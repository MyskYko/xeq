//
// Conformal-LEC Version 20.10-d132 (30-Jun-2020)
//
module top(RIc0c7950_66,RIc0c9750_2,RIc0c96d8_3,RIc0c9660_4,RIc0c78d8_67,RIc0c95e8_5,RIc0c9570_6,RIc0c7860_68,RIc0c77e8_69,
        RIc0c94f8_7,RIc0c9480_8,RIc0c7770_70,RIc0c76f8_71,RIc0c9408_9,RIc0c9390_10,RIc0c7680_72,RIc0c7608_73,RIc0c9318_11,RIc0c92a0_12,
        RIc0c7590_74,RIc0c7518_75,RIc0c9228_13,RIc0c91b0_14,RIc0c74a0_76,RIc0c7428_77,RIc0c9138_15,RIc0c90c0_16,RIc0c73b0_78,RIc0c7338_79,
        RIc0c9048_17,RIc0c8fd0_18,RIc0c72c0_80,RIc0c7248_81,RIc0c8f58_19,RIc0c8ee0_20,RIc0c71d0_82,RIc0c8e68_21,RIc0c8df0_22,RIc0c7158_83,
        RIc0c70e0_84,RIc0c7068_85,RIc0c8d78_23,RIc0c8d00_24,RIc0c6ff0_86,RIc0c6f78_87,RIc0c8c88_25,RIc0c8c10_26,RIc0c6f00_88,RIc0c6e88_89,
        RIc0c8b98_27,RIc0c8b20_28,RIc0c6e10_90,RIc0c6d98_91,RIc0c8aa8_29,RIc0c8a30_30,RIc0c6d20_92,RIc0c6ca8_93,RIc0c89b8_31,RIc0c8940_32,
        RIc0c6c30_94,RIc0c6bb8_95,RIc0c88c8_33,RIc0c8850_34,RIc0c6b40_96,RIc0c6ac8_97,RIc0c87d8_35,RIc0c8760_36,RIc0c6a50_98,RIc0c69d8_99,
        RIc0c86e8_37,RIc0c8670_38,RIc0c6960_100,RIc0c85f8_39,RIc0c8580_40,RIc0c68e8_101,RIc0c6870_102,RIc0c67f8_103,RIc0c8508_41,RIc0c8490_42,
        RIc0c6780_104,RIc0c6708_105,RIc0c8418_43,RIc0c83a0_44,RIc0c6690_106,RIc0c6618_107,RIc0c8328_45,RIc0c82b0_46,RIc0c65a0_108,RIc0c6528_109,
        RIc0c8238_47,RIc0c81c0_48,RIc0c64b0_110,RIc0c6438_111,RIc0c8148_49,RIc0c80d0_50,RIc0c63c0_112,RIc0c6348_113,RIc0c8058_51,RIc0c7fe0_52,
        RIc0c62d0_114,RIc0c6258_115,RIc0c7f68_53,RIc0c7ef0_54,RIc0c61e0_116,RIc0c6168_117,RIc0c7e78_55,RIc0c7e00_56,RIc0c60f0_118,RIc0c7d88_57,
        RIc0c7d10_58,RIc0c6078_119,RIc0c6000_120,RIc0c5f88_121,RIc0c7c98_59,RIc0c7c20_60,RIc0c5f10_122,RIc0c5e98_123,RIc0c7ba8_61,RIc0c7b30_62,
        RIc0c5e20_124,RIc0c5da8_125,RIc0c7ab8_63,RIc0c7a40_64,RIc0c5d30_126,RIc340530_127,RIc3405a8_128,RIc0c79c8_65,RIc340620_129,RIc340698_130,
        RIc340710_131,RIc340788_132,RIc340800_133,RIc340878_134,RIc3408f0_135,RIc340968_136,RIc3409e0_137,RIc340a58_138,RIc340ad0_139,RIc340b48_140,
        RIc340bc0_141,RIc340c38_142,RIc340cb0_143,RIc340d28_144,RIc340da0_145,RIc340e18_146,RIc340e90_147,RIc340f08_148,RIc340f80_149,RIc340ff8_150,
        RIc341070_151,RIc3410e8_152,RIc341160_153,RIc3411d8_154,RIc341250_155,RIc3412c8_156,RIc341340_157,RIc3413b8_158,RIc341430_159,RIc3414a8_160,
        RIc341520_161,RIc341598_162,RIc341610_163,RIc341688_164,RIc341700_165,RIc341778_166,RIc3417f0_167,RIc341868_168,RIc3418e0_169,RIc341958_170,
        RIc3419d0_171,RIc341a48_172,RIc341ac0_173,RIc341b38_174,RIc341bb0_175,RIc341c28_176,RIc341ca0_177,RIc341d18_178,RIc341d90_179,RIc341e08_180,
        RIc341e80_181,RIc341ef8_182,RIc341f70_183,RIc341fe8_184,RIc342060_185,RIc3420d8_186,RIc342150_187,RIc3421c8_188,RIc342240_189,RIc3422b8_190,
        RIc342330_191,RIc3423a8_192,RIc342420_193,RIc0c97c8_1,R_c2_9969708,R_c3_99697b0,R_c4_9969858,R_c5_9969900,R_c6_99699a8,R_c7_9969a50,
        R_c8_9969af8,R_c9_9969ba0,R_ca_9969c48,R_cb_9969cf0,R_cc_9969d98,R_cd_9969e40,R_ce_9969ee8,R_cf_9969f90,R_d0_996a038,R_d1_996a0e0,
        R_d2_996a188,R_d3_996a230,R_d4_996a2d8,R_d5_996a380,R_d6_996a428,R_d7_996a4d0,R_d8_996a578,R_d9_996a620,R_da_996a6c8,R_db_996a770,
        R_dc_996a818,R_dd_996a8c0,R_de_996a968,R_df_996aa10,R_e0_996aab8,R_e1_996ab60,R_e2_996ac08,R_e3_996acb0,R_e4_996ad58,R_e5_996ae00,
        R_e6_996aea8,R_e7_996af50,R_e8_996aff8,R_e9_996b0a0,R_ea_996b148,R_eb_996b1f0,R_ec_996b298,R_ed_996b340,R_ee_996b3e8,R_ef_996b490,
        R_f0_996b538,R_f1_996b5e0,R_f2_996b688,R_f3_996b730,R_f4_996b7d8,R_f5_996b880,R_f6_996b928,R_f7_996b9d0,R_f8_996ba78,R_f9_996bb20,
        R_fa_996bbc8,R_fb_996bc70,R_fc_996bd18,R_fd_996bdc0,R_fe_996be68,R_ff_996bf10,R_100_996bfb8,R_101_996c060,R_102_996c108,R_103_996c1b0,
        R_104_996c258,R_105_996c300,R_106_996c3a8,R_107_996c450,R_108_996c4f8,R_109_996c5a0,R_10a_996c648,R_10b_996c6f0,R_10c_996c798,R_10d_996c840,
        R_10e_996c8e8,R_10f_996c990,R_110_996ca38,R_111_996cae0,R_112_996cb88,R_113_996cc30,R_114_996ccd8,R_115_996cd80,R_116_996ce28,R_117_996ced0,
        R_118_996cf78,R_119_996d020,R_11a_996d0c8,R_11b_996d170,R_11c_996d218,R_11d_996d2c0,R_11e_996d368,R_11f_996d410,R_120_996d4b8,R_121_996d560,
        R_122_996d608,R_123_996d6b0,R_124_996d758,R_125_996d800,R_126_996d8a8,R_127_996d950,R_128_996d9f8,R_129_996daa0,R_12a_996db48,R_12b_996dbf0,
        R_12c_996dc98,R_12d_996dd40,R_12e_996dde8,R_12f_996de90,R_130_996df38,R_131_996dfe0,R_132_996e088,R_133_996e130,R_134_996e1d8,R_135_996e280,
        R_136_996e328,R_137_996e3d0,R_138_996e478,R_139_996e520);
input RIc0c7950_66,RIc0c9750_2,RIc0c96d8_3,RIc0c9660_4,RIc0c78d8_67,RIc0c95e8_5,RIc0c9570_6,RIc0c7860_68,RIc0c77e8_69,
        RIc0c94f8_7,RIc0c9480_8,RIc0c7770_70,RIc0c76f8_71,RIc0c9408_9,RIc0c9390_10,RIc0c7680_72,RIc0c7608_73,RIc0c9318_11,RIc0c92a0_12,
        RIc0c7590_74,RIc0c7518_75,RIc0c9228_13,RIc0c91b0_14,RIc0c74a0_76,RIc0c7428_77,RIc0c9138_15,RIc0c90c0_16,RIc0c73b0_78,RIc0c7338_79,
        RIc0c9048_17,RIc0c8fd0_18,RIc0c72c0_80,RIc0c7248_81,RIc0c8f58_19,RIc0c8ee0_20,RIc0c71d0_82,RIc0c8e68_21,RIc0c8df0_22,RIc0c7158_83,
        RIc0c70e0_84,RIc0c7068_85,RIc0c8d78_23,RIc0c8d00_24,RIc0c6ff0_86,RIc0c6f78_87,RIc0c8c88_25,RIc0c8c10_26,RIc0c6f00_88,RIc0c6e88_89,
        RIc0c8b98_27,RIc0c8b20_28,RIc0c6e10_90,RIc0c6d98_91,RIc0c8aa8_29,RIc0c8a30_30,RIc0c6d20_92,RIc0c6ca8_93,RIc0c89b8_31,RIc0c8940_32,
        RIc0c6c30_94,RIc0c6bb8_95,RIc0c88c8_33,RIc0c8850_34,RIc0c6b40_96,RIc0c6ac8_97,RIc0c87d8_35,RIc0c8760_36,RIc0c6a50_98,RIc0c69d8_99,
        RIc0c86e8_37,RIc0c8670_38,RIc0c6960_100,RIc0c85f8_39,RIc0c8580_40,RIc0c68e8_101,RIc0c6870_102,RIc0c67f8_103,RIc0c8508_41,RIc0c8490_42,
        RIc0c6780_104,RIc0c6708_105,RIc0c8418_43,RIc0c83a0_44,RIc0c6690_106,RIc0c6618_107,RIc0c8328_45,RIc0c82b0_46,RIc0c65a0_108,RIc0c6528_109,
        RIc0c8238_47,RIc0c81c0_48,RIc0c64b0_110,RIc0c6438_111,RIc0c8148_49,RIc0c80d0_50,RIc0c63c0_112,RIc0c6348_113,RIc0c8058_51,RIc0c7fe0_52,
        RIc0c62d0_114,RIc0c6258_115,RIc0c7f68_53,RIc0c7ef0_54,RIc0c61e0_116,RIc0c6168_117,RIc0c7e78_55,RIc0c7e00_56,RIc0c60f0_118,RIc0c7d88_57,
        RIc0c7d10_58,RIc0c6078_119,RIc0c6000_120,RIc0c5f88_121,RIc0c7c98_59,RIc0c7c20_60,RIc0c5f10_122,RIc0c5e98_123,RIc0c7ba8_61,RIc0c7b30_62,
        RIc0c5e20_124,RIc0c5da8_125,RIc0c7ab8_63,RIc0c7a40_64,RIc0c5d30_126,RIc340530_127,RIc3405a8_128,RIc0c79c8_65,RIc340620_129,RIc340698_130,
        RIc340710_131,RIc340788_132,RIc340800_133,RIc340878_134,RIc3408f0_135,RIc340968_136,RIc3409e0_137,RIc340a58_138,RIc340ad0_139,RIc340b48_140,
        RIc340bc0_141,RIc340c38_142,RIc340cb0_143,RIc340d28_144,RIc340da0_145,RIc340e18_146,RIc340e90_147,RIc340f08_148,RIc340f80_149,RIc340ff8_150,
        RIc341070_151,RIc3410e8_152,RIc341160_153,RIc3411d8_154,RIc341250_155,RIc3412c8_156,RIc341340_157,RIc3413b8_158,RIc341430_159,RIc3414a8_160,
        RIc341520_161,RIc341598_162,RIc341610_163,RIc341688_164,RIc341700_165,RIc341778_166,RIc3417f0_167,RIc341868_168,RIc3418e0_169,RIc341958_170,
        RIc3419d0_171,RIc341a48_172,RIc341ac0_173,RIc341b38_174,RIc341bb0_175,RIc341c28_176,RIc341ca0_177,RIc341d18_178,RIc341d90_179,RIc341e08_180,
        RIc341e80_181,RIc341ef8_182,RIc341f70_183,RIc341fe8_184,RIc342060_185,RIc3420d8_186,RIc342150_187,RIc3421c8_188,RIc342240_189,RIc3422b8_190,
        RIc342330_191,RIc3423a8_192,RIc342420_193,RIc0c97c8_1;
output R_c2_9969708,R_c3_99697b0,R_c4_9969858,R_c5_9969900,R_c6_99699a8,R_c7_9969a50,R_c8_9969af8,R_c9_9969ba0,R_ca_9969c48,
        R_cb_9969cf0,R_cc_9969d98,R_cd_9969e40,R_ce_9969ee8,R_cf_9969f90,R_d0_996a038,R_d1_996a0e0,R_d2_996a188,R_d3_996a230,R_d4_996a2d8,
        R_d5_996a380,R_d6_996a428,R_d7_996a4d0,R_d8_996a578,R_d9_996a620,R_da_996a6c8,R_db_996a770,R_dc_996a818,R_dd_996a8c0,R_de_996a968,
        R_df_996aa10,R_e0_996aab8,R_e1_996ab60,R_e2_996ac08,R_e3_996acb0,R_e4_996ad58,R_e5_996ae00,R_e6_996aea8,R_e7_996af50,R_e8_996aff8,
        R_e9_996b0a0,R_ea_996b148,R_eb_996b1f0,R_ec_996b298,R_ed_996b340,R_ee_996b3e8,R_ef_996b490,R_f0_996b538,R_f1_996b5e0,R_f2_996b688,
        R_f3_996b730,R_f4_996b7d8,R_f5_996b880,R_f6_996b928,R_f7_996b9d0,R_f8_996ba78,R_f9_996bb20,R_fa_996bbc8,R_fb_996bc70,R_fc_996bd18,
        R_fd_996bdc0,R_fe_996be68,R_ff_996bf10,R_100_996bfb8,R_101_996c060,R_102_996c108,R_103_996c1b0,R_104_996c258,R_105_996c300,R_106_996c3a8,
        R_107_996c450,R_108_996c4f8,R_109_996c5a0,R_10a_996c648,R_10b_996c6f0,R_10c_996c798,R_10d_996c840,R_10e_996c8e8,R_10f_996c990,R_110_996ca38,
        R_111_996cae0,R_112_996cb88,R_113_996cc30,R_114_996ccd8,R_115_996cd80,R_116_996ce28,R_117_996ced0,R_118_996cf78,R_119_996d020,R_11a_996d0c8,
        R_11b_996d170,R_11c_996d218,R_11d_996d2c0,R_11e_996d368,R_11f_996d410,R_120_996d4b8,R_121_996d560,R_122_996d608,R_123_996d6b0,R_124_996d758,
        R_125_996d800,R_126_996d8a8,R_127_996d950,R_128_996d9f8,R_129_996daa0,R_12a_996db48,R_12b_996dbf0,R_12c_996dc98,R_12d_996dd40,R_12e_996dde8,
        R_12f_996de90,R_130_996df38,R_131_996dfe0,R_132_996e088,R_133_996e130,R_134_996e1d8,R_135_996e280,R_136_996e328,R_137_996e3d0,R_138_996e478,
        R_139_996e520;

wire \314_ZERO , \315_ONE , \316 , \317 , \318 , \319 , \320 , \321 , \322 ,
         \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 ,
         \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 ,
         \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 ,
         \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 ,
         \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 ,
         \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 ,
         \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 ,
         \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 ,
         \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 ,
         \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 ,
         \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 ,
         \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 ,
         \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 ,
         \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 ,
         \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 ,
         \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 ,
         \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 ,
         \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 ,
         \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 ,
         \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 ,
         \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 ,
         \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 ,
         \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 ,
         \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 ,
         \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 ,
         \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 ,
         \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 ,
         \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 ,
         \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 ,
         \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 ,
         \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 ,
         \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 ,
         \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 ,
         \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 ,
         \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 ,
         \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 ,
         \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 ,
         \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 ,
         \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 ,
         \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 ,
         \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 ,
         \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 ,
         \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 ,
         \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 ,
         \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 ,
         \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 ,
         \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 ,
         \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 ,
         \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 ,
         \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 ,
         \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 ,
         \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 ,
         \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 ,
         \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 ,
         \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 ,
         \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 ,
         \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 ,
         \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 ,
         \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 ,
         \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 ,
         \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 ,
         \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 ,
         \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 ,
         \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 ,
         \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 ,
         \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 ,
         \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 ,
         \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 ,
         \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 ,
         \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 ,
         \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 ,
         \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 ,
         \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 ,
         \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 ,
         \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 ,
         \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 ,
         \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 ,
         \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 ,
         \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 ,
         \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 ,
         \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 ,
         \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 ,
         \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 ,
         \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 ,
         \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 ,
         \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 ,
         \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 ,
         \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 ,
         \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 ,
         \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 ,
         \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 ,
         \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 ,
         \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 ,
         \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 ,
         \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 ,
         \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 ,
         \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 ,
         \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 ,
         \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 ,
         \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 ,
         \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 ,
         \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 ,
         \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 ,
         \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 ,
         \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 ,
         \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 ,
         \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 ,
         \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 ,
         \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 ,
         \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 ,
         \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 ,
         \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 ,
         \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 ,
         \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 ,
         \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 ,
         \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 ,
         \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 ,
         \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 ,
         \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 ,
         \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 ,
         \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 ,
         \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 ,
         \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 ,
         \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 ,
         \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 ,
         \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 ,
         \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 ,
         \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 ,
         \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 ,
         \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 ,
         \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 ,
         \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 ,
         \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 ,
         \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 ,
         \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 ,
         \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 ,
         \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 ,
         \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 ,
         \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 ,
         \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 ,
         \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 ,
         \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 ,
         \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 ,
         \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 ,
         \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 ,
         \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 ,
         \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 ,
         \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 ,
         \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 ,
         \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 ,
         \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 ,
         \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 ,
         \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 ,
         \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 ,
         \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 ,
         \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 ,
         \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 ,
         \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 ,
         \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 ,
         \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 ,
         \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 ,
         \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 ,
         \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 ,
         \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 ,
         \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 ,
         \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 ,
         \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 ,
         \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 ,
         \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 ,
         \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 ,
         \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 ,
         \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 ,
         \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 ,
         \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 ,
         \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 ,
         \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 ,
         \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 ,
         \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 ,
         \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 ,
         \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 ,
         \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 ,
         \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 ,
         \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 ,
         \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 ,
         \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 ,
         \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 ,
         \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 ,
         \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 ,
         \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 ,
         \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 ,
         \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 ,
         \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 ,
         \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 ,
         \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 ,
         \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 ,
         \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 ,
         \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 ,
         \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 ,
         \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 ,
         \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 ,
         \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 ,
         \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 ,
         \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 ,
         \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 ,
         \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 ,
         \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 ,
         \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 ,
         \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 ,
         \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 ,
         \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 ,
         \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 ,
         \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 ,
         \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 ,
         \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 ,
         \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 ,
         \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 ,
         \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 ,
         \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 ,
         \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 ,
         \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 ,
         \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 ,
         \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 ,
         \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 ,
         \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 ,
         \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 ,
         \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 ,
         \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 ,
         \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 ,
         \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 ,
         \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 ,
         \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 ,
         \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 ,
         \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 ,
         \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 ,
         \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 ,
         \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 ,
         \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 ,
         \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 ,
         \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 ,
         \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 ,
         \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 ,
         \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 ,
         \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 ,
         \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 ,
         \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 ,
         \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 ,
         \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 ,
         \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 ,
         \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 ,
         \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 ,
         \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 ,
         \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 ,
         \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 ,
         \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 ,
         \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 ,
         \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 ,
         \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 ,
         \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 ,
         \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 ,
         \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 ,
         \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 ,
         \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 ,
         \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 ,
         \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 ,
         \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 ,
         \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 ,
         \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 ,
         \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 ,
         \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 ,
         \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 ,
         \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 ,
         \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 ,
         \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 ,
         \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 ,
         \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 ,
         \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 ,
         \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 ,
         \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 ,
         \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 ,
         \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 ,
         \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 ,
         \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 ,
         \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 ,
         \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 ,
         \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 ,
         \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 ,
         \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 ,
         \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 ,
         \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 ,
         \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 ,
         \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 ,
         \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 ,
         \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 ,
         \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 ,
         \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 ,
         \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 ,
         \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 ,
         \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 ,
         \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 ,
         \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 ,
         \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 ,
         \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 ,
         \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 ,
         \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 ,
         \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 ,
         \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 ,
         \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 ,
         \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 ,
         \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 ,
         \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 ,
         \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 ,
         \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 ,
         \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 ,
         \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 ,
         \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 ,
         \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 ,
         \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 ,
         \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 ,
         \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 ,
         \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 ,
         \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 ,
         \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 ,
         \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 ,
         \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 ,
         \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 ,
         \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 ,
         \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 ,
         \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 ,
         \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 ,
         \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 ,
         \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 ,
         \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 ,
         \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 ,
         \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 ,
         \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 ,
         \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 ,
         \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 ,
         \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 ,
         \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 ,
         \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 ,
         \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 ,
         \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 ,
         \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 ,
         \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 ,
         \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 ,
         \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 ,
         \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 ,
         \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 ,
         \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 ,
         \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 ,
         \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 ,
         \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 ,
         \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 ,
         \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 ,
         \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 ,
         \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 ,
         \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 ,
         \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 ,
         \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 ,
         \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 ,
         \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 ,
         \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 ,
         \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 ,
         \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 ,
         \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 ,
         \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 ,
         \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 ,
         \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 ,
         \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 ,
         \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 ,
         \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 ,
         \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 ,
         \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 ,
         \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 ,
         \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 ,
         \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 ,
         \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 ,
         \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 ,
         \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 ,
         \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 ,
         \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 ,
         \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 ,
         \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 ,
         \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 ,
         \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 ,
         \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 ,
         \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 ,
         \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 ,
         \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 ,
         \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 ,
         \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 ,
         \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 ,
         \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 ,
         \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 ,
         \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 ,
         \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 ,
         \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 ,
         \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 ,
         \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 ,
         \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 ,
         \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 ,
         \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 ,
         \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 ,
         \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 ,
         \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 ,
         \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 ,
         \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 ,
         \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 ,
         \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 ,
         \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 ,
         \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 ,
         \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 ,
         \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 ,
         \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 ,
         \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 ,
         \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 ,
         \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 ,
         \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 ,
         \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 ,
         \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 ,
         \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 ,
         \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 ,
         \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 ,
         \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 ,
         \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 ,
         \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 ,
         \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 ,
         \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 ,
         \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 ,
         \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 ,
         \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 ,
         \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 ,
         \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 ,
         \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 ,
         \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 ,
         \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 ,
         \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 ,
         \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 ,
         \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 ,
         \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 ,
         \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 ,
         \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 ,
         \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 ,
         \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 ,
         \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 ,
         \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 ,
         \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 ,
         \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 ,
         \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 ,
         \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 ,
         \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 ,
         \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 ,
         \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 ,
         \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 ,
         \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 ,
         \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 ,
         \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 ,
         \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 ,
         \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 ,
         \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 ,
         \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 ,
         \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 ,
         \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 ,
         \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 ,
         \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 ,
         \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 ,
         \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 ,
         \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 ,
         \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 ,
         \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 ,
         \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 ,
         \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 ,
         \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 ,
         \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 ,
         \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 ,
         \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 ,
         \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 ,
         \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 ,
         \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 ,
         \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 ,
         \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 ,
         \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 ,
         \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 ,
         \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 ,
         \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 ,
         \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 ,
         \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 ,
         \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 ,
         \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 ,
         \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 ,
         \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 ,
         \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 ,
         \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 ,
         \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 ,
         \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 ,
         \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 ,
         \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 ,
         \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 ,
         \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 ,
         \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 ,
         \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 ,
         \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 ,
         \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 ,
         \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 ,
         \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 ,
         \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 ,
         \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 ,
         \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 ,
         \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 ,
         \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 ,
         \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 ,
         \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 ,
         \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 ,
         \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 ,
         \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 ,
         \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 ,
         \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 ,
         \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 ,
         \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 ,
         \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 ,
         \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 ,
         \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 ,
         \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 ,
         \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 ,
         \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 ,
         \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 ,
         \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 ,
         \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 ,
         \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 ,
         \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 ,
         \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 ,
         \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 ,
         \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 ,
         \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 ,
         \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 ,
         \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 ,
         \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 ,
         \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 ,
         \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 ,
         \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 ,
         \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 ,
         \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 ,
         \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 ,
         \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 ,
         \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 ,
         \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 ,
         \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 ,
         \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 ,
         \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 ,
         \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 ,
         \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 ,
         \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 ,
         \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 ,
         \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 ,
         \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 ,
         \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 ,
         \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 ,
         \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 ,
         \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 ,
         \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 ,
         \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 ,
         \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 ,
         \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 ,
         \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 ,
         \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 ,
         \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 ,
         \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 ,
         \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 ,
         \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 ,
         \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 ,
         \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 ,
         \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 ,
         \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 ,
         \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 ,
         \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 ,
         \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 ,
         \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 ,
         \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 ,
         \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 ,
         \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 ,
         \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 ,
         \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 ,
         \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 ,
         \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 ,
         \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 ,
         \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 ,
         \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 ,
         \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 ,
         \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 ,
         \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 ,
         \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 ,
         \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 ,
         \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 ,
         \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 ,
         \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 ,
         \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 ,
         \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 ,
         \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 ,
         \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 ,
         \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 ,
         \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 ,
         \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 ,
         \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 ,
         \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 ,
         \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 ,
         \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 ,
         \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 ,
         \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 ,
         \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 ,
         \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 ,
         \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 ,
         \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 ,
         \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 ,
         \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 ,
         \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 ,
         \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 ,
         \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 ,
         \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 ,
         \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 ,
         \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 ,
         \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 ,
         \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 ,
         \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 ,
         \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 ,
         \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 ,
         \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 ,
         \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 ,
         \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 ,
         \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 ,
         \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 ,
         \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 ,
         \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 ,
         \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 ,
         \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 ,
         \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 ,
         \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 ,
         \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 ,
         \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 ,
         \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 ,
         \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 ,
         \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 ,
         \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 ,
         \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 ,
         \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 ,
         \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 ,
         \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 ,
         \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 ,
         \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 ,
         \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 ,
         \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 ,
         \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 ,
         \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 ,
         \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 ,
         \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 ,
         \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 ,
         \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 ,
         \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 ,
         \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 ,
         \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 ,
         \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 ,
         \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 ,
         \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 ,
         \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 ,
         \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 ,
         \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 ,
         \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 ,
         \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 ,
         \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 ,
         \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 ,
         \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 ,
         \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 ,
         \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 ,
         \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 ,
         \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 ,
         \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 ,
         \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 ,
         \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 ,
         \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 ,
         \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 ,
         \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 ,
         \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 ,
         \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 ,
         \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 ,
         \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 ,
         \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 ,
         \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 ,
         \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 ,
         \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 ,
         \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 ,
         \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 ,
         \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 ,
         \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 ,
         \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 ,
         \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 ,
         \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 ,
         \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 ,
         \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 ,
         \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 ,
         \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 ,
         \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 ,
         \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 ,
         \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 ,
         \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 ,
         \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 ,
         \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 ,
         \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 ,
         \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 ,
         \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 ,
         \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 ,
         \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 ,
         \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 ,
         \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 ,
         \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 ,
         \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 ,
         \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 ,
         \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 ,
         \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 ,
         \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 ,
         \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 ,
         \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 ,
         \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 ,
         \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 ,
         \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 ,
         \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 ,
         \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 ,
         \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 ,
         \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 ,
         \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 ,
         \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 ,
         \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 ,
         \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 ,
         \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 ,
         \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 ,
         \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 ,
         \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 ,
         \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 ,
         \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 ,
         \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 ,
         \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 ,
         \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 ,
         \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 ,
         \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 ,
         \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 ,
         \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 ,
         \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 ,
         \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 ,
         \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 ,
         \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 ,
         \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 ,
         \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 ,
         \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 ,
         \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 ,
         \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 ,
         \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 ,
         \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 ,
         \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 ,
         \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 ,
         \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 ,
         \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 ,
         \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 ,
         \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 ,
         \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 ,
         \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 ,
         \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 ,
         \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 ,
         \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 ,
         \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 ,
         \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 ,
         \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 ,
         \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 ,
         \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 ,
         \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 ,
         \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 ,
         \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 ,
         \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 ,
         \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 ,
         \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 ,
         \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 ,
         \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 ,
         \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 ,
         \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 ,
         \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 ,
         \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 ,
         \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 ,
         \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 ,
         \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 ,
         \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 ,
         \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 ,
         \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 ,
         \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 ,
         \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 ,
         \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 ,
         \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 ,
         \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 ,
         \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 ,
         \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 ,
         \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 ,
         \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 ,
         \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 ,
         \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 ,
         \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 ,
         \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 ,
         \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 ,
         \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 ,
         \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 ,
         \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 ,
         \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 ,
         \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 ,
         \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 ,
         \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 ,
         \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 ,
         \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 ,
         \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 ,
         \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 ,
         \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 ,
         \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 ,
         \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 ,
         \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 ,
         \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 ,
         \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 ,
         \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 ,
         \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 ,
         \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 ,
         \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 ,
         \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 ,
         \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 ,
         \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 ,
         \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 ,
         \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 ,
         \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 ,
         \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 ,
         \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 ,
         \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 ,
         \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 ,
         \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 ,
         \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 ,
         \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 ,
         \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 ,
         \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 ,
         \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 ,
         \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 ,
         \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 ,
         \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 ,
         \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 ,
         \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 ,
         \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 ,
         \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 ,
         \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 ,
         \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 ,
         \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 ,
         \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 ,
         \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 ,
         \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 ,
         \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 ,
         \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 ,
         \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 ,
         \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 ,
         \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 ,
         \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 ,
         \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 ,
         \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 ,
         \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 ,
         \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 ,
         \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 ,
         \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 ,
         \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 ,
         \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 ,
         \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 ,
         \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 ,
         \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 ,
         \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 ,
         \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 ,
         \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 ,
         \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 ,
         \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 ,
         \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 ,
         \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 ,
         \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 ,
         \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 ,
         \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 ,
         \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 ,
         \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 ,
         \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 ,
         \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 ,
         \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 ,
         \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 ,
         \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 ,
         \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 ,
         \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 ,
         \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 ,
         \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 ,
         \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 ,
         \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 ,
         \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 ,
         \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 ,
         \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 ,
         \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 ,
         \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 ,
         \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 ,
         \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 ,
         \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 ,
         \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 ,
         \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 ,
         \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 ,
         \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 ,
         \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 ,
         \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 ,
         \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 ,
         \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 ,
         \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 ,
         \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 ,
         \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 ,
         \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 ,
         \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 ,
         \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 ,
         \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 ,
         \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 ,
         \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 ,
         \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 ,
         \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 ,
         \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 ,
         \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 ,
         \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 ,
         \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 ,
         \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 ,
         \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 ,
         \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 ,
         \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 ,
         \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 ,
         \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 ,
         \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 ,
         \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 ,
         \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 ,
         \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 ,
         \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 ,
         \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 ,
         \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 ,
         \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 ,
         \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 ,
         \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 ,
         \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 ,
         \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 ,
         \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 ,
         \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 ,
         \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 ,
         \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 ,
         \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 ,
         \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 ,
         \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 ,
         \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 ,
         \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 ,
         \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 ,
         \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 ,
         \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 ,
         \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 ,
         \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 ,
         \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 ,
         \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 ,
         \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 ,
         \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 ,
         \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 ,
         \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 ,
         \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 ,
         \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 ,
         \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 ,
         \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 ,
         \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 ,
         \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 ,
         \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 ,
         \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 ,
         \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 ,
         \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 ,
         \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 ,
         \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 ,
         \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 ,
         \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 ,
         \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 ,
         \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 ,
         \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 ,
         \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 ,
         \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 ,
         \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 ,
         \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 ,
         \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 ,
         \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 ,
         \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 ,
         \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 ,
         \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 ,
         \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 ,
         \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 ,
         \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 ,
         \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 ,
         \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 ,
         \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 ,
         \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 ,
         \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 ,
         \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 ,
         \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 ,
         \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 ,
         \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 ,
         \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 ,
         \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 ,
         \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 ,
         \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 ,
         \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 ,
         \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 ,
         \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 ,
         \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 ,
         \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 ,
         \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 ,
         \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 ,
         \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 ,
         \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 ,
         \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 ,
         \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 ,
         \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 ,
         \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 ,
         \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 ,
         \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 ,
         \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 ,
         \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 ,
         \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 ,
         \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 ,
         \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 ,
         \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 ,
         \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 ,
         \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 ,
         \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 ,
         \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 ,
         \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 ,
         \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 ,
         \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 ,
         \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 ,
         \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 ,
         \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 ,
         \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 ,
         \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 ,
         \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 ,
         \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 ,
         \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 ,
         \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 ,
         \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 ,
         \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 ,
         \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 ,
         \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 ,
         \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 ,
         \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 ,
         \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 ,
         \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 ,
         \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 ,
         \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 ,
         \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 ,
         \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 ,
         \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 ,
         \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 ,
         \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 ,
         \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 ,
         \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 ,
         \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 ,
         \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 ,
         \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 ,
         \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 ,
         \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 ,
         \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 ,
         \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 ,
         \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 ,
         \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 ,
         \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 ,
         \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 ,
         \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 ,
         \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 ,
         \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 ,
         \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 ,
         \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 ,
         \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 ,
         \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 ,
         \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 ,
         \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 ,
         \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 ,
         \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 ,
         \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 ,
         \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 ,
         \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 ,
         \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 ,
         \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 ,
         \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 ,
         \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 ,
         \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 ,
         \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 ,
         \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 ,
         \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 ,
         \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 ,
         \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 ,
         \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 ,
         \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 ,
         \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 ,
         \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 ,
         \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 ,
         \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 ,
         \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 ,
         \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 ,
         \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 ,
         \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 ,
         \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 ,
         \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 ,
         \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 ,
         \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 ,
         \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 ,
         \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 ,
         \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 ,
         \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 ,
         \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 ,
         \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 ,
         \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 ,
         \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 ,
         \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 ,
         \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 ,
         \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 ,
         \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 ,
         \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 ,
         \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 ,
         \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 ,
         \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 ,
         \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 ,
         \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 ,
         \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 ,
         \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 ,
         \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 ,
         \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 ,
         \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 ,
         \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 ,
         \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 ,
         \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 ,
         \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 ,
         \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 ,
         \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 ,
         \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 ,
         \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 ,
         \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 ,
         \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 ,
         \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 ,
         \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 ,
         \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 ,
         \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 ,
         \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 ,
         \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 ,
         \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 ,
         \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 ,
         \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 ,
         \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 ,
         \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 ,
         \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 ,
         \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 ,
         \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 ,
         \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 ,
         \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 ,
         \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 ,
         \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 ,
         \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 ,
         \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 ,
         \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 ,
         \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 ,
         \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 ,
         \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 ,
         \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 ,
         \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 ,
         \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 ,
         \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 ,
         \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 ,
         \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 ,
         \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 ,
         \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 ,
         \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 ,
         \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 ,
         \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 ,
         \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 ,
         \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 ,
         \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 ,
         \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 ,
         \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 ,
         \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 ,
         \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 ,
         \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 ,
         \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 ,
         \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 ,
         \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 ,
         \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 ,
         \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 ,
         \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 ,
         \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 ,
         \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 ,
         \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 ,
         \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 ,
         \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 ,
         \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 ,
         \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 ,
         \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 ,
         \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 ,
         \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 ,
         \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 ,
         \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 ,
         \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 ,
         \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 ,
         \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 ,
         \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 ,
         \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 ,
         \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 ,
         \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 ,
         \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 ,
         \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 ,
         \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 ,
         \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 ,
         \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 ,
         \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 ,
         \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 ,
         \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 ,
         \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 ,
         \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 ,
         \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 ,
         \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 ,
         \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 ,
         \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 ,
         \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 ,
         \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 ,
         \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 ,
         \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 ,
         \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 ,
         \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 ,
         \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 ,
         \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 ,
         \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 ,
         \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 ,
         \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 ,
         \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 ,
         \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 ,
         \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 ,
         \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 ,
         \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 ,
         \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 ,
         \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 ,
         \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 ,
         \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 ,
         \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 ,
         \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 ,
         \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 ,
         \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 ,
         \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 ,
         \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 ,
         \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 ,
         \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 ,
         \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 ,
         \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 ,
         \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 ,
         \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 ,
         \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 ,
         \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 ,
         \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 ,
         \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 ,
         \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 ,
         \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 ,
         \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 ,
         \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 ,
         \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 ,
         \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 ,
         \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 ,
         \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 ,
         \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 ,
         \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 ,
         \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 ,
         \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 ,
         \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 ,
         \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 ,
         \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 ,
         \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 ,
         \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 ,
         \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 ,
         \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 ,
         \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 ,
         \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 ,
         \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 ,
         \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 ,
         \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 ,
         \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 ,
         \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 ,
         \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 ,
         \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 ,
         \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 ,
         \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 ,
         \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 ,
         \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 ,
         \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 ,
         \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 ,
         \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 ,
         \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 ,
         \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 ,
         \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 ,
         \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 ,
         \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 ,
         \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 ,
         \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 ,
         \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 ,
         \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 ,
         \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 ,
         \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 ,
         \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 ,
         \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 ,
         \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 ,
         \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 ,
         \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 ,
         \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 ,
         \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 ,
         \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 ,
         \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 ,
         \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 ,
         \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 ,
         \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 ,
         \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 ,
         \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 ,
         \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 ,
         \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 ,
         \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 ,
         \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 ,
         \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 ,
         \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 ,
         \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 ,
         \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 ,
         \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 ,
         \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 ,
         \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 ,
         \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 ,
         \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 ,
         \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 ,
         \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 ,
         \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 ,
         \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 ,
         \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 ,
         \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 ,
         \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 ,
         \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 ,
         \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 ,
         \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 ,
         \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 ,
         \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 ,
         \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 ,
         \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 ,
         \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 ,
         \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 ,
         \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 ,
         \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 ,
         \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 ,
         \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 ,
         \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 ,
         \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 ,
         \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 ,
         \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 ,
         \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 ,
         \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 ,
         \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 ,
         \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 ,
         \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 ,
         \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 ,
         \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 ,
         \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 ,
         \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 ,
         \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 ,
         \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 ,
         \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 ,
         \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 ,
         \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 ,
         \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 ,
         \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 ,
         \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 ,
         \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 ,
         \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 ,
         \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 ,
         \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 ,
         \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 ,
         \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 ,
         \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 ,
         \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 ,
         \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 ,
         \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 ,
         \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 ,
         \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 ,
         \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 ,
         \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 ,
         \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 ,
         \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 ,
         \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 ,
         \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 ,
         \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 ,
         \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 ,
         \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 ,
         \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 ,
         \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 ,
         \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 ,
         \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 ,
         \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 ,
         \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 ,
         \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 ,
         \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 ,
         \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 ,
         \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 ,
         \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 ,
         \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 ,
         \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 ,
         \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 ,
         \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 ,
         \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 ,
         \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 ,
         \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 ,
         \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 ,
         \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 ,
         \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 ,
         \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 ,
         \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 ,
         \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 ,
         \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 ,
         \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 ,
         \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 ,
         \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 ,
         \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 ,
         \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 ,
         \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 ,
         \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 ,
         \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 ,
         \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 ,
         \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 ,
         \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 ,
         \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 ,
         \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 ,
         \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 ,
         \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 ,
         \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 ,
         \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 ,
         \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 ,
         \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 ,
         \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 ,
         \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 ,
         \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 ,
         \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 ,
         \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 ,
         \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 ,
         \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 ,
         \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 ,
         \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 ,
         \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 ,
         \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 ,
         \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 ,
         \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 ,
         \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 ,
         \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 ,
         \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 ,
         \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 ,
         \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 ,
         \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 ,
         \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 ,
         \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 ,
         \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 ,
         \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 ,
         \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 ,
         \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 ,
         \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 ,
         \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 ,
         \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 ,
         \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 ,
         \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 ,
         \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 ,
         \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 ,
         \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 ,
         \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 ,
         \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 ,
         \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 ,
         \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 ,
         \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 ,
         \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 ,
         \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 ,
         \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 ,
         \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 ,
         \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 ,
         \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 ,
         \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 ,
         \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 ,
         \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 ,
         \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 ,
         \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 ,
         \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 ,
         \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 ,
         \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 ,
         \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 ,
         \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 ,
         \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 ,
         \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 ,
         \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 ,
         \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 ,
         \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 ,
         \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 ,
         \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 ,
         \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 ,
         \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 ,
         \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 ,
         \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 ,
         \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 ,
         \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 ,
         \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 ,
         \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 ,
         \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 ,
         \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 ,
         \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 ,
         \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 ,
         \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 ,
         \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 ,
         \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 ,
         \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 ,
         \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 ,
         \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 ,
         \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 ,
         \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 ,
         \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 ,
         \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 ,
         \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 ,
         \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 ,
         \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 ,
         \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 ,
         \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 ,
         \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 ,
         \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 ,
         \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 ,
         \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 ,
         \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 ,
         \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 ,
         \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 ,
         \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 ,
         \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 ,
         \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 ,
         \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 ,
         \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 ,
         \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 ,
         \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 ,
         \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 ,
         \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 ,
         \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 ,
         \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 ,
         \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 ,
         \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 ,
         \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 ,
         \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 ,
         \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 ,
         \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 ,
         \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 ,
         \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 ,
         \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 ,
         \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 ,
         \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 ,
         \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 ,
         \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 ,
         \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 ,
         \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 ,
         \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 ,
         \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 ,
         \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 ,
         \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 ,
         \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 ,
         \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 ,
         \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 ,
         \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 ,
         \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 ,
         \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 ,
         \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 ,
         \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 ,
         \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 ,
         \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 ,
         \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 ,
         \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 ,
         \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 ,
         \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 ,
         \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 ,
         \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 ,
         \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 ,
         \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 ,
         \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 ,
         \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 ,
         \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 ,
         \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 ,
         \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 ,
         \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 ,
         \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 ,
         \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 ,
         \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 ,
         \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 ,
         \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 ,
         \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 ,
         \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 ,
         \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 ,
         \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 ,
         \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 ,
         \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 ,
         \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 ,
         \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 ,
         \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 ,
         \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 ,
         \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 ,
         \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 ,
         \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 ,
         \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 ,
         \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 ,
         \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 ,
         \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 ,
         \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 ,
         \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 ,
         \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 ,
         \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 ,
         \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 ,
         \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 ,
         \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 ,
         \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 ,
         \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 ,
         \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 ,
         \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 ,
         \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 ,
         \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 ,
         \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 ,
         \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 ,
         \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 ,
         \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 ,
         \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 ,
         \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 ,
         \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 ,
         \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 ,
         \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 ,
         \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 ,
         \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 ,
         \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 ,
         \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 ,
         \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 ,
         \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 ,
         \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 ,
         \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 ,
         \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 ,
         \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 ,
         \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 ,
         \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 ,
         \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 ,
         \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 ,
         \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 ,
         \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 ,
         \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 ,
         \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 ,
         \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 ,
         \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 ,
         \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 ,
         \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 ,
         \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 ,
         \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 ,
         \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 ,
         \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 ,
         \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 ,
         \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 ,
         \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 ,
         \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 ,
         \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 ,
         \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 ,
         \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 ,
         \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 ,
         \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 ,
         \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 ,
         \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 ,
         \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 ,
         \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 ,
         \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 ,
         \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 ,
         \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 ,
         \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 ,
         \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 ,
         \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 ,
         \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 ,
         \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 ,
         \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 ,
         \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 ,
         \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 ,
         \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 ,
         \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 ,
         \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 ,
         \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 ,
         \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 ,
         \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 ,
         \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 ,
         \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 ,
         \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 ,
         \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 ,
         \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 ,
         \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 ,
         \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 ,
         \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 ,
         \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 ,
         \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 ,
         \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 ,
         \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 ,
         \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 ,
         \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 ,
         \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 ,
         \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 ,
         \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 ,
         \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 ,
         \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 ,
         \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 ,
         \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 ,
         \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 ,
         \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 ,
         \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 ,
         \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 ,
         \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 ,
         \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 ,
         \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 ,
         \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 ,
         \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 ,
         \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 ,
         \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 ,
         \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 ,
         \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 ,
         \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 ,
         \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 ,
         \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 ,
         \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 ,
         \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 ,
         \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 ,
         \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 ,
         \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 ,
         \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 ,
         \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 ,
         \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 ,
         \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 ,
         \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 ,
         \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 ,
         \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 ,
         \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 ,
         \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 ,
         \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 ,
         \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 ,
         \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 ,
         \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 ,
         \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 ,
         \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 ,
         \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 ,
         \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 ,
         \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 ,
         \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 ,
         \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 ,
         \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 ,
         \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 ,
         \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 ,
         \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 ,
         \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 ,
         \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 ,
         \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 ,
         \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 ,
         \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 ,
         \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 ,
         \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 ,
         \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 ,
         \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 ,
         \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 ,
         \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 ,
         \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 ,
         \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 ,
         \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 ,
         \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 ,
         \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 ,
         \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 ,
         \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 ,
         \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 ,
         \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 ,
         \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 ,
         \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 ,
         \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 ,
         \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 ,
         \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 ,
         \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 ,
         \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 ,
         \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 ,
         \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 ,
         \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 ,
         \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 ,
         \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 ,
         \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 ,
         \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 ,
         \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 ,
         \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 ,
         \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 ,
         \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 ,
         \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 ,
         \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 ,
         \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 ,
         \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 ,
         \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 ,
         \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 ,
         \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 ,
         \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 ,
         \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 ,
         \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 ,
         \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 ,
         \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 ,
         \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 ,
         \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 ,
         \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 ,
         \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 ,
         \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 ,
         \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 ,
         \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 ,
         \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 ,
         \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 ,
         \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 ,
         \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 ,
         \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 ,
         \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 ,
         \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 ,
         \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 ,
         \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 ,
         \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 ,
         \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 ,
         \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 ,
         \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 ,
         \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 ,
         \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 ,
         \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 ,
         \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 ,
         \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 ,
         \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 ,
         \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 ,
         \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 ,
         \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 ,
         \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 ,
         \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 ,
         \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 ,
         \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 ,
         \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 ,
         \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 ,
         \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 ,
         \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 ,
         \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 ,
         \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 ,
         \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 ,
         \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 ,
         \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 ,
         \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 ,
         \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 ,
         \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 ,
         \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 ,
         \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 ,
         \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 ,
         \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 ,
         \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 ,
         \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 ,
         \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 ,
         \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 ,
         \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 ,
         \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 ,
         \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 ,
         \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 ,
         \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 ,
         \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 ,
         \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 ,
         \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 ,
         \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 ,
         \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 ,
         \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 ,
         \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 ,
         \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 ,
         \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 ,
         \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 ,
         \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 ,
         \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 ,
         \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 ,
         \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 ,
         \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 ,
         \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 ,
         \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 ,
         \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 ,
         \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 ,
         \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 ,
         \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 ,
         \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 ,
         \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 ,
         \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 ,
         \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 ,
         \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 ,
         \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 ,
         \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 ,
         \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 ,
         \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 ,
         \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 ,
         \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 ,
         \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 ,
         \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 ,
         \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 ,
         \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 ,
         \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 ,
         \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 ,
         \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 ,
         \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 ,
         \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 ,
         \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 ,
         \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 ,
         \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 ,
         \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 ,
         \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 ,
         \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 ,
         \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 ,
         \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 ,
         \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 ,
         \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 ,
         \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 ,
         \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 ,
         \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 ,
         \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 ,
         \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 ,
         \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 ,
         \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 ,
         \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 ,
         \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 ,
         \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 ,
         \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 ,
         \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 ,
         \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 ,
         \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 ,
         \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 ,
         \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 ,
         \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 ,
         \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 ,
         \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 ,
         \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 ,
         \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 ,
         \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 ,
         \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 ,
         \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 ,
         \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 ,
         \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 ,
         \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 ,
         \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 ,
         \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 ,
         \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 ,
         \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 ,
         \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 ,
         \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 ,
         \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 ,
         \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 ,
         \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 ,
         \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 ,
         \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 ,
         \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 ,
         \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 ,
         \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 ,
         \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 ,
         \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 ,
         \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 ,
         \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 ,
         \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 ,
         \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 ,
         \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 ,
         \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 ,
         \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 ,
         \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 ,
         \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 ,
         \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 ,
         \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 ,
         \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 ,
         \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 ,
         \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 ,
         \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 ,
         \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 ,
         \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 ,
         \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 ,
         \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 ,
         \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 ,
         \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 ,
         \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 ,
         \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 ,
         \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 ,
         \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 ,
         \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 ,
         \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 ,
         \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 ,
         \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 ,
         \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 ,
         \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 ,
         \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 ,
         \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 ,
         \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 ,
         \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 ,
         \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 ,
         \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 ,
         \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 ,
         \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 ,
         \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 ,
         \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 ,
         \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 ,
         \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 ,
         \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 ,
         \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 ,
         \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 ,
         \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 ,
         \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 ,
         \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 ,
         \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 ,
         \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 ,
         \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 ,
         \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 ,
         \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 ,
         \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 ,
         \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 ,
         \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 ,
         \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 ,
         \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 ,
         \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 ,
         \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 ,
         \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 ,
         \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 ,
         \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 ,
         \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 ,
         \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 ,
         \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 ,
         \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 ,
         \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 ,
         \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 ,
         \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 ,
         \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 ,
         \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 ,
         \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 ,
         \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 ,
         \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 ,
         \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 ,
         \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 ,
         \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 ,
         \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 ,
         \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 ,
         \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 ,
         \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 ,
         \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 ,
         \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 ,
         \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 ,
         \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 ,
         \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 ,
         \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 ,
         \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 ,
         \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 ,
         \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 ,
         \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 ,
         \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 ,
         \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 ,
         \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 ,
         \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 ,
         \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 ,
         \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 ,
         \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 ,
         \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 ,
         \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 ,
         \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 ,
         \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 ,
         \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 ,
         \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 ,
         \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 ,
         \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 ,
         \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 ,
         \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 ,
         \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 ,
         \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 ,
         \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 ,
         \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 ,
         \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 ,
         \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 ,
         \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 ,
         \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 ,
         \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 ,
         \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 ,
         \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 ,
         \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 ,
         \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 ,
         \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 ,
         \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 ,
         \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 ,
         \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 ,
         \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 ,
         \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 ,
         \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 ,
         \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 ,
         \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 ,
         \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 ,
         \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 ,
         \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 ,
         \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 ,
         \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 ,
         \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 ,
         \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 ,
         \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 ,
         \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 ,
         \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 ,
         \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 ,
         \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 ,
         \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 ,
         \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 ,
         \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 ,
         \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 ,
         \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 ,
         \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 ,
         \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 ,
         \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 ,
         \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 ,
         \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 ,
         \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 ,
         \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 ,
         \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 ,
         \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 ,
         \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 ,
         \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 ,
         \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 ,
         \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 ,
         \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 ,
         \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 ,
         \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 ,
         \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 ,
         \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 ,
         \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 ,
         \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 ,
         \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 ,
         \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 ,
         \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 ,
         \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 ,
         \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 ,
         \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 ,
         \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 ,
         \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 ,
         \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 ,
         \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 ,
         \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 ,
         \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 ,
         \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 ,
         \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 ,
         \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 ,
         \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 ,
         \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 ,
         \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 ,
         \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 ,
         \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 ,
         \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 ,
         \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 ,
         \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 ,
         \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 ,
         \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 ,
         \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 ,
         \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 ,
         \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 ,
         \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 ,
         \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 ,
         \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 ,
         \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 ,
         \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 ,
         \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 ,
         \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 ,
         \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 ,
         \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 ,
         \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 ,
         \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 ,
         \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 ,
         \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 ,
         \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 ,
         \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 ,
         \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 ,
         \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 ,
         \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 ,
         \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 ,
         \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 ,
         \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 ,
         \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 ,
         \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 ,
         \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 ,
         \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 ,
         \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 ,
         \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 ,
         \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 ,
         \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 ,
         \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 ,
         \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 ,
         \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 ,
         \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 ,
         \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 ,
         \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 ,
         \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 ,
         \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 ,
         \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 ,
         \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 ,
         \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 ,
         \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 ,
         \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 ,
         \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 ,
         \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 ,
         \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 ,
         \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 ,
         \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 ,
         \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 ,
         \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 ,
         \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 ,
         \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 ,
         \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 ,
         \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 ,
         \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 ,
         \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 ,
         \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 ,
         \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 ,
         \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 ,
         \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 ,
         \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 ,
         \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 ,
         \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 ,
         \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 ,
         \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 ,
         \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 ,
         \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 ,
         \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 ,
         \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 ,
         \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 ,
         \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 ,
         \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 ,
         \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 ,
         \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 ,
         \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 ,
         \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 ,
         \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 ,
         \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 ,
         \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 ,
         \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 ,
         \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 ,
         \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 ,
         \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 ,
         \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 ,
         \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 ,
         \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 ,
         \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 ,
         \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 ,
         \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 ,
         \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 ,
         \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 ,
         \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 ,
         \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 ,
         \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 ,
         \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 ,
         \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 ,
         \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 ,
         \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 ,
         \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 ,
         \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 ,
         \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 ,
         \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 ,
         \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 ,
         \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 ,
         \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 ,
         \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 ,
         \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 ,
         \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 ,
         \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 ,
         \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 ,
         \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 ,
         \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 ,
         \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 ,
         \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 ,
         \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 ,
         \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 ,
         \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 ,
         \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 ,
         \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 ,
         \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 ,
         \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 ,
         \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 ,
         \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 ,
         \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 ,
         \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 ,
         \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 ,
         \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 ,
         \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 ,
         \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 ,
         \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 ,
         \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 ,
         \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 ,
         \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 ,
         \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 ,
         \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 ,
         \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 ,
         \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 ,
         \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 ,
         \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 ,
         \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 ,
         \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 ,
         \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 ,
         \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 ,
         \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 ,
         \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 ,
         \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 ,
         \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 ,
         \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 ,
         \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 ,
         \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 ,
         \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 ,
         \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 ,
         \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 ,
         \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 ,
         \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 ,
         \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 ,
         \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 ,
         \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 ,
         \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 ,
         \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 ,
         \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 ,
         \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 ,
         \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 ,
         \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 ,
         \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 ,
         \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 ,
         \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 ,
         \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 ,
         \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 ,
         \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 ,
         \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 ,
         \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 ,
         \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 ,
         \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 ,
         \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 ,
         \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 ,
         \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 ,
         \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 ,
         \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 ,
         \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 ,
         \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 ,
         \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 ,
         \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 ,
         \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 ,
         \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 ,
         \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 ,
         \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 ,
         \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 ,
         \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 ,
         \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 ,
         \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 ,
         \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 ,
         \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 ,
         \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 ,
         \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 ,
         \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 ,
         \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 ,
         \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 ,
         \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 ,
         \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 ,
         \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 ,
         \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 ,
         \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 ,
         \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 ,
         \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 ,
         \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 ,
         \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 ,
         \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 ,
         \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 ,
         \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 ,
         \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 ,
         \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 ,
         \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 ,
         \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 ,
         \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 ,
         \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 ,
         \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 ,
         \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 ,
         \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 ,
         \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 ,
         \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 ,
         \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 ,
         \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 ,
         \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 ,
         \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 ,
         \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 ,
         \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 ,
         \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 ,
         \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 ,
         \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 ,
         \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 ,
         \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 ,
         \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 ,
         \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 ,
         \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 ,
         \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 ,
         \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 ,
         \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 ,
         \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 ,
         \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 ,
         \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 ,
         \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 ,
         \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 ,
         \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 ,
         \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 ,
         \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 ,
         \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 ,
         \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 ,
         \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 ,
         \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 ,
         \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 ,
         \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 ,
         \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 ,
         \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 ,
         \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 ,
         \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 ,
         \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 ,
         \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 ,
         \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 ,
         \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 ,
         \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 ,
         \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 ,
         \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 ,
         \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 ,
         \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 ,
         \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 ,
         \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 ,
         \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 ,
         \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 ,
         \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 ,
         \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 ,
         \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 ,
         \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 ,
         \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 ,
         \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 ,
         \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 ,
         \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 ,
         \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 ,
         \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 ,
         \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 ,
         \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 ,
         \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 ,
         \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 ,
         \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 ,
         \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 ,
         \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 ,
         \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 ,
         \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 ,
         \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 ,
         \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 ,
         \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 ,
         \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 ,
         \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 ,
         \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 ,
         \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 ,
         \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 ,
         \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 ,
         \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 ,
         \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 ,
         \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 ,
         \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 ,
         \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 ,
         \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 ,
         \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 ,
         \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 ,
         \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 ,
         \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 ,
         \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 ,
         \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 ,
         \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 ,
         \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 ,
         \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 ,
         \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 ,
         \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 ,
         \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 ,
         \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 ,
         \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 ,
         \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 ,
         \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 ,
         \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 ,
         \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 ,
         \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 ,
         \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 ,
         \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 ,
         \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 ,
         \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 ,
         \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 ,
         \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 ,
         \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 ,
         \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 ,
         \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 ,
         \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 ,
         \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 ,
         \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 ,
         \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 ,
         \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 ,
         \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 ,
         \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 ,
         \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 ,
         \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 ,
         \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 ,
         \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 ,
         \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 ,
         \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 ,
         \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 ,
         \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 ,
         \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 ,
         \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 ,
         \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 ,
         \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 ,
         \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 ,
         \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 ,
         \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 ,
         \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 ,
         \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 ,
         \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 ,
         \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 ,
         \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 ,
         \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 ,
         \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 ,
         \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 ,
         \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 ,
         \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 ,
         \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 ,
         \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 ,
         \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 ,
         \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 ,
         \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 ,
         \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 ,
         \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 ,
         \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 ,
         \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 ,
         \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 ,
         \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 ,
         \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 ,
         \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 ,
         \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 ,
         \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 ,
         \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 ,
         \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 ,
         \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 ,
         \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 ,
         \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 ,
         \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 ,
         \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 ,
         \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 ,
         \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 ,
         \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 ,
         \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 ,
         \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 ,
         \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 ,
         \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 ,
         \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 ,
         \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 ,
         \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 ,
         \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 ,
         \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 ,
         \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 ,
         \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 ,
         \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 ,
         \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 ,
         \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 ,
         \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 ,
         \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 ,
         \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 ,
         \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 ,
         \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 ,
         \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 ,
         \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 ,
         \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 ,
         \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 ,
         \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 ,
         \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 ,
         \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 ,
         \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 ,
         \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 ,
         \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 ,
         \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 ,
         \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 ,
         \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 ,
         \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 ,
         \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 ,
         \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 ,
         \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 ,
         \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 ,
         \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 ,
         \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 ,
         \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 ,
         \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 ,
         \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 ,
         \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 ,
         \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 ,
         \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 ,
         \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 ,
         \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 ,
         \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 ,
         \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 ,
         \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 ,
         \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 ,
         \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 ,
         \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 ,
         \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 ,
         \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 ,
         \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 ,
         \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 ,
         \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 ,
         \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 ,
         \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 ,
         \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 ,
         \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 ,
         \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 ,
         \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 ,
         \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 ,
         \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 ,
         \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 ,
         \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 ,
         \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 ,
         \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 ,
         \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 ,
         \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 ,
         \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 ,
         \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 ,
         \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 ,
         \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 ,
         \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 ,
         \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 ,
         \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 ,
         \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 ,
         \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 ,
         \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 ,
         \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 ,
         \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 ,
         \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 ,
         \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 ,
         \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 ,
         \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 ,
         \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 ,
         \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 ,
         \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 ,
         \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 ,
         \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 ,
         \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 ,
         \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 ,
         \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 ,
         \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 ,
         \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 ,
         \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 ,
         \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 ,
         \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 ,
         \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 ,
         \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 ,
         \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 ,
         \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 ,
         \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 ,
         \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 ,
         \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 ,
         \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 ,
         \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 ,
         \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 ,
         \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 ,
         \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 ,
         \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 ,
         \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 ,
         \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 ,
         \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 ,
         \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 ,
         \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 ,
         \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 ,
         \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 ,
         \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 ,
         \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 ,
         \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 ,
         \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 ,
         \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 ,
         \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 ,
         \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 ,
         \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 ,
         \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 ,
         \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 ,
         \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 ,
         \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 ,
         \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 ,
         \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 ,
         \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 ,
         \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 ,
         \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 ,
         \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 ,
         \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 ,
         \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 ,
         \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 ,
         \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 ,
         \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 ,
         \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 ,
         \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 ,
         \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 ,
         \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 ,
         \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 ,
         \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 ,
         \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 ,
         \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 ,
         \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 ,
         \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 ,
         \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 ,
         \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 ,
         \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 ,
         \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 ,
         \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 ,
         \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 ,
         \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 ,
         \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 ,
         \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 ,
         \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 ,
         \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 ,
         \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 ,
         \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 ,
         \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 ,
         \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 ,
         \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 ,
         \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 ,
         \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 ,
         \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 ,
         \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 ,
         \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 ,
         \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 ,
         \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 ,
         \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 ,
         \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 ,
         \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 ,
         \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 ,
         \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 ,
         \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 ,
         \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 ,
         \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 ,
         \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 ,
         \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 ,
         \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 ,
         \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 ,
         \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 ,
         \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 ,
         \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 ,
         \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 ,
         \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 ,
         \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 ,
         \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 ,
         \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 ,
         \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 ,
         \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 ,
         \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 ,
         \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 ,
         \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 ,
         \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 ,
         \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 ,
         \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 ,
         \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 ,
         \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 ,
         \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 ,
         \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 ,
         \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 ,
         \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 ,
         \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 ,
         \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 ,
         \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 ,
         \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 ,
         \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 ,
         \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 ,
         \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 ,
         \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 ,
         \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 ,
         \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 ,
         \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 ,
         \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 ,
         \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 ,
         \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 ,
         \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 ,
         \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 ,
         \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 ,
         \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 ,
         \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 ,
         \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 ,
         \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 ,
         \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 ,
         \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 ,
         \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 ,
         \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 ,
         \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 ,
         \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 ,
         \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 ,
         \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 ,
         \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 ,
         \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 ,
         \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 ,
         \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 ,
         \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 ,
         \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 ,
         \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 ,
         \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 ,
         \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 ,
         \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 ,
         \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 ,
         \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 ,
         \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 ,
         \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 ,
         \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 ,
         \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 ,
         \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 ,
         \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 ,
         \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 ,
         \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 ,
         \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 ,
         \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 ,
         \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 ,
         \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 ,
         \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 ,
         \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 ,
         \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 ,
         \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 ,
         \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 ,
         \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 ,
         \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 ,
         \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 ,
         \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 ,
         \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 ,
         \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 ,
         \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 ,
         \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 ,
         \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 ,
         \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 ,
         \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 ,
         \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 ,
         \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 ,
         \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 ,
         \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 ,
         \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 ,
         \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 ,
         \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 ,
         \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 ,
         \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 ,
         \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 ,
         \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 ,
         \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 ,
         \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 ,
         \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 ,
         \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 ,
         \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 ,
         \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 ,
         \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 ,
         \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 ,
         \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 ,
         \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 ,
         \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 ,
         \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 ,
         \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 ,
         \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 ,
         \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 ,
         \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 ,
         \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 ,
         \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 ,
         \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 ,
         \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 ,
         \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 ,
         \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 ,
         \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 ,
         \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 ,
         \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 ,
         \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 ,
         \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 ,
         \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 ,
         \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 ,
         \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 ,
         \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 ,
         \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 ,
         \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 ,
         \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 ,
         \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 ,
         \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 ,
         \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 ,
         \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 ,
         \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 ,
         \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 ,
         \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 ,
         \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 ,
         \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 ,
         \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 ,
         \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 ,
         \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 ,
         \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 ,
         \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 ,
         \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 ,
         \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 ,
         \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 ,
         \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 ,
         \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 ,
         \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 ,
         \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 ,
         \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 ,
         \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 ,
         \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 ,
         \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 ,
         \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 ,
         \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 ,
         \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 ,
         \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 ,
         \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 ,
         \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 ,
         \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 ,
         \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 ,
         \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 ,
         \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 ,
         \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 ,
         \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 ,
         \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 ,
         \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 ,
         \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 ,
         \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 ,
         \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 ,
         \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 ,
         \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 ,
         \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 ,
         \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 ,
         \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 ,
         \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 ,
         \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 ,
         \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 ,
         \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 ,
         \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 ,
         \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 ,
         \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 ,
         \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 ,
         \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 ,
         \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 ,
         \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 ,
         \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 ,
         \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 ,
         \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 ,
         \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 ,
         \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 ,
         \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 ,
         \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 ,
         \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 ,
         \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 ,
         \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 ,
         \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 ,
         \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 ,
         \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 ,
         \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 ,
         \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 ,
         \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 ,
         \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 ,
         \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 ,
         \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 ,
         \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 ,
         \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 ,
         \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 ,
         \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 ,
         \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 ,
         \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 ,
         \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 ,
         \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 ,
         \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 ,
         \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 ,
         \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 ,
         \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 ,
         \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 ,
         \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 ,
         \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 ,
         \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 ,
         \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 ,
         \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 ,
         \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 ,
         \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 ,
         \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 ,
         \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 ,
         \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 ,
         \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 ,
         \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 ,
         \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 ,
         \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 ,
         \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 ,
         \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 ,
         \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 ,
         \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 ,
         \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 ,
         \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 ,
         \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 ,
         \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 ,
         \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 ,
         \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 ,
         \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 ,
         \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 ,
         \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 ,
         \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 ,
         \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 ,
         \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 ,
         \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 ,
         \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 ,
         \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 ,
         \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 ,
         \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 ,
         \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 ,
         \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 ,
         \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 ,
         \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 ,
         \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 ,
         \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 ,
         \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 ,
         \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 ,
         \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 ,
         \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 ,
         \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 ,
         \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 ,
         \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 ,
         \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 ,
         \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 ,
         \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 ,
         \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 ,
         \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 ,
         \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 ,
         \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 ,
         \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 ,
         \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 ,
         \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 ,
         \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 ,
         \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 ,
         \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 ,
         \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 ,
         \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 ,
         \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 ,
         \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 ,
         \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 ,
         \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 ,
         \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 ,
         \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 ,
         \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 ,
         \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 ,
         \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 ,
         \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 ,
         \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 ,
         \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 ,
         \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 ,
         \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 ,
         \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 ,
         \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 ,
         \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 ,
         \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 ,
         \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 ,
         \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 ,
         \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 ,
         \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 ,
         \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 ,
         \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 ,
         \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 ,
         \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 ,
         \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 ,
         \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 ,
         \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 ,
         \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 ,
         \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 ,
         \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 ,
         \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 ,
         \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 ,
         \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 ,
         \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 ,
         \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 ,
         \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 ,
         \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 ,
         \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 ,
         \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 ,
         \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 ,
         \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 ,
         \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 ,
         \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 ,
         \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 ,
         \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 ,
         \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 ,
         \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 ,
         \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 ,
         \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 ,
         \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 ,
         \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 ,
         \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 ,
         \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 ,
         \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 ,
         \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 ,
         \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 ,
         \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 ,
         \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 ,
         \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 ,
         \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 ,
         \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 ,
         \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 ,
         \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 ,
         \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 ,
         \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 ,
         \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 ,
         \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 ,
         \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 ,
         \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 ,
         \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 ,
         \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 ,
         \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 ,
         \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 ,
         \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 ,
         \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 ,
         \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 ,
         \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 ,
         \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 ,
         \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 ,
         \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 ,
         \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 ,
         \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 ,
         \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 ,
         \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 ,
         \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 ,
         \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 ,
         \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 ,
         \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 ,
         \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 ,
         \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 ,
         \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 ,
         \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 ,
         \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 ,
         \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 ,
         \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 ,
         \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 ,
         \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 ,
         \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 ,
         \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 ,
         \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 ,
         \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 ,
         \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 ,
         \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 ,
         \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 ,
         \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 ,
         \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 ,
         \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 ,
         \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 ,
         \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 ,
         \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 ,
         \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 ,
         \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 ,
         \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 ,
         \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 ,
         \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 ,
         \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 ,
         \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 ,
         \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 ,
         \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 ,
         \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 ,
         \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 ,
         \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 ,
         \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 ,
         \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 ,
         \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 ,
         \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 ,
         \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 ,
         \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 ,
         \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 ,
         \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 ,
         \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 ,
         \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 ,
         \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 ,
         \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 ,
         \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 ,
         \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 ,
         \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 ,
         \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 ,
         \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 ,
         \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 ,
         \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 ,
         \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 ,
         \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 ,
         \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 ,
         \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 ,
         \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 ,
         \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 ,
         \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 ,
         \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 ,
         \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 ,
         \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 ,
         \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 ,
         \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 ,
         \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 ,
         \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 ,
         \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 ,
         \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 ,
         \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 ,
         \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 ,
         \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 ,
         \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 ,
         \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 ,
         \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 ,
         \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 ,
         \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 ,
         \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 ,
         \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 ,
         \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 ,
         \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 ,
         \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 ,
         \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 ,
         \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 ,
         \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 ,
         \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 ,
         \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 ,
         \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 ,
         \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 ,
         \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 ,
         \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 ,
         \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 ,
         \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 ,
         \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 ,
         \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 ,
         \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 ,
         \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 ,
         \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 ,
         \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 ,
         \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 ,
         \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 ,
         \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 ,
         \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 ,
         \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 ,
         \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 ,
         \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 ,
         \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 ,
         \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 ,
         \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 ,
         \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 ,
         \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 ,
         \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 ,
         \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 ,
         \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 ,
         \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 ,
         \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 ,
         \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 ,
         \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 ,
         \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 ,
         \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 ,
         \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 ,
         \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 ,
         \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 ,
         \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 ,
         \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 ,
         \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 ,
         \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 ,
         \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 ,
         \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 ,
         \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 ,
         \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 ,
         \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 ,
         \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 ,
         \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 ,
         \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 ,
         \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 ,
         \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 ,
         \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 ,
         \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 ,
         \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 ,
         \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 ,
         \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 ,
         \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 ,
         \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 ,
         \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 ,
         \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 ,
         \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 ,
         \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 ,
         \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 ,
         \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 ,
         \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 ,
         \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 ,
         \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 ,
         \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 ,
         \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 ,
         \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 ,
         \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 ,
         \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 ,
         \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 ,
         \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 ,
         \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 ,
         \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 ,
         \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 ,
         \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 ,
         \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 ,
         \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 ,
         \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 ,
         \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 ,
         \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 ,
         \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 ,
         \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 ,
         \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 ,
         \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 ,
         \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 ,
         \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 ,
         \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 ,
         \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 ,
         \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 ,
         \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 ,
         \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 ,
         \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 ,
         \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 ,
         \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 ,
         \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 ,
         \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 ,
         \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 ,
         \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 ,
         \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 ,
         \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 ,
         \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 ,
         \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 ,
         \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 ,
         \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 ,
         \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 ,
         \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 ,
         \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 ,
         \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 ,
         \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 ,
         \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 ,
         \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 ,
         \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 ,
         \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 ,
         \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 ,
         \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 ,
         \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 ,
         \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 ,
         \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 ,
         \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 ,
         \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 ,
         \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 ,
         \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 ,
         \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 ,
         \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 ,
         \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 ,
         \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 ,
         \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 ,
         \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 ,
         \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 ,
         \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 ,
         \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 ,
         \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 ,
         \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 ,
         \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 ,
         \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 ,
         \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 ,
         \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 ,
         \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 ,
         \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 ,
         \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 ,
         \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 ,
         \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 ,
         \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 ,
         \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 ,
         \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 ,
         \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 ,
         \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 ,
         \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 ,
         \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 ,
         \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 ,
         \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 ,
         \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 ,
         \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 ,
         \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 ,
         \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 ,
         \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 ,
         \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 ,
         \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 ,
         \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 ,
         \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 ,
         \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 ,
         \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 ,
         \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 ,
         \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 ,
         \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 ,
         \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 ,
         \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 ,
         \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 ,
         \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 ,
         \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 ,
         \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 ,
         \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 ,
         \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 ,
         \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 ,
         \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 ,
         \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 ,
         \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 ,
         \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 ,
         \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 ,
         \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 ,
         \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 ,
         \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 ,
         \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 ,
         \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 ,
         \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 ,
         \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 ,
         \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 ,
         \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 ,
         \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 ,
         \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 ,
         \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 ,
         \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 ,
         \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 ,
         \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 ,
         \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 ,
         \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 ,
         \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 ,
         \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 ,
         \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 ,
         \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 ,
         \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 ,
         \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 ,
         \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 ,
         \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 ,
         \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 ,
         \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 ,
         \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 ,
         \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 ,
         \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 ,
         \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 ,
         \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 ,
         \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 ,
         \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 ,
         \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 ,
         \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 ,
         \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 ,
         \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 ,
         \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 ,
         \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 ,
         \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 ,
         \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 ,
         \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 ,
         \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 ,
         \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 ,
         \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 ,
         \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 ,
         \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 ,
         \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 ,
         \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 ,
         \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 ,
         \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 ,
         \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 ,
         \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 ,
         \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 ,
         \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 ,
         \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 ,
         \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 ,
         \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 ,
         \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 ,
         \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 ,
         \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 ,
         \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 ,
         \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 ,
         \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 ,
         \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 ,
         \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 ,
         \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 ,
         \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 ,
         \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 ,
         \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 ,
         \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 ,
         \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 ,
         \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 ,
         \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 ,
         \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 ,
         \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 ,
         \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 ,
         \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 ,
         \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 ,
         \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 ,
         \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 ,
         \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 ,
         \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 ,
         \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 ,
         \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 ,
         \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 ,
         \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 ,
         \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 ,
         \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 ,
         \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 ,
         \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 ,
         \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 ,
         \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 ,
         \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 ,
         \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 ,
         \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 ,
         \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 ,
         \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 ,
         \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 ,
         \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 ,
         \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 ,
         \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 ,
         \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 ,
         \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 ,
         \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 ,
         \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 ,
         \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 ,
         \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 ,
         \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 ,
         \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 ,
         \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 ,
         \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 ,
         \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 ,
         \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 ,
         \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 ,
         \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 ,
         \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 ,
         \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 ,
         \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 ,
         \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 ,
         \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 ,
         \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 ,
         \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 ,
         \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 ,
         \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 ,
         \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 ,
         \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 ,
         \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 ,
         \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 ,
         \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 ,
         \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 ,
         \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 ,
         \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 ,
         \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 ,
         \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 ,
         \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 ,
         \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 ,
         \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 ,
         \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 ,
         \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 ,
         \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 ,
         \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 ,
         \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 ,
         \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 ,
         \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 ,
         \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 ,
         \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 ,
         \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 ,
         \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 ,
         \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 ,
         \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 ,
         \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 ,
         \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 ,
         \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 ,
         \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 ,
         \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 ,
         \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 ,
         \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 ,
         \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 ,
         \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 ,
         \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 ,
         \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 ,
         \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 ,
         \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 ,
         \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 ,
         \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 ,
         \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 ,
         \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 ,
         \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 ,
         \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 ,
         \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 ,
         \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 ,
         \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 ,
         \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 ,
         \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 ,
         \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 ,
         \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 ,
         \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 ,
         \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 ,
         \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 ,
         \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 ,
         \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 ,
         \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 ,
         \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 ,
         \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 ,
         \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 ,
         \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 ,
         \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 ,
         \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 ,
         \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 ,
         \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 ,
         \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 ,
         \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 ,
         \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 ,
         \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 ,
         \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 ,
         \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 ,
         \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 ,
         \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 ,
         \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 ,
         \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 ,
         \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 ,
         \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 ,
         \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 ,
         \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 ,
         \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 ,
         \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 ,
         \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 ,
         \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 ,
         \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 ,
         \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 ,
         \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 ,
         \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 ,
         \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 ,
         \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 ,
         \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 ,
         \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 ,
         \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 ,
         \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 ,
         \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 ,
         \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 ,
         \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 ,
         \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 ,
         \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 ,
         \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 ,
         \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 ,
         \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 ,
         \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 ,
         \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 ,
         \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 ,
         \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 ,
         \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 ,
         \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 ,
         \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 ,
         \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 ,
         \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 ,
         \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 ,
         \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 ,
         \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 ,
         \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 ,
         \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 ,
         \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 ,
         \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 ,
         \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 ,
         \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 ,
         \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 ,
         \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 ,
         \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 ,
         \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 ,
         \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 ,
         \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 ,
         \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 ,
         \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 ,
         \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 ,
         \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 ,
         \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 ,
         \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 ,
         \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 ,
         \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 ,
         \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 ,
         \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 ,
         \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 ,
         \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 ,
         \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 ,
         \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 ,
         \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 ,
         \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 ,
         \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 ,
         \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 ,
         \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 ,
         \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 ,
         \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 ,
         \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 ,
         \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 ,
         \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 ,
         \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 ,
         \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 ,
         \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 ,
         \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 ,
         \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 ,
         \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 ,
         \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 ,
         \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 ,
         \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 ,
         \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 ,
         \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 ,
         \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 ,
         \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 ,
         \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 ,
         \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 ,
         \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 ,
         \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 ,
         \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 ,
         \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 ,
         \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 ,
         \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 ,
         \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 ,
         \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 ,
         \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 ,
         \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 ,
         \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 ,
         \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 ,
         \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 ,
         \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 ,
         \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 ,
         \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 ,
         \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 ,
         \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 ,
         \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 ,
         \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 ,
         \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 ,
         \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 ,
         \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 ,
         \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 ,
         \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 ,
         \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 ,
         \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 ,
         \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 ,
         \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 ,
         \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 ,
         \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 ,
         \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 ,
         \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 ,
         \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 ,
         \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 ,
         \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 ,
         \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 ,
         \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 ,
         \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 ,
         \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 ,
         \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 ,
         \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 ,
         \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 ,
         \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 ,
         \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 ,
         \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 ,
         \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 ,
         \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 ,
         \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 ,
         \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 ,
         \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 ,
         \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 ,
         \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 ,
         \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 ,
         \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 ,
         \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 ,
         \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 ,
         \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 ,
         \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 ,
         \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 ,
         \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 ,
         \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 ,
         \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 ,
         \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 ,
         \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 ,
         \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 ,
         \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 ,
         \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 ,
         \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 ,
         \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 ,
         \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 ,
         \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 ,
         \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 ,
         \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 ,
         \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 ,
         \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 ,
         \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 ,
         \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 ,
         \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 ,
         \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 ,
         \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 ,
         \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 ,
         \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 ,
         \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 ,
         \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 ,
         \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 ,
         \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 ,
         \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 ,
         \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 ,
         \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 ,
         \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 ,
         \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 ,
         \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 ,
         \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 ,
         \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 ,
         \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 ,
         \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 ,
         \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 ,
         \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 ,
         \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 ,
         \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 ,
         \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 ,
         \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 ,
         \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 ,
         \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 ,
         \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 ,
         \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 ,
         \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 ,
         \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 ,
         \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 ,
         \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 ,
         \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 ,
         \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 ,
         \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 ,
         \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 ,
         \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 ,
         \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 ,
         \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 ,
         \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 ,
         \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 ,
         \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 ,
         \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 ,
         \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 ,
         \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 ,
         \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 ,
         \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 ,
         \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 ,
         \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 ,
         \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 ,
         \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 ,
         \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 ,
         \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 ,
         \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 ,
         \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 ,
         \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 ,
         \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 ,
         \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 ,
         \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 ,
         \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 ,
         \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 ,
         \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 ,
         \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 ,
         \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 ,
         \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 ,
         \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 ,
         \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 ,
         \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 ,
         \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 ,
         \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 ,
         \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 ,
         \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 ,
         \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 ,
         \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 ,
         \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 ,
         \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 ,
         \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 ,
         \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 ,
         \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 ,
         \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 ,
         \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 ,
         \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 ,
         \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 ,
         \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 ,
         \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 ,
         \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 ,
         \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 ,
         \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 ,
         \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 ,
         \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 ,
         \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 ,
         \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 ,
         \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 ,
         \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 ,
         \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 ,
         \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 ,
         \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 ,
         \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 ,
         \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 ,
         \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 ,
         \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 ,
         \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 ,
         \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 ,
         \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 ,
         \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 ,
         \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 ,
         \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 ,
         \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 ,
         \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 ,
         \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 ,
         \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 ,
         \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 ,
         \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 ,
         \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 ,
         \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 ,
         \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 ,
         \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 ,
         \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 ,
         \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 ,
         \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 ,
         \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 ,
         \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 ,
         \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 ,
         \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 ,
         \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 ,
         \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 ,
         \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 ,
         \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 ,
         \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 ,
         \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 ,
         \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 ,
         \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 ,
         \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 ,
         \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 ,
         \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 ,
         \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 ,
         \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 ,
         \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 ,
         \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 ,
         \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 ,
         \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 ,
         \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 ,
         \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 ,
         \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 ,
         \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 ,
         \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 ,
         \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 ,
         \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 ,
         \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 ,
         \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 ,
         \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 ,
         \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 ,
         \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 ,
         \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 ,
         \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 ,
         \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 ,
         \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 ,
         \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 ,
         \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 ,
         \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 ,
         \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 ,
         \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 ,
         \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 ,
         \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 ,
         \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 ,
         \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 ,
         \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 ,
         \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 ,
         \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 ,
         \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 ,
         \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 ,
         \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 ,
         \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 ,
         \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 ,
         \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 ,
         \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 ,
         \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 ,
         \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 ,
         \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 ,
         \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 ,
         \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 ,
         \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 ,
         \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 ,
         \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 ,
         \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 ,
         \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 ,
         \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 ,
         \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 ,
         \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 ,
         \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 ,
         \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 ,
         \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 ,
         \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 ,
         \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 ,
         \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 ,
         \42393 , \42394 , \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 ,
         \42403 , \42404 , \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 ,
         \42413 , \42414 , \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 ,
         \42423 , \42424 , \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 ,
         \42433 , \42434 , \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 ,
         \42443 , \42444 , \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 ,
         \42453 , \42454 , \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 ,
         \42463 , \42464 , \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 ,
         \42473 , \42474 , \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 ,
         \42483 , \42484 , \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 ,
         \42493 , \42494 , \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 ,
         \42503 , \42504 , \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 ,
         \42513 , \42514 , \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 ,
         \42523 , \42524 , \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 ,
         \42533 , \42534 , \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 ,
         \42543 , \42544 , \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 ,
         \42553 , \42554 , \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 ,
         \42563 , \42564 , \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 ,
         \42573 , \42574 , \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 ,
         \42583 , \42584 , \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 ,
         \42593 , \42594 , \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 ,
         \42603 , \42604 , \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 ,
         \42613 , \42614 , \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 ,
         \42623 , \42624 , \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 ,
         \42633 , \42634 , \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 ,
         \42643 , \42644 , \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 ,
         \42653 , \42654 , \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 ,
         \42663 , \42664 , \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 ,
         \42673 , \42674 , \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 ,
         \42683 , \42684 , \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 ,
         \42693 , \42694 , \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 ,
         \42703 , \42704 , \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 ,
         \42713 , \42714 , \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 ,
         \42723 , \42724 , \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 ,
         \42733 , \42734 , \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 ,
         \42743 , \42744 , \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 ,
         \42753 , \42754 , \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 ,
         \42763 , \42764 , \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 ,
         \42773 , \42774 , \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 ,
         \42783 , \42784 , \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 ,
         \42793 , \42794 , \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 ,
         \42803 , \42804 , \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 ,
         \42813 , \42814 , \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 ,
         \42823 , \42824 , \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 ,
         \42833 , \42834 , \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 ,
         \42843 , \42844 , \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 ,
         \42853 , \42854 , \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 ,
         \42863 , \42864 , \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 ,
         \42873 , \42874 , \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 ,
         \42883 , \42884 , \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 ,
         \42893 , \42894 , \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 ,
         \42903 , \42904 , \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 ,
         \42913 , \42914 , \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 ,
         \42923 , \42924 , \42925 , \42926 , \42927 , \42928 , \42929 , \42930 , \42931 , \42932 ,
         \42933 , \42934 , \42935 , \42936 , \42937 , \42938 , \42939 , \42940 , \42941 , \42942 ,
         \42943 , \42944 , \42945 , \42946 , \42947 , \42948 , \42949 , \42950 , \42951 , \42952 ,
         \42953 , \42954 , \42955 , \42956 , \42957 , \42958 , \42959 , \42960 , \42961 , \42962 ,
         \42963 , \42964 , \42965 , \42966 , \42967 , \42968 , \42969 , \42970 , \42971 , \42972 ,
         \42973 , \42974 , \42975 , \42976 , \42977 , \42978 , \42979 , \42980 , \42981 , \42982 ,
         \42983 , \42984 , \42985 , \42986 , \42987 , \42988 , \42989 , \42990 , \42991 , \42992 ,
         \42993 , \42994 , \42995 , \42996 , \42997 , \42998 , \42999 , \43000 , \43001 , \43002 ,
         \43003 , \43004 , \43005 , \43006 , \43007 , \43008 , \43009 , \43010 , \43011 , \43012 ,
         \43013 , \43014 , \43015 , \43016 , \43017 , \43018 , \43019 , \43020 , \43021 , \43022 ,
         \43023 , \43024 , \43025 , \43026 , \43027 , \43028 , \43029 , \43030 , \43031 , \43032 ,
         \43033 , \43034 , \43035 , \43036 , \43037 , \43038 , \43039 , \43040 , \43041 , \43042 ,
         \43043 , \43044 , \43045 , \43046 , \43047 , \43048 , \43049 , \43050 , \43051 , \43052 ,
         \43053 , \43054 , \43055 , \43056 , \43057 , \43058 , \43059 , \43060 , \43061 , \43062 ,
         \43063 , \43064 , \43065 , \43066 , \43067 , \43068 , \43069 , \43070 , \43071 , \43072 ,
         \43073 , \43074 , \43075 , \43076 , \43077 , \43078 , \43079 , \43080 , \43081 , \43082 ,
         \43083 , \43084 , \43085 , \43086 , \43087 , \43088 , \43089 , \43090 , \43091 , \43092 ,
         \43093 , \43094 , \43095 , \43096 , \43097 , \43098 , \43099 , \43100 , \43101 , \43102 ,
         \43103 , \43104 , \43105 , \43106 , \43107 , \43108 , \43109 , \43110 , \43111 , \43112 ,
         \43113 , \43114 , \43115 , \43116 , \43117 , \43118 , \43119 , \43120 , \43121 , \43122 ,
         \43123 , \43124 , \43125 , \43126 , \43127 , \43128 , \43129 , \43130 , \43131 , \43132 ,
         \43133 , \43134 , \43135 , \43136 , \43137 , \43138 , \43139 , \43140 , \43141 , \43142 ,
         \43143 , \43144 , \43145 , \43146 , \43147 , \43148 , \43149 , \43150 , \43151 , \43152 ,
         \43153 , \43154 , \43155 , \43156 , \43157 , \43158 , \43159 , \43160 , \43161 , \43162 ,
         \43163 , \43164 , \43165 , \43166 , \43167 , \43168 , \43169 , \43170 , \43171 , \43172 ,
         \43173 , \43174 , \43175 , \43176 , \43177 , \43178 , \43179 , \43180 , \43181 , \43182 ,
         \43183 , \43184 , \43185 , \43186 , \43187 , \43188 , \43189 , \43190 , \43191 , \43192 ,
         \43193 , \43194 , \43195 , \43196 , \43197 , \43198 , \43199 , \43200 , \43201 , \43202 ,
         \43203 , \43204 , \43205 , \43206 , \43207 , \43208 , \43209 , \43210 , \43211 , \43212 ,
         \43213 , \43214 , \43215 , \43216 , \43217 , \43218 , \43219 , \43220 , \43221 , \43222 ,
         \43223 , \43224 , \43225 , \43226 , \43227 , \43228 , \43229 , \43230 , \43231 , \43232 ,
         \43233 , \43234 , \43235 , \43236 , \43237 , \43238 , \43239 , \43240 , \43241 , \43242 ,
         \43243 , \43244 , \43245 , \43246 , \43247 , \43248 , \43249 , \43250 , \43251 , \43252 ,
         \43253 , \43254 , \43255 , \43256 , \43257 , \43258 , \43259 , \43260 , \43261 , \43262 ,
         \43263 , \43264 , \43265 , \43266 , \43267 , \43268 , \43269 , \43270 , \43271 , \43272 ,
         \43273 , \43274 , \43275 , \43276 , \43277 , \43278 , \43279 , \43280 , \43281 , \43282 ,
         \43283 , \43284 , \43285 , \43286 , \43287 , \43288 , \43289 , \43290 , \43291 , \43292 ,
         \43293 , \43294 , \43295 , \43296 , \43297 , \43298 , \43299 , \43300 , \43301 , \43302 ,
         \43303 , \43304 , \43305 , \43306 , \43307 , \43308 , \43309 , \43310 , \43311 , \43312 ,
         \43313 , \43314 , \43315 , \43316 , \43317 , \43318 , \43319 , \43320 , \43321 , \43322 ,
         \43323 , \43324 , \43325 , \43326 , \43327 , \43328 , \43329 , \43330 , \43331 , \43332 ,
         \43333 , \43334 , \43335 , \43336 , \43337 , \43338 , \43339 , \43340 , \43341 , \43342 ,
         \43343 , \43344 , \43345 , \43346 , \43347 , \43348 , \43349 , \43350 , \43351 , \43352 ,
         \43353 , \43354 , \43355 , \43356 , \43357 , \43358 , \43359 , \43360 , \43361 , \43362 ,
         \43363 , \43364 , \43365 , \43366 , \43367 , \43368 , \43369 , \43370 , \43371 , \43372 ,
         \43373 , \43374 , \43375 , \43376 , \43377 , \43378 , \43379 , \43380 , \43381 , \43382 ,
         \43383 , \43384 , \43385 , \43386 , \43387 , \43388 , \43389 , \43390 , \43391 , \43392 ,
         \43393 , \43394 , \43395 , \43396 , \43397 , \43398 , \43399 , \43400 , \43401 , \43402 ,
         \43403 , \43404 , \43405 , \43406 , \43407 , \43408 , \43409 , \43410 , \43411 , \43412 ,
         \43413 , \43414 , \43415 , \43416 , \43417 , \43418 , \43419 , \43420 , \43421 , \43422 ,
         \43423 , \43424 , \43425 , \43426 , \43427 , \43428 , \43429 , \43430 , \43431 , \43432 ,
         \43433 , \43434 , \43435 , \43436 , \43437 , \43438 , \43439 , \43440 , \43441 , \43442 ,
         \43443 , \43444 , \43445 , \43446 , \43447 , \43448 , \43449 , \43450 , \43451 , \43452 ,
         \43453 , \43454 , \43455 , \43456 , \43457 , \43458 , \43459 , \43460 , \43461 , \43462 ,
         \43463 , \43464 , \43465 , \43466 , \43467 , \43468 , \43469 , \43470 , \43471 , \43472 ,
         \43473 , \43474 , \43475 , \43476 , \43477 , \43478 , \43479 , \43480 , \43481 , \43482 ,
         \43483 , \43484 , \43485 , \43486 , \43487 , \43488 , \43489 , \43490 , \43491 , \43492 ,
         \43493 , \43494 , \43495 , \43496 , \43497 , \43498 , \43499 , \43500 , \43501 , \43502 ,
         \43503 , \43504 , \43505 , \43506 , \43507 , \43508 , \43509 , \43510 , \43511 , \43512 ,
         \43513 , \43514 , \43515 , \43516 , \43517 , \43518 , \43519 , \43520 , \43521 , \43522 ,
         \43523 , \43524 , \43525 , \43526 , \43527 , \43528 , \43529 , \43530 , \43531 , \43532 ,
         \43533 , \43534 , \43535 , \43536 , \43537 , \43538 , \43539 , \43540 , \43541 , \43542 ,
         \43543 , \43544 , \43545 , \43546 , \43547 , \43548 , \43549 , \43550 , \43551 , \43552 ,
         \43553 , \43554 , \43555 , \43556 , \43557 , \43558 , \43559 , \43560 , \43561 , \43562 ,
         \43563 , \43564 , \43565 , \43566 , \43567 , \43568 , \43569 , \43570 , \43571 , \43572 ,
         \43573 , \43574 , \43575 , \43576 , \43577 , \43578 , \43579 , \43580 , \43581 , \43582 ,
         \43583 , \43584 , \43585 , \43586 , \43587 , \43588 , \43589 , \43590 , \43591 , \43592 ,
         \43593 , \43594 , \43595 , \43596 , \43597 , \43598 , \43599 , \43600 , \43601 , \43602 ,
         \43603 , \43604 , \43605 , \43606 , \43607 , \43608 , \43609 , \43610 , \43611 , \43612 ,
         \43613 , \43614 , \43615 , \43616 , \43617 , \43618 , \43619 , \43620 , \43621 , \43622 ,
         \43623 , \43624 , \43625 , \43626 , \43627 , \43628 , \43629 , \43630 , \43631 , \43632 ,
         \43633 , \43634 , \43635 , \43636 , \43637 , \43638 , \43639 , \43640 , \43641 , \43642 ,
         \43643 , \43644 , \43645 , \43646 , \43647 , \43648 , \43649 , \43650 , \43651 , \43652 ,
         \43653 , \43654 , \43655 , \43656 , \43657 , \43658 , \43659 , \43660 , \43661 , \43662 ,
         \43663 , \43664 , \43665 , \43666 , \43667 , \43668 , \43669 , \43670 , \43671 , \43672 ,
         \43673 , \43674 , \43675 , \43676 , \43677 , \43678 , \43679 , \43680 , \43681 , \43682 ,
         \43683 , \43684 , \43685 , \43686 , \43687 , \43688 , \43689 , \43690 , \43691 , \43692 ,
         \43693 , \43694 , \43695 , \43696 , \43697 , \43698 , \43699 , \43700 , \43701 , \43702 ,
         \43703 , \43704 , \43705 , \43706 , \43707 , \43708 , \43709 , \43710 , \43711 , \43712 ,
         \43713 , \43714 , \43715 , \43716 , \43717 , \43718 , \43719 , \43720 , \43721 , \43722 ,
         \43723 , \43724 , \43725 , \43726 , \43727 , \43728 , \43729 , \43730 , \43731 , \43732 ,
         \43733 , \43734 , \43735 , \43736 , \43737 , \43738 , \43739 , \43740 , \43741 , \43742 ,
         \43743 , \43744 , \43745 , \43746 , \43747 , \43748 , \43749 , \43750 , \43751 , \43752 ,
         \43753 , \43754 , \43755 , \43756 , \43757 , \43758 , \43759 , \43760 , \43761 , \43762 ,
         \43763 , \43764 , \43765 , \43766 , \43767 , \43768 , \43769 , \43770 , \43771 , \43772 ,
         \43773 , \43774 , \43775 , \43776 , \43777 , \43778 , \43779 , \43780 , \43781 , \43782 ,
         \43783 , \43784 , \43785 , \43786 , \43787 , \43788 , \43789 , \43790 , \43791 , \43792 ,
         \43793 , \43794 , \43795 , \43796 , \43797 , \43798 , \43799 , \43800 , \43801 , \43802 ,
         \43803 , \43804 , \43805 , \43806 , \43807 , \43808 , \43809 , \43810 , \43811 , \43812 ,
         \43813 , \43814 , \43815 , \43816 , \43817 , \43818 , \43819 , \43820 , \43821 , \43822 ,
         \43823 , \43824 , \43825 , \43826 , \43827 , \43828 , \43829 , \43830 , \43831 , \43832 ,
         \43833 , \43834 , \43835 , \43836 , \43837 , \43838 , \43839 , \43840 , \43841 , \43842 ,
         \43843 , \43844 , \43845 , \43846 , \43847 , \43848 , \43849 , \43850 , \43851 , \43852 ,
         \43853 , \43854 , \43855 , \43856 , \43857 , \43858 , \43859 , \43860 , \43861 , \43862 ,
         \43863 , \43864 , \43865 , \43866_nRb622 , \43867 , \43868 , \43869 , \43870 , \43871 , \43872 ,
         \43873 , \43874 , \43875 , \43876 , \43877 , \43878 , \43879 , \43880 , \43881 , \43882 ,
         \43883 , \43884 , \43885 , \43886 , \43887 , \43888 , \43889 , \43890 , \43891 , \43892 ,
         \43893 , \43894 , \43895 , \43896 , \43897 , \43898 , \43899 , \43900 , \43901 , \43902 ,
         \43903 , \43904 , \43905 , \43906 , \43907 , \43908 , \43909 , \43910 , \43911 , \43912 ,
         \43913 , \43914 , \43915 , \43916 , \43917 , \43918 , \43919 , \43920 , \43921 , \43922 ,
         \43923 , \43924 , \43925 , \43926 , \43927 , \43928 , \43929 , \43930 , \43931 , \43932 ,
         \43933 , \43934 , \43935 , \43936 , \43937 , \43938 , \43939 , \43940 , \43941 , \43942 ,
         \43943 , \43944 , \43945 , \43946 , \43947 , \43948 , \43949 , \43950 , \43951 , \43952 ,
         \43953 , \43954 , \43955 , \43956 , \43957 , \43958 , \43959 , \43960 , \43961 , \43962 ,
         \43963 , \43964 , \43965 , \43966 , \43967 , \43968 , \43969 , \43970 , \43971 , \43972 ,
         \43973 , \43974 , \43975 , \43976 , \43977 , \43978 , \43979 , \43980 , \43981 , \43982 ,
         \43983 , \43984 , \43985 , \43986 , \43987 , \43988 , \43989 , \43990 , \43991 , \43992 ,
         \43993 , \43994 , \43995 , \43996 , \43997 , \43998 , \43999 , \44000 , \44001 , \44002 ,
         \44003 , \44004 , \44005 , \44006 , \44007 , \44008 , \44009 , \44010 , \44011 , \44012 ,
         \44013 , \44014 , \44015 , \44016 , \44017 , \44018 , \44019 , \44020 , \44021 , \44022 ,
         \44023 , \44024 , \44025 , \44026 , \44027 , \44028 , \44029 , \44030 , \44031 , \44032 ,
         \44033 , \44034 , \44035 , \44036 , \44037 , \44038 , \44039 , \44040 , \44041 , \44042 ,
         \44043 , \44044 , \44045 , \44046 , \44047 , \44048 , \44049 , \44050 , \44051 , \44052 ,
         \44053 , \44054 , \44055 , \44056 , \44057 , \44058 , \44059 , \44060 , \44061 , \44062 ,
         \44063 , \44064 , \44065 , \44066 , \44067 , \44068 , \44069 , \44070 , \44071 , \44072 ,
         \44073 , \44074 , \44075 , \44076 , \44077 , \44078 , \44079 , \44080 , \44081 , \44082 ,
         \44083 , \44084 , \44085 , \44086 , \44087 , \44088 , \44089 , \44090 , \44091 , \44092 ,
         \44093 , \44094 , \44095 , \44096 , \44097 , \44098 , \44099 , \44100 , \44101 , \44102 ,
         \44103 , \44104 , \44105 , \44106 , \44107 , \44108 , \44109 , \44110 , \44111 , \44112 ,
         \44113 , \44114 , \44115 , \44116 , \44117 , \44118 , \44119 , \44120 , \44121 , \44122 ,
         \44123 , \44124 , \44125 , \44126 , \44127 , \44128 , \44129 , \44130 , \44131 , \44132 ,
         \44133 , \44134 , \44135 , \44136 , \44137 , \44138 , \44139 , \44140 , \44141 , \44142 ,
         \44143 , \44144 , \44145 , \44146 , \44147 , \44148 , \44149 , \44150 , \44151 , \44152 ,
         \44153 , \44154 , \44155 , \44156 , \44157 , \44158 , \44159 , \44160 , \44161 , \44162 ,
         \44163 , \44164 , \44165 , \44166 , \44167 , \44168 , \44169 , \44170 , \44171 , \44172 ,
         \44173 , \44174 , \44175 , \44176 , \44177 , \44178 , \44179 , \44180 , \44181 , \44182 ,
         \44183 , \44184 , \44185 , \44186 , \44187 , \44188 , \44189 , \44190 , \44191 , \44192 ,
         \44193 , \44194 , \44195 , \44196 , \44197 , \44198 , \44199 , \44200 , \44201 , \44202 ,
         \44203 , \44204 , \44205 , \44206 , \44207 , \44208 , \44209 , \44210 , \44211 , \44212 ,
         \44213 , \44214 , \44215 , \44216 , \44217 , \44218 , \44219 , \44220 , \44221 , \44222 ,
         \44223 , \44224 , \44225 , \44226 , \44227 , \44228 , \44229 , \44230 , \44231 , \44232 ,
         \44233 , \44234 , \44235 , \44236 , \44237 , \44238 , \44239 , \44240 , \44241 , \44242_nRb5ec ,
         \44243 , \44244 , \44245 , \44246 , \44247 , \44248 , \44249 , \44250 , \44251 , \44252 ,
         \44253 , \44254 , \44255 , \44256 , \44257 , \44258 , \44259 , \44260 , \44261 , \44262 ,
         \44263 , \44264 , \44265 , \44266 , \44267 , \44268 , \44269 , \44270 , \44271 , \44272 ,
         \44273 , \44274 , \44275 , \44276 , \44277 , \44278 , \44279 , \44280 , \44281 , \44282 ,
         \44283 , \44284 , \44285 , \44286 , \44287 , \44288 , \44289 , \44290 , \44291 , \44292 ,
         \44293 , \44294 , \44295 , \44296 , \44297 , \44298 , \44299 , \44300 , \44301 , \44302 ,
         \44303 , \44304 , \44305 , \44306 , \44307 , \44308 , \44309 , \44310 , \44311 , \44312 ,
         \44313 , \44314 , \44315 , \44316 , \44317 , \44318 , \44319 , \44320 , \44321 , \44322 ,
         \44323 , \44324 , \44325 , \44326 , \44327 , \44328 , \44329 , \44330 , \44331 , \44332 ,
         \44333 , \44334 , \44335 , \44336 , \44337 , \44338 , \44339 , \44340 , \44341 , \44342 ,
         \44343 , \44344 , \44345 , \44346 , \44347 , \44348 , \44349 , \44350 , \44351 , \44352 ,
         \44353 , \44354 , \44355 , \44356 , \44357 , \44358 , \44359 , \44360 , \44361 , \44362 ,
         \44363 , \44364 , \44365 , \44366 , \44367 , \44368 , \44369 , \44370 , \44371 , \44372 ,
         \44373 , \44374 , \44375 , \44376 , \44377 , \44378 , \44379 , \44380 , \44381 , \44382 ,
         \44383 , \44384 , \44385 , \44386 , \44387 , \44388 , \44389 , \44390 , \44391 , \44392 ,
         \44393 , \44394 , \44395 , \44396 , \44397 , \44398 , \44399 , \44400 , \44401 , \44402 ,
         \44403 , \44404 , \44405 , \44406 , \44407 , \44408 , \44409 , \44410 , \44411 , \44412 ,
         \44413 , \44414 , \44415 , \44416 , \44417 , \44418 , \44419 , \44420 , \44421 , \44422 ,
         \44423 , \44424 , \44425 , \44426 , \44427 , \44428 , \44429 , \44430_nRb5a9 , \44431 , \44432 ,
         \44433 , \44434 , \44435 , \44436 , \44437 , \44438 , \44439 , \44440 , \44441 , \44442 ,
         \44443 , \44444 , \44445 , \44446 , \44447 , \44448 , \44449 , \44450 , \44451 , \44452 ,
         \44453 , \44454 , \44455 , \44456 , \44457 , \44458 , \44459 , \44460 , \44461 , \44462 ,
         \44463 , \44464 , \44465 , \44466 , \44467 , \44468 , \44469 , \44470 , \44471 , \44472 ,
         \44473 , \44474 , \44475 , \44476 , \44477 , \44478 , \44479 , \44480 , \44481 , \44482 ,
         \44483 , \44484 , \44485 , \44486 , \44487 , \44488 , \44489 , \44490 , \44491 , \44492 ,
         \44493 , \44494 , \44495 , \44496 , \44497 , \44498 , \44499 , \44500 , \44501 , \44502 ,
         \44503 , \44504 , \44505 , \44506 , \44507 , \44508 , \44509 , \44510 , \44511 , \44512 ,
         \44513 , \44514 , \44515 , \44516 , \44517 , \44518 , \44519 , \44520 , \44521 , \44522 ,
         \44523 , \44524 , \44525 , \44526 , \44527 , \44528 , \44529 , \44530 , \44531 , \44532 ,
         \44533 , \44534 , \44535 , \44536 , \44537 , \44538 , \44539 , \44540 , \44541 , \44542 ,
         \44543 , \44544 , \44545 , \44546 , \44547 , \44548 , \44549 , \44550 , \44551 , \44552 ,
         \44553 , \44554 , \44555 , \44556 , \44557 , \44558 , \44559 , \44560 , \44561 , \44562 ,
         \44563 , \44564 , \44565 , \44566 , \44567 , \44568 , \44569 , \44570 , \44571 , \44572 ,
         \44573 , \44574 , \44575 , \44576 , \44577 , \44578 , \44579 , \44580 , \44581 , \44582 ,
         \44583 , \44584 , \44585 , \44586 , \44587 , \44588 , \44589 , \44590 , \44591 , \44592 ,
         \44593 , \44594 , \44595 , \44596 , \44597 , \44598 , \44599 , \44600 , \44601 , \44602 ,
         \44603 , \44604 , \44605 , \44606 , \44607 , \44608 , \44609 , \44610 , \44611 , \44612 ,
         \44613 , \44614 , \44615 , \44616 , \44617 , \44618 , \44619_nRb55a , \44620 , \44621 , \44622 ,
         \44623 , \44624 , \44625 , \44626 , \44627 , \44628 , \44629 , \44630 , \44631 , \44632 ,
         \44633 , \44634 , \44635 , \44636 , \44637 , \44638 , \44639 , \44640 , \44641 , \44642 ,
         \44643 , \44644 , \44645 , \44646 , \44647 , \44648 , \44649 , \44650 , \44651 , \44652 ,
         \44653 , \44654 , \44655 , \44656 , \44657 , \44658 , \44659 , \44660 , \44661 , \44662 ,
         \44663 , \44664 , \44665 , \44666 , \44667 , \44668 , \44669 , \44670 , \44671 , \44672 ,
         \44673 , \44674 , \44675 , \44676 , \44677 , \44678 , \44679 , \44680 , \44681 , \44682 ,
         \44683 , \44684 , \44685 , \44686 , \44687 , \44688 , \44689 , \44690 , \44691 , \44692 ,
         \44693 , \44694 , \44695 , \44696 , \44697 , \44698 , \44699 , \44700 , \44701 , \44702 ,
         \44703 , \44704 , \44705 , \44706 , \44707 , \44708 , \44709 , \44710 , \44711 , \44712 ,
         \44713 , \44714_nRb500 , \44715 , \44716 , \44717 , \44718 , \44719 , \44720 , \44721 , \44722 ,
         \44723 , \44724 , \44725 , \44726 , \44727 , \44728 , \44729 , \44730 , \44731 , \44732 ,
         \44733 , \44734 , \44735 , \44736 , \44737 , \44738 , \44739 , \44740 , \44741 , \44742 ,
         \44743 , \44744 , \44745 , \44746 , \44747 , \44748 , \44749 , \44750 , \44751 , \44752 ,
         \44753 , \44754 , \44755 , \44756 , \44757 , \44758 , \44759 , \44760 , \44761 , \44762 ,
         \44763 , \44764 , \44765 , \44766 , \44767 , \44768 , \44769 , \44770 , \44771 , \44772 ,
         \44773 , \44774 , \44775 , \44776 , \44777 , \44778 , \44779 , \44780 , \44781 , \44782 ,
         \44783 , \44784 , \44785 , \44786 , \44787 , \44788 , \44789 , \44790 , \44791 , \44792 ,
         \44793 , \44794 , \44795 , \44796 , \44797 , \44798 , \44799 , \44800 , \44801 , \44802 ,
         \44803 , \44804 , \44805 , \44806 , \44807 , \44808 , \44809_nRb49d , \44810 , \44811 , \44812 ,
         \44813 , \44814 , \44815 , \44816 , \44817 , \44818 , \44819 , \44820 , \44821 , \44822 ,
         \44823 , \44824 , \44825 , \44826 , \44827 , \44828 , \44829 , \44830 , \44831 , \44832 ,
         \44833 , \44834 , \44835 , \44836 , \44837 , \44838 , \44839 , \44840 , \44841 , \44842 ,
         \44843 , \44844 , \44845 , \44846 , \44847 , \44848 , \44849 , \44850 , \44851 , \44852 ,
         \44853 , \44854 , \44855 , \44856 , \44857 , \44858 , \44859 , \44860 , \44861 , \44862 ,
         \44863 , \44864 , \44865 , \44866 , \44867 , \44868 , \44869 , \44870 , \44871 , \44872 ,
         \44873 , \44874 , \44875 , \44876 , \44877 , \44878 , \44879 , \44880 , \44881 , \44882 ,
         \44883 , \44884 , \44885 , \44886 , \44887 , \44888 , \44889 , \44890 , \44891 , \44892 ,
         \44893 , \44894 , \44895 , \44896 , \44897 , \44898 , \44899 , \44900 , \44901 , \44902_nRb432 ,
         \44903 , \44904 , \44905 , \44906 , \44907 , \44908 , \44909 , \44910 , \44911 , \44912 ,
         \44913 , \44914 , \44915 , \44916 , \44917 , \44918 , \44919 , \44920 , \44921 , \44922 ,
         \44923 , \44924 , \44925 , \44926 , \44927 , \44928 , \44929 , \44930 , \44931 , \44932 ,
         \44933 , \44934 , \44935 , \44936 , \44937 , \44938 , \44939 , \44940 , \44941 , \44942 ,
         \44943 , \44944 , \44945 , \44946 , \44947 , \44948 , \44949 , \44950 , \44951 , \44952 ,
         \44953 , \44954 , \44955 , \44956 , \44957 , \44958 , \44959 , \44960 , \44961 , \44962 ,
         \44963 , \44964 , \44965 , \44966 , \44967 , \44968 , \44969 , \44970 , \44971 , \44972 ,
         \44973 , \44974 , \44975 , \44976 , \44977 , \44978 , \44979 , \44980 , \44981 , \44982 ,
         \44983 , \44984 , \44985 , \44986 , \44987 , \44988 , \44989 , \44990 , \44991 , \44992 ,
         \44993 , \44994 , \44995_nRb3bb , \44996 , \44997 , \44998 , \44999 , \45000 , \45001 , \45002 ,
         \45003 , \45004 , \45005 , \45006 , \45007 , \45008 , \45009 , \45010 , \45011 , \45012 ,
         \45013 , \45014 , \45015 , \45016 , \45017 , \45018 , \45019 , \45020 , \45021 , \45022 ,
         \45023 , \45024 , \45025 , \45026 , \45027 , \45028 , \45029 , \45030 , \45031 , \45032 ,
         \45033 , \45034 , \45035 , \45036 , \45037 , \45038 , \45039 , \45040 , \45041 , \45042 ,
         \45043 , \45044_nRb33b , \45045 , \45046 , \45047 , \45048 , \45049 , \45050 , \45051 , \45052 ,
         \45053 , \45054 , \45055 , \45056 , \45057 , \45058 , \45059 , \45060 , \45061 , \45062 ,
         \45063 , \45064 , \45065 , \45066 , \45067 , \45068 , \45069 , \45070 , \45071 , \45072 ,
         \45073 , \45074 , \45075 , \45076 , \45077 , \45078 , \45079 , \45080 , \45081 , \45082 ,
         \45083 , \45084 , \45085 , \45086 , \45087 , \45088 , \45089 , \45090 , \45091 , \45092 ,
         \45093_nRb2b1 , \45094 , \45095 , \45096 , \45097 , \45098 , \45099 , \45100 , \45101 , \45102 ,
         \45103 , \45104 , \45105 , \45106 , \45107 , \45108 , \45109 , \45110 , \45111 , \45112 ,
         \45113 , \45114 , \45115 , \45116 , \45117 , \45118 , \45119 , \45120 , \45121 , \45122 ,
         \45123 , \45124 , \45125 , \45126 , \45127 , \45128 , \45129 , \45130 , \45131 , \45132 ,
         \45133 , \45134 , \45135 , \45136 , \45137 , \45138 , \45139 , \45140 , \45141_nRb21b , \45142 ,
         \45143 , \45144 , \45145 , \45146 , \45147 , \45148 , \45149 , \45150 , \45151 , \45152 ,
         \45153 , \45154 , \45155 , \45156 , \45157 , \45158 , \45159 , \45160 , \45161 , \45162 ,
         \45163 , \45164 , \45165 , \45166 , \45167 , \45168 , \45169 , \45170 , \45171 , \45172 ,
         \45173 , \45174 , \45175 , \45176 , \45177 , \45178 , \45179 , \45180 , \45181 , \45182 ,
         \45183 , \45184 , \45185 , \45186 , \45187 , \45188 , \45189_nRb17c , \45190 , \45191 , \45192 ,
         \45193 , \45194 , \45195 , \45196 , \45197 , \45198 , \45199 , \45200 , \45201 , \45202 ,
         \45203 , \45204 , \45205 , \45206 , \45207 , \45208 , \45209 , \45210 , \45211 , \45212 ,
         \45213 , \45214 , \45215 , \45216 , \45217 , \45218 , \45219 , \45220 , \45221 , \45222 ,
         \45223 , \45224 , \45225 , \45226 , \45227 , \45228 , \45229 , \45230 , \45231 , \45232 ,
         \45233 , \45234 , \45235 , \45236 , \45237_nRb0d5 , \45238 , \45239 , \45240 , \45241 , \45242 ,
         \45243 , \45244 , \45245 , \45246 , \45247 , \45248 , \45249 , \45250 , \45251 , \45252 ,
         \45253 , \45254 , \45255 , \45256 , \45257 , \45258 , \45259 , \45260 , \45261 , \45262 ,
         \45263 , \45264 , \45265 , \45266 , \45267 , \45268 , \45269 , \45270 , \45271 , \45272 ,
         \45273 , \45274 , \45275 , \45276 , \45277 , \45278 , \45279 , \45280 , \45281 , \45282 ,
         \45283 , \45284 , \45285_nRb022 , \45286 , \45287 , \45288 , \45289 , \45290 , \45291 , \45292 ,
         \45293 , \45294 , \45295 , \45296 , \45297 , \45298 , \45299 , \45300 , \45301 , \45302 ,
         \45303 , \45304 , \45305 , \45306 , \45307 , \45308 , \45309 , \45310 , \45311 , \45312 ,
         \45313 , \45314 , \45315 , \45316 , \45317 , \45318 , \45319 , \45320 , \45321 , \45322 ,
         \45323 , \45324 , \45325 , \45326 , \45327 , \45328 , \45329 , \45330 , \45331_nRaf66 , \45332 ,
         \45333 , \45334 , \45335 , \45336 , \45337 , \45338 , \45339 , \45340 , \45341 , \45342 ,
         \45343 , \45344 , \45345 , \45346 , \45347 , \45348 , \45349 , \45350 , \45351 , \45352 ,
         \45353 , \45354 , \45355 , \45356 , \45357 , \45358 , \45359 , \45360 , \45361 , \45362 ,
         \45363 , \45364 , \45365 , \45366 , \45367 , \45368 , \45369 , \45370 , \45371 , \45372 ,
         \45373 , \45374 , \45375 , \45376 , \45377_nRaea0 , \45378 , \45379 , \45380 , \45381 , \45382 ,
         \45383 , \45384 , \45385 , \45386 , \45387 , \45388 , \45389 , \45390 , \45391 , \45392 ,
         \45393 , \45394 , \45395 , \45396 , \45397 , \45398 , \45399 , \45400 , \45401 , \45402 ,
         \45403_nRadd0 , \45404 , \45405 , \45406 , \45407 , \45408 , \45409 , \45410 , \45411 , \45412 ,
         \45413 , \45414 , \45415 , \45416 , \45417 , \45418 , \45419 , \45420 , \45421 , \45422 ,
         \45423 , \45424 , \45425 , \45426 , \45427 , \45428 , \45429_nRacf6 , \45430 , \45431 , \45432 ,
         \45433 , \45434 , \45435 , \45436 , \45437 , \45438 , \45439 , \45440 , \45441 , \45442 ,
         \45443 , \45444 , \45445 , \45446 , \45447 , \45448 , \45449 , \45450 , \45451 , \45452 ,
         \45453 , \45454 , \45455_nRac12 , \45456 , \45457 , \45458 , \45459 , \45460 , \45461 , \45462 ,
         \45463 , \45464 , \45465 , \45466 , \45467 , \45468 , \45469 , \45470 , \45471 , \45472 ,
         \45473 , \45474 , \45475 , \45476 , \45477 , \45478 , \45479 , \45480 , \45481_nRab27 , \45482 ,
         \45483 , \45484 , \45485 , \45486 , \45487 , \45488 , \45489 , \45490 , \45491 , \45492 ,
         \45493 , \45494 , \45495 , \45496 , \45497 , \45498 , \45499 , \45500 , \45501 , \45502 ,
         \45503 , \45504 , \45505 , \45506 , \45507_nRaa31 , \45508 , \45509 , \45510 , \45511 , \45512 ,
         \45513 , \45514 , \45515 , \45516 , \45517 , \45518 , \45519 , \45520 , \45521 , \45522 ,
         \45523 , \45524 , \45525 , \45526 , \45527 , \45528 , \45529 , \45530 , \45531 , \45532 ,
         \45533_nRa92e , \45534 , \45535 , \45536 , \45537 , \45538 , \45539 , \45540 , \45541 , \45542 ,
         \45543 , \45544 , \45545 , \45546 , \45547 , \45548 , \45549 , \45550 , \45551 , \45552 ,
         \45553 , \45554 , \45555 , \45556 , \45557 , \45558_nRa820 , \45559 , \45560 , \45561 , \45562 ,
         \45563 , \45564 , \45565 , \45566 , \45567 , \45568 , \45569 , \45570 , \45571 , \45572 ,
         \45573 , \45574 , \45575 , \45576 , \45577 , \45578 , \45579 , \45580 , \45581 , \45582 ,
         \45583_nRa706 , \45584 , \45585 , \45586 , \45587 , \45588 , \45589 , \45590 , \45591 , \45592 ,
         \45593 , \45594 , \45595 , \45596 , \45597 , \45598 , \45599 , \45600 , \45601 , \45602 ,
         \45603 , \45604 , \45605 , \45606 , \45607 , \45608_nRa5e5 , \45609 , \45610 , \45611 , \45612 ,
         \45613 , \45614 , \45615 , \45616 , \45617 , \45618 , \45619 , \45620 , \45621 , \45622 ,
         \45623 , \45624 , \45625 , \45626 , \45627 , \45628 , \45629 , \45630 , \45631 , \45632 ,
         \45633_nRa4bb , \45634 , \45635 , \45636 , \45637 , \45638 , \45639 , \45640 , \45641 , \45642 ,
         \45643 , \45644 , \45645 , \45646 , \45647 , \45648 , \45649 , \45650 , \45651 , \45652 ,
         \45653 , \45654 , \45655 , \45656 , \45657 , \45658_nRa384 , \45659 , \45660 , \45661 , \45662 ,
         \45663 , \45664 , \45665 , \45666 , \45667 , \45668 , \45669 , \45670 , \45671 , \45672 ,
         \45673 , \45674 , \45675 , \45676 , \45677 , \45678 , \45679 , \45680 , \45681 , \45682 ,
         \45683_nRa241 , \45684 , \45685 , \45686 , \45687 , \45688 , \45689 , \45690 , \45691 , \45692 ,
         \45693 , \45694 , \45695 , \45696 , \45697 , \45698 , \45699 , \45700 , \45701 , \45702 ,
         \45703 , \45704 , \45705 , \45706 , \45707 , \45708_nRa0f3 , \45709 , \45710 , \45711 , \45712 ,
         \45713 , \45714 , \45715 , \45716 , \45717 , \45718 , \45719 , \45720 , \45721 , \45722 ,
         \45723 , \45724 , \45725 , \45726 , \45727 , \45728 , \45729 , \45730 , \45731 , \45732 ,
         \45733_nR9f9c , \45734 , \45735 , \45736 , \45737 , \45738 , \45739 , \45740 , \45741 , \45742 ,
         \45743 , \45744 , \45745 , \45746 , \45747 , \45748 , \45749 , \45750 , \45751 , \45752 ,
         \45753 , \45754 , \45755 , \45756_nR9e40 , \45757 , \45758 , \45759 , \45760 , \45761 , \45762 ,
         \45763 , \45764 , \45765 , \45766 , \45767 , \45768 , \45769 , \45770 , \45771 , \45772 ,
         \45773 , \45774 , \45775 , \45776 , \45777 , \45778 , \45779_nR9cdd , \45780 , \45781 , \45782 ,
         \45783 , \45784 , \45785 , \45786 , \45787 , \45788 , \45789 , \45790 , \45791 , \45792 ,
         \45793 , \45794_nR9b72 , \45795 , \45796 , \45797 , \45798 , \45799 , \45800 , \45801 , \45802 ,
         \45803 , \45804 , \45805 , \45806 , \45807 , \45808 , \45809_nR99fc , \45810 , \45811 , \45812 ,
         \45813 , \45814 , \45815 , \45816 , \45817 , \45818 , \45819 , \45820 , \45821 , \45822 ,
         \45823 , \45824_nR9879 , \45825 , \45826 , \45827 , \45828 , \45829 , \45830 , \45831 , \45832 ,
         \45833 , \45834 , \45835 , \45836 , \45837 , \45838 , \45839_nR96ea , \45840 , \45841 , \45842 ,
         \45843 , \45844 , \45845 , \45846 , \45847 , \45848 , \45849 , \45850 , \45851 , \45852 ,
         \45853 , \45854_nR9552 , \45855 , \45856 , \45857 , \45858 , \45859 , \45860 , \45861 , \45862 ,
         \45863 , \45864 , \45865 , \45866 , \45867 , \45868 , \45869_nR93b0 , \45870 , \45871 , \45872 ,
         \45873 , \45874 , \45875 , \45876 , \45877 , \45878 , \45879 , \45880 , \45881 , \45882 ,
         \45883 , \45884_nR9204 , \45885 , \45886 , \45887 , \45888 , \45889 , \45890 , \45891 , \45892 ,
         \45893 , \45894 , \45895 , \45896 , \45897 , \45898 , \45899_nR904e , \45900 , \45901 , \45902 ,
         \45903 , \45904 , \45905 , \45906 , \45907 , \45908 , \45909 , \45910 , \45911 , \45912 ,
         \45913 , \45914_nR8e8c , \45915 , \45916 , \45917 , \45918 , \45919 , \45920 , \45921 , \45922 ,
         \45923 , \45924 , \45925 , \45926 , \45927 , \45928 , \45929_nR8cbe , \45930 , \45931 , \45932 ,
         \45933 , \45934 , \45935 , \45936 , \45937 , \45938 , \45939 , \45940 , \45941 , \45942 ,
         \45943 , \45944_nR8ae6 , \45945 , \45946 , \45947 , \45948 , \45949 , \45950 , \45951 , \45952 ,
         \45953 , \45954 , \45955 , \45956 , \45957 , \45958 , \45959_nR8903 , \45960 , \45961 , \45962 ,
         \45963 , \45964 , \45965 , \45966 , \45967 , \45968 , \45969 , \45970 , \45971 , \45972 ,
         \45973 , \45974_nR8717 , \45975 , \45976 , \45977 , \45978 , \45979 , \45980 , \45981 , \45982 ,
         \45983 , \45984 , \45985 , \45986 , \45987 , \45988 , \45989_nR8521 , \45990 , \45991 , \45992 ,
         \45993 , \45994 , \45995 , \45996 , \45997 , \45998 , \45999 , \46000 , \46001 , \46002 ,
         \46003_nR831f , \46004 , \46005 , \46006 , \46007 , \46008 , \46009 , \46010 , \46011 , \46012 ,
         \46013 , \46014 , \46015 , \46016 , \46017_nR8114 , \46018 , \46019 , \46020 , \46021 , \46022 ,
         \46023 , \46024 , \46025 , \46026 , \46027 , \46028 , \46029 , \46030 , \46031_nR7f04 , \46032 ,
         \46033 , \46034 , \46035 , \46036 , \46037 , \46038 , \46039 , \46040 , \46041 , \46042 ,
         \46043 , \46044 , \46045_nR7ced , \46046 , \46047 , \46048 , \46049 , \46050 , \46051 , \46052 ,
         \46053 , \46054 , \46055 , \46056 , \46057 , \46058 , \46059_nR7acb , \46060 , \46061 , \46062 ,
         \46063 , \46064 , \46065 , \46066 , \46067 , \46068 , \46069 , \46070 , \46071 , \46072 ,
         \46073_nR789f , \46074 , \46075 , \46076 , \46077 , \46078 , \46079 , \46080 , \46081 , \46082 ,
         \46083 , \46084 , \46085 , \46086 , \46087_nR766c , \46088 , \46089 , \46090 , \46091 , \46092 ,
         \46093 , \46094 , \46095 , \46096 , \46097 , \46098 , \46099 , \46100 , \46101_nR742e , \46102 ,
         \46103 , \46104 , \46105 , \46106 , \46107 , \46108 , \46109 , \46110 , \46111 , \46112 ,
         \46113 , \46114 , \46115_nR71e6 , \46116 , \46117 , \46118 , \46119 , \46120 , \46121 , \46122 ,
         \46123 , \46124 , \46125 , \46126 , \46127 , \46128 , \46129_nR6f94 , \46130 , \46131 , \46132 ,
         \46133 , \46134 , \46135 , \46136 , \46137 , \46138 , \46139 , \46140 , \46141 , \46142 ,
         \46143_nR6d35 , \46144 , \46145 , \46146 , \46147 , \46148 , \46149 , \46150 , \46151 , \46152 ,
         \46153 , \46154 , \46155 , \46156 , \46157_nR6aca , \46158 , \46159 , \46160 , \46161 , \46162 ,
         \46163 , \46164 , \46165 , \46166 , \46167 , \46168 , \46169 , \46170 , \46171_nR6854 , \46172 ,
         \46173 , \46174 , \46175 , \46176 , \46177 , \46178 , \46179 , \46180 , \46181 , \46182 ,
         \46183 , \46184 , \46185_nR65d5 , \46186 , \46187 , \46188 , \46189 , \46190 , \46191 , \46192 ,
         \46193 , \46194 , \46195 , \46196 , \46197 , \46198 , \46199_nR634e , \46200 , \46201 , \46202 ,
         \46203 , \46204 , \46205 , \46206 , \46207 , \46208 , \46209 , \46210 , \46211 , \46212 ,
         \46213_nR60c1 , \46214 , \46215 , \46216 , \46217 , \46218 , \46219 , \46220 , \46221 , \46222 ,
         \46223_nR5e2f , \46224 , \46225 , \46226 , \46227 , \46228 , \46229 , \46230 , \46231 , \46232 ,
         \46233_nR5ba1 , \46234 , \46235 , \46236 , \46237 , \46238 , \46239 , \46240 , \46241_nR590c , \46242 ,
         \46243 , \46244 , \46245 , \46246 , \46247 , \46248 , \46249_nR5671 , \46250 , \46251 , \46252 ,
         \46253 , \46254 , \46255 , \46256 , \46257_nR53dc , \46258 , \46259 , \46260 , \46261 , \46262 ,
         \46263 , \46264 , \46265_nR5155 , \46266 , \46267 , \46268 , \46269 , \46270 , \46271 , \46272 ,
         \46273_nR4ed4 , \46274 , \46275 , \46276 , \46277 , \46278 , \46279 , \46280 , \46281_nR4c61 , \46282 ,
         \46283 , \46284 , \46285 , \46286 , \46287 , \46288 , \46289_nR49f4 , \46290 , \46291 , \46292 ,
         \46293 , \46294 , \46295 , \46296 , \46297_nR4795 , \46298 , \46299 , \46300 , \46301 , \46302 ,
         \46303 , \46304 , \46305_nR453c , \46306 , \46307 , \46308 , \46309 , \46310 , \46311 , \46312 ,
         \46313_nR42f1 , \46314 , \46315 , \46316 , \46317 , \46318 , \46319 , \46320 , \46321_nR40ac , \46322 ,
         \46323 , \46324 , \46325 , \46326 , \46327 , \46328 , \46329_nR3e75 , \46330 , \46331 , \46332 ,
         \46333 , \46334 , \46335 , \46336 , \46337_nR3c44 , \46338 , \46339 , \46340 , \46341 , \46342 ,
         \46343 , \46344 , \46345_nR3a21 , \46346 , \46347 , \46348 , \46349 , \46350 , \46351 , \46352 ,
         \46353_nR3804 , \46354 , \46355 , \46356 , \46357 , \46358 , \46359 , \46360 , \46361_nR35f4 , \46362 ,
         \46363 , \46364 , \46365 , \46366 , \46367 , \46368 , \46369_nR33ea , \46370 , \46371 , \46372 ,
         \46373 , \46374 , \46375 , \46376 , \46377_nR31ee , \46378 , \46379 , \46380 , \46381 , \46382 ,
         \46383 , \46384 , \46385_nR2ff8 , \46386 , \46387 , \46388 , \46389 , \46390 , \46391 , \46392 ,
         \46393_nR2e10 , \46394 , \46395 , \46396 , \46397 , \46398 , \46399 , \46400 , \46401_nR2c28 , \46402 ,
         \46403 , \46404 , \46405 , \46406 , \46407 , \46408 , \46409_nR2a56 , \46410 , \46411 , \46412 ,
         \46413 , \46414 , \46415 , \46416 , \46417_nR2888 , \46418 , \46419 , \46420 , \46421 , \46422 ,
         \46423 , \46424 , \46425_nR26c9 , \46426 , \46427 , \46428 , \46429 , \46430 , \46431 , \46432 ,
         \46433_nR2510 , \46434 , \46435 , \46436 , \46437 , \46438 , \46439 , \46440 , \46441_nR2365 , \46442 ,
         \46443 , \46444 , \46445 , \46446 , \46447 , \46448 , \46449_nR21c0 , \46450 , \46451 , \46452 ,
         \46453 , \46454 , \46455 , \46456 , \46457_nR2029 , \46458 , \46459 , \46460 , \46461 , \46462 ,
         \46463 , \46464 , \46465_nR1e98 , \46466 , \46467 , \46468 , \46469 , \46470 , \46471 , \46472 ,
         \46473_nR1d15 , \46474 , \46475 , \46476 , \46477 , \46478 , \46479 , \46480 , \46481_nR1b98 , \46482 ,
         \46483 , \46484 , \46485 , \46486 , \46487 , \46488 , \46489_nR1a2b , \46490 , \46491 , \46492 ,
         \46493 , \46494 , \46495 , \46496 , \46497_nR18c4 , \46498 , \46499 , \46500 , \46501 , \46502 ,
         \46503 , \46504 , \46505_nR176b , \46506 , \46507 , \46508 , \46509 , \46510 , \46511 , \46512 ,
         \46513_nR1618 , \46514 , \46515 , \46516 , \46517 , \46518 , \46519 , \46520 , \46521_nR14d3 , \46522 ,
         \46523 , \46524 , \46525 , \46526 , \46527 , \46528 , \46529_nR1394 , \46530 , \46531 , \46532 ,
         \46533 , \46534 , \46535 , \46536 , \46537_nR1263 , \46538 , \46539 , \46540 , \46541 , \46542 ,
         \46543 , \46544 , \46545_nR1138 , \46546 , \46547 , \46548 , \46549 , \46550 , \46551 , \46552 ,
         \46553_nR101b , \46554 , \46555 , \46556 , \46557 , \46558 , \46559 , \46560 , \46561_nRf04 , \46562 ,
         \46563 , \46564 , \46565 , \46566 , \46567 , \46568 , \46569_nRdfb , \46570 , \46571 , \46572 ,
         \46573 , \46574 , \46575 , \46576 , \46577_nRcf8 , \46578 , \46579 , \46580 , \46581 , \46582 ,
         \46583 , \46584 , \46585_nRc03 , \46586 , \46587 , \46588 , \46589 , \46590 , \46591 , \46592 ,
         \46593_nRb14 , \46594 , \46595 , \46596 , \46597 , \46598 , \46599 , \46600 , \46601_nRa33 , \46602 ,
         \46603 , \46604 , \46605 , \46606 , \46607 , \46608 , \46609_nR958 , \46610 , \46611 , \46612 ,
         \46613 , \46614 , \46615 , \46616 , \46617_nR88f , \46618 , \46619 , \46620 , \46621 , \46622 ,
         \46623 , \46624 , \46625_nR7cc , \46626 , \46627 , \46628 , \46629 , \46630 , \46631 , \46632 ,
         \46633_nR717 , \46634 , \46635 , \46636 , \46637 , \46638 , \46639 , \46640 , \46641_nR668 , \46642 ,
         \46643 , \46644 , \46645 , \46646 , \46647 , \46648 , \46649_nR5c6 , \46650 , \46651 , \46652 ,
         \46653 , \46654 , \46655 , \46656 , \46657_nR52a , \46658 , \46659 , \46660 , \46661 , \46662 ,
         \46663 , \46664 , \46665_nR49d , \46666 , \46667 , \46668 , \46669 , \46670 , \46671 , \46672 ,
         \46673_nR416 , \46674 , \46675 , \46676 , \46677 , \46678 , \46679 , \46680 , \46681_nR39f , \46682 ;
buf \U$labaj4707 ( R_c2_9969708, \43867 );
buf \U$labaj4708 ( R_c3_99697b0, \44243 );
buf \U$labaj4709 ( R_c4_9969858, \44431 );
buf \U$labaj4710 ( R_c5_9969900, \44620 );
buf \U$labaj4711 ( R_c6_99699a8, \44715 );
buf \U$labaj4712 ( R_c7_9969a50, \44810 );
buf \U$labaj4713 ( R_c8_9969af8, \44903 );
buf \U$labaj4714 ( R_c9_9969ba0, \44996 );
buf \U$labaj4715 ( R_ca_9969c48, \45045 );
buf \U$labaj4716 ( R_cb_9969cf0, \45094 );
buf \U$labaj4717 ( R_cc_9969d98, \45142 );
buf \U$labaj4718 ( R_cd_9969e40, \45190 );
buf \U$labaj4719 ( R_ce_9969ee8, \45238 );
buf \U$labaj4720 ( R_cf_9969f90, \45286 );
buf \U$labaj4721 ( R_d0_996a038, \45332 );
buf \U$labaj4722 ( R_d1_996a0e0, \45378 );
buf \U$labaj4723 ( R_d2_996a188, \45404 );
buf \U$labaj4724 ( R_d3_996a230, \45430 );
buf \U$labaj4725 ( R_d4_996a2d8, \45456 );
buf \U$labaj4726 ( R_d5_996a380, \45482 );
buf \U$labaj4727 ( R_d6_996a428, \45508 );
buf \U$labaj4728 ( R_d7_996a4d0, \45534 );
buf \U$labaj4729 ( R_d8_996a578, \45559 );
buf \U$labaj4730 ( R_d9_996a620, \45584 );
buf \U$labaj4731 ( R_da_996a6c8, \45609 );
buf \U$labaj4732 ( R_db_996a770, \45634 );
buf \U$labaj4733 ( R_dc_996a818, \45659 );
buf \U$labaj4734 ( R_dd_996a8c0, \45684 );
buf \U$labaj4735 ( R_de_996a968, \45709 );
buf \U$labaj4736 ( R_df_996aa10, \45734 );
buf \U$labaj4737 ( R_e0_996aab8, \45757 );
buf \U$labaj4738 ( R_e1_996ab60, \45780 );
buf \U$labaj4739 ( R_e2_996ac08, \45795 );
buf \U$labaj4740 ( R_e3_996acb0, \45810 );
buf \U$labaj4741 ( R_e4_996ad58, \45825 );
buf \U$labaj4742 ( R_e5_996ae00, \45840 );
buf \U$labaj4743 ( R_e6_996aea8, \45855 );
buf \U$labaj4744 ( R_e7_996af50, \45870 );
buf \U$labaj4745 ( R_e8_996aff8, \45885 );
buf \U$labaj4746 ( R_e9_996b0a0, \45900 );
buf \U$labaj4747 ( R_ea_996b148, \45915 );
buf \U$labaj4748 ( R_eb_996b1f0, \45930 );
buf \U$labaj4749 ( R_ec_996b298, \45945 );
buf \U$labaj4750 ( R_ed_996b340, \45960 );
buf \U$labaj4751 ( R_ee_996b3e8, \45975 );
buf \U$labaj4752 ( R_ef_996b490, \45990 );
buf \U$labaj4753 ( R_f0_996b538, \46004 );
buf \U$labaj4754 ( R_f1_996b5e0, \46018 );
buf \U$labaj4755 ( R_f2_996b688, \46032 );
buf \U$labaj4756 ( R_f3_996b730, \46046 );
buf \U$labaj4757 ( R_f4_996b7d8, \46060 );
buf \U$labaj4758 ( R_f5_996b880, \46074 );
buf \U$labaj4759 ( R_f6_996b928, \46088 );
buf \U$labaj4760 ( R_f7_996b9d0, \46102 );
buf \U$labaj4761 ( R_f8_996ba78, \46116 );
buf \U$labaj4762 ( R_f9_996bb20, \46130 );
buf \U$labaj4763 ( R_fa_996bbc8, \46144 );
buf \U$labaj4764 ( R_fb_996bc70, \46158 );
buf \U$labaj4765 ( R_fc_996bd18, \46172 );
buf \U$labaj4766 ( R_fd_996bdc0, \46186 );
buf \U$labaj4767 ( R_fe_996be68, \46200 );
buf \U$labaj4768 ( R_ff_996bf10, \46214 );
buf \U$labaj4769 ( R_100_996bfb8, \46224 );
buf \U$labaj4770 ( R_101_996c060, \46234 );
buf \U$labaj4771 ( R_102_996c108, \46242 );
buf \U$labaj4772 ( R_103_996c1b0, \46250 );
buf \U$labaj4773 ( R_104_996c258, \46258 );
buf \U$labaj4774 ( R_105_996c300, \46266 );
buf \U$labaj4775 ( R_106_996c3a8, \46274 );
buf \U$labaj4776 ( R_107_996c450, \46282 );
buf \U$labaj4777 ( R_108_996c4f8, \46290 );
buf \U$labaj4778 ( R_109_996c5a0, \46298 );
buf \U$labaj4779 ( R_10a_996c648, \46306 );
buf \U$labaj4780 ( R_10b_996c6f0, \46314 );
buf \U$labaj4781 ( R_10c_996c798, \46322 );
buf \U$labaj4782 ( R_10d_996c840, \46330 );
buf \U$labaj4783 ( R_10e_996c8e8, \46338 );
buf \U$labaj4784 ( R_10f_996c990, \46346 );
buf \U$labaj4785 ( R_110_996ca38, \46354 );
buf \U$labaj4786 ( R_111_996cae0, \46362 );
buf \U$labaj4787 ( R_112_996cb88, \46370 );
buf \U$labaj4788 ( R_113_996cc30, \46378 );
buf \U$labaj4789 ( R_114_996ccd8, \46386 );
buf \U$labaj4790 ( R_115_996cd80, \46394 );
buf \U$labaj4791 ( R_116_996ce28, \46402 );
buf \U$labaj4792 ( R_117_996ced0, \46410 );
buf \U$labaj4793 ( R_118_996cf78, \46418 );
buf \U$labaj4794 ( R_119_996d020, \46426 );
buf \U$labaj4795 ( R_11a_996d0c8, \46434 );
buf \U$labaj4796 ( R_11b_996d170, \46442 );
buf \U$labaj4797 ( R_11c_996d218, \46450 );
buf \U$labaj4798 ( R_11d_996d2c0, \46458 );
buf \U$labaj4799 ( R_11e_996d368, \46466 );
buf \U$labaj4800 ( R_11f_996d410, \46474 );
buf \U$labaj4801 ( R_120_996d4b8, \46482 );
buf \U$labaj4802 ( R_121_996d560, \46490 );
buf \U$labaj4803 ( R_122_996d608, \46498 );
buf \U$labaj4804 ( R_123_996d6b0, \46506 );
buf \U$labaj4805 ( R_124_996d758, \46514 );
buf \U$labaj4806 ( R_125_996d800, \46522 );
buf \U$labaj4807 ( R_126_996d8a8, \46530 );
buf \U$labaj4808 ( R_127_996d950, \46538 );
buf \U$labaj4809 ( R_128_996d9f8, \46546 );
buf \U$labaj4810 ( R_129_996daa0, \46554 );
buf \U$labaj4811 ( R_12a_996db48, \46562 );
buf \U$labaj4812 ( R_12b_996dbf0, \46570 );
buf \U$labaj4813 ( R_12c_996dc98, \46578 );
buf \U$labaj4814 ( R_12d_996dd40, \46586 );
buf \U$labaj4815 ( R_12e_996dde8, \46594 );
buf \U$labaj4816 ( R_12f_996de90, \46602 );
buf \U$labaj4817 ( R_130_996df38, \46610 );
buf \U$labaj4818 ( R_131_996dfe0, \46618 );
buf \U$labaj4819 ( R_132_996e088, \46626 );
buf \U$labaj4820 ( R_133_996e130, \46634 );
buf \U$labaj4821 ( R_134_996e1d8, \46642 );
buf \U$labaj4822 ( R_135_996e280, \46650 );
buf \U$labaj4823 ( R_136_996e328, \46658 );
buf \U$labaj4824 ( R_137_996e3d0, \46666 );
buf \U$labaj4825 ( R_138_996e478, \46674 );
buf \U$labaj4826 ( R_139_996e520, \46682 );
buf \U$1 ( \316 , RIc0c7950_66);
buf \U$2 ( \317 , RIc0c9750_2);
buf \U$3 ( \318 , RIc0c96d8_3);
xor \U$4 ( \319 , \317 , \318 );
buf \U$5 ( \320 , RIc0c9660_4);
xor \U$6 ( \321 , \318 , \320 );
not \U$7 ( \322 , \321 );
and \U$8 ( \323 , \319 , \322 );
and \U$9 ( \324 , \316 , \323 );
not \U$10 ( \325 , \324 );
and \U$11 ( \326 , \318 , \320 );
not \U$12 ( \327 , \326 );
and \U$13 ( \328 , \317 , \327 );
xnor \U$14 ( \329 , \325 , \328 );
buf \U$15 ( \330 , RIc0c78d8_67);
and \U$16 ( \331 , \330 , \317 );
or \U$17 ( \332 , \329 , \331 );
not \U$18 ( \333 , \328 );
xor \U$19 ( \334 , \332 , \333 );
and \U$20 ( \335 , \316 , \317 );
xor \U$21 ( \336 , \334 , \335 );
buf \U$22 ( \337 , RIc0c95e8_5);
buf \U$23 ( \338 , RIc0c9570_6);
and \U$24 ( \339 , \337 , \338 );
not \U$25 ( \340 , \339 );
and \U$26 ( \341 , \320 , \340 );
not \U$27 ( \342 , \341 );
and \U$28 ( \343 , \330 , \323 );
and \U$29 ( \344 , \316 , \321 );
nor \U$30 ( \345 , \343 , \344 );
xnor \U$31 ( \346 , \345 , \328 );
and \U$32 ( \347 , \342 , \346 );
buf \U$33 ( \348 , RIc0c7860_68);
and \U$34 ( \349 , \348 , \317 );
and \U$35 ( \350 , \346 , \349 );
and \U$36 ( \351 , \342 , \349 );
or \U$37 ( \352 , \347 , \350 , \351 );
xnor \U$38 ( \353 , \329 , \331 );
and \U$39 ( \354 , \352 , \353 );
xor \U$40 ( \355 , \336 , \354 );
xor \U$41 ( \356 , \352 , \353 );
xor \U$42 ( \357 , \320 , \337 );
xor \U$43 ( \358 , \337 , \338 );
not \U$44 ( \359 , \358 );
and \U$45 ( \360 , \357 , \359 );
and \U$46 ( \361 , \316 , \360 );
not \U$47 ( \362 , \361 );
xnor \U$48 ( \363 , \362 , \341 );
and \U$49 ( \364 , \348 , \323 );
and \U$50 ( \365 , \330 , \321 );
nor \U$51 ( \366 , \364 , \365 );
xnor \U$52 ( \367 , \366 , \328 );
and \U$53 ( \368 , \363 , \367 );
buf \U$54 ( \369 , RIc0c77e8_69);
and \U$55 ( \370 , \369 , \317 );
and \U$56 ( \371 , \367 , \370 );
and \U$57 ( \372 , \363 , \370 );
or \U$58 ( \373 , \368 , \371 , \372 );
buf \U$59 ( \374 , RIc0c94f8_7);
buf \U$60 ( \375 , RIc0c9480_8);
and \U$61 ( \376 , \374 , \375 );
not \U$62 ( \377 , \376 );
and \U$63 ( \378 , \338 , \377 );
not \U$64 ( \379 , \378 );
and \U$65 ( \380 , \330 , \360 );
and \U$66 ( \381 , \316 , \358 );
nor \U$67 ( \382 , \380 , \381 );
xnor \U$68 ( \383 , \382 , \341 );
and \U$69 ( \384 , \379 , \383 );
and \U$70 ( \385 , \369 , \323 );
and \U$71 ( \386 , \348 , \321 );
nor \U$72 ( \387 , \385 , \386 );
xnor \U$73 ( \388 , \387 , \328 );
and \U$74 ( \389 , \383 , \388 );
and \U$75 ( \390 , \379 , \388 );
or \U$76 ( \391 , \384 , \389 , \390 );
xor \U$77 ( \392 , \363 , \367 );
xor \U$78 ( \393 , \392 , \370 );
or \U$79 ( \394 , \391 , \393 );
and \U$80 ( \395 , \373 , \394 );
xor \U$81 ( \396 , \342 , \346 );
xor \U$82 ( \397 , \396 , \349 );
and \U$83 ( \398 , \394 , \397 );
and \U$84 ( \399 , \373 , \397 );
or \U$85 ( \400 , \395 , \398 , \399 );
and \U$86 ( \401 , \356 , \400 );
xor \U$87 ( \402 , \356 , \400 );
xor \U$88 ( \403 , \373 , \394 );
xor \U$89 ( \404 , \403 , \397 );
xor \U$90 ( \405 , \338 , \374 );
xor \U$91 ( \406 , \374 , \375 );
not \U$92 ( \407 , \406 );
and \U$93 ( \408 , \405 , \407 );
and \U$94 ( \409 , \316 , \408 );
not \U$95 ( \410 , \409 );
xnor \U$96 ( \411 , \410 , \378 );
and \U$97 ( \412 , \348 , \360 );
and \U$98 ( \413 , \330 , \358 );
nor \U$99 ( \414 , \412 , \413 );
xnor \U$100 ( \415 , \414 , \341 );
and \U$101 ( \416 , \411 , \415 );
buf \U$102 ( \417 , RIc0c7770_70);
and \U$103 ( \418 , \417 , \323 );
and \U$104 ( \419 , \369 , \321 );
nor \U$105 ( \420 , \418 , \419 );
xnor \U$106 ( \421 , \420 , \328 );
and \U$107 ( \422 , \415 , \421 );
and \U$108 ( \423 , \411 , \421 );
or \U$109 ( \424 , \416 , \422 , \423 );
buf \U$110 ( \425 , RIc0c76f8_71);
and \U$111 ( \426 , \425 , \317 );
buf \U$112 ( \427 , \426 );
and \U$113 ( \428 , \424 , \427 );
and \U$114 ( \429 , \417 , \317 );
and \U$115 ( \430 , \427 , \429 );
and \U$116 ( \431 , \424 , \429 );
or \U$117 ( \432 , \428 , \430 , \431 );
buf \U$118 ( \433 , RIc0c9408_9);
buf \U$119 ( \434 , RIc0c9390_10);
and \U$120 ( \435 , \433 , \434 );
not \U$121 ( \436 , \435 );
and \U$122 ( \437 , \375 , \436 );
not \U$123 ( \438 , \437 );
and \U$124 ( \439 , \330 , \408 );
and \U$125 ( \440 , \316 , \406 );
nor \U$126 ( \441 , \439 , \440 );
xnor \U$127 ( \442 , \441 , \378 );
and \U$128 ( \443 , \438 , \442 );
and \U$129 ( \444 , \369 , \360 );
and \U$130 ( \445 , \348 , \358 );
nor \U$131 ( \446 , \444 , \445 );
xnor \U$132 ( \447 , \446 , \341 );
and \U$133 ( \448 , \442 , \447 );
and \U$134 ( \449 , \438 , \447 );
or \U$135 ( \450 , \443 , \448 , \449 );
xor \U$136 ( \451 , \411 , \415 );
xor \U$137 ( \452 , \451 , \421 );
and \U$138 ( \453 , \450 , \452 );
not \U$139 ( \454 , \426 );
and \U$140 ( \455 , \452 , \454 );
and \U$141 ( \456 , \450 , \454 );
or \U$142 ( \457 , \453 , \455 , \456 );
xor \U$143 ( \458 , \379 , \383 );
xor \U$144 ( \459 , \458 , \388 );
and \U$145 ( \460 , \457 , \459 );
xor \U$146 ( \461 , \424 , \427 );
xor \U$147 ( \462 , \461 , \429 );
and \U$148 ( \463 , \459 , \462 );
and \U$149 ( \464 , \457 , \462 );
or \U$150 ( \465 , \460 , \463 , \464 );
and \U$151 ( \466 , \432 , \465 );
xnor \U$152 ( \467 , \391 , \393 );
and \U$153 ( \468 , \465 , \467 );
and \U$154 ( \469 , \432 , \467 );
or \U$155 ( \470 , \466 , \468 , \469 );
and \U$156 ( \471 , \404 , \470 );
xor \U$157 ( \472 , \404 , \470 );
xor \U$158 ( \473 , \432 , \465 );
xor \U$159 ( \474 , \473 , \467 );
xor \U$160 ( \475 , \375 , \433 );
xor \U$161 ( \476 , \433 , \434 );
not \U$162 ( \477 , \476 );
and \U$163 ( \478 , \475 , \477 );
and \U$164 ( \479 , \316 , \478 );
not \U$165 ( \480 , \479 );
xnor \U$166 ( \481 , \480 , \437 );
and \U$167 ( \482 , \348 , \408 );
and \U$168 ( \483 , \330 , \406 );
nor \U$169 ( \484 , \482 , \483 );
xnor \U$170 ( \485 , \484 , \378 );
and \U$171 ( \486 , \481 , \485 );
and \U$172 ( \487 , \417 , \360 );
and \U$173 ( \488 , \369 , \358 );
nor \U$174 ( \489 , \487 , \488 );
xnor \U$175 ( \490 , \489 , \341 );
and \U$176 ( \491 , \485 , \490 );
and \U$177 ( \492 , \481 , \490 );
or \U$178 ( \493 , \486 , \491 , \492 );
buf \U$179 ( \494 , RIc0c7680_72);
and \U$180 ( \495 , \494 , \323 );
and \U$181 ( \496 , \425 , \321 );
nor \U$182 ( \497 , \495 , \496 );
xnor \U$183 ( \498 , \497 , \328 );
buf \U$184 ( \499 , RIc0c7608_73);
and \U$185 ( \500 , \499 , \317 );
or \U$186 ( \501 , \498 , \500 );
and \U$187 ( \502 , \493 , \501 );
and \U$188 ( \503 , \425 , \323 );
and \U$189 ( \504 , \417 , \321 );
nor \U$190 ( \505 , \503 , \504 );
xnor \U$191 ( \506 , \505 , \328 );
and \U$192 ( \507 , \501 , \506 );
and \U$193 ( \508 , \493 , \506 );
or \U$194 ( \509 , \502 , \507 , \508 );
and \U$195 ( \510 , \494 , \317 );
xor \U$196 ( \511 , \438 , \442 );
xor \U$197 ( \512 , \511 , \447 );
and \U$198 ( \513 , \510 , \512 );
and \U$199 ( \514 , \509 , \513 );
xor \U$200 ( \515 , \450 , \452 );
xor \U$201 ( \516 , \515 , \454 );
and \U$202 ( \517 , \513 , \516 );
and \U$203 ( \518 , \509 , \516 );
or \U$204 ( \519 , \514 , \517 , \518 );
xor \U$205 ( \520 , \457 , \459 );
xor \U$206 ( \521 , \520 , \462 );
and \U$207 ( \522 , \519 , \521 );
and \U$208 ( \523 , \474 , \522 );
xor \U$209 ( \524 , \474 , \522 );
xor \U$210 ( \525 , \519 , \521 );
buf \U$211 ( \526 , RIc0c9318_11);
buf \U$212 ( \527 , RIc0c92a0_12);
and \U$213 ( \528 , \526 , \527 );
not \U$214 ( \529 , \528 );
and \U$215 ( \530 , \434 , \529 );
not \U$216 ( \531 , \530 );
and \U$217 ( \532 , \330 , \478 );
and \U$218 ( \533 , \316 , \476 );
nor \U$219 ( \534 , \532 , \533 );
xnor \U$220 ( \535 , \534 , \437 );
and \U$221 ( \536 , \531 , \535 );
and \U$222 ( \537 , \369 , \408 );
and \U$223 ( \538 , \348 , \406 );
nor \U$224 ( \539 , \537 , \538 );
xnor \U$225 ( \540 , \539 , \378 );
and \U$226 ( \541 , \535 , \540 );
and \U$227 ( \542 , \531 , \540 );
or \U$228 ( \543 , \536 , \541 , \542 );
and \U$229 ( \544 , \425 , \360 );
and \U$230 ( \545 , \417 , \358 );
nor \U$231 ( \546 , \544 , \545 );
xnor \U$232 ( \547 , \546 , \341 );
and \U$233 ( \548 , \499 , \323 );
and \U$234 ( \549 , \494 , \321 );
nor \U$235 ( \550 , \548 , \549 );
xnor \U$236 ( \551 , \550 , \328 );
and \U$237 ( \552 , \547 , \551 );
buf \U$238 ( \553 , RIc0c7590_74);
and \U$239 ( \554 , \553 , \317 );
and \U$240 ( \555 , \551 , \554 );
and \U$241 ( \556 , \547 , \554 );
or \U$242 ( \557 , \552 , \555 , \556 );
and \U$243 ( \558 , \543 , \557 );
xnor \U$244 ( \559 , \498 , \500 );
and \U$245 ( \560 , \557 , \559 );
and \U$246 ( \561 , \543 , \559 );
or \U$247 ( \562 , \558 , \560 , \561 );
xor \U$248 ( \563 , \493 , \501 );
xor \U$249 ( \564 , \563 , \506 );
and \U$250 ( \565 , \562 , \564 );
xor \U$251 ( \566 , \510 , \512 );
and \U$252 ( \567 , \564 , \566 );
and \U$253 ( \568 , \562 , \566 );
or \U$254 ( \569 , \565 , \567 , \568 );
xor \U$255 ( \570 , \509 , \513 );
xor \U$256 ( \571 , \570 , \516 );
and \U$257 ( \572 , \569 , \571 );
and \U$258 ( \573 , \525 , \572 );
xor \U$259 ( \574 , \525 , \572 );
xor \U$260 ( \575 , \569 , \571 );
xor \U$261 ( \576 , \434 , \526 );
xor \U$262 ( \577 , \526 , \527 );
not \U$263 ( \578 , \577 );
and \U$264 ( \579 , \576 , \578 );
and \U$265 ( \580 , \316 , \579 );
not \U$266 ( \581 , \580 );
xnor \U$267 ( \582 , \581 , \530 );
and \U$268 ( \583 , \348 , \478 );
and \U$269 ( \584 , \330 , \476 );
nor \U$270 ( \585 , \583 , \584 );
xnor \U$271 ( \586 , \585 , \437 );
and \U$272 ( \587 , \582 , \586 );
and \U$273 ( \588 , \417 , \408 );
and \U$274 ( \589 , \369 , \406 );
nor \U$275 ( \590 , \588 , \589 );
xnor \U$276 ( \591 , \590 , \378 );
and \U$277 ( \592 , \586 , \591 );
and \U$278 ( \593 , \582 , \591 );
or \U$279 ( \594 , \587 , \592 , \593 );
and \U$280 ( \595 , \494 , \360 );
and \U$281 ( \596 , \425 , \358 );
nor \U$282 ( \597 , \595 , \596 );
xnor \U$283 ( \598 , \597 , \341 );
and \U$284 ( \599 , \553 , \323 );
and \U$285 ( \600 , \499 , \321 );
nor \U$286 ( \601 , \599 , \600 );
xnor \U$287 ( \602 , \601 , \328 );
and \U$288 ( \603 , \598 , \602 );
buf \U$289 ( \604 , RIc0c7518_75);
and \U$290 ( \605 , \604 , \317 );
and \U$291 ( \606 , \602 , \605 );
and \U$292 ( \607 , \598 , \605 );
or \U$293 ( \608 , \603 , \606 , \607 );
and \U$294 ( \609 , \594 , \608 );
xor \U$295 ( \610 , \547 , \551 );
xor \U$296 ( \611 , \610 , \554 );
and \U$297 ( \612 , \608 , \611 );
and \U$298 ( \613 , \594 , \611 );
or \U$299 ( \614 , \609 , \612 , \613 );
xor \U$300 ( \615 , \481 , \485 );
xor \U$301 ( \616 , \615 , \490 );
and \U$302 ( \617 , \614 , \616 );
xor \U$303 ( \618 , \543 , \557 );
xor \U$304 ( \619 , \618 , \559 );
and \U$305 ( \620 , \616 , \619 );
and \U$306 ( \621 , \614 , \619 );
or \U$307 ( \622 , \617 , \620 , \621 );
xor \U$308 ( \623 , \562 , \564 );
xor \U$309 ( \624 , \623 , \566 );
and \U$310 ( \625 , \622 , \624 );
and \U$311 ( \626 , \575 , \625 );
xor \U$312 ( \627 , \575 , \625 );
xor \U$313 ( \628 , \622 , \624 );
and \U$314 ( \629 , \425 , \408 );
and \U$315 ( \630 , \417 , \406 );
nor \U$316 ( \631 , \629 , \630 );
xnor \U$317 ( \632 , \631 , \378 );
and \U$318 ( \633 , \499 , \360 );
and \U$319 ( \634 , \494 , \358 );
nor \U$320 ( \635 , \633 , \634 );
xnor \U$321 ( \636 , \635 , \341 );
and \U$322 ( \637 , \632 , \636 );
and \U$323 ( \638 , \604 , \323 );
and \U$324 ( \639 , \553 , \321 );
nor \U$325 ( \640 , \638 , \639 );
xnor \U$326 ( \641 , \640 , \328 );
and \U$327 ( \642 , \636 , \641 );
and \U$328 ( \643 , \632 , \641 );
or \U$329 ( \644 , \637 , \642 , \643 );
buf \U$330 ( \645 , RIc0c9228_13);
buf \U$331 ( \646 , RIc0c91b0_14);
and \U$332 ( \647 , \645 , \646 );
not \U$333 ( \648 , \647 );
and \U$334 ( \649 , \527 , \648 );
not \U$335 ( \650 , \649 );
and \U$336 ( \651 , \330 , \579 );
and \U$337 ( \652 , \316 , \577 );
nor \U$338 ( \653 , \651 , \652 );
xnor \U$339 ( \654 , \653 , \530 );
and \U$340 ( \655 , \650 , \654 );
and \U$341 ( \656 , \369 , \478 );
and \U$342 ( \657 , \348 , \476 );
nor \U$343 ( \658 , \656 , \657 );
xnor \U$344 ( \659 , \658 , \437 );
and \U$345 ( \660 , \654 , \659 );
and \U$346 ( \661 , \650 , \659 );
or \U$347 ( \662 , \655 , \660 , \661 );
or \U$348 ( \663 , \644 , \662 );
xor \U$349 ( \664 , \531 , \535 );
xor \U$350 ( \665 , \664 , \540 );
and \U$351 ( \666 , \663 , \665 );
xor \U$352 ( \667 , \594 , \608 );
xor \U$353 ( \668 , \667 , \611 );
and \U$354 ( \669 , \665 , \668 );
and \U$355 ( \670 , \663 , \668 );
or \U$356 ( \671 , \666 , \669 , \670 );
and \U$357 ( \672 , \494 , \408 );
and \U$358 ( \673 , \425 , \406 );
nor \U$359 ( \674 , \672 , \673 );
xnor \U$360 ( \675 , \674 , \378 );
and \U$361 ( \676 , \553 , \360 );
and \U$362 ( \677 , \499 , \358 );
nor \U$363 ( \678 , \676 , \677 );
xnor \U$364 ( \679 , \678 , \341 );
and \U$365 ( \680 , \675 , \679 );
buf \U$366 ( \681 , RIc0c74a0_76);
and \U$367 ( \682 , \681 , \323 );
and \U$368 ( \683 , \604 , \321 );
nor \U$369 ( \684 , \682 , \683 );
xnor \U$370 ( \685 , \684 , \328 );
and \U$371 ( \686 , \679 , \685 );
and \U$372 ( \687 , \675 , \685 );
or \U$373 ( \688 , \680 , \686 , \687 );
xor \U$374 ( \689 , \527 , \645 );
xor \U$375 ( \690 , \645 , \646 );
not \U$376 ( \691 , \690 );
and \U$377 ( \692 , \689 , \691 );
and \U$378 ( \693 , \316 , \692 );
not \U$379 ( \694 , \693 );
xnor \U$380 ( \695 , \694 , \649 );
and \U$381 ( \696 , \348 , \579 );
and \U$382 ( \697 , \330 , \577 );
nor \U$383 ( \698 , \696 , \697 );
xnor \U$384 ( \699 , \698 , \530 );
and \U$385 ( \700 , \695 , \699 );
and \U$386 ( \701 , \417 , \478 );
and \U$387 ( \702 , \369 , \476 );
nor \U$388 ( \703 , \701 , \702 );
xnor \U$389 ( \704 , \703 , \437 );
and \U$390 ( \705 , \699 , \704 );
and \U$391 ( \706 , \695 , \704 );
or \U$392 ( \707 , \700 , \705 , \706 );
and \U$393 ( \708 , \688 , \707 );
buf \U$394 ( \709 , RIc0c7428_77);
and \U$395 ( \710 , \709 , \317 );
buf \U$396 ( \711 , \710 );
and \U$397 ( \712 , \707 , \711 );
and \U$398 ( \713 , \688 , \711 );
or \U$399 ( \714 , \708 , \712 , \713 );
and \U$400 ( \715 , \681 , \317 );
xor \U$401 ( \716 , \632 , \636 );
xor \U$402 ( \717 , \716 , \641 );
and \U$403 ( \718 , \715 , \717 );
xor \U$404 ( \719 , \650 , \654 );
xor \U$405 ( \720 , \719 , \659 );
and \U$406 ( \721 , \717 , \720 );
and \U$407 ( \722 , \715 , \720 );
or \U$408 ( \723 , \718 , \721 , \722 );
and \U$409 ( \724 , \714 , \723 );
xor \U$410 ( \725 , \598 , \602 );
xor \U$411 ( \726 , \725 , \605 );
and \U$412 ( \727 , \723 , \726 );
and \U$413 ( \728 , \714 , \726 );
or \U$414 ( \729 , \724 , \727 , \728 );
xor \U$415 ( \730 , \582 , \586 );
xor \U$416 ( \731 , \730 , \591 );
xnor \U$417 ( \732 , \644 , \662 );
and \U$418 ( \733 , \731 , \732 );
and \U$419 ( \734 , \729 , \733 );
xor \U$420 ( \735 , \663 , \665 );
xor \U$421 ( \736 , \735 , \668 );
and \U$422 ( \737 , \733 , \736 );
and \U$423 ( \738 , \729 , \736 );
or \U$424 ( \739 , \734 , \737 , \738 );
and \U$425 ( \740 , \671 , \739 );
xor \U$426 ( \741 , \614 , \616 );
xor \U$427 ( \742 , \741 , \619 );
and \U$428 ( \743 , \739 , \742 );
and \U$429 ( \744 , \671 , \742 );
or \U$430 ( \745 , \740 , \743 , \744 );
and \U$431 ( \746 , \628 , \745 );
xor \U$432 ( \747 , \628 , \745 );
xor \U$433 ( \748 , \671 , \739 );
xor \U$434 ( \749 , \748 , \742 );
buf \U$435 ( \750 , RIc0c9138_15);
buf \U$436 ( \751 , RIc0c90c0_16);
and \U$437 ( \752 , \750 , \751 );
not \U$438 ( \753 , \752 );
and \U$439 ( \754 , \646 , \753 );
not \U$440 ( \755 , \754 );
and \U$441 ( \756 , \330 , \692 );
and \U$442 ( \757 , \316 , \690 );
nor \U$443 ( \758 , \756 , \757 );
xnor \U$444 ( \759 , \758 , \649 );
and \U$445 ( \760 , \755 , \759 );
and \U$446 ( \761 , \369 , \579 );
and \U$447 ( \762 , \348 , \577 );
nor \U$448 ( \763 , \761 , \762 );
xnor \U$449 ( \764 , \763 , \530 );
and \U$450 ( \765 , \759 , \764 );
and \U$451 ( \766 , \755 , \764 );
or \U$452 ( \767 , \760 , \765 , \766 );
and \U$453 ( \768 , \425 , \478 );
and \U$454 ( \769 , \417 , \476 );
nor \U$455 ( \770 , \768 , \769 );
xnor \U$456 ( \771 , \770 , \437 );
and \U$457 ( \772 , \499 , \408 );
and \U$458 ( \773 , \494 , \406 );
nor \U$459 ( \774 , \772 , \773 );
xnor \U$460 ( \775 , \774 , \378 );
and \U$461 ( \776 , \771 , \775 );
and \U$462 ( \777 , \604 , \360 );
and \U$463 ( \778 , \553 , \358 );
nor \U$464 ( \779 , \777 , \778 );
xnor \U$465 ( \780 , \779 , \341 );
and \U$466 ( \781 , \775 , \780 );
and \U$467 ( \782 , \771 , \780 );
or \U$468 ( \783 , \776 , \781 , \782 );
and \U$469 ( \784 , \767 , \783 );
and \U$470 ( \785 , \709 , \323 );
and \U$471 ( \786 , \681 , \321 );
nor \U$472 ( \787 , \785 , \786 );
xnor \U$473 ( \788 , \787 , \328 );
buf \U$474 ( \789 , RIc0c73b0_78);
and \U$475 ( \790 , \789 , \317 );
and \U$476 ( \791 , \788 , \790 );
and \U$477 ( \792 , \783 , \791 );
and \U$478 ( \793 , \767 , \791 );
or \U$479 ( \794 , \784 , \792 , \793 );
xor \U$480 ( \795 , \675 , \679 );
xor \U$481 ( \796 , \795 , \685 );
xor \U$482 ( \797 , \695 , \699 );
xor \U$483 ( \798 , \797 , \704 );
and \U$484 ( \799 , \796 , \798 );
not \U$485 ( \800 , \710 );
and \U$486 ( \801 , \798 , \800 );
and \U$487 ( \802 , \796 , \800 );
or \U$488 ( \803 , \799 , \801 , \802 );
and \U$489 ( \804 , \794 , \803 );
xor \U$490 ( \805 , \715 , \717 );
xor \U$491 ( \806 , \805 , \720 );
and \U$492 ( \807 , \803 , \806 );
and \U$493 ( \808 , \794 , \806 );
or \U$494 ( \809 , \804 , \807 , \808 );
xor \U$495 ( \810 , \714 , \723 );
xor \U$496 ( \811 , \810 , \726 );
and \U$497 ( \812 , \809 , \811 );
xor \U$498 ( \813 , \731 , \732 );
and \U$499 ( \814 , \811 , \813 );
and \U$500 ( \815 , \809 , \813 );
or \U$501 ( \816 , \812 , \814 , \815 );
xor \U$502 ( \817 , \729 , \733 );
xor \U$503 ( \818 , \817 , \736 );
and \U$504 ( \819 , \816 , \818 );
and \U$505 ( \820 , \749 , \819 );
xor \U$506 ( \821 , \749 , \819 );
xor \U$507 ( \822 , \816 , \818 );
xor \U$508 ( \823 , \646 , \750 );
xor \U$509 ( \824 , \750 , \751 );
not \U$510 ( \825 , \824 );
and \U$511 ( \826 , \823 , \825 );
and \U$512 ( \827 , \316 , \826 );
not \U$513 ( \828 , \827 );
xnor \U$514 ( \829 , \828 , \754 );
and \U$515 ( \830 , \348 , \692 );
and \U$516 ( \831 , \330 , \690 );
nor \U$517 ( \832 , \830 , \831 );
xnor \U$518 ( \833 , \832 , \649 );
and \U$519 ( \834 , \829 , \833 );
and \U$520 ( \835 , \417 , \579 );
and \U$521 ( \836 , \369 , \577 );
nor \U$522 ( \837 , \835 , \836 );
xnor \U$523 ( \838 , \837 , \530 );
and \U$524 ( \839 , \833 , \838 );
and \U$525 ( \840 , \829 , \838 );
or \U$526 ( \841 , \834 , \839 , \840 );
and \U$527 ( \842 , \494 , \478 );
and \U$528 ( \843 , \425 , \476 );
nor \U$529 ( \844 , \842 , \843 );
xnor \U$530 ( \845 , \844 , \437 );
and \U$531 ( \846 , \553 , \408 );
and \U$532 ( \847 , \499 , \406 );
nor \U$533 ( \848 , \846 , \847 );
xnor \U$534 ( \849 , \848 , \378 );
and \U$535 ( \850 , \845 , \849 );
and \U$536 ( \851 , \681 , \360 );
and \U$537 ( \852 , \604 , \358 );
nor \U$538 ( \853 , \851 , \852 );
xnor \U$539 ( \854 , \853 , \341 );
and \U$540 ( \855 , \849 , \854 );
and \U$541 ( \856 , \845 , \854 );
or \U$542 ( \857 , \850 , \855 , \856 );
and \U$543 ( \858 , \841 , \857 );
and \U$544 ( \859 , \789 , \323 );
and \U$545 ( \860 , \709 , \321 );
nor \U$546 ( \861 , \859 , \860 );
xnor \U$547 ( \862 , \861 , \328 );
buf \U$548 ( \863 , RIc0c7338_79);
and \U$549 ( \864 , \863 , \317 );
or \U$550 ( \865 , \862 , \864 );
and \U$551 ( \866 , \857 , \865 );
and \U$552 ( \867 , \841 , \865 );
or \U$553 ( \868 , \858 , \866 , \867 );
xor \U$554 ( \869 , \755 , \759 );
xor \U$555 ( \870 , \869 , \764 );
xor \U$556 ( \871 , \771 , \775 );
xor \U$557 ( \872 , \871 , \780 );
and \U$558 ( \873 , \870 , \872 );
xor \U$559 ( \874 , \788 , \790 );
and \U$560 ( \875 , \872 , \874 );
and \U$561 ( \876 , \870 , \874 );
or \U$562 ( \877 , \873 , \875 , \876 );
and \U$563 ( \878 , \868 , \877 );
xor \U$564 ( \879 , \796 , \798 );
xor \U$565 ( \880 , \879 , \800 );
and \U$566 ( \881 , \877 , \880 );
and \U$567 ( \882 , \868 , \880 );
or \U$568 ( \883 , \878 , \881 , \882 );
xor \U$569 ( \884 , \688 , \707 );
xor \U$570 ( \885 , \884 , \711 );
and \U$571 ( \886 , \883 , \885 );
xor \U$572 ( \887 , \794 , \803 );
xor \U$573 ( \888 , \887 , \806 );
and \U$574 ( \889 , \885 , \888 );
and \U$575 ( \890 , \883 , \888 );
or \U$576 ( \891 , \886 , \889 , \890 );
xor \U$577 ( \892 , \809 , \811 );
xor \U$578 ( \893 , \892 , \813 );
and \U$579 ( \894 , \891 , \893 );
and \U$580 ( \895 , \822 , \894 );
xor \U$581 ( \896 , \822 , \894 );
xor \U$582 ( \897 , \891 , \893 );
buf \U$583 ( \898 , RIc0c9048_17);
buf \U$584 ( \899 , RIc0c8fd0_18);
and \U$585 ( \900 , \898 , \899 );
not \U$586 ( \901 , \900 );
and \U$587 ( \902 , \751 , \901 );
not \U$588 ( \903 , \902 );
and \U$589 ( \904 , \330 , \826 );
and \U$590 ( \905 , \316 , \824 );
nor \U$591 ( \906 , \904 , \905 );
xnor \U$592 ( \907 , \906 , \754 );
and \U$593 ( \908 , \903 , \907 );
and \U$594 ( \909 , \369 , \692 );
and \U$595 ( \910 , \348 , \690 );
nor \U$596 ( \911 , \909 , \910 );
xnor \U$597 ( \912 , \911 , \649 );
and \U$598 ( \913 , \907 , \912 );
and \U$599 ( \914 , \903 , \912 );
or \U$600 ( \915 , \908 , \913 , \914 );
and \U$601 ( \916 , \709 , \360 );
and \U$602 ( \917 , \681 , \358 );
nor \U$603 ( \918 , \916 , \917 );
xnor \U$604 ( \919 , \918 , \341 );
and \U$605 ( \920 , \863 , \323 );
and \U$606 ( \921 , \789 , \321 );
nor \U$607 ( \922 , \920 , \921 );
xnor \U$608 ( \923 , \922 , \328 );
and \U$609 ( \924 , \919 , \923 );
buf \U$610 ( \925 , RIc0c72c0_80);
and \U$611 ( \926 , \925 , \317 );
and \U$612 ( \927 , \923 , \926 );
and \U$613 ( \928 , \919 , \926 );
or \U$614 ( \929 , \924 , \927 , \928 );
and \U$615 ( \930 , \915 , \929 );
and \U$616 ( \931 , \425 , \579 );
and \U$617 ( \932 , \417 , \577 );
nor \U$618 ( \933 , \931 , \932 );
xnor \U$619 ( \934 , \933 , \530 );
and \U$620 ( \935 , \499 , \478 );
and \U$621 ( \936 , \494 , \476 );
nor \U$622 ( \937 , \935 , \936 );
xnor \U$623 ( \938 , \937 , \437 );
and \U$624 ( \939 , \934 , \938 );
and \U$625 ( \940 , \604 , \408 );
and \U$626 ( \941 , \553 , \406 );
nor \U$627 ( \942 , \940 , \941 );
xnor \U$628 ( \943 , \942 , \378 );
and \U$629 ( \944 , \938 , \943 );
and \U$630 ( \945 , \934 , \943 );
or \U$631 ( \946 , \939 , \944 , \945 );
and \U$632 ( \947 , \929 , \946 );
and \U$633 ( \948 , \915 , \946 );
or \U$634 ( \949 , \930 , \947 , \948 );
xor \U$635 ( \950 , \829 , \833 );
xor \U$636 ( \951 , \950 , \838 );
xor \U$637 ( \952 , \845 , \849 );
xor \U$638 ( \953 , \952 , \854 );
and \U$639 ( \954 , \951 , \953 );
xnor \U$640 ( \955 , \862 , \864 );
and \U$641 ( \956 , \953 , \955 );
and \U$642 ( \957 , \951 , \955 );
or \U$643 ( \958 , \954 , \956 , \957 );
and \U$644 ( \959 , \949 , \958 );
xor \U$645 ( \960 , \870 , \872 );
xor \U$646 ( \961 , \960 , \874 );
and \U$647 ( \962 , \958 , \961 );
and \U$648 ( \963 , \949 , \961 );
or \U$649 ( \964 , \959 , \962 , \963 );
xor \U$650 ( \965 , \767 , \783 );
xor \U$651 ( \966 , \965 , \791 );
and \U$652 ( \967 , \964 , \966 );
xor \U$653 ( \968 , \868 , \877 );
xor \U$654 ( \969 , \968 , \880 );
and \U$655 ( \970 , \966 , \969 );
and \U$656 ( \971 , \964 , \969 );
or \U$657 ( \972 , \967 , \970 , \971 );
xor \U$658 ( \973 , \883 , \885 );
xor \U$659 ( \974 , \973 , \888 );
and \U$660 ( \975 , \972 , \974 );
and \U$661 ( \976 , \897 , \975 );
xor \U$662 ( \977 , \897 , \975 );
xor \U$663 ( \978 , \972 , \974 );
and \U$664 ( \979 , \789 , \360 );
and \U$665 ( \980 , \709 , \358 );
nor \U$666 ( \981 , \979 , \980 );
xnor \U$667 ( \982 , \981 , \341 );
and \U$668 ( \983 , \925 , \323 );
and \U$669 ( \984 , \863 , \321 );
nor \U$670 ( \985 , \983 , \984 );
xnor \U$671 ( \986 , \985 , \328 );
and \U$672 ( \987 , \982 , \986 );
buf \U$673 ( \988 , RIc0c7248_81);
and \U$674 ( \989 , \988 , \317 );
and \U$675 ( \990 , \986 , \989 );
and \U$676 ( \991 , \982 , \989 );
or \U$677 ( \992 , \987 , \990 , \991 );
xor \U$678 ( \993 , \751 , \898 );
xor \U$679 ( \994 , \898 , \899 );
not \U$680 ( \995 , \994 );
and \U$681 ( \996 , \993 , \995 );
and \U$682 ( \997 , \316 , \996 );
not \U$683 ( \998 , \997 );
xnor \U$684 ( \999 , \998 , \902 );
and \U$685 ( \1000 , \348 , \826 );
and \U$686 ( \1001 , \330 , \824 );
nor \U$687 ( \1002 , \1000 , \1001 );
xnor \U$688 ( \1003 , \1002 , \754 );
and \U$689 ( \1004 , \999 , \1003 );
and \U$690 ( \1005 , \417 , \692 );
and \U$691 ( \1006 , \369 , \690 );
nor \U$692 ( \1007 , \1005 , \1006 );
xnor \U$693 ( \1008 , \1007 , \649 );
and \U$694 ( \1009 , \1003 , \1008 );
and \U$695 ( \1010 , \999 , \1008 );
or \U$696 ( \1011 , \1004 , \1009 , \1010 );
and \U$697 ( \1012 , \992 , \1011 );
and \U$698 ( \1013 , \494 , \579 );
and \U$699 ( \1014 , \425 , \577 );
nor \U$700 ( \1015 , \1013 , \1014 );
xnor \U$701 ( \1016 , \1015 , \530 );
and \U$702 ( \1017 , \553 , \478 );
and \U$703 ( \1018 , \499 , \476 );
nor \U$704 ( \1019 , \1017 , \1018 );
xnor \U$705 ( \1020 , \1019 , \437 );
and \U$706 ( \1021 , \1016 , \1020 );
and \U$707 ( \1022 , \681 , \408 );
and \U$708 ( \1023 , \604 , \406 );
nor \U$709 ( \1024 , \1022 , \1023 );
xnor \U$710 ( \1025 , \1024 , \378 );
and \U$711 ( \1026 , \1020 , \1025 );
and \U$712 ( \1027 , \1016 , \1025 );
or \U$713 ( \1028 , \1021 , \1026 , \1027 );
and \U$714 ( \1029 , \1011 , \1028 );
and \U$715 ( \1030 , \992 , \1028 );
or \U$716 ( \1031 , \1012 , \1029 , \1030 );
xor \U$717 ( \1032 , \903 , \907 );
xor \U$718 ( \1033 , \1032 , \912 );
xor \U$719 ( \1034 , \919 , \923 );
xor \U$720 ( \1035 , \1034 , \926 );
and \U$721 ( \1036 , \1033 , \1035 );
xor \U$722 ( \1037 , \934 , \938 );
xor \U$723 ( \1038 , \1037 , \943 );
and \U$724 ( \1039 , \1035 , \1038 );
and \U$725 ( \1040 , \1033 , \1038 );
or \U$726 ( \1041 , \1036 , \1039 , \1040 );
and \U$727 ( \1042 , \1031 , \1041 );
xor \U$728 ( \1043 , \951 , \953 );
xor \U$729 ( \1044 , \1043 , \955 );
and \U$730 ( \1045 , \1041 , \1044 );
and \U$731 ( \1046 , \1031 , \1044 );
or \U$732 ( \1047 , \1042 , \1045 , \1046 );
xor \U$733 ( \1048 , \841 , \857 );
xor \U$734 ( \1049 , \1048 , \865 );
and \U$735 ( \1050 , \1047 , \1049 );
xor \U$736 ( \1051 , \949 , \958 );
xor \U$737 ( \1052 , \1051 , \961 );
and \U$738 ( \1053 , \1049 , \1052 );
and \U$739 ( \1054 , \1047 , \1052 );
or \U$740 ( \1055 , \1050 , \1053 , \1054 );
xor \U$741 ( \1056 , \964 , \966 );
xor \U$742 ( \1057 , \1056 , \969 );
and \U$743 ( \1058 , \1055 , \1057 );
and \U$744 ( \1059 , \978 , \1058 );
xor \U$745 ( \1060 , \978 , \1058 );
xor \U$746 ( \1061 , \1055 , \1057 );
and \U$747 ( \1062 , \425 , \692 );
and \U$748 ( \1063 , \417 , \690 );
nor \U$749 ( \1064 , \1062 , \1063 );
xnor \U$750 ( \1065 , \1064 , \649 );
and \U$751 ( \1066 , \499 , \579 );
and \U$752 ( \1067 , \494 , \577 );
nor \U$753 ( \1068 , \1066 , \1067 );
xnor \U$754 ( \1069 , \1068 , \530 );
and \U$755 ( \1070 , \1065 , \1069 );
and \U$756 ( \1071 , \604 , \478 );
and \U$757 ( \1072 , \553 , \476 );
nor \U$758 ( \1073 , \1071 , \1072 );
xnor \U$759 ( \1074 , \1073 , \437 );
and \U$760 ( \1075 , \1069 , \1074 );
and \U$761 ( \1076 , \1065 , \1074 );
or \U$762 ( \1077 , \1070 , \1075 , \1076 );
buf \U$763 ( \1078 , RIc0c8f58_19);
buf \U$764 ( \1079 , RIc0c8ee0_20);
and \U$765 ( \1080 , \1078 , \1079 );
not \U$766 ( \1081 , \1080 );
and \U$767 ( \1082 , \899 , \1081 );
not \U$768 ( \1083 , \1082 );
and \U$769 ( \1084 , \330 , \996 );
and \U$770 ( \1085 , \316 , \994 );
nor \U$771 ( \1086 , \1084 , \1085 );
xnor \U$772 ( \1087 , \1086 , \902 );
and \U$773 ( \1088 , \1083 , \1087 );
and \U$774 ( \1089 , \369 , \826 );
and \U$775 ( \1090 , \348 , \824 );
nor \U$776 ( \1091 , \1089 , \1090 );
xnor \U$777 ( \1092 , \1091 , \754 );
and \U$778 ( \1093 , \1087 , \1092 );
and \U$779 ( \1094 , \1083 , \1092 );
or \U$780 ( \1095 , \1088 , \1093 , \1094 );
and \U$781 ( \1096 , \1077 , \1095 );
and \U$782 ( \1097 , \709 , \408 );
and \U$783 ( \1098 , \681 , \406 );
nor \U$784 ( \1099 , \1097 , \1098 );
xnor \U$785 ( \1100 , \1099 , \378 );
and \U$786 ( \1101 , \863 , \360 );
and \U$787 ( \1102 , \789 , \358 );
nor \U$788 ( \1103 , \1101 , \1102 );
xnor \U$789 ( \1104 , \1103 , \341 );
and \U$790 ( \1105 , \1100 , \1104 );
and \U$791 ( \1106 , \988 , \323 );
and \U$792 ( \1107 , \925 , \321 );
nor \U$793 ( \1108 , \1106 , \1107 );
xnor \U$794 ( \1109 , \1108 , \328 );
and \U$795 ( \1110 , \1104 , \1109 );
and \U$796 ( \1111 , \1100 , \1109 );
or \U$797 ( \1112 , \1105 , \1110 , \1111 );
and \U$798 ( \1113 , \1095 , \1112 );
and \U$799 ( \1114 , \1077 , \1112 );
or \U$800 ( \1115 , \1096 , \1113 , \1114 );
xor \U$801 ( \1116 , \982 , \986 );
xor \U$802 ( \1117 , \1116 , \989 );
xor \U$803 ( \1118 , \1016 , \1020 );
xor \U$804 ( \1119 , \1118 , \1025 );
or \U$805 ( \1120 , \1117 , \1119 );
and \U$806 ( \1121 , \1115 , \1120 );
xor \U$807 ( \1122 , \1033 , \1035 );
xor \U$808 ( \1123 , \1122 , \1038 );
and \U$809 ( \1124 , \1120 , \1123 );
and \U$810 ( \1125 , \1115 , \1123 );
or \U$811 ( \1126 , \1121 , \1124 , \1125 );
xor \U$812 ( \1127 , \915 , \929 );
xor \U$813 ( \1128 , \1127 , \946 );
and \U$814 ( \1129 , \1126 , \1128 );
xor \U$815 ( \1130 , \1031 , \1041 );
xor \U$816 ( \1131 , \1130 , \1044 );
and \U$817 ( \1132 , \1128 , \1131 );
and \U$818 ( \1133 , \1126 , \1131 );
or \U$819 ( \1134 , \1129 , \1132 , \1133 );
xor \U$820 ( \1135 , \1047 , \1049 );
xor \U$821 ( \1136 , \1135 , \1052 );
and \U$822 ( \1137 , \1134 , \1136 );
and \U$823 ( \1138 , \1061 , \1137 );
xor \U$824 ( \1139 , \1061 , \1137 );
xor \U$825 ( \1140 , \1134 , \1136 );
and \U$826 ( \1141 , \494 , \692 );
and \U$827 ( \1142 , \425 , \690 );
nor \U$828 ( \1143 , \1141 , \1142 );
xnor \U$829 ( \1144 , \1143 , \649 );
and \U$830 ( \1145 , \553 , \579 );
and \U$831 ( \1146 , \499 , \577 );
nor \U$832 ( \1147 , \1145 , \1146 );
xnor \U$833 ( \1148 , \1147 , \530 );
and \U$834 ( \1149 , \1144 , \1148 );
and \U$835 ( \1150 , \681 , \478 );
and \U$836 ( \1151 , \604 , \476 );
nor \U$837 ( \1152 , \1150 , \1151 );
xnor \U$838 ( \1153 , \1152 , \437 );
and \U$839 ( \1154 , \1148 , \1153 );
and \U$840 ( \1155 , \1144 , \1153 );
or \U$841 ( \1156 , \1149 , \1154 , \1155 );
xor \U$842 ( \1157 , \899 , \1078 );
xor \U$843 ( \1158 , \1078 , \1079 );
not \U$844 ( \1159 , \1158 );
and \U$845 ( \1160 , \1157 , \1159 );
and \U$846 ( \1161 , \316 , \1160 );
not \U$847 ( \1162 , \1161 );
xnor \U$848 ( \1163 , \1162 , \1082 );
and \U$849 ( \1164 , \348 , \996 );
and \U$850 ( \1165 , \330 , \994 );
nor \U$851 ( \1166 , \1164 , \1165 );
xnor \U$852 ( \1167 , \1166 , \902 );
and \U$853 ( \1168 , \1163 , \1167 );
and \U$854 ( \1169 , \417 , \826 );
and \U$855 ( \1170 , \369 , \824 );
nor \U$856 ( \1171 , \1169 , \1170 );
xnor \U$857 ( \1172 , \1171 , \754 );
and \U$858 ( \1173 , \1167 , \1172 );
and \U$859 ( \1174 , \1163 , \1172 );
or \U$860 ( \1175 , \1168 , \1173 , \1174 );
and \U$861 ( \1176 , \1156 , \1175 );
and \U$862 ( \1177 , \789 , \408 );
and \U$863 ( \1178 , \709 , \406 );
nor \U$864 ( \1179 , \1177 , \1178 );
xnor \U$865 ( \1180 , \1179 , \378 );
and \U$866 ( \1181 , \925 , \360 );
and \U$867 ( \1182 , \863 , \358 );
nor \U$868 ( \1183 , \1181 , \1182 );
xnor \U$869 ( \1184 , \1183 , \341 );
and \U$870 ( \1185 , \1180 , \1184 );
buf \U$871 ( \1186 , RIc0c71d0_82);
and \U$872 ( \1187 , \1186 , \323 );
and \U$873 ( \1188 , \988 , \321 );
nor \U$874 ( \1189 , \1187 , \1188 );
xnor \U$875 ( \1190 , \1189 , \328 );
and \U$876 ( \1191 , \1184 , \1190 );
and \U$877 ( \1192 , \1180 , \1190 );
or \U$878 ( \1193 , \1185 , \1191 , \1192 );
and \U$879 ( \1194 , \1175 , \1193 );
and \U$880 ( \1195 , \1156 , \1193 );
or \U$881 ( \1196 , \1176 , \1194 , \1195 );
and \U$882 ( \1197 , \1186 , \317 );
xor \U$883 ( \1198 , \1065 , \1069 );
xor \U$884 ( \1199 , \1198 , \1074 );
and \U$885 ( \1200 , \1197 , \1199 );
xor \U$886 ( \1201 , \1100 , \1104 );
xor \U$887 ( \1202 , \1201 , \1109 );
and \U$888 ( \1203 , \1199 , \1202 );
and \U$889 ( \1204 , \1197 , \1202 );
or \U$890 ( \1205 , \1200 , \1203 , \1204 );
and \U$891 ( \1206 , \1196 , \1205 );
xor \U$892 ( \1207 , \999 , \1003 );
xor \U$893 ( \1208 , \1207 , \1008 );
and \U$894 ( \1209 , \1205 , \1208 );
and \U$895 ( \1210 , \1196 , \1208 );
or \U$896 ( \1211 , \1206 , \1209 , \1210 );
xor \U$897 ( \1212 , \992 , \1011 );
xor \U$898 ( \1213 , \1212 , \1028 );
and \U$899 ( \1214 , \1211 , \1213 );
xor \U$900 ( \1215 , \1115 , \1120 );
xor \U$901 ( \1216 , \1215 , \1123 );
and \U$902 ( \1217 , \1213 , \1216 );
and \U$903 ( \1218 , \1211 , \1216 );
or \U$904 ( \1219 , \1214 , \1217 , \1218 );
buf \U$905 ( \1220 , RIc0c8e68_21);
buf \U$906 ( \1221 , RIc0c8df0_22);
and \U$907 ( \1222 , \1220 , \1221 );
not \U$908 ( \1223 , \1222 );
and \U$909 ( \1224 , \1079 , \1223 );
not \U$910 ( \1225 , \1224 );
and \U$911 ( \1226 , \330 , \1160 );
and \U$912 ( \1227 , \316 , \1158 );
nor \U$913 ( \1228 , \1226 , \1227 );
xnor \U$914 ( \1229 , \1228 , \1082 );
and \U$915 ( \1230 , \1225 , \1229 );
and \U$916 ( \1231 , \369 , \996 );
and \U$917 ( \1232 , \348 , \994 );
nor \U$918 ( \1233 , \1231 , \1232 );
xnor \U$919 ( \1234 , \1233 , \902 );
and \U$920 ( \1235 , \1229 , \1234 );
and \U$921 ( \1236 , \1225 , \1234 );
or \U$922 ( \1237 , \1230 , \1235 , \1236 );
and \U$923 ( \1238 , \425 , \826 );
and \U$924 ( \1239 , \417 , \824 );
nor \U$925 ( \1240 , \1238 , \1239 );
xnor \U$926 ( \1241 , \1240 , \754 );
and \U$927 ( \1242 , \499 , \692 );
and \U$928 ( \1243 , \494 , \690 );
nor \U$929 ( \1244 , \1242 , \1243 );
xnor \U$930 ( \1245 , \1244 , \649 );
and \U$931 ( \1246 , \1241 , \1245 );
and \U$932 ( \1247 , \604 , \579 );
and \U$933 ( \1248 , \553 , \577 );
nor \U$934 ( \1249 , \1247 , \1248 );
xnor \U$935 ( \1250 , \1249 , \530 );
and \U$936 ( \1251 , \1245 , \1250 );
and \U$937 ( \1252 , \1241 , \1250 );
or \U$938 ( \1253 , \1246 , \1251 , \1252 );
and \U$939 ( \1254 , \1237 , \1253 );
and \U$940 ( \1255 , \709 , \478 );
and \U$941 ( \1256 , \681 , \476 );
nor \U$942 ( \1257 , \1255 , \1256 );
xnor \U$943 ( \1258 , \1257 , \437 );
and \U$944 ( \1259 , \863 , \408 );
and \U$945 ( \1260 , \789 , \406 );
nor \U$946 ( \1261 , \1259 , \1260 );
xnor \U$947 ( \1262 , \1261 , \378 );
and \U$948 ( \1263 , \1258 , \1262 );
and \U$949 ( \1264 , \988 , \360 );
and \U$950 ( \1265 , \925 , \358 );
nor \U$951 ( \1266 , \1264 , \1265 );
xnor \U$952 ( \1267 , \1266 , \341 );
and \U$953 ( \1268 , \1262 , \1267 );
and \U$954 ( \1269 , \1258 , \1267 );
or \U$955 ( \1270 , \1263 , \1268 , \1269 );
and \U$956 ( \1271 , \1253 , \1270 );
and \U$957 ( \1272 , \1237 , \1270 );
or \U$958 ( \1273 , \1254 , \1271 , \1272 );
buf \U$959 ( \1274 , RIc0c7158_83);
and \U$960 ( \1275 , \1274 , \317 );
xor \U$961 ( \1276 , \1180 , \1184 );
xor \U$962 ( \1277 , \1276 , \1190 );
or \U$963 ( \1278 , \1275 , \1277 );
and \U$964 ( \1279 , \1273 , \1278 );
xor \U$965 ( \1280 , \1144 , \1148 );
xor \U$966 ( \1281 , \1280 , \1153 );
xor \U$967 ( \1282 , \1163 , \1167 );
xor \U$968 ( \1283 , \1282 , \1172 );
and \U$969 ( \1284 , \1281 , \1283 );
and \U$970 ( \1285 , \1278 , \1284 );
and \U$971 ( \1286 , \1273 , \1284 );
or \U$972 ( \1287 , \1279 , \1285 , \1286 );
xor \U$973 ( \1288 , \1083 , \1087 );
xor \U$974 ( \1289 , \1288 , \1092 );
xor \U$975 ( \1290 , \1156 , \1175 );
xor \U$976 ( \1291 , \1290 , \1193 );
and \U$977 ( \1292 , \1289 , \1291 );
xor \U$978 ( \1293 , \1197 , \1199 );
xor \U$979 ( \1294 , \1293 , \1202 );
and \U$980 ( \1295 , \1291 , \1294 );
and \U$981 ( \1296 , \1289 , \1294 );
or \U$982 ( \1297 , \1292 , \1295 , \1296 );
and \U$983 ( \1298 , \1287 , \1297 );
xnor \U$984 ( \1299 , \1117 , \1119 );
and \U$985 ( \1300 , \1297 , \1299 );
and \U$986 ( \1301 , \1287 , \1299 );
or \U$987 ( \1302 , \1298 , \1300 , \1301 );
xor \U$988 ( \1303 , \1077 , \1095 );
xor \U$989 ( \1304 , \1303 , \1112 );
xor \U$990 ( \1305 , \1196 , \1205 );
xor \U$991 ( \1306 , \1305 , \1208 );
and \U$992 ( \1307 , \1304 , \1306 );
and \U$993 ( \1308 , \1302 , \1307 );
xor \U$994 ( \1309 , \1211 , \1213 );
xor \U$995 ( \1310 , \1309 , \1216 );
and \U$996 ( \1311 , \1307 , \1310 );
and \U$997 ( \1312 , \1302 , \1310 );
or \U$998 ( \1313 , \1308 , \1311 , \1312 );
and \U$999 ( \1314 , \1219 , \1313 );
xor \U$1000 ( \1315 , \1126 , \1128 );
xor \U$1001 ( \1316 , \1315 , \1131 );
and \U$1002 ( \1317 , \1313 , \1316 );
and \U$1003 ( \1318 , \1219 , \1316 );
or \U$1004 ( \1319 , \1314 , \1317 , \1318 );
and \U$1005 ( \1320 , \1140 , \1319 );
xor \U$1006 ( \1321 , \1140 , \1319 );
xor \U$1007 ( \1322 , \1219 , \1313 );
xor \U$1008 ( \1323 , \1322 , \1316 );
and \U$1009 ( \1324 , \789 , \478 );
and \U$1010 ( \1325 , \709 , \476 );
nor \U$1011 ( \1326 , \1324 , \1325 );
xnor \U$1012 ( \1327 , \1326 , \437 );
and \U$1013 ( \1328 , \925 , \408 );
and \U$1014 ( \1329 , \863 , \406 );
nor \U$1015 ( \1330 , \1328 , \1329 );
xnor \U$1016 ( \1331 , \1330 , \378 );
and \U$1017 ( \1332 , \1327 , \1331 );
and \U$1018 ( \1333 , \1186 , \360 );
and \U$1019 ( \1334 , \988 , \358 );
nor \U$1020 ( \1335 , \1333 , \1334 );
xnor \U$1021 ( \1336 , \1335 , \341 );
and \U$1022 ( \1337 , \1331 , \1336 );
and \U$1023 ( \1338 , \1327 , \1336 );
or \U$1024 ( \1339 , \1332 , \1337 , \1338 );
and \U$1025 ( \1340 , \494 , \826 );
and \U$1026 ( \1341 , \425 , \824 );
nor \U$1027 ( \1342 , \1340 , \1341 );
xnor \U$1028 ( \1343 , \1342 , \754 );
and \U$1029 ( \1344 , \553 , \692 );
and \U$1030 ( \1345 , \499 , \690 );
nor \U$1031 ( \1346 , \1344 , \1345 );
xnor \U$1032 ( \1347 , \1346 , \649 );
and \U$1033 ( \1348 , \1343 , \1347 );
and \U$1034 ( \1349 , \681 , \579 );
and \U$1035 ( \1350 , \604 , \577 );
nor \U$1036 ( \1351 , \1349 , \1350 );
xnor \U$1037 ( \1352 , \1351 , \530 );
and \U$1038 ( \1353 , \1347 , \1352 );
and \U$1039 ( \1354 , \1343 , \1352 );
or \U$1040 ( \1355 , \1348 , \1353 , \1354 );
and \U$1041 ( \1356 , \1339 , \1355 );
xor \U$1042 ( \1357 , \1079 , \1220 );
xor \U$1043 ( \1358 , \1220 , \1221 );
not \U$1044 ( \1359 , \1358 );
and \U$1045 ( \1360 , \1357 , \1359 );
and \U$1046 ( \1361 , \316 , \1360 );
not \U$1047 ( \1362 , \1361 );
xnor \U$1048 ( \1363 , \1362 , \1224 );
and \U$1049 ( \1364 , \348 , \1160 );
and \U$1050 ( \1365 , \330 , \1158 );
nor \U$1051 ( \1366 , \1364 , \1365 );
xnor \U$1052 ( \1367 , \1366 , \1082 );
and \U$1053 ( \1368 , \1363 , \1367 );
and \U$1054 ( \1369 , \417 , \996 );
and \U$1055 ( \1370 , \369 , \994 );
nor \U$1056 ( \1371 , \1369 , \1370 );
xnor \U$1057 ( \1372 , \1371 , \902 );
and \U$1058 ( \1373 , \1367 , \1372 );
and \U$1059 ( \1374 , \1363 , \1372 );
or \U$1060 ( \1375 , \1368 , \1373 , \1374 );
and \U$1061 ( \1376 , \1355 , \1375 );
and \U$1062 ( \1377 , \1339 , \1375 );
or \U$1063 ( \1378 , \1356 , \1376 , \1377 );
buf \U$1064 ( \1379 , RIc0c70e0_84);
and \U$1065 ( \1380 , \1379 , \323 );
and \U$1066 ( \1381 , \1274 , \321 );
nor \U$1067 ( \1382 , \1380 , \1381 );
xnor \U$1068 ( \1383 , \1382 , \328 );
buf \U$1069 ( \1384 , RIc0c7068_85);
and \U$1070 ( \1385 , \1384 , \317 );
or \U$1071 ( \1386 , \1383 , \1385 );
and \U$1072 ( \1387 , \1274 , \323 );
and \U$1073 ( \1388 , \1186 , \321 );
nor \U$1074 ( \1389 , \1387 , \1388 );
xnor \U$1075 ( \1390 , \1389 , \328 );
and \U$1076 ( \1391 , \1386 , \1390 );
and \U$1077 ( \1392 , \1379 , \317 );
and \U$1078 ( \1393 , \1390 , \1392 );
and \U$1079 ( \1394 , \1386 , \1392 );
or \U$1080 ( \1395 , \1391 , \1393 , \1394 );
and \U$1081 ( \1396 , \1378 , \1395 );
xor \U$1082 ( \1397 , \1225 , \1229 );
xor \U$1083 ( \1398 , \1397 , \1234 );
xor \U$1084 ( \1399 , \1241 , \1245 );
xor \U$1085 ( \1400 , \1399 , \1250 );
and \U$1086 ( \1401 , \1398 , \1400 );
xor \U$1087 ( \1402 , \1258 , \1262 );
xor \U$1088 ( \1403 , \1402 , \1267 );
and \U$1089 ( \1404 , \1400 , \1403 );
and \U$1090 ( \1405 , \1398 , \1403 );
or \U$1091 ( \1406 , \1401 , \1404 , \1405 );
and \U$1092 ( \1407 , \1395 , \1406 );
and \U$1093 ( \1408 , \1378 , \1406 );
or \U$1094 ( \1409 , \1396 , \1407 , \1408 );
xor \U$1095 ( \1410 , \1237 , \1253 );
xor \U$1096 ( \1411 , \1410 , \1270 );
xnor \U$1097 ( \1412 , \1275 , \1277 );
and \U$1098 ( \1413 , \1411 , \1412 );
xor \U$1099 ( \1414 , \1281 , \1283 );
and \U$1100 ( \1415 , \1412 , \1414 );
and \U$1101 ( \1416 , \1411 , \1414 );
or \U$1102 ( \1417 , \1413 , \1415 , \1416 );
and \U$1103 ( \1418 , \1409 , \1417 );
xor \U$1104 ( \1419 , \1289 , \1291 );
xor \U$1105 ( \1420 , \1419 , \1294 );
and \U$1106 ( \1421 , \1417 , \1420 );
and \U$1107 ( \1422 , \1409 , \1420 );
or \U$1108 ( \1423 , \1418 , \1421 , \1422 );
xor \U$1109 ( \1424 , \1287 , \1297 );
xor \U$1110 ( \1425 , \1424 , \1299 );
and \U$1111 ( \1426 , \1423 , \1425 );
xor \U$1112 ( \1427 , \1304 , \1306 );
and \U$1113 ( \1428 , \1425 , \1427 );
and \U$1114 ( \1429 , \1423 , \1427 );
or \U$1115 ( \1430 , \1426 , \1428 , \1429 );
xor \U$1116 ( \1431 , \1302 , \1307 );
xor \U$1117 ( \1432 , \1431 , \1310 );
and \U$1118 ( \1433 , \1430 , \1432 );
and \U$1119 ( \1434 , \1323 , \1433 );
xor \U$1120 ( \1435 , \1323 , \1433 );
xor \U$1121 ( \1436 , \1430 , \1432 );
buf \U$1122 ( \1437 , RIc0c8d78_23);
buf \U$1123 ( \1438 , RIc0c8d00_24);
and \U$1124 ( \1439 , \1437 , \1438 );
not \U$1125 ( \1440 , \1439 );
and \U$1126 ( \1441 , \1221 , \1440 );
not \U$1127 ( \1442 , \1441 );
and \U$1128 ( \1443 , \330 , \1360 );
and \U$1129 ( \1444 , \316 , \1358 );
nor \U$1130 ( \1445 , \1443 , \1444 );
xnor \U$1131 ( \1446 , \1445 , \1224 );
and \U$1132 ( \1447 , \1442 , \1446 );
and \U$1133 ( \1448 , \369 , \1160 );
and \U$1134 ( \1449 , \348 , \1158 );
nor \U$1135 ( \1450 , \1448 , \1449 );
xnor \U$1136 ( \1451 , \1450 , \1082 );
and \U$1137 ( \1452 , \1446 , \1451 );
and \U$1138 ( \1453 , \1442 , \1451 );
or \U$1139 ( \1454 , \1447 , \1452 , \1453 );
and \U$1140 ( \1455 , \709 , \579 );
and \U$1141 ( \1456 , \681 , \577 );
nor \U$1142 ( \1457 , \1455 , \1456 );
xnor \U$1143 ( \1458 , \1457 , \530 );
and \U$1144 ( \1459 , \863 , \478 );
and \U$1145 ( \1460 , \789 , \476 );
nor \U$1146 ( \1461 , \1459 , \1460 );
xnor \U$1147 ( \1462 , \1461 , \437 );
and \U$1148 ( \1463 , \1458 , \1462 );
and \U$1149 ( \1464 , \988 , \408 );
and \U$1150 ( \1465 , \925 , \406 );
nor \U$1151 ( \1466 , \1464 , \1465 );
xnor \U$1152 ( \1467 , \1466 , \378 );
and \U$1153 ( \1468 , \1462 , \1467 );
and \U$1154 ( \1469 , \1458 , \1467 );
or \U$1155 ( \1470 , \1463 , \1468 , \1469 );
and \U$1156 ( \1471 , \1454 , \1470 );
and \U$1157 ( \1472 , \425 , \996 );
and \U$1158 ( \1473 , \417 , \994 );
nor \U$1159 ( \1474 , \1472 , \1473 );
xnor \U$1160 ( \1475 , \1474 , \902 );
and \U$1161 ( \1476 , \499 , \826 );
and \U$1162 ( \1477 , \494 , \824 );
nor \U$1163 ( \1478 , \1476 , \1477 );
xnor \U$1164 ( \1479 , \1478 , \754 );
and \U$1165 ( \1480 , \1475 , \1479 );
and \U$1166 ( \1481 , \604 , \692 );
and \U$1167 ( \1482 , \553 , \690 );
nor \U$1168 ( \1483 , \1481 , \1482 );
xnor \U$1169 ( \1484 , \1483 , \649 );
and \U$1170 ( \1485 , \1479 , \1484 );
and \U$1171 ( \1486 , \1475 , \1484 );
or \U$1172 ( \1487 , \1480 , \1485 , \1486 );
and \U$1173 ( \1488 , \1470 , \1487 );
and \U$1174 ( \1489 , \1454 , \1487 );
or \U$1175 ( \1490 , \1471 , \1488 , \1489 );
and \U$1176 ( \1491 , \1274 , \360 );
and \U$1177 ( \1492 , \1186 , \358 );
nor \U$1178 ( \1493 , \1491 , \1492 );
xnor \U$1179 ( \1494 , \1493 , \341 );
and \U$1180 ( \1495 , \1384 , \323 );
and \U$1181 ( \1496 , \1379 , \321 );
nor \U$1182 ( \1497 , \1495 , \1496 );
xnor \U$1183 ( \1498 , \1497 , \328 );
and \U$1184 ( \1499 , \1494 , \1498 );
buf \U$1185 ( \1500 , RIc0c6ff0_86);
and \U$1186 ( \1501 , \1500 , \317 );
and \U$1187 ( \1502 , \1498 , \1501 );
and \U$1188 ( \1503 , \1494 , \1501 );
or \U$1189 ( \1504 , \1499 , \1502 , \1503 );
xor \U$1190 ( \1505 , \1327 , \1331 );
xor \U$1191 ( \1506 , \1505 , \1336 );
and \U$1192 ( \1507 , \1504 , \1506 );
xnor \U$1193 ( \1508 , \1383 , \1385 );
and \U$1194 ( \1509 , \1506 , \1508 );
and \U$1195 ( \1510 , \1504 , \1508 );
or \U$1196 ( \1511 , \1507 , \1509 , \1510 );
and \U$1197 ( \1512 , \1490 , \1511 );
xor \U$1198 ( \1513 , \1343 , \1347 );
xor \U$1199 ( \1514 , \1513 , \1352 );
xor \U$1200 ( \1515 , \1363 , \1367 );
xor \U$1201 ( \1516 , \1515 , \1372 );
and \U$1202 ( \1517 , \1514 , \1516 );
and \U$1203 ( \1518 , \1511 , \1517 );
and \U$1204 ( \1519 , \1490 , \1517 );
or \U$1205 ( \1520 , \1512 , \1518 , \1519 );
xor \U$1206 ( \1521 , \1339 , \1355 );
xor \U$1207 ( \1522 , \1521 , \1375 );
xor \U$1208 ( \1523 , \1386 , \1390 );
xor \U$1209 ( \1524 , \1523 , \1392 );
and \U$1210 ( \1525 , \1522 , \1524 );
xor \U$1211 ( \1526 , \1398 , \1400 );
xor \U$1212 ( \1527 , \1526 , \1403 );
and \U$1213 ( \1528 , \1524 , \1527 );
and \U$1214 ( \1529 , \1522 , \1527 );
or \U$1215 ( \1530 , \1525 , \1528 , \1529 );
and \U$1216 ( \1531 , \1520 , \1530 );
xor \U$1217 ( \1532 , \1411 , \1412 );
xor \U$1218 ( \1533 , \1532 , \1414 );
and \U$1219 ( \1534 , \1530 , \1533 );
and \U$1220 ( \1535 , \1520 , \1533 );
or \U$1221 ( \1536 , \1531 , \1534 , \1535 );
xor \U$1222 ( \1537 , \1273 , \1278 );
xor \U$1223 ( \1538 , \1537 , \1284 );
and \U$1224 ( \1539 , \1536 , \1538 );
xor \U$1225 ( \1540 , \1409 , \1417 );
xor \U$1226 ( \1541 , \1540 , \1420 );
and \U$1227 ( \1542 , \1538 , \1541 );
and \U$1228 ( \1543 , \1536 , \1541 );
or \U$1229 ( \1544 , \1539 , \1542 , \1543 );
xor \U$1230 ( \1545 , \1423 , \1425 );
xor \U$1231 ( \1546 , \1545 , \1427 );
and \U$1232 ( \1547 , \1544 , \1546 );
and \U$1233 ( \1548 , \1436 , \1547 );
xor \U$1234 ( \1549 , \1436 , \1547 );
xor \U$1235 ( \1550 , \1544 , \1546 );
xor \U$1236 ( \1551 , \1221 , \1437 );
xor \U$1237 ( \1552 , \1437 , \1438 );
not \U$1238 ( \1553 , \1552 );
and \U$1239 ( \1554 , \1551 , \1553 );
and \U$1240 ( \1555 , \316 , \1554 );
not \U$1241 ( \1556 , \1555 );
xnor \U$1242 ( \1557 , \1556 , \1441 );
and \U$1243 ( \1558 , \348 , \1360 );
and \U$1244 ( \1559 , \330 , \1358 );
nor \U$1245 ( \1560 , \1558 , \1559 );
xnor \U$1246 ( \1561 , \1560 , \1224 );
and \U$1247 ( \1562 , \1557 , \1561 );
and \U$1248 ( \1563 , \417 , \1160 );
and \U$1249 ( \1564 , \369 , \1158 );
nor \U$1250 ( \1565 , \1563 , \1564 );
xnor \U$1251 ( \1566 , \1565 , \1082 );
and \U$1252 ( \1567 , \1561 , \1566 );
and \U$1253 ( \1568 , \1557 , \1566 );
or \U$1254 ( \1569 , \1562 , \1567 , \1568 );
and \U$1255 ( \1570 , \789 , \579 );
and \U$1256 ( \1571 , \709 , \577 );
nor \U$1257 ( \1572 , \1570 , \1571 );
xnor \U$1258 ( \1573 , \1572 , \530 );
and \U$1259 ( \1574 , \925 , \478 );
and \U$1260 ( \1575 , \863 , \476 );
nor \U$1261 ( \1576 , \1574 , \1575 );
xnor \U$1262 ( \1577 , \1576 , \437 );
and \U$1263 ( \1578 , \1573 , \1577 );
and \U$1264 ( \1579 , \1186 , \408 );
and \U$1265 ( \1580 , \988 , \406 );
nor \U$1266 ( \1581 , \1579 , \1580 );
xnor \U$1267 ( \1582 , \1581 , \378 );
and \U$1268 ( \1583 , \1577 , \1582 );
and \U$1269 ( \1584 , \1573 , \1582 );
or \U$1270 ( \1585 , \1578 , \1583 , \1584 );
and \U$1271 ( \1586 , \1569 , \1585 );
and \U$1272 ( \1587 , \494 , \996 );
and \U$1273 ( \1588 , \425 , \994 );
nor \U$1274 ( \1589 , \1587 , \1588 );
xnor \U$1275 ( \1590 , \1589 , \902 );
and \U$1276 ( \1591 , \553 , \826 );
and \U$1277 ( \1592 , \499 , \824 );
nor \U$1278 ( \1593 , \1591 , \1592 );
xnor \U$1279 ( \1594 , \1593 , \754 );
and \U$1280 ( \1595 , \1590 , \1594 );
and \U$1281 ( \1596 , \681 , \692 );
and \U$1282 ( \1597 , \604 , \690 );
nor \U$1283 ( \1598 , \1596 , \1597 );
xnor \U$1284 ( \1599 , \1598 , \649 );
and \U$1285 ( \1600 , \1594 , \1599 );
and \U$1286 ( \1601 , \1590 , \1599 );
or \U$1287 ( \1602 , \1595 , \1600 , \1601 );
and \U$1288 ( \1603 , \1585 , \1602 );
and \U$1289 ( \1604 , \1569 , \1602 );
or \U$1290 ( \1605 , \1586 , \1603 , \1604 );
and \U$1291 ( \1606 , \1379 , \360 );
and \U$1292 ( \1607 , \1274 , \358 );
nor \U$1293 ( \1608 , \1606 , \1607 );
xnor \U$1294 ( \1609 , \1608 , \341 );
and \U$1295 ( \1610 , \1500 , \323 );
and \U$1296 ( \1611 , \1384 , \321 );
nor \U$1297 ( \1612 , \1610 , \1611 );
xnor \U$1298 ( \1613 , \1612 , \328 );
and \U$1299 ( \1614 , \1609 , \1613 );
buf \U$1300 ( \1615 , RIc0c6f78_87);
and \U$1301 ( \1616 , \1615 , \317 );
and \U$1302 ( \1617 , \1613 , \1616 );
and \U$1303 ( \1618 , \1609 , \1616 );
or \U$1304 ( \1619 , \1614 , \1617 , \1618 );
xor \U$1305 ( \1620 , \1494 , \1498 );
xor \U$1306 ( \1621 , \1620 , \1501 );
and \U$1307 ( \1622 , \1619 , \1621 );
xor \U$1308 ( \1623 , \1458 , \1462 );
xor \U$1309 ( \1624 , \1623 , \1467 );
and \U$1310 ( \1625 , \1621 , \1624 );
and \U$1311 ( \1626 , \1619 , \1624 );
or \U$1312 ( \1627 , \1622 , \1625 , \1626 );
and \U$1313 ( \1628 , \1605 , \1627 );
xor \U$1314 ( \1629 , \1442 , \1446 );
xor \U$1315 ( \1630 , \1629 , \1451 );
xor \U$1316 ( \1631 , \1475 , \1479 );
xor \U$1317 ( \1632 , \1631 , \1484 );
and \U$1318 ( \1633 , \1630 , \1632 );
and \U$1319 ( \1634 , \1627 , \1633 );
and \U$1320 ( \1635 , \1605 , \1633 );
or \U$1321 ( \1636 , \1628 , \1634 , \1635 );
xor \U$1322 ( \1637 , \1454 , \1470 );
xor \U$1323 ( \1638 , \1637 , \1487 );
xor \U$1324 ( \1639 , \1504 , \1506 );
xor \U$1325 ( \1640 , \1639 , \1508 );
and \U$1326 ( \1641 , \1638 , \1640 );
xor \U$1327 ( \1642 , \1514 , \1516 );
and \U$1328 ( \1643 , \1640 , \1642 );
and \U$1329 ( \1644 , \1638 , \1642 );
or \U$1330 ( \1645 , \1641 , \1643 , \1644 );
and \U$1331 ( \1646 , \1636 , \1645 );
xor \U$1332 ( \1647 , \1522 , \1524 );
xor \U$1333 ( \1648 , \1647 , \1527 );
and \U$1334 ( \1649 , \1645 , \1648 );
and \U$1335 ( \1650 , \1636 , \1648 );
or \U$1336 ( \1651 , \1646 , \1649 , \1650 );
xor \U$1337 ( \1652 , \1378 , \1395 );
xor \U$1338 ( \1653 , \1652 , \1406 );
and \U$1339 ( \1654 , \1651 , \1653 );
xor \U$1340 ( \1655 , \1520 , \1530 );
xor \U$1341 ( \1656 , \1655 , \1533 );
and \U$1342 ( \1657 , \1653 , \1656 );
and \U$1343 ( \1658 , \1651 , \1656 );
or \U$1344 ( \1659 , \1654 , \1657 , \1658 );
xor \U$1345 ( \1660 , \1536 , \1538 );
xor \U$1346 ( \1661 , \1660 , \1541 );
and \U$1347 ( \1662 , \1659 , \1661 );
and \U$1348 ( \1663 , \1550 , \1662 );
xor \U$1349 ( \1664 , \1550 , \1662 );
xor \U$1350 ( \1665 , \1659 , \1661 );
buf \U$1351 ( \1666 , RIc0c8c88_25);
buf \U$1352 ( \1667 , RIc0c8c10_26);
and \U$1353 ( \1668 , \1666 , \1667 );
not \U$1354 ( \1669 , \1668 );
and \U$1355 ( \1670 , \1438 , \1669 );
not \U$1356 ( \1671 , \1670 );
and \U$1357 ( \1672 , \330 , \1554 );
and \U$1358 ( \1673 , \316 , \1552 );
nor \U$1359 ( \1674 , \1672 , \1673 );
xnor \U$1360 ( \1675 , \1674 , \1441 );
and \U$1361 ( \1676 , \1671 , \1675 );
and \U$1362 ( \1677 , \369 , \1360 );
and \U$1363 ( \1678 , \348 , \1358 );
nor \U$1364 ( \1679 , \1677 , \1678 );
xnor \U$1365 ( \1680 , \1679 , \1224 );
and \U$1366 ( \1681 , \1675 , \1680 );
and \U$1367 ( \1682 , \1671 , \1680 );
or \U$1368 ( \1683 , \1676 , \1681 , \1682 );
and \U$1369 ( \1684 , \425 , \1160 );
and \U$1370 ( \1685 , \417 , \1158 );
nor \U$1371 ( \1686 , \1684 , \1685 );
xnor \U$1372 ( \1687 , \1686 , \1082 );
and \U$1373 ( \1688 , \499 , \996 );
and \U$1374 ( \1689 , \494 , \994 );
nor \U$1375 ( \1690 , \1688 , \1689 );
xnor \U$1376 ( \1691 , \1690 , \902 );
and \U$1377 ( \1692 , \1687 , \1691 );
and \U$1378 ( \1693 , \604 , \826 );
and \U$1379 ( \1694 , \553 , \824 );
nor \U$1380 ( \1695 , \1693 , \1694 );
xnor \U$1381 ( \1696 , \1695 , \754 );
and \U$1382 ( \1697 , \1691 , \1696 );
and \U$1383 ( \1698 , \1687 , \1696 );
or \U$1384 ( \1699 , \1692 , \1697 , \1698 );
and \U$1385 ( \1700 , \1683 , \1699 );
and \U$1386 ( \1701 , \709 , \692 );
and \U$1387 ( \1702 , \681 , \690 );
nor \U$1388 ( \1703 , \1701 , \1702 );
xnor \U$1389 ( \1704 , \1703 , \649 );
and \U$1390 ( \1705 , \863 , \579 );
and \U$1391 ( \1706 , \789 , \577 );
nor \U$1392 ( \1707 , \1705 , \1706 );
xnor \U$1393 ( \1708 , \1707 , \530 );
and \U$1394 ( \1709 , \1704 , \1708 );
and \U$1395 ( \1710 , \988 , \478 );
and \U$1396 ( \1711 , \925 , \476 );
nor \U$1397 ( \1712 , \1710 , \1711 );
xnor \U$1398 ( \1713 , \1712 , \437 );
and \U$1399 ( \1714 , \1708 , \1713 );
and \U$1400 ( \1715 , \1704 , \1713 );
or \U$1401 ( \1716 , \1709 , \1714 , \1715 );
and \U$1402 ( \1717 , \1699 , \1716 );
and \U$1403 ( \1718 , \1683 , \1716 );
or \U$1404 ( \1719 , \1700 , \1717 , \1718 );
xor \U$1405 ( \1720 , \1557 , \1561 );
xor \U$1406 ( \1721 , \1720 , \1566 );
xor \U$1407 ( \1722 , \1573 , \1577 );
xor \U$1408 ( \1723 , \1722 , \1582 );
and \U$1409 ( \1724 , \1721 , \1723 );
xor \U$1410 ( \1725 , \1590 , \1594 );
xor \U$1411 ( \1726 , \1725 , \1599 );
and \U$1412 ( \1727 , \1723 , \1726 );
and \U$1413 ( \1728 , \1721 , \1726 );
or \U$1414 ( \1729 , \1724 , \1727 , \1728 );
and \U$1415 ( \1730 , \1719 , \1729 );
and \U$1416 ( \1731 , \1274 , \408 );
and \U$1417 ( \1732 , \1186 , \406 );
nor \U$1418 ( \1733 , \1731 , \1732 );
xnor \U$1419 ( \1734 , \1733 , \378 );
and \U$1420 ( \1735 , \1384 , \360 );
and \U$1421 ( \1736 , \1379 , \358 );
nor \U$1422 ( \1737 , \1735 , \1736 );
xnor \U$1423 ( \1738 , \1737 , \341 );
and \U$1424 ( \1739 , \1734 , \1738 );
and \U$1425 ( \1740 , \1615 , \323 );
and \U$1426 ( \1741 , \1500 , \321 );
nor \U$1427 ( \1742 , \1740 , \1741 );
xnor \U$1428 ( \1743 , \1742 , \328 );
and \U$1429 ( \1744 , \1738 , \1743 );
and \U$1430 ( \1745 , \1734 , \1743 );
or \U$1431 ( \1746 , \1739 , \1744 , \1745 );
xor \U$1432 ( \1747 , \1609 , \1613 );
xor \U$1433 ( \1748 , \1747 , \1616 );
or \U$1434 ( \1749 , \1746 , \1748 );
and \U$1435 ( \1750 , \1729 , \1749 );
and \U$1436 ( \1751 , \1719 , \1749 );
or \U$1437 ( \1752 , \1730 , \1750 , \1751 );
xor \U$1438 ( \1753 , \1569 , \1585 );
xor \U$1439 ( \1754 , \1753 , \1602 );
xor \U$1440 ( \1755 , \1619 , \1621 );
xor \U$1441 ( \1756 , \1755 , \1624 );
and \U$1442 ( \1757 , \1754 , \1756 );
xor \U$1443 ( \1758 , \1630 , \1632 );
and \U$1444 ( \1759 , \1756 , \1758 );
and \U$1445 ( \1760 , \1754 , \1758 );
or \U$1446 ( \1761 , \1757 , \1759 , \1760 );
and \U$1447 ( \1762 , \1752 , \1761 );
xor \U$1448 ( \1763 , \1638 , \1640 );
xor \U$1449 ( \1764 , \1763 , \1642 );
and \U$1450 ( \1765 , \1761 , \1764 );
and \U$1451 ( \1766 , \1752 , \1764 );
or \U$1452 ( \1767 , \1762 , \1765 , \1766 );
xor \U$1453 ( \1768 , \1490 , \1511 );
xor \U$1454 ( \1769 , \1768 , \1517 );
and \U$1455 ( \1770 , \1767 , \1769 );
xor \U$1456 ( \1771 , \1636 , \1645 );
xor \U$1457 ( \1772 , \1771 , \1648 );
and \U$1458 ( \1773 , \1769 , \1772 );
and \U$1459 ( \1774 , \1767 , \1772 );
or \U$1460 ( \1775 , \1770 , \1773 , \1774 );
xor \U$1461 ( \1776 , \1651 , \1653 );
xor \U$1462 ( \1777 , \1776 , \1656 );
and \U$1463 ( \1778 , \1775 , \1777 );
and \U$1464 ( \1779 , \1665 , \1778 );
xor \U$1465 ( \1780 , \1665 , \1778 );
xor \U$1466 ( \1781 , \1775 , \1777 );
and \U$1467 ( \1782 , \1379 , \408 );
and \U$1468 ( \1783 , \1274 , \406 );
nor \U$1469 ( \1784 , \1782 , \1783 );
xnor \U$1470 ( \1785 , \1784 , \378 );
and \U$1471 ( \1786 , \1500 , \360 );
and \U$1472 ( \1787 , \1384 , \358 );
nor \U$1473 ( \1788 , \1786 , \1787 );
xnor \U$1474 ( \1789 , \1788 , \341 );
and \U$1475 ( \1790 , \1785 , \1789 );
buf \U$1476 ( \1791 , RIc0c6f00_88);
and \U$1477 ( \1792 , \1791 , \323 );
and \U$1478 ( \1793 , \1615 , \321 );
nor \U$1479 ( \1794 , \1792 , \1793 );
xnor \U$1480 ( \1795 , \1794 , \328 );
and \U$1481 ( \1796 , \1789 , \1795 );
and \U$1482 ( \1797 , \1785 , \1795 );
or \U$1483 ( \1798 , \1790 , \1796 , \1797 );
buf \U$1484 ( \1799 , RIc0c6e88_89);
and \U$1485 ( \1800 , \1799 , \317 );
buf \U$1486 ( \1801 , \1800 );
and \U$1487 ( \1802 , \1798 , \1801 );
and \U$1488 ( \1803 , \1791 , \317 );
and \U$1489 ( \1804 , \1801 , \1803 );
and \U$1490 ( \1805 , \1798 , \1803 );
or \U$1491 ( \1806 , \1802 , \1804 , \1805 );
and \U$1492 ( \1807 , \494 , \1160 );
and \U$1493 ( \1808 , \425 , \1158 );
nor \U$1494 ( \1809 , \1807 , \1808 );
xnor \U$1495 ( \1810 , \1809 , \1082 );
and \U$1496 ( \1811 , \553 , \996 );
and \U$1497 ( \1812 , \499 , \994 );
nor \U$1498 ( \1813 , \1811 , \1812 );
xnor \U$1499 ( \1814 , \1813 , \902 );
and \U$1500 ( \1815 , \1810 , \1814 );
and \U$1501 ( \1816 , \681 , \826 );
and \U$1502 ( \1817 , \604 , \824 );
nor \U$1503 ( \1818 , \1816 , \1817 );
xnor \U$1504 ( \1819 , \1818 , \754 );
and \U$1505 ( \1820 , \1814 , \1819 );
and \U$1506 ( \1821 , \1810 , \1819 );
or \U$1507 ( \1822 , \1815 , \1820 , \1821 );
xor \U$1508 ( \1823 , \1438 , \1666 );
xor \U$1509 ( \1824 , \1666 , \1667 );
not \U$1510 ( \1825 , \1824 );
and \U$1511 ( \1826 , \1823 , \1825 );
and \U$1512 ( \1827 , \316 , \1826 );
not \U$1513 ( \1828 , \1827 );
xnor \U$1514 ( \1829 , \1828 , \1670 );
and \U$1515 ( \1830 , \348 , \1554 );
and \U$1516 ( \1831 , \330 , \1552 );
nor \U$1517 ( \1832 , \1830 , \1831 );
xnor \U$1518 ( \1833 , \1832 , \1441 );
and \U$1519 ( \1834 , \1829 , \1833 );
and \U$1520 ( \1835 , \417 , \1360 );
and \U$1521 ( \1836 , \369 , \1358 );
nor \U$1522 ( \1837 , \1835 , \1836 );
xnor \U$1523 ( \1838 , \1837 , \1224 );
and \U$1524 ( \1839 , \1833 , \1838 );
and \U$1525 ( \1840 , \1829 , \1838 );
or \U$1526 ( \1841 , \1834 , \1839 , \1840 );
and \U$1527 ( \1842 , \1822 , \1841 );
and \U$1528 ( \1843 , \789 , \692 );
and \U$1529 ( \1844 , \709 , \690 );
nor \U$1530 ( \1845 , \1843 , \1844 );
xnor \U$1531 ( \1846 , \1845 , \649 );
and \U$1532 ( \1847 , \925 , \579 );
and \U$1533 ( \1848 , \863 , \577 );
nor \U$1534 ( \1849 , \1847 , \1848 );
xnor \U$1535 ( \1850 , \1849 , \530 );
and \U$1536 ( \1851 , \1846 , \1850 );
and \U$1537 ( \1852 , \1186 , \478 );
and \U$1538 ( \1853 , \988 , \476 );
nor \U$1539 ( \1854 , \1852 , \1853 );
xnor \U$1540 ( \1855 , \1854 , \437 );
and \U$1541 ( \1856 , \1850 , \1855 );
and \U$1542 ( \1857 , \1846 , \1855 );
or \U$1543 ( \1858 , \1851 , \1856 , \1857 );
and \U$1544 ( \1859 , \1841 , \1858 );
and \U$1545 ( \1860 , \1822 , \1858 );
or \U$1546 ( \1861 , \1842 , \1859 , \1860 );
and \U$1547 ( \1862 , \1806 , \1861 );
xor \U$1548 ( \1863 , \1687 , \1691 );
xor \U$1549 ( \1864 , \1863 , \1696 );
xor \U$1550 ( \1865 , \1734 , \1738 );
xor \U$1551 ( \1866 , \1865 , \1743 );
and \U$1552 ( \1867 , \1864 , \1866 );
xor \U$1553 ( \1868 , \1704 , \1708 );
xor \U$1554 ( \1869 , \1868 , \1713 );
and \U$1555 ( \1870 , \1866 , \1869 );
and \U$1556 ( \1871 , \1864 , \1869 );
or \U$1557 ( \1872 , \1867 , \1870 , \1871 );
and \U$1558 ( \1873 , \1861 , \1872 );
and \U$1559 ( \1874 , \1806 , \1872 );
or \U$1560 ( \1875 , \1862 , \1873 , \1874 );
xor \U$1561 ( \1876 , \1683 , \1699 );
xor \U$1562 ( \1877 , \1876 , \1716 );
xor \U$1563 ( \1878 , \1721 , \1723 );
xor \U$1564 ( \1879 , \1878 , \1726 );
and \U$1565 ( \1880 , \1877 , \1879 );
xnor \U$1566 ( \1881 , \1746 , \1748 );
and \U$1567 ( \1882 , \1879 , \1881 );
and \U$1568 ( \1883 , \1877 , \1881 );
or \U$1569 ( \1884 , \1880 , \1882 , \1883 );
and \U$1570 ( \1885 , \1875 , \1884 );
xor \U$1571 ( \1886 , \1754 , \1756 );
xor \U$1572 ( \1887 , \1886 , \1758 );
and \U$1573 ( \1888 , \1884 , \1887 );
and \U$1574 ( \1889 , \1875 , \1887 );
or \U$1575 ( \1890 , \1885 , \1888 , \1889 );
xor \U$1576 ( \1891 , \1605 , \1627 );
xor \U$1577 ( \1892 , \1891 , \1633 );
and \U$1578 ( \1893 , \1890 , \1892 );
xor \U$1579 ( \1894 , \1752 , \1761 );
xor \U$1580 ( \1895 , \1894 , \1764 );
and \U$1581 ( \1896 , \1892 , \1895 );
and \U$1582 ( \1897 , \1890 , \1895 );
or \U$1583 ( \1898 , \1893 , \1896 , \1897 );
xor \U$1584 ( \1899 , \1767 , \1769 );
xor \U$1585 ( \1900 , \1899 , \1772 );
and \U$1586 ( \1901 , \1898 , \1900 );
and \U$1587 ( \1902 , \1781 , \1901 );
xor \U$1588 ( \1903 , \1781 , \1901 );
xor \U$1589 ( \1904 , \1898 , \1900 );
and \U$1590 ( \1905 , \709 , \826 );
and \U$1591 ( \1906 , \681 , \824 );
nor \U$1592 ( \1907 , \1905 , \1906 );
xnor \U$1593 ( \1908 , \1907 , \754 );
and \U$1594 ( \1909 , \863 , \692 );
and \U$1595 ( \1910 , \789 , \690 );
nor \U$1596 ( \1911 , \1909 , \1910 );
xnor \U$1597 ( \1912 , \1911 , \649 );
and \U$1598 ( \1913 , \1908 , \1912 );
and \U$1599 ( \1914 , \988 , \579 );
and \U$1600 ( \1915 , \925 , \577 );
nor \U$1601 ( \1916 , \1914 , \1915 );
xnor \U$1602 ( \1917 , \1916 , \530 );
and \U$1603 ( \1918 , \1912 , \1917 );
and \U$1604 ( \1919 , \1908 , \1917 );
or \U$1605 ( \1920 , \1913 , \1918 , \1919 );
and \U$1606 ( \1921 , \425 , \1360 );
and \U$1607 ( \1922 , \417 , \1358 );
nor \U$1608 ( \1923 , \1921 , \1922 );
xnor \U$1609 ( \1924 , \1923 , \1224 );
and \U$1610 ( \1925 , \499 , \1160 );
and \U$1611 ( \1926 , \494 , \1158 );
nor \U$1612 ( \1927 , \1925 , \1926 );
xnor \U$1613 ( \1928 , \1927 , \1082 );
and \U$1614 ( \1929 , \1924 , \1928 );
and \U$1615 ( \1930 , \604 , \996 );
and \U$1616 ( \1931 , \553 , \994 );
nor \U$1617 ( \1932 , \1930 , \1931 );
xnor \U$1618 ( \1933 , \1932 , \902 );
and \U$1619 ( \1934 , \1928 , \1933 );
and \U$1620 ( \1935 , \1924 , \1933 );
or \U$1621 ( \1936 , \1929 , \1934 , \1935 );
and \U$1622 ( \1937 , \1920 , \1936 );
buf \U$1623 ( \1938 , RIc0c8b98_27);
buf \U$1624 ( \1939 , RIc0c8b20_28);
and \U$1625 ( \1940 , \1938 , \1939 );
not \U$1626 ( \1941 , \1940 );
and \U$1627 ( \1942 , \1667 , \1941 );
not \U$1628 ( \1943 , \1942 );
and \U$1629 ( \1944 , \330 , \1826 );
and \U$1630 ( \1945 , \316 , \1824 );
nor \U$1631 ( \1946 , \1944 , \1945 );
xnor \U$1632 ( \1947 , \1946 , \1670 );
and \U$1633 ( \1948 , \1943 , \1947 );
and \U$1634 ( \1949 , \369 , \1554 );
and \U$1635 ( \1950 , \348 , \1552 );
nor \U$1636 ( \1951 , \1949 , \1950 );
xnor \U$1637 ( \1952 , \1951 , \1441 );
and \U$1638 ( \1953 , \1947 , \1952 );
and \U$1639 ( \1954 , \1943 , \1952 );
or \U$1640 ( \1955 , \1948 , \1953 , \1954 );
and \U$1641 ( \1956 , \1936 , \1955 );
and \U$1642 ( \1957 , \1920 , \1955 );
or \U$1643 ( \1958 , \1937 , \1956 , \1957 );
xor \U$1644 ( \1959 , \1810 , \1814 );
xor \U$1645 ( \1960 , \1959 , \1819 );
xor \U$1646 ( \1961 , \1829 , \1833 );
xor \U$1647 ( \1962 , \1961 , \1838 );
and \U$1648 ( \1963 , \1960 , \1962 );
xor \U$1649 ( \1964 , \1846 , \1850 );
xor \U$1650 ( \1965 , \1964 , \1855 );
and \U$1651 ( \1966 , \1962 , \1965 );
and \U$1652 ( \1967 , \1960 , \1965 );
or \U$1653 ( \1968 , \1963 , \1966 , \1967 );
and \U$1654 ( \1969 , \1958 , \1968 );
and \U$1655 ( \1970 , \1274 , \478 );
and \U$1656 ( \1971 , \1186 , \476 );
nor \U$1657 ( \1972 , \1970 , \1971 );
xnor \U$1658 ( \1973 , \1972 , \437 );
and \U$1659 ( \1974 , \1384 , \408 );
and \U$1660 ( \1975 , \1379 , \406 );
nor \U$1661 ( \1976 , \1974 , \1975 );
xnor \U$1662 ( \1977 , \1976 , \378 );
and \U$1663 ( \1978 , \1973 , \1977 );
and \U$1664 ( \1979 , \1615 , \360 );
and \U$1665 ( \1980 , \1500 , \358 );
nor \U$1666 ( \1981 , \1979 , \1980 );
xnor \U$1667 ( \1982 , \1981 , \341 );
and \U$1668 ( \1983 , \1977 , \1982 );
and \U$1669 ( \1984 , \1973 , \1982 );
or \U$1670 ( \1985 , \1978 , \1983 , \1984 );
xor \U$1671 ( \1986 , \1785 , \1789 );
xor \U$1672 ( \1987 , \1986 , \1795 );
and \U$1673 ( \1988 , \1985 , \1987 );
not \U$1674 ( \1989 , \1800 );
and \U$1675 ( \1990 , \1987 , \1989 );
and \U$1676 ( \1991 , \1985 , \1989 );
or \U$1677 ( \1992 , \1988 , \1990 , \1991 );
and \U$1678 ( \1993 , \1968 , \1992 );
and \U$1679 ( \1994 , \1958 , \1992 );
or \U$1680 ( \1995 , \1969 , \1993 , \1994 );
xor \U$1681 ( \1996 , \1671 , \1675 );
xor \U$1682 ( \1997 , \1996 , \1680 );
xor \U$1683 ( \1998 , \1798 , \1801 );
xor \U$1684 ( \1999 , \1998 , \1803 );
and \U$1685 ( \2000 , \1997 , \1999 );
xor \U$1686 ( \2001 , \1864 , \1866 );
xor \U$1687 ( \2002 , \2001 , \1869 );
and \U$1688 ( \2003 , \1999 , \2002 );
and \U$1689 ( \2004 , \1997 , \2002 );
or \U$1690 ( \2005 , \2000 , \2003 , \2004 );
and \U$1691 ( \2006 , \1995 , \2005 );
xor \U$1692 ( \2007 , \1877 , \1879 );
xor \U$1693 ( \2008 , \2007 , \1881 );
and \U$1694 ( \2009 , \2005 , \2008 );
and \U$1695 ( \2010 , \1995 , \2008 );
or \U$1696 ( \2011 , \2006 , \2009 , \2010 );
xor \U$1697 ( \2012 , \1719 , \1729 );
xor \U$1698 ( \2013 , \2012 , \1749 );
and \U$1699 ( \2014 , \2011 , \2013 );
xor \U$1700 ( \2015 , \1875 , \1884 );
xor \U$1701 ( \2016 , \2015 , \1887 );
and \U$1702 ( \2017 , \2013 , \2016 );
and \U$1703 ( \2018 , \2011 , \2016 );
or \U$1704 ( \2019 , \2014 , \2017 , \2018 );
xor \U$1705 ( \2020 , \1890 , \1892 );
xor \U$1706 ( \2021 , \2020 , \1895 );
and \U$1707 ( \2022 , \2019 , \2021 );
and \U$1708 ( \2023 , \1904 , \2022 );
xor \U$1709 ( \2024 , \1904 , \2022 );
xor \U$1710 ( \2025 , \2019 , \2021 );
and \U$1711 ( \2026 , \1379 , \478 );
and \U$1712 ( \2027 , \1274 , \476 );
nor \U$1713 ( \2028 , \2026 , \2027 );
xnor \U$1714 ( \2029 , \2028 , \437 );
and \U$1715 ( \2030 , \1500 , \408 );
and \U$1716 ( \2031 , \1384 , \406 );
nor \U$1717 ( \2032 , \2030 , \2031 );
xnor \U$1718 ( \2033 , \2032 , \378 );
and \U$1719 ( \2034 , \2029 , \2033 );
and \U$1720 ( \2035 , \1791 , \360 );
and \U$1721 ( \2036 , \1615 , \358 );
nor \U$1722 ( \2037 , \2035 , \2036 );
xnor \U$1723 ( \2038 , \2037 , \341 );
and \U$1724 ( \2039 , \2033 , \2038 );
and \U$1725 ( \2040 , \2029 , \2038 );
or \U$1726 ( \2041 , \2034 , \2039 , \2040 );
buf \U$1727 ( \2042 , RIc0c6e10_90);
and \U$1728 ( \2043 , \2042 , \323 );
and \U$1729 ( \2044 , \1799 , \321 );
nor \U$1730 ( \2045 , \2043 , \2044 );
xnor \U$1731 ( \2046 , \2045 , \328 );
buf \U$1732 ( \2047 , RIc0c6d98_91);
and \U$1733 ( \2048 , \2047 , \317 );
or \U$1734 ( \2049 , \2046 , \2048 );
and \U$1735 ( \2050 , \2041 , \2049 );
and \U$1736 ( \2051 , \1799 , \323 );
and \U$1737 ( \2052 , \1791 , \321 );
nor \U$1738 ( \2053 , \2051 , \2052 );
xnor \U$1739 ( \2054 , \2053 , \328 );
and \U$1740 ( \2055 , \2049 , \2054 );
and \U$1741 ( \2056 , \2041 , \2054 );
or \U$1742 ( \2057 , \2050 , \2055 , \2056 );
and \U$1743 ( \2058 , \789 , \826 );
and \U$1744 ( \2059 , \709 , \824 );
nor \U$1745 ( \2060 , \2058 , \2059 );
xnor \U$1746 ( \2061 , \2060 , \754 );
and \U$1747 ( \2062 , \925 , \692 );
and \U$1748 ( \2063 , \863 , \690 );
nor \U$1749 ( \2064 , \2062 , \2063 );
xnor \U$1750 ( \2065 , \2064 , \649 );
and \U$1751 ( \2066 , \2061 , \2065 );
and \U$1752 ( \2067 , \1186 , \579 );
and \U$1753 ( \2068 , \988 , \577 );
nor \U$1754 ( \2069 , \2067 , \2068 );
xnor \U$1755 ( \2070 , \2069 , \530 );
and \U$1756 ( \2071 , \2065 , \2070 );
and \U$1757 ( \2072 , \2061 , \2070 );
or \U$1758 ( \2073 , \2066 , \2071 , \2072 );
and \U$1759 ( \2074 , \494 , \1360 );
and \U$1760 ( \2075 , \425 , \1358 );
nor \U$1761 ( \2076 , \2074 , \2075 );
xnor \U$1762 ( \2077 , \2076 , \1224 );
and \U$1763 ( \2078 , \553 , \1160 );
and \U$1764 ( \2079 , \499 , \1158 );
nor \U$1765 ( \2080 , \2078 , \2079 );
xnor \U$1766 ( \2081 , \2080 , \1082 );
and \U$1767 ( \2082 , \2077 , \2081 );
and \U$1768 ( \2083 , \681 , \996 );
and \U$1769 ( \2084 , \604 , \994 );
nor \U$1770 ( \2085 , \2083 , \2084 );
xnor \U$1771 ( \2086 , \2085 , \902 );
and \U$1772 ( \2087 , \2081 , \2086 );
and \U$1773 ( \2088 , \2077 , \2086 );
or \U$1774 ( \2089 , \2082 , \2087 , \2088 );
and \U$1775 ( \2090 , \2073 , \2089 );
xor \U$1776 ( \2091 , \1667 , \1938 );
xor \U$1777 ( \2092 , \1938 , \1939 );
not \U$1778 ( \2093 , \2092 );
and \U$1779 ( \2094 , \2091 , \2093 );
and \U$1780 ( \2095 , \316 , \2094 );
not \U$1781 ( \2096 , \2095 );
xnor \U$1782 ( \2097 , \2096 , \1942 );
and \U$1783 ( \2098 , \348 , \1826 );
and \U$1784 ( \2099 , \330 , \1824 );
nor \U$1785 ( \2100 , \2098 , \2099 );
xnor \U$1786 ( \2101 , \2100 , \1670 );
and \U$1787 ( \2102 , \2097 , \2101 );
and \U$1788 ( \2103 , \417 , \1554 );
and \U$1789 ( \2104 , \369 , \1552 );
nor \U$1790 ( \2105 , \2103 , \2104 );
xnor \U$1791 ( \2106 , \2105 , \1441 );
and \U$1792 ( \2107 , \2101 , \2106 );
and \U$1793 ( \2108 , \2097 , \2106 );
or \U$1794 ( \2109 , \2102 , \2107 , \2108 );
and \U$1795 ( \2110 , \2089 , \2109 );
and \U$1796 ( \2111 , \2073 , \2109 );
or \U$1797 ( \2112 , \2090 , \2110 , \2111 );
and \U$1798 ( \2113 , \2057 , \2112 );
and \U$1799 ( \2114 , \2042 , \317 );
xor \U$1800 ( \2115 , \1908 , \1912 );
xor \U$1801 ( \2116 , \2115 , \1917 );
and \U$1802 ( \2117 , \2114 , \2116 );
xor \U$1803 ( \2118 , \1973 , \1977 );
xor \U$1804 ( \2119 , \2118 , \1982 );
and \U$1805 ( \2120 , \2116 , \2119 );
and \U$1806 ( \2121 , \2114 , \2119 );
or \U$1807 ( \2122 , \2117 , \2120 , \2121 );
and \U$1808 ( \2123 , \2112 , \2122 );
and \U$1809 ( \2124 , \2057 , \2122 );
or \U$1810 ( \2125 , \2113 , \2123 , \2124 );
xor \U$1811 ( \2126 , \1920 , \1936 );
xor \U$1812 ( \2127 , \2126 , \1955 );
xor \U$1813 ( \2128 , \1960 , \1962 );
xor \U$1814 ( \2129 , \2128 , \1965 );
and \U$1815 ( \2130 , \2127 , \2129 );
xor \U$1816 ( \2131 , \1985 , \1987 );
xor \U$1817 ( \2132 , \2131 , \1989 );
and \U$1818 ( \2133 , \2129 , \2132 );
and \U$1819 ( \2134 , \2127 , \2132 );
or \U$1820 ( \2135 , \2130 , \2133 , \2134 );
and \U$1821 ( \2136 , \2125 , \2135 );
xor \U$1822 ( \2137 , \1822 , \1841 );
xor \U$1823 ( \2138 , \2137 , \1858 );
and \U$1824 ( \2139 , \2135 , \2138 );
and \U$1825 ( \2140 , \2125 , \2138 );
or \U$1826 ( \2141 , \2136 , \2139 , \2140 );
xor \U$1827 ( \2142 , \1958 , \1968 );
xor \U$1828 ( \2143 , \2142 , \1992 );
xor \U$1829 ( \2144 , \1997 , \1999 );
xor \U$1830 ( \2145 , \2144 , \2002 );
and \U$1831 ( \2146 , \2143 , \2145 );
and \U$1832 ( \2147 , \2141 , \2146 );
xor \U$1833 ( \2148 , \1806 , \1861 );
xor \U$1834 ( \2149 , \2148 , \1872 );
and \U$1835 ( \2150 , \2146 , \2149 );
and \U$1836 ( \2151 , \2141 , \2149 );
or \U$1837 ( \2152 , \2147 , \2150 , \2151 );
xor \U$1838 ( \2153 , \2011 , \2013 );
xor \U$1839 ( \2154 , \2153 , \2016 );
and \U$1840 ( \2155 , \2152 , \2154 );
and \U$1841 ( \2156 , \2025 , \2155 );
xor \U$1842 ( \2157 , \2025 , \2155 );
xor \U$1843 ( \2158 , \2152 , \2154 );
buf \U$1844 ( \2159 , RIc0c8aa8_29);
buf \U$1845 ( \2160 , RIc0c8a30_30);
and \U$1846 ( \2161 , \2159 , \2160 );
not \U$1847 ( \2162 , \2161 );
and \U$1848 ( \2163 , \1939 , \2162 );
not \U$1849 ( \2164 , \2163 );
and \U$1850 ( \2165 , \330 , \2094 );
and \U$1851 ( \2166 , \316 , \2092 );
nor \U$1852 ( \2167 , \2165 , \2166 );
xnor \U$1853 ( \2168 , \2167 , \1942 );
and \U$1854 ( \2169 , \2164 , \2168 );
and \U$1855 ( \2170 , \369 , \1826 );
and \U$1856 ( \2171 , \348 , \1824 );
nor \U$1857 ( \2172 , \2170 , \2171 );
xnor \U$1858 ( \2173 , \2172 , \1670 );
and \U$1859 ( \2174 , \2168 , \2173 );
and \U$1860 ( \2175 , \2164 , \2173 );
or \U$1861 ( \2176 , \2169 , \2174 , \2175 );
and \U$1862 ( \2177 , \425 , \1554 );
and \U$1863 ( \2178 , \417 , \1552 );
nor \U$1864 ( \2179 , \2177 , \2178 );
xnor \U$1865 ( \2180 , \2179 , \1441 );
and \U$1866 ( \2181 , \499 , \1360 );
and \U$1867 ( \2182 , \494 , \1358 );
nor \U$1868 ( \2183 , \2181 , \2182 );
xnor \U$1869 ( \2184 , \2183 , \1224 );
and \U$1870 ( \2185 , \2180 , \2184 );
and \U$1871 ( \2186 , \604 , \1160 );
and \U$1872 ( \2187 , \553 , \1158 );
nor \U$1873 ( \2188 , \2186 , \2187 );
xnor \U$1874 ( \2189 , \2188 , \1082 );
and \U$1875 ( \2190 , \2184 , \2189 );
and \U$1876 ( \2191 , \2180 , \2189 );
or \U$1877 ( \2192 , \2185 , \2190 , \2191 );
and \U$1878 ( \2193 , \2176 , \2192 );
and \U$1879 ( \2194 , \709 , \996 );
and \U$1880 ( \2195 , \681 , \994 );
nor \U$1881 ( \2196 , \2194 , \2195 );
xnor \U$1882 ( \2197 , \2196 , \902 );
and \U$1883 ( \2198 , \863 , \826 );
and \U$1884 ( \2199 , \789 , \824 );
nor \U$1885 ( \2200 , \2198 , \2199 );
xnor \U$1886 ( \2201 , \2200 , \754 );
and \U$1887 ( \2202 , \2197 , \2201 );
and \U$1888 ( \2203 , \988 , \692 );
and \U$1889 ( \2204 , \925 , \690 );
nor \U$1890 ( \2205 , \2203 , \2204 );
xnor \U$1891 ( \2206 , \2205 , \649 );
and \U$1892 ( \2207 , \2201 , \2206 );
and \U$1893 ( \2208 , \2197 , \2206 );
or \U$1894 ( \2209 , \2202 , \2207 , \2208 );
and \U$1895 ( \2210 , \2192 , \2209 );
and \U$1896 ( \2211 , \2176 , \2209 );
or \U$1897 ( \2212 , \2193 , \2210 , \2211 );
xor \U$1898 ( \2213 , \2061 , \2065 );
xor \U$1899 ( \2214 , \2213 , \2070 );
xor \U$1900 ( \2215 , \2077 , \2081 );
xor \U$1901 ( \2216 , \2215 , \2086 );
and \U$1902 ( \2217 , \2214 , \2216 );
xor \U$1903 ( \2218 , \2029 , \2033 );
xor \U$1904 ( \2219 , \2218 , \2038 );
and \U$1905 ( \2220 , \2216 , \2219 );
and \U$1906 ( \2221 , \2214 , \2219 );
or \U$1907 ( \2222 , \2217 , \2220 , \2221 );
and \U$1908 ( \2223 , \2212 , \2222 );
and \U$1909 ( \2224 , \1799 , \360 );
and \U$1910 ( \2225 , \1791 , \358 );
nor \U$1911 ( \2226 , \2224 , \2225 );
xnor \U$1912 ( \2227 , \2226 , \341 );
and \U$1913 ( \2228 , \2047 , \323 );
and \U$1914 ( \2229 , \2042 , \321 );
nor \U$1915 ( \2230 , \2228 , \2229 );
xnor \U$1916 ( \2231 , \2230 , \328 );
and \U$1917 ( \2232 , \2227 , \2231 );
buf \U$1918 ( \2233 , RIc0c6d20_92);
and \U$1919 ( \2234 , \2233 , \317 );
and \U$1920 ( \2235 , \2231 , \2234 );
and \U$1921 ( \2236 , \2227 , \2234 );
or \U$1922 ( \2237 , \2232 , \2235 , \2236 );
and \U$1923 ( \2238 , \1274 , \579 );
and \U$1924 ( \2239 , \1186 , \577 );
nor \U$1925 ( \2240 , \2238 , \2239 );
xnor \U$1926 ( \2241 , \2240 , \530 );
and \U$1927 ( \2242 , \1384 , \478 );
and \U$1928 ( \2243 , \1379 , \476 );
nor \U$1929 ( \2244 , \2242 , \2243 );
xnor \U$1930 ( \2245 , \2244 , \437 );
and \U$1931 ( \2246 , \2241 , \2245 );
and \U$1932 ( \2247 , \1615 , \408 );
and \U$1933 ( \2248 , \1500 , \406 );
nor \U$1934 ( \2249 , \2247 , \2248 );
xnor \U$1935 ( \2250 , \2249 , \378 );
and \U$1936 ( \2251 , \2245 , \2250 );
and \U$1937 ( \2252 , \2241 , \2250 );
or \U$1938 ( \2253 , \2246 , \2251 , \2252 );
and \U$1939 ( \2254 , \2237 , \2253 );
xnor \U$1940 ( \2255 , \2046 , \2048 );
and \U$1941 ( \2256 , \2253 , \2255 );
and \U$1942 ( \2257 , \2237 , \2255 );
or \U$1943 ( \2258 , \2254 , \2256 , \2257 );
and \U$1944 ( \2259 , \2222 , \2258 );
and \U$1945 ( \2260 , \2212 , \2258 );
or \U$1946 ( \2261 , \2223 , \2259 , \2260 );
xor \U$1947 ( \2262 , \1924 , \1928 );
xor \U$1948 ( \2263 , \2262 , \1933 );
xor \U$1949 ( \2264 , \1943 , \1947 );
xor \U$1950 ( \2265 , \2264 , \1952 );
and \U$1951 ( \2266 , \2263 , \2265 );
xor \U$1952 ( \2267 , \2114 , \2116 );
xor \U$1953 ( \2268 , \2267 , \2119 );
and \U$1954 ( \2269 , \2265 , \2268 );
and \U$1955 ( \2270 , \2263 , \2268 );
or \U$1956 ( \2271 , \2266 , \2269 , \2270 );
and \U$1957 ( \2272 , \2261 , \2271 );
xor \U$1958 ( \2273 , \2127 , \2129 );
xor \U$1959 ( \2274 , \2273 , \2132 );
and \U$1960 ( \2275 , \2271 , \2274 );
and \U$1961 ( \2276 , \2261 , \2274 );
or \U$1962 ( \2277 , \2272 , \2275 , \2276 );
xor \U$1963 ( \2278 , \2125 , \2135 );
xor \U$1964 ( \2279 , \2278 , \2138 );
and \U$1965 ( \2280 , \2277 , \2279 );
xor \U$1966 ( \2281 , \2143 , \2145 );
and \U$1967 ( \2282 , \2279 , \2281 );
and \U$1968 ( \2283 , \2277 , \2281 );
or \U$1969 ( \2284 , \2280 , \2282 , \2283 );
xor \U$1970 ( \2285 , \2141 , \2146 );
xor \U$1971 ( \2286 , \2285 , \2149 );
and \U$1972 ( \2287 , \2284 , \2286 );
xor \U$1973 ( \2288 , \1995 , \2005 );
xor \U$1974 ( \2289 , \2288 , \2008 );
and \U$1975 ( \2290 , \2286 , \2289 );
and \U$1976 ( \2291 , \2284 , \2289 );
or \U$1977 ( \2292 , \2287 , \2290 , \2291 );
and \U$1978 ( \2293 , \2158 , \2292 );
xor \U$1979 ( \2294 , \2158 , \2292 );
xor \U$1980 ( \2295 , \2284 , \2286 );
xor \U$1981 ( \2296 , \2295 , \2289 );
xor \U$1982 ( \2297 , \1939 , \2159 );
xor \U$1983 ( \2298 , \2159 , \2160 );
not \U$1984 ( \2299 , \2298 );
and \U$1985 ( \2300 , \2297 , \2299 );
and \U$1986 ( \2301 , \316 , \2300 );
not \U$1987 ( \2302 , \2301 );
xnor \U$1988 ( \2303 , \2302 , \2163 );
and \U$1989 ( \2304 , \348 , \2094 );
and \U$1990 ( \2305 , \330 , \2092 );
nor \U$1991 ( \2306 , \2304 , \2305 );
xnor \U$1992 ( \2307 , \2306 , \1942 );
and \U$1993 ( \2308 , \2303 , \2307 );
and \U$1994 ( \2309 , \417 , \1826 );
and \U$1995 ( \2310 , \369 , \1824 );
nor \U$1996 ( \2311 , \2309 , \2310 );
xnor \U$1997 ( \2312 , \2311 , \1670 );
and \U$1998 ( \2313 , \2307 , \2312 );
and \U$1999 ( \2314 , \2303 , \2312 );
or \U$2000 ( \2315 , \2308 , \2313 , \2314 );
and \U$2001 ( \2316 , \494 , \1554 );
and \U$2002 ( \2317 , \425 , \1552 );
nor \U$2003 ( \2318 , \2316 , \2317 );
xnor \U$2004 ( \2319 , \2318 , \1441 );
and \U$2005 ( \2320 , \553 , \1360 );
and \U$2006 ( \2321 , \499 , \1358 );
nor \U$2007 ( \2322 , \2320 , \2321 );
xnor \U$2008 ( \2323 , \2322 , \1224 );
and \U$2009 ( \2324 , \2319 , \2323 );
and \U$2010 ( \2325 , \681 , \1160 );
and \U$2011 ( \2326 , \604 , \1158 );
nor \U$2012 ( \2327 , \2325 , \2326 );
xnor \U$2013 ( \2328 , \2327 , \1082 );
and \U$2014 ( \2329 , \2323 , \2328 );
and \U$2015 ( \2330 , \2319 , \2328 );
or \U$2016 ( \2331 , \2324 , \2329 , \2330 );
and \U$2017 ( \2332 , \2315 , \2331 );
and \U$2018 ( \2333 , \789 , \996 );
and \U$2019 ( \2334 , \709 , \994 );
nor \U$2020 ( \2335 , \2333 , \2334 );
xnor \U$2021 ( \2336 , \2335 , \902 );
and \U$2022 ( \2337 , \925 , \826 );
and \U$2023 ( \2338 , \863 , \824 );
nor \U$2024 ( \2339 , \2337 , \2338 );
xnor \U$2025 ( \2340 , \2339 , \754 );
and \U$2026 ( \2341 , \2336 , \2340 );
and \U$2027 ( \2342 , \1186 , \692 );
and \U$2028 ( \2343 , \988 , \690 );
nor \U$2029 ( \2344 , \2342 , \2343 );
xnor \U$2030 ( \2345 , \2344 , \649 );
and \U$2031 ( \2346 , \2340 , \2345 );
and \U$2032 ( \2347 , \2336 , \2345 );
or \U$2033 ( \2348 , \2341 , \2346 , \2347 );
and \U$2034 ( \2349 , \2331 , \2348 );
and \U$2035 ( \2350 , \2315 , \2348 );
or \U$2036 ( \2351 , \2332 , \2349 , \2350 );
and \U$2037 ( \2352 , \1379 , \579 );
and \U$2038 ( \2353 , \1274 , \577 );
nor \U$2039 ( \2354 , \2352 , \2353 );
xnor \U$2040 ( \2355 , \2354 , \530 );
and \U$2041 ( \2356 , \1500 , \478 );
and \U$2042 ( \2357 , \1384 , \476 );
nor \U$2043 ( \2358 , \2356 , \2357 );
xnor \U$2044 ( \2359 , \2358 , \437 );
and \U$2045 ( \2360 , \2355 , \2359 );
and \U$2046 ( \2361 , \1791 , \408 );
and \U$2047 ( \2362 , \1615 , \406 );
nor \U$2048 ( \2363 , \2361 , \2362 );
xnor \U$2049 ( \2364 , \2363 , \378 );
and \U$2050 ( \2365 , \2359 , \2364 );
and \U$2051 ( \2366 , \2355 , \2364 );
or \U$2052 ( \2367 , \2360 , \2365 , \2366 );
and \U$2053 ( \2368 , \2042 , \360 );
and \U$2054 ( \2369 , \1799 , \358 );
nor \U$2055 ( \2370 , \2368 , \2369 );
xnor \U$2056 ( \2371 , \2370 , \341 );
and \U$2057 ( \2372 , \2233 , \323 );
and \U$2058 ( \2373 , \2047 , \321 );
nor \U$2059 ( \2374 , \2372 , \2373 );
xnor \U$2060 ( \2375 , \2374 , \328 );
and \U$2061 ( \2376 , \2371 , \2375 );
buf \U$2062 ( \2377 , RIc0c6ca8_93);
and \U$2063 ( \2378 , \2377 , \317 );
and \U$2064 ( \2379 , \2375 , \2378 );
and \U$2065 ( \2380 , \2371 , \2378 );
or \U$2066 ( \2381 , \2376 , \2379 , \2380 );
and \U$2067 ( \2382 , \2367 , \2381 );
xor \U$2068 ( \2383 , \2227 , \2231 );
xor \U$2069 ( \2384 , \2383 , \2234 );
and \U$2070 ( \2385 , \2381 , \2384 );
and \U$2071 ( \2386 , \2367 , \2384 );
or \U$2072 ( \2387 , \2382 , \2385 , \2386 );
and \U$2073 ( \2388 , \2351 , \2387 );
xor \U$2074 ( \2389 , \2180 , \2184 );
xor \U$2075 ( \2390 , \2389 , \2189 );
xor \U$2076 ( \2391 , \2241 , \2245 );
xor \U$2077 ( \2392 , \2391 , \2250 );
and \U$2078 ( \2393 , \2390 , \2392 );
xor \U$2079 ( \2394 , \2197 , \2201 );
xor \U$2080 ( \2395 , \2394 , \2206 );
and \U$2081 ( \2396 , \2392 , \2395 );
and \U$2082 ( \2397 , \2390 , \2395 );
or \U$2083 ( \2398 , \2393 , \2396 , \2397 );
and \U$2084 ( \2399 , \2387 , \2398 );
and \U$2085 ( \2400 , \2351 , \2398 );
or \U$2086 ( \2401 , \2388 , \2399 , \2400 );
xor \U$2087 ( \2402 , \2097 , \2101 );
xor \U$2088 ( \2403 , \2402 , \2106 );
xor \U$2089 ( \2404 , \2214 , \2216 );
xor \U$2090 ( \2405 , \2404 , \2219 );
and \U$2091 ( \2406 , \2403 , \2405 );
xor \U$2092 ( \2407 , \2237 , \2253 );
xor \U$2093 ( \2408 , \2407 , \2255 );
and \U$2094 ( \2409 , \2405 , \2408 );
and \U$2095 ( \2410 , \2403 , \2408 );
or \U$2096 ( \2411 , \2406 , \2409 , \2410 );
and \U$2097 ( \2412 , \2401 , \2411 );
xor \U$2098 ( \2413 , \2041 , \2049 );
xor \U$2099 ( \2414 , \2413 , \2054 );
and \U$2100 ( \2415 , \2411 , \2414 );
and \U$2101 ( \2416 , \2401 , \2414 );
or \U$2102 ( \2417 , \2412 , \2415 , \2416 );
xor \U$2103 ( \2418 , \2073 , \2089 );
xor \U$2104 ( \2419 , \2418 , \2109 );
xor \U$2105 ( \2420 , \2212 , \2222 );
xor \U$2106 ( \2421 , \2420 , \2258 );
and \U$2107 ( \2422 , \2419 , \2421 );
xor \U$2108 ( \2423 , \2263 , \2265 );
xor \U$2109 ( \2424 , \2423 , \2268 );
and \U$2110 ( \2425 , \2421 , \2424 );
and \U$2111 ( \2426 , \2419 , \2424 );
or \U$2112 ( \2427 , \2422 , \2425 , \2426 );
and \U$2113 ( \2428 , \2417 , \2427 );
xor \U$2114 ( \2429 , \2057 , \2112 );
xor \U$2115 ( \2430 , \2429 , \2122 );
and \U$2116 ( \2431 , \2427 , \2430 );
and \U$2117 ( \2432 , \2417 , \2430 );
or \U$2118 ( \2433 , \2428 , \2431 , \2432 );
and \U$2119 ( \2434 , \425 , \1826 );
and \U$2120 ( \2435 , \417 , \1824 );
nor \U$2121 ( \2436 , \2434 , \2435 );
xnor \U$2122 ( \2437 , \2436 , \1670 );
and \U$2123 ( \2438 , \499 , \1554 );
and \U$2124 ( \2439 , \494 , \1552 );
nor \U$2125 ( \2440 , \2438 , \2439 );
xnor \U$2126 ( \2441 , \2440 , \1441 );
and \U$2127 ( \2442 , \2437 , \2441 );
and \U$2128 ( \2443 , \604 , \1360 );
and \U$2129 ( \2444 , \553 , \1358 );
nor \U$2130 ( \2445 , \2443 , \2444 );
xnor \U$2131 ( \2446 , \2445 , \1224 );
and \U$2132 ( \2447 , \2441 , \2446 );
and \U$2133 ( \2448 , \2437 , \2446 );
or \U$2134 ( \2449 , \2442 , \2447 , \2448 );
buf \U$2135 ( \2450 , RIc0c89b8_31);
buf \U$2136 ( \2451 , RIc0c8940_32);
and \U$2137 ( \2452 , \2450 , \2451 );
not \U$2138 ( \2453 , \2452 );
and \U$2139 ( \2454 , \2160 , \2453 );
not \U$2140 ( \2455 , \2454 );
and \U$2141 ( \2456 , \330 , \2300 );
and \U$2142 ( \2457 , \316 , \2298 );
nor \U$2143 ( \2458 , \2456 , \2457 );
xnor \U$2144 ( \2459 , \2458 , \2163 );
and \U$2145 ( \2460 , \2455 , \2459 );
and \U$2146 ( \2461 , \369 , \2094 );
and \U$2147 ( \2462 , \348 , \2092 );
nor \U$2148 ( \2463 , \2461 , \2462 );
xnor \U$2149 ( \2464 , \2463 , \1942 );
and \U$2150 ( \2465 , \2459 , \2464 );
and \U$2151 ( \2466 , \2455 , \2464 );
or \U$2152 ( \2467 , \2460 , \2465 , \2466 );
and \U$2153 ( \2468 , \2449 , \2467 );
and \U$2154 ( \2469 , \709 , \1160 );
and \U$2155 ( \2470 , \681 , \1158 );
nor \U$2156 ( \2471 , \2469 , \2470 );
xnor \U$2157 ( \2472 , \2471 , \1082 );
and \U$2158 ( \2473 , \863 , \996 );
and \U$2159 ( \2474 , \789 , \994 );
nor \U$2160 ( \2475 , \2473 , \2474 );
xnor \U$2161 ( \2476 , \2475 , \902 );
and \U$2162 ( \2477 , \2472 , \2476 );
and \U$2163 ( \2478 , \988 , \826 );
and \U$2164 ( \2479 , \925 , \824 );
nor \U$2165 ( \2480 , \2478 , \2479 );
xnor \U$2166 ( \2481 , \2480 , \754 );
and \U$2167 ( \2482 , \2476 , \2481 );
and \U$2168 ( \2483 , \2472 , \2481 );
or \U$2169 ( \2484 , \2477 , \2482 , \2483 );
and \U$2170 ( \2485 , \2467 , \2484 );
and \U$2171 ( \2486 , \2449 , \2484 );
or \U$2172 ( \2487 , \2468 , \2485 , \2486 );
xor \U$2173 ( \2488 , \2355 , \2359 );
xor \U$2174 ( \2489 , \2488 , \2364 );
xor \U$2175 ( \2490 , \2371 , \2375 );
xor \U$2176 ( \2491 , \2490 , \2378 );
and \U$2177 ( \2492 , \2489 , \2491 );
xor \U$2178 ( \2493 , \2336 , \2340 );
xor \U$2179 ( \2494 , \2493 , \2345 );
and \U$2180 ( \2495 , \2491 , \2494 );
and \U$2181 ( \2496 , \2489 , \2494 );
or \U$2182 ( \2497 , \2492 , \2495 , \2496 );
and \U$2183 ( \2498 , \2487 , \2497 );
and \U$2184 ( \2499 , \1799 , \408 );
and \U$2185 ( \2500 , \1791 , \406 );
nor \U$2186 ( \2501 , \2499 , \2500 );
xnor \U$2187 ( \2502 , \2501 , \378 );
and \U$2188 ( \2503 , \2047 , \360 );
and \U$2189 ( \2504 , \2042 , \358 );
nor \U$2190 ( \2505 , \2503 , \2504 );
xnor \U$2191 ( \2506 , \2505 , \341 );
and \U$2192 ( \2507 , \2502 , \2506 );
and \U$2193 ( \2508 , \2377 , \323 );
and \U$2194 ( \2509 , \2233 , \321 );
nor \U$2195 ( \2510 , \2508 , \2509 );
xnor \U$2196 ( \2511 , \2510 , \328 );
and \U$2197 ( \2512 , \2506 , \2511 );
and \U$2198 ( \2513 , \2502 , \2511 );
or \U$2199 ( \2514 , \2507 , \2512 , \2513 );
and \U$2200 ( \2515 , \1274 , \692 );
and \U$2201 ( \2516 , \1186 , \690 );
nor \U$2202 ( \2517 , \2515 , \2516 );
xnor \U$2203 ( \2518 , \2517 , \649 );
and \U$2204 ( \2519 , \1384 , \579 );
and \U$2205 ( \2520 , \1379 , \577 );
nor \U$2206 ( \2521 , \2519 , \2520 );
xnor \U$2207 ( \2522 , \2521 , \530 );
and \U$2208 ( \2523 , \2518 , \2522 );
and \U$2209 ( \2524 , \1615 , \478 );
and \U$2210 ( \2525 , \1500 , \476 );
nor \U$2211 ( \2526 , \2524 , \2525 );
xnor \U$2212 ( \2527 , \2526 , \437 );
and \U$2213 ( \2528 , \2522 , \2527 );
and \U$2214 ( \2529 , \2518 , \2527 );
or \U$2215 ( \2530 , \2523 , \2528 , \2529 );
or \U$2216 ( \2531 , \2514 , \2530 );
and \U$2217 ( \2532 , \2497 , \2531 );
and \U$2218 ( \2533 , \2487 , \2531 );
or \U$2219 ( \2534 , \2498 , \2532 , \2533 );
xor \U$2220 ( \2535 , \2164 , \2168 );
xor \U$2221 ( \2536 , \2535 , \2173 );
xor \U$2222 ( \2537 , \2367 , \2381 );
xor \U$2223 ( \2538 , \2537 , \2384 );
and \U$2224 ( \2539 , \2536 , \2538 );
xor \U$2225 ( \2540 , \2390 , \2392 );
xor \U$2226 ( \2541 , \2540 , \2395 );
and \U$2227 ( \2542 , \2538 , \2541 );
and \U$2228 ( \2543 , \2536 , \2541 );
or \U$2229 ( \2544 , \2539 , \2542 , \2543 );
and \U$2230 ( \2545 , \2534 , \2544 );
xor \U$2231 ( \2546 , \2176 , \2192 );
xor \U$2232 ( \2547 , \2546 , \2209 );
and \U$2233 ( \2548 , \2544 , \2547 );
and \U$2234 ( \2549 , \2534 , \2547 );
or \U$2235 ( \2550 , \2545 , \2548 , \2549 );
xor \U$2236 ( \2551 , \2401 , \2411 );
xor \U$2237 ( \2552 , \2551 , \2414 );
and \U$2238 ( \2553 , \2550 , \2552 );
xor \U$2239 ( \2554 , \2419 , \2421 );
xor \U$2240 ( \2555 , \2554 , \2424 );
and \U$2241 ( \2556 , \2552 , \2555 );
and \U$2242 ( \2557 , \2550 , \2555 );
or \U$2243 ( \2558 , \2553 , \2556 , \2557 );
xor \U$2244 ( \2559 , \2417 , \2427 );
xor \U$2245 ( \2560 , \2559 , \2430 );
and \U$2246 ( \2561 , \2558 , \2560 );
xor \U$2247 ( \2562 , \2261 , \2271 );
xor \U$2248 ( \2563 , \2562 , \2274 );
and \U$2249 ( \2564 , \2560 , \2563 );
and \U$2250 ( \2565 , \2558 , \2563 );
or \U$2251 ( \2566 , \2561 , \2564 , \2565 );
and \U$2252 ( \2567 , \2433 , \2566 );
xor \U$2253 ( \2568 , \2277 , \2279 );
xor \U$2254 ( \2569 , \2568 , \2281 );
and \U$2255 ( \2570 , \2566 , \2569 );
and \U$2256 ( \2571 , \2433 , \2569 );
or \U$2257 ( \2572 , \2567 , \2570 , \2571 );
and \U$2258 ( \2573 , \2296 , \2572 );
xor \U$2259 ( \2574 , \2296 , \2572 );
xor \U$2260 ( \2575 , \2433 , \2566 );
xor \U$2261 ( \2576 , \2575 , \2569 );
and \U$2262 ( \2577 , \494 , \1826 );
and \U$2263 ( \2578 , \425 , \1824 );
nor \U$2264 ( \2579 , \2577 , \2578 );
xnor \U$2265 ( \2580 , \2579 , \1670 );
and \U$2266 ( \2581 , \553 , \1554 );
and \U$2267 ( \2582 , \499 , \1552 );
nor \U$2268 ( \2583 , \2581 , \2582 );
xnor \U$2269 ( \2584 , \2583 , \1441 );
and \U$2270 ( \2585 , \2580 , \2584 );
and \U$2271 ( \2586 , \681 , \1360 );
and \U$2272 ( \2587 , \604 , \1358 );
nor \U$2273 ( \2588 , \2586 , \2587 );
xnor \U$2274 ( \2589 , \2588 , \1224 );
and \U$2275 ( \2590 , \2584 , \2589 );
and \U$2276 ( \2591 , \2580 , \2589 );
or \U$2277 ( \2592 , \2585 , \2590 , \2591 );
xor \U$2278 ( \2593 , \2160 , \2450 );
xor \U$2279 ( \2594 , \2450 , \2451 );
not \U$2280 ( \2595 , \2594 );
and \U$2281 ( \2596 , \2593 , \2595 );
and \U$2282 ( \2597 , \316 , \2596 );
not \U$2283 ( \2598 , \2597 );
xnor \U$2284 ( \2599 , \2598 , \2454 );
and \U$2285 ( \2600 , \348 , \2300 );
and \U$2286 ( \2601 , \330 , \2298 );
nor \U$2287 ( \2602 , \2600 , \2601 );
xnor \U$2288 ( \2603 , \2602 , \2163 );
and \U$2289 ( \2604 , \2599 , \2603 );
and \U$2290 ( \2605 , \417 , \2094 );
and \U$2291 ( \2606 , \369 , \2092 );
nor \U$2292 ( \2607 , \2605 , \2606 );
xnor \U$2293 ( \2608 , \2607 , \1942 );
and \U$2294 ( \2609 , \2603 , \2608 );
and \U$2295 ( \2610 , \2599 , \2608 );
or \U$2296 ( \2611 , \2604 , \2609 , \2610 );
and \U$2297 ( \2612 , \2592 , \2611 );
and \U$2298 ( \2613 , \789 , \1160 );
and \U$2299 ( \2614 , \709 , \1158 );
nor \U$2300 ( \2615 , \2613 , \2614 );
xnor \U$2301 ( \2616 , \2615 , \1082 );
and \U$2302 ( \2617 , \925 , \996 );
and \U$2303 ( \2618 , \863 , \994 );
nor \U$2304 ( \2619 , \2617 , \2618 );
xnor \U$2305 ( \2620 , \2619 , \902 );
and \U$2306 ( \2621 , \2616 , \2620 );
and \U$2307 ( \2622 , \1186 , \826 );
and \U$2308 ( \2623 , \988 , \824 );
nor \U$2309 ( \2624 , \2622 , \2623 );
xnor \U$2310 ( \2625 , \2624 , \754 );
and \U$2311 ( \2626 , \2620 , \2625 );
and \U$2312 ( \2627 , \2616 , \2625 );
or \U$2313 ( \2628 , \2621 , \2626 , \2627 );
and \U$2314 ( \2629 , \2611 , \2628 );
and \U$2315 ( \2630 , \2592 , \2628 );
or \U$2316 ( \2631 , \2612 , \2629 , \2630 );
and \U$2317 ( \2632 , \2042 , \408 );
and \U$2318 ( \2633 , \1799 , \406 );
nor \U$2319 ( \2634 , \2632 , \2633 );
xnor \U$2320 ( \2635 , \2634 , \378 );
and \U$2321 ( \2636 , \2233 , \360 );
and \U$2322 ( \2637 , \2047 , \358 );
nor \U$2323 ( \2638 , \2636 , \2637 );
xnor \U$2324 ( \2639 , \2638 , \341 );
and \U$2325 ( \2640 , \2635 , \2639 );
buf \U$2326 ( \2641 , RIc0c6c30_94);
and \U$2327 ( \2642 , \2641 , \323 );
and \U$2328 ( \2643 , \2377 , \321 );
nor \U$2329 ( \2644 , \2642 , \2643 );
xnor \U$2330 ( \2645 , \2644 , \328 );
and \U$2331 ( \2646 , \2639 , \2645 );
and \U$2332 ( \2647 , \2635 , \2645 );
or \U$2333 ( \2648 , \2640 , \2646 , \2647 );
and \U$2334 ( \2649 , \1379 , \692 );
and \U$2335 ( \2650 , \1274 , \690 );
nor \U$2336 ( \2651 , \2649 , \2650 );
xnor \U$2337 ( \2652 , \2651 , \649 );
and \U$2338 ( \2653 , \1500 , \579 );
and \U$2339 ( \2654 , \1384 , \577 );
nor \U$2340 ( \2655 , \2653 , \2654 );
xnor \U$2341 ( \2656 , \2655 , \530 );
and \U$2342 ( \2657 , \2652 , \2656 );
and \U$2343 ( \2658 , \1791 , \478 );
and \U$2344 ( \2659 , \1615 , \476 );
nor \U$2345 ( \2660 , \2658 , \2659 );
xnor \U$2346 ( \2661 , \2660 , \437 );
and \U$2347 ( \2662 , \2656 , \2661 );
and \U$2348 ( \2663 , \2652 , \2661 );
or \U$2349 ( \2664 , \2657 , \2662 , \2663 );
and \U$2350 ( \2665 , \2648 , \2664 );
buf \U$2351 ( \2666 , RIc0c6bb8_95);
and \U$2352 ( \2667 , \2666 , \317 );
buf \U$2353 ( \2668 , \2667 );
and \U$2354 ( \2669 , \2664 , \2668 );
and \U$2355 ( \2670 , \2648 , \2668 );
or \U$2356 ( \2671 , \2665 , \2669 , \2670 );
and \U$2357 ( \2672 , \2631 , \2671 );
and \U$2358 ( \2673 , \2641 , \317 );
xor \U$2359 ( \2674 , \2502 , \2506 );
xor \U$2360 ( \2675 , \2674 , \2511 );
and \U$2361 ( \2676 , \2673 , \2675 );
xor \U$2362 ( \2677 , \2518 , \2522 );
xor \U$2363 ( \2678 , \2677 , \2527 );
and \U$2364 ( \2679 , \2675 , \2678 );
and \U$2365 ( \2680 , \2673 , \2678 );
or \U$2366 ( \2681 , \2676 , \2679 , \2680 );
and \U$2367 ( \2682 , \2671 , \2681 );
and \U$2368 ( \2683 , \2631 , \2681 );
or \U$2369 ( \2684 , \2672 , \2682 , \2683 );
xor \U$2370 ( \2685 , \2437 , \2441 );
xor \U$2371 ( \2686 , \2685 , \2446 );
xor \U$2372 ( \2687 , \2455 , \2459 );
xor \U$2373 ( \2688 , \2687 , \2464 );
and \U$2374 ( \2689 , \2686 , \2688 );
xor \U$2375 ( \2690 , \2472 , \2476 );
xor \U$2376 ( \2691 , \2690 , \2481 );
and \U$2377 ( \2692 , \2688 , \2691 );
and \U$2378 ( \2693 , \2686 , \2691 );
or \U$2379 ( \2694 , \2689 , \2692 , \2693 );
xor \U$2380 ( \2695 , \2303 , \2307 );
xor \U$2381 ( \2696 , \2695 , \2312 );
and \U$2382 ( \2697 , \2694 , \2696 );
xor \U$2383 ( \2698 , \2319 , \2323 );
xor \U$2384 ( \2699 , \2698 , \2328 );
and \U$2385 ( \2700 , \2696 , \2699 );
and \U$2386 ( \2701 , \2694 , \2699 );
or \U$2387 ( \2702 , \2697 , \2700 , \2701 );
and \U$2388 ( \2703 , \2684 , \2702 );
xor \U$2389 ( \2704 , \2449 , \2467 );
xor \U$2390 ( \2705 , \2704 , \2484 );
xor \U$2391 ( \2706 , \2489 , \2491 );
xor \U$2392 ( \2707 , \2706 , \2494 );
and \U$2393 ( \2708 , \2705 , \2707 );
xnor \U$2394 ( \2709 , \2514 , \2530 );
and \U$2395 ( \2710 , \2707 , \2709 );
and \U$2396 ( \2711 , \2705 , \2709 );
or \U$2397 ( \2712 , \2708 , \2710 , \2711 );
and \U$2398 ( \2713 , \2702 , \2712 );
and \U$2399 ( \2714 , \2684 , \2712 );
or \U$2400 ( \2715 , \2703 , \2713 , \2714 );
xor \U$2401 ( \2716 , \2315 , \2331 );
xor \U$2402 ( \2717 , \2716 , \2348 );
xor \U$2403 ( \2718 , \2487 , \2497 );
xor \U$2404 ( \2719 , \2718 , \2531 );
and \U$2405 ( \2720 , \2717 , \2719 );
xor \U$2406 ( \2721 , \2536 , \2538 );
xor \U$2407 ( \2722 , \2721 , \2541 );
and \U$2408 ( \2723 , \2719 , \2722 );
and \U$2409 ( \2724 , \2717 , \2722 );
or \U$2410 ( \2725 , \2720 , \2723 , \2724 );
and \U$2411 ( \2726 , \2715 , \2725 );
xor \U$2412 ( \2727 , \2403 , \2405 );
xor \U$2413 ( \2728 , \2727 , \2408 );
and \U$2414 ( \2729 , \2725 , \2728 );
and \U$2415 ( \2730 , \2715 , \2728 );
or \U$2416 ( \2731 , \2726 , \2729 , \2730 );
xor \U$2417 ( \2732 , \2351 , \2387 );
xor \U$2418 ( \2733 , \2732 , \2398 );
xor \U$2419 ( \2734 , \2534 , \2544 );
xor \U$2420 ( \2735 , \2734 , \2547 );
and \U$2421 ( \2736 , \2733 , \2735 );
and \U$2422 ( \2737 , \2731 , \2736 );
xor \U$2423 ( \2738 , \2550 , \2552 );
xor \U$2424 ( \2739 , \2738 , \2555 );
and \U$2425 ( \2740 , \2736 , \2739 );
and \U$2426 ( \2741 , \2731 , \2739 );
or \U$2427 ( \2742 , \2737 , \2740 , \2741 );
xor \U$2428 ( \2743 , \2558 , \2560 );
xor \U$2429 ( \2744 , \2743 , \2563 );
and \U$2430 ( \2745 , \2742 , \2744 );
and \U$2431 ( \2746 , \2576 , \2745 );
xor \U$2432 ( \2747 , \2576 , \2745 );
xor \U$2433 ( \2748 , \2742 , \2744 );
and \U$2434 ( \2749 , \709 , \1360 );
and \U$2435 ( \2750 , \681 , \1358 );
nor \U$2436 ( \2751 , \2749 , \2750 );
xnor \U$2437 ( \2752 , \2751 , \1224 );
and \U$2438 ( \2753 , \863 , \1160 );
and \U$2439 ( \2754 , \789 , \1158 );
nor \U$2440 ( \2755 , \2753 , \2754 );
xnor \U$2441 ( \2756 , \2755 , \1082 );
and \U$2442 ( \2757 , \2752 , \2756 );
and \U$2443 ( \2758 , \988 , \996 );
and \U$2444 ( \2759 , \925 , \994 );
nor \U$2445 ( \2760 , \2758 , \2759 );
xnor \U$2446 ( \2761 , \2760 , \902 );
and \U$2447 ( \2762 , \2756 , \2761 );
and \U$2448 ( \2763 , \2752 , \2761 );
or \U$2449 ( \2764 , \2757 , \2762 , \2763 );
buf \U$2450 ( \2765 , RIc0c88c8_33);
buf \U$2451 ( \2766 , RIc0c8850_34);
and \U$2452 ( \2767 , \2765 , \2766 );
not \U$2453 ( \2768 , \2767 );
and \U$2454 ( \2769 , \2451 , \2768 );
not \U$2455 ( \2770 , \2769 );
and \U$2456 ( \2771 , \330 , \2596 );
and \U$2457 ( \2772 , \316 , \2594 );
nor \U$2458 ( \2773 , \2771 , \2772 );
xnor \U$2459 ( \2774 , \2773 , \2454 );
and \U$2460 ( \2775 , \2770 , \2774 );
and \U$2461 ( \2776 , \369 , \2300 );
and \U$2462 ( \2777 , \348 , \2298 );
nor \U$2463 ( \2778 , \2776 , \2777 );
xnor \U$2464 ( \2779 , \2778 , \2163 );
and \U$2465 ( \2780 , \2774 , \2779 );
and \U$2466 ( \2781 , \2770 , \2779 );
or \U$2467 ( \2782 , \2775 , \2780 , \2781 );
and \U$2468 ( \2783 , \2764 , \2782 );
and \U$2469 ( \2784 , \425 , \2094 );
and \U$2470 ( \2785 , \417 , \2092 );
nor \U$2471 ( \2786 , \2784 , \2785 );
xnor \U$2472 ( \2787 , \2786 , \1942 );
and \U$2473 ( \2788 , \499 , \1826 );
and \U$2474 ( \2789 , \494 , \1824 );
nor \U$2475 ( \2790 , \2788 , \2789 );
xnor \U$2476 ( \2791 , \2790 , \1670 );
and \U$2477 ( \2792 , \2787 , \2791 );
and \U$2478 ( \2793 , \604 , \1554 );
and \U$2479 ( \2794 , \553 , \1552 );
nor \U$2480 ( \2795 , \2793 , \2794 );
xnor \U$2481 ( \2796 , \2795 , \1441 );
and \U$2482 ( \2797 , \2791 , \2796 );
and \U$2483 ( \2798 , \2787 , \2796 );
or \U$2484 ( \2799 , \2792 , \2797 , \2798 );
and \U$2485 ( \2800 , \2782 , \2799 );
and \U$2486 ( \2801 , \2764 , \2799 );
or \U$2487 ( \2802 , \2783 , \2800 , \2801 );
and \U$2488 ( \2803 , \1799 , \478 );
and \U$2489 ( \2804 , \1791 , \476 );
nor \U$2490 ( \2805 , \2803 , \2804 );
xnor \U$2491 ( \2806 , \2805 , \437 );
and \U$2492 ( \2807 , \2047 , \408 );
and \U$2493 ( \2808 , \2042 , \406 );
nor \U$2494 ( \2809 , \2807 , \2808 );
xnor \U$2495 ( \2810 , \2809 , \378 );
and \U$2496 ( \2811 , \2806 , \2810 );
and \U$2497 ( \2812 , \2377 , \360 );
and \U$2498 ( \2813 , \2233 , \358 );
nor \U$2499 ( \2814 , \2812 , \2813 );
xnor \U$2500 ( \2815 , \2814 , \341 );
and \U$2501 ( \2816 , \2810 , \2815 );
and \U$2502 ( \2817 , \2806 , \2815 );
or \U$2503 ( \2818 , \2811 , \2816 , \2817 );
and \U$2504 ( \2819 , \1274 , \826 );
and \U$2505 ( \2820 , \1186 , \824 );
nor \U$2506 ( \2821 , \2819 , \2820 );
xnor \U$2507 ( \2822 , \2821 , \754 );
and \U$2508 ( \2823 , \1384 , \692 );
and \U$2509 ( \2824 , \1379 , \690 );
nor \U$2510 ( \2825 , \2823 , \2824 );
xnor \U$2511 ( \2826 , \2825 , \649 );
and \U$2512 ( \2827 , \2822 , \2826 );
and \U$2513 ( \2828 , \1615 , \579 );
and \U$2514 ( \2829 , \1500 , \577 );
nor \U$2515 ( \2830 , \2828 , \2829 );
xnor \U$2516 ( \2831 , \2830 , \530 );
and \U$2517 ( \2832 , \2826 , \2831 );
and \U$2518 ( \2833 , \2822 , \2831 );
or \U$2519 ( \2834 , \2827 , \2832 , \2833 );
and \U$2520 ( \2835 , \2818 , \2834 );
and \U$2521 ( \2836 , \2666 , \323 );
and \U$2522 ( \2837 , \2641 , \321 );
nor \U$2523 ( \2838 , \2836 , \2837 );
xnor \U$2524 ( \2839 , \2838 , \328 );
buf \U$2525 ( \2840 , RIc0c6b40_96);
and \U$2526 ( \2841 , \2840 , \317 );
and \U$2527 ( \2842 , \2839 , \2841 );
and \U$2528 ( \2843 , \2834 , \2842 );
and \U$2529 ( \2844 , \2818 , \2842 );
or \U$2530 ( \2845 , \2835 , \2843 , \2844 );
and \U$2531 ( \2846 , \2802 , \2845 );
xor \U$2532 ( \2847 , \2635 , \2639 );
xor \U$2533 ( \2848 , \2847 , \2645 );
xor \U$2534 ( \2849 , \2652 , \2656 );
xor \U$2535 ( \2850 , \2849 , \2661 );
and \U$2536 ( \2851 , \2848 , \2850 );
not \U$2537 ( \2852 , \2667 );
and \U$2538 ( \2853 , \2850 , \2852 );
and \U$2539 ( \2854 , \2848 , \2852 );
or \U$2540 ( \2855 , \2851 , \2853 , \2854 );
and \U$2541 ( \2856 , \2845 , \2855 );
and \U$2542 ( \2857 , \2802 , \2855 );
or \U$2543 ( \2858 , \2846 , \2856 , \2857 );
xor \U$2544 ( \2859 , \2580 , \2584 );
xor \U$2545 ( \2860 , \2859 , \2589 );
xor \U$2546 ( \2861 , \2599 , \2603 );
xor \U$2547 ( \2862 , \2861 , \2608 );
and \U$2548 ( \2863 , \2860 , \2862 );
xor \U$2549 ( \2864 , \2616 , \2620 );
xor \U$2550 ( \2865 , \2864 , \2625 );
and \U$2551 ( \2866 , \2862 , \2865 );
and \U$2552 ( \2867 , \2860 , \2865 );
or \U$2553 ( \2868 , \2863 , \2866 , \2867 );
xor \U$2554 ( \2869 , \2686 , \2688 );
xor \U$2555 ( \2870 , \2869 , \2691 );
and \U$2556 ( \2871 , \2868 , \2870 );
xor \U$2557 ( \2872 , \2673 , \2675 );
xor \U$2558 ( \2873 , \2872 , \2678 );
and \U$2559 ( \2874 , \2870 , \2873 );
and \U$2560 ( \2875 , \2868 , \2873 );
or \U$2561 ( \2876 , \2871 , \2874 , \2875 );
and \U$2562 ( \2877 , \2858 , \2876 );
xor \U$2563 ( \2878 , \2592 , \2611 );
xor \U$2564 ( \2879 , \2878 , \2628 );
xor \U$2565 ( \2880 , \2648 , \2664 );
xor \U$2566 ( \2881 , \2880 , \2668 );
and \U$2567 ( \2882 , \2879 , \2881 );
and \U$2568 ( \2883 , \2876 , \2882 );
and \U$2569 ( \2884 , \2858 , \2882 );
or \U$2570 ( \2885 , \2877 , \2883 , \2884 );
xor \U$2571 ( \2886 , \2631 , \2671 );
xor \U$2572 ( \2887 , \2886 , \2681 );
xor \U$2573 ( \2888 , \2694 , \2696 );
xor \U$2574 ( \2889 , \2888 , \2699 );
and \U$2575 ( \2890 , \2887 , \2889 );
xor \U$2576 ( \2891 , \2705 , \2707 );
xor \U$2577 ( \2892 , \2891 , \2709 );
and \U$2578 ( \2893 , \2889 , \2892 );
and \U$2579 ( \2894 , \2887 , \2892 );
or \U$2580 ( \2895 , \2890 , \2893 , \2894 );
and \U$2581 ( \2896 , \2885 , \2895 );
xor \U$2582 ( \2897 , \2717 , \2719 );
xor \U$2583 ( \2898 , \2897 , \2722 );
and \U$2584 ( \2899 , \2895 , \2898 );
and \U$2585 ( \2900 , \2885 , \2898 );
or \U$2586 ( \2901 , \2896 , \2899 , \2900 );
xor \U$2587 ( \2902 , \2715 , \2725 );
xor \U$2588 ( \2903 , \2902 , \2728 );
and \U$2589 ( \2904 , \2901 , \2903 );
xor \U$2590 ( \2905 , \2733 , \2735 );
and \U$2591 ( \2906 , \2903 , \2905 );
and \U$2592 ( \2907 , \2901 , \2905 );
or \U$2593 ( \2908 , \2904 , \2906 , \2907 );
xor \U$2594 ( \2909 , \2731 , \2736 );
xor \U$2595 ( \2910 , \2909 , \2739 );
and \U$2596 ( \2911 , \2908 , \2910 );
and \U$2597 ( \2912 , \2748 , \2911 );
xor \U$2598 ( \2913 , \2748 , \2911 );
xor \U$2599 ( \2914 , \2908 , \2910 );
xor \U$2600 ( \2915 , \2451 , \2765 );
xor \U$2601 ( \2916 , \2765 , \2766 );
not \U$2602 ( \2917 , \2916 );
and \U$2603 ( \2918 , \2915 , \2917 );
and \U$2604 ( \2919 , \316 , \2918 );
not \U$2605 ( \2920 , \2919 );
xnor \U$2606 ( \2921 , \2920 , \2769 );
and \U$2607 ( \2922 , \348 , \2596 );
and \U$2608 ( \2923 , \330 , \2594 );
nor \U$2609 ( \2924 , \2922 , \2923 );
xnor \U$2610 ( \2925 , \2924 , \2454 );
and \U$2611 ( \2926 , \2921 , \2925 );
and \U$2612 ( \2927 , \417 , \2300 );
and \U$2613 ( \2928 , \369 , \2298 );
nor \U$2614 ( \2929 , \2927 , \2928 );
xnor \U$2615 ( \2930 , \2929 , \2163 );
and \U$2616 ( \2931 , \2925 , \2930 );
and \U$2617 ( \2932 , \2921 , \2930 );
or \U$2618 ( \2933 , \2926 , \2931 , \2932 );
and \U$2619 ( \2934 , \789 , \1360 );
and \U$2620 ( \2935 , \709 , \1358 );
nor \U$2621 ( \2936 , \2934 , \2935 );
xnor \U$2622 ( \2937 , \2936 , \1224 );
and \U$2623 ( \2938 , \925 , \1160 );
and \U$2624 ( \2939 , \863 , \1158 );
nor \U$2625 ( \2940 , \2938 , \2939 );
xnor \U$2626 ( \2941 , \2940 , \1082 );
and \U$2627 ( \2942 , \2937 , \2941 );
and \U$2628 ( \2943 , \1186 , \996 );
and \U$2629 ( \2944 , \988 , \994 );
nor \U$2630 ( \2945 , \2943 , \2944 );
xnor \U$2631 ( \2946 , \2945 , \902 );
and \U$2632 ( \2947 , \2941 , \2946 );
and \U$2633 ( \2948 , \2937 , \2946 );
or \U$2634 ( \2949 , \2942 , \2947 , \2948 );
and \U$2635 ( \2950 , \2933 , \2949 );
and \U$2636 ( \2951 , \494 , \2094 );
and \U$2637 ( \2952 , \425 , \2092 );
nor \U$2638 ( \2953 , \2951 , \2952 );
xnor \U$2639 ( \2954 , \2953 , \1942 );
and \U$2640 ( \2955 , \553 , \1826 );
and \U$2641 ( \2956 , \499 , \1824 );
nor \U$2642 ( \2957 , \2955 , \2956 );
xnor \U$2643 ( \2958 , \2957 , \1670 );
and \U$2644 ( \2959 , \2954 , \2958 );
and \U$2645 ( \2960 , \681 , \1554 );
and \U$2646 ( \2961 , \604 , \1552 );
nor \U$2647 ( \2962 , \2960 , \2961 );
xnor \U$2648 ( \2963 , \2962 , \1441 );
and \U$2649 ( \2964 , \2958 , \2963 );
and \U$2650 ( \2965 , \2954 , \2963 );
or \U$2651 ( \2966 , \2959 , \2964 , \2965 );
and \U$2652 ( \2967 , \2949 , \2966 );
and \U$2653 ( \2968 , \2933 , \2966 );
or \U$2654 ( \2969 , \2950 , \2967 , \2968 );
and \U$2655 ( \2970 , \2042 , \478 );
and \U$2656 ( \2971 , \1799 , \476 );
nor \U$2657 ( \2972 , \2970 , \2971 );
xnor \U$2658 ( \2973 , \2972 , \437 );
and \U$2659 ( \2974 , \2233 , \408 );
and \U$2660 ( \2975 , \2047 , \406 );
nor \U$2661 ( \2976 , \2974 , \2975 );
xnor \U$2662 ( \2977 , \2976 , \378 );
and \U$2663 ( \2978 , \2973 , \2977 );
and \U$2664 ( \2979 , \2641 , \360 );
and \U$2665 ( \2980 , \2377 , \358 );
nor \U$2666 ( \2981 , \2979 , \2980 );
xnor \U$2667 ( \2982 , \2981 , \341 );
and \U$2668 ( \2983 , \2977 , \2982 );
and \U$2669 ( \2984 , \2973 , \2982 );
or \U$2670 ( \2985 , \2978 , \2983 , \2984 );
and \U$2671 ( \2986 , \1379 , \826 );
and \U$2672 ( \2987 , \1274 , \824 );
nor \U$2673 ( \2988 , \2986 , \2987 );
xnor \U$2674 ( \2989 , \2988 , \754 );
and \U$2675 ( \2990 , \1500 , \692 );
and \U$2676 ( \2991 , \1384 , \690 );
nor \U$2677 ( \2992 , \2990 , \2991 );
xnor \U$2678 ( \2993 , \2992 , \649 );
and \U$2679 ( \2994 , \2989 , \2993 );
and \U$2680 ( \2995 , \1791 , \579 );
and \U$2681 ( \2996 , \1615 , \577 );
nor \U$2682 ( \2997 , \2995 , \2996 );
xnor \U$2683 ( \2998 , \2997 , \530 );
and \U$2684 ( \2999 , \2993 , \2998 );
and \U$2685 ( \3000 , \2989 , \2998 );
or \U$2686 ( \3001 , \2994 , \2999 , \3000 );
and \U$2687 ( \3002 , \2985 , \3001 );
and \U$2688 ( \3003 , \2840 , \323 );
and \U$2689 ( \3004 , \2666 , \321 );
nor \U$2690 ( \3005 , \3003 , \3004 );
xnor \U$2691 ( \3006 , \3005 , \328 );
buf \U$2692 ( \3007 , RIc0c6ac8_97);
and \U$2693 ( \3008 , \3007 , \317 );
or \U$2694 ( \3009 , \3006 , \3008 );
and \U$2695 ( \3010 , \3001 , \3009 );
and \U$2696 ( \3011 , \2985 , \3009 );
or \U$2697 ( \3012 , \3002 , \3010 , \3011 );
and \U$2698 ( \3013 , \2969 , \3012 );
xor \U$2699 ( \3014 , \2806 , \2810 );
xor \U$2700 ( \3015 , \3014 , \2815 );
xor \U$2701 ( \3016 , \2822 , \2826 );
xor \U$2702 ( \3017 , \3016 , \2831 );
and \U$2703 ( \3018 , \3015 , \3017 );
xor \U$2704 ( \3019 , \2839 , \2841 );
and \U$2705 ( \3020 , \3017 , \3019 );
and \U$2706 ( \3021 , \3015 , \3019 );
or \U$2707 ( \3022 , \3018 , \3020 , \3021 );
and \U$2708 ( \3023 , \3012 , \3022 );
and \U$2709 ( \3024 , \2969 , \3022 );
or \U$2710 ( \3025 , \3013 , \3023 , \3024 );
xor \U$2711 ( \3026 , \2752 , \2756 );
xor \U$2712 ( \3027 , \3026 , \2761 );
xor \U$2713 ( \3028 , \2770 , \2774 );
xor \U$2714 ( \3029 , \3028 , \2779 );
and \U$2715 ( \3030 , \3027 , \3029 );
xor \U$2716 ( \3031 , \2787 , \2791 );
xor \U$2717 ( \3032 , \3031 , \2796 );
and \U$2718 ( \3033 , \3029 , \3032 );
and \U$2719 ( \3034 , \3027 , \3032 );
or \U$2720 ( \3035 , \3030 , \3033 , \3034 );
xor \U$2721 ( \3036 , \2860 , \2862 );
xor \U$2722 ( \3037 , \3036 , \2865 );
and \U$2723 ( \3038 , \3035 , \3037 );
xor \U$2724 ( \3039 , \2848 , \2850 );
xor \U$2725 ( \3040 , \3039 , \2852 );
and \U$2726 ( \3041 , \3037 , \3040 );
and \U$2727 ( \3042 , \3035 , \3040 );
or \U$2728 ( \3043 , \3038 , \3041 , \3042 );
and \U$2729 ( \3044 , \3025 , \3043 );
xor \U$2730 ( \3045 , \2764 , \2782 );
xor \U$2731 ( \3046 , \3045 , \2799 );
xor \U$2732 ( \3047 , \2818 , \2834 );
xor \U$2733 ( \3048 , \3047 , \2842 );
and \U$2734 ( \3049 , \3046 , \3048 );
and \U$2735 ( \3050 , \3043 , \3049 );
and \U$2736 ( \3051 , \3025 , \3049 );
or \U$2737 ( \3052 , \3044 , \3050 , \3051 );
xor \U$2738 ( \3053 , \2802 , \2845 );
xor \U$2739 ( \3054 , \3053 , \2855 );
xor \U$2740 ( \3055 , \2868 , \2870 );
xor \U$2741 ( \3056 , \3055 , \2873 );
and \U$2742 ( \3057 , \3054 , \3056 );
xor \U$2743 ( \3058 , \2879 , \2881 );
and \U$2744 ( \3059 , \3056 , \3058 );
and \U$2745 ( \3060 , \3054 , \3058 );
or \U$2746 ( \3061 , \3057 , \3059 , \3060 );
and \U$2747 ( \3062 , \3052 , \3061 );
xor \U$2748 ( \3063 , \2887 , \2889 );
xor \U$2749 ( \3064 , \3063 , \2892 );
and \U$2750 ( \3065 , \3061 , \3064 );
and \U$2751 ( \3066 , \3052 , \3064 );
or \U$2752 ( \3067 , \3062 , \3065 , \3066 );
xor \U$2753 ( \3068 , \2684 , \2702 );
xor \U$2754 ( \3069 , \3068 , \2712 );
and \U$2755 ( \3070 , \3067 , \3069 );
xor \U$2756 ( \3071 , \2885 , \2895 );
xor \U$2757 ( \3072 , \3071 , \2898 );
and \U$2758 ( \3073 , \3069 , \3072 );
and \U$2759 ( \3074 , \3067 , \3072 );
or \U$2760 ( \3075 , \3070 , \3073 , \3074 );
xor \U$2761 ( \3076 , \2901 , \2903 );
xor \U$2762 ( \3077 , \3076 , \2905 );
and \U$2763 ( \3078 , \3075 , \3077 );
and \U$2764 ( \3079 , \2914 , \3078 );
xor \U$2765 ( \3080 , \2914 , \3078 );
xor \U$2766 ( \3081 , \3075 , \3077 );
and \U$2767 ( \3082 , \425 , \2300 );
and \U$2768 ( \3083 , \417 , \2298 );
nor \U$2769 ( \3084 , \3082 , \3083 );
xnor \U$2770 ( \3085 , \3084 , \2163 );
and \U$2771 ( \3086 , \499 , \2094 );
and \U$2772 ( \3087 , \494 , \2092 );
nor \U$2773 ( \3088 , \3086 , \3087 );
xnor \U$2774 ( \3089 , \3088 , \1942 );
and \U$2775 ( \3090 , \3085 , \3089 );
and \U$2776 ( \3091 , \604 , \1826 );
and \U$2777 ( \3092 , \553 , \1824 );
nor \U$2778 ( \3093 , \3091 , \3092 );
xnor \U$2779 ( \3094 , \3093 , \1670 );
and \U$2780 ( \3095 , \3089 , \3094 );
and \U$2781 ( \3096 , \3085 , \3094 );
or \U$2782 ( \3097 , \3090 , \3095 , \3096 );
and \U$2783 ( \3098 , \709 , \1554 );
and \U$2784 ( \3099 , \681 , \1552 );
nor \U$2785 ( \3100 , \3098 , \3099 );
xnor \U$2786 ( \3101 , \3100 , \1441 );
and \U$2787 ( \3102 , \863 , \1360 );
and \U$2788 ( \3103 , \789 , \1358 );
nor \U$2789 ( \3104 , \3102 , \3103 );
xnor \U$2790 ( \3105 , \3104 , \1224 );
and \U$2791 ( \3106 , \3101 , \3105 );
and \U$2792 ( \3107 , \988 , \1160 );
and \U$2793 ( \3108 , \925 , \1158 );
nor \U$2794 ( \3109 , \3107 , \3108 );
xnor \U$2795 ( \3110 , \3109 , \1082 );
and \U$2796 ( \3111 , \3105 , \3110 );
and \U$2797 ( \3112 , \3101 , \3110 );
or \U$2798 ( \3113 , \3106 , \3111 , \3112 );
and \U$2799 ( \3114 , \3097 , \3113 );
buf \U$2800 ( \3115 , RIc0c87d8_35);
buf \U$2801 ( \3116 , RIc0c8760_36);
and \U$2802 ( \3117 , \3115 , \3116 );
not \U$2803 ( \3118 , \3117 );
and \U$2804 ( \3119 , \2766 , \3118 );
not \U$2805 ( \3120 , \3119 );
and \U$2806 ( \3121 , \330 , \2918 );
and \U$2807 ( \3122 , \316 , \2916 );
nor \U$2808 ( \3123 , \3121 , \3122 );
xnor \U$2809 ( \3124 , \3123 , \2769 );
and \U$2810 ( \3125 , \3120 , \3124 );
and \U$2811 ( \3126 , \369 , \2596 );
and \U$2812 ( \3127 , \348 , \2594 );
nor \U$2813 ( \3128 , \3126 , \3127 );
xnor \U$2814 ( \3129 , \3128 , \2454 );
and \U$2815 ( \3130 , \3124 , \3129 );
and \U$2816 ( \3131 , \3120 , \3129 );
or \U$2817 ( \3132 , \3125 , \3130 , \3131 );
and \U$2818 ( \3133 , \3113 , \3132 );
and \U$2819 ( \3134 , \3097 , \3132 );
or \U$2820 ( \3135 , \3114 , \3133 , \3134 );
and \U$2821 ( \3136 , \2666 , \360 );
and \U$2822 ( \3137 , \2641 , \358 );
nor \U$2823 ( \3138 , \3136 , \3137 );
xnor \U$2824 ( \3139 , \3138 , \341 );
and \U$2825 ( \3140 , \3007 , \323 );
and \U$2826 ( \3141 , \2840 , \321 );
nor \U$2827 ( \3142 , \3140 , \3141 );
xnor \U$2828 ( \3143 , \3142 , \328 );
and \U$2829 ( \3144 , \3139 , \3143 );
buf \U$2830 ( \3145 , RIc0c6a50_98);
and \U$2831 ( \3146 , \3145 , \317 );
and \U$2832 ( \3147 , \3143 , \3146 );
and \U$2833 ( \3148 , \3139 , \3146 );
or \U$2834 ( \3149 , \3144 , \3147 , \3148 );
and \U$2835 ( \3150 , \1799 , \579 );
and \U$2836 ( \3151 , \1791 , \577 );
nor \U$2837 ( \3152 , \3150 , \3151 );
xnor \U$2838 ( \3153 , \3152 , \530 );
and \U$2839 ( \3154 , \2047 , \478 );
and \U$2840 ( \3155 , \2042 , \476 );
nor \U$2841 ( \3156 , \3154 , \3155 );
xnor \U$2842 ( \3157 , \3156 , \437 );
and \U$2843 ( \3158 , \3153 , \3157 );
and \U$2844 ( \3159 , \2377 , \408 );
and \U$2845 ( \3160 , \2233 , \406 );
nor \U$2846 ( \3161 , \3159 , \3160 );
xnor \U$2847 ( \3162 , \3161 , \378 );
and \U$2848 ( \3163 , \3157 , \3162 );
and \U$2849 ( \3164 , \3153 , \3162 );
or \U$2850 ( \3165 , \3158 , \3163 , \3164 );
and \U$2851 ( \3166 , \3149 , \3165 );
and \U$2852 ( \3167 , \1274 , \996 );
and \U$2853 ( \3168 , \1186 , \994 );
nor \U$2854 ( \3169 , \3167 , \3168 );
xnor \U$2855 ( \3170 , \3169 , \902 );
and \U$2856 ( \3171 , \1384 , \826 );
and \U$2857 ( \3172 , \1379 , \824 );
nor \U$2858 ( \3173 , \3171 , \3172 );
xnor \U$2859 ( \3174 , \3173 , \754 );
and \U$2860 ( \3175 , \3170 , \3174 );
and \U$2861 ( \3176 , \1615 , \692 );
and \U$2862 ( \3177 , \1500 , \690 );
nor \U$2863 ( \3178 , \3176 , \3177 );
xnor \U$2864 ( \3179 , \3178 , \649 );
and \U$2865 ( \3180 , \3174 , \3179 );
and \U$2866 ( \3181 , \3170 , \3179 );
or \U$2867 ( \3182 , \3175 , \3180 , \3181 );
and \U$2868 ( \3183 , \3165 , \3182 );
and \U$2869 ( \3184 , \3149 , \3182 );
or \U$2870 ( \3185 , \3166 , \3183 , \3184 );
and \U$2871 ( \3186 , \3135 , \3185 );
xor \U$2872 ( \3187 , \2973 , \2977 );
xor \U$2873 ( \3188 , \3187 , \2982 );
xor \U$2874 ( \3189 , \2989 , \2993 );
xor \U$2875 ( \3190 , \3189 , \2998 );
and \U$2876 ( \3191 , \3188 , \3190 );
xnor \U$2877 ( \3192 , \3006 , \3008 );
and \U$2878 ( \3193 , \3190 , \3192 );
and \U$2879 ( \3194 , \3188 , \3192 );
or \U$2880 ( \3195 , \3191 , \3193 , \3194 );
and \U$2881 ( \3196 , \3185 , \3195 );
and \U$2882 ( \3197 , \3135 , \3195 );
or \U$2883 ( \3198 , \3186 , \3196 , \3197 );
xor \U$2884 ( \3199 , \2921 , \2925 );
xor \U$2885 ( \3200 , \3199 , \2930 );
xor \U$2886 ( \3201 , \2937 , \2941 );
xor \U$2887 ( \3202 , \3201 , \2946 );
and \U$2888 ( \3203 , \3200 , \3202 );
xor \U$2889 ( \3204 , \2954 , \2958 );
xor \U$2890 ( \3205 , \3204 , \2963 );
and \U$2891 ( \3206 , \3202 , \3205 );
and \U$2892 ( \3207 , \3200 , \3205 );
or \U$2893 ( \3208 , \3203 , \3206 , \3207 );
xor \U$2894 ( \3209 , \3027 , \3029 );
xor \U$2895 ( \3210 , \3209 , \3032 );
and \U$2896 ( \3211 , \3208 , \3210 );
xor \U$2897 ( \3212 , \3015 , \3017 );
xor \U$2898 ( \3213 , \3212 , \3019 );
and \U$2899 ( \3214 , \3210 , \3213 );
and \U$2900 ( \3215 , \3208 , \3213 );
or \U$2901 ( \3216 , \3211 , \3214 , \3215 );
and \U$2902 ( \3217 , \3198 , \3216 );
xor \U$2903 ( \3218 , \2933 , \2949 );
xor \U$2904 ( \3219 , \3218 , \2966 );
xor \U$2905 ( \3220 , \2985 , \3001 );
xor \U$2906 ( \3221 , \3220 , \3009 );
and \U$2907 ( \3222 , \3219 , \3221 );
and \U$2908 ( \3223 , \3216 , \3222 );
and \U$2909 ( \3224 , \3198 , \3222 );
or \U$2910 ( \3225 , \3217 , \3223 , \3224 );
xor \U$2911 ( \3226 , \2969 , \3012 );
xor \U$2912 ( \3227 , \3226 , \3022 );
xor \U$2913 ( \3228 , \3035 , \3037 );
xor \U$2914 ( \3229 , \3228 , \3040 );
and \U$2915 ( \3230 , \3227 , \3229 );
xor \U$2916 ( \3231 , \3046 , \3048 );
and \U$2917 ( \3232 , \3229 , \3231 );
and \U$2918 ( \3233 , \3227 , \3231 );
or \U$2919 ( \3234 , \3230 , \3232 , \3233 );
and \U$2920 ( \3235 , \3225 , \3234 );
xor \U$2921 ( \3236 , \3054 , \3056 );
xor \U$2922 ( \3237 , \3236 , \3058 );
and \U$2923 ( \3238 , \3234 , \3237 );
and \U$2924 ( \3239 , \3225 , \3237 );
or \U$2925 ( \3240 , \3235 , \3238 , \3239 );
xor \U$2926 ( \3241 , \2858 , \2876 );
xor \U$2927 ( \3242 , \3241 , \2882 );
and \U$2928 ( \3243 , \3240 , \3242 );
xor \U$2929 ( \3244 , \3052 , \3061 );
xor \U$2930 ( \3245 , \3244 , \3064 );
and \U$2931 ( \3246 , \3242 , \3245 );
and \U$2932 ( \3247 , \3240 , \3245 );
or \U$2933 ( \3248 , \3243 , \3246 , \3247 );
xor \U$2934 ( \3249 , \3067 , \3069 );
xor \U$2935 ( \3250 , \3249 , \3072 );
and \U$2936 ( \3251 , \3248 , \3250 );
and \U$2937 ( \3252 , \3081 , \3251 );
xor \U$2938 ( \3253 , \3081 , \3251 );
xor \U$2939 ( \3254 , \3248 , \3250 );
and \U$2940 ( \3255 , \2840 , \360 );
and \U$2941 ( \3256 , \2666 , \358 );
nor \U$2942 ( \3257 , \3255 , \3256 );
xnor \U$2943 ( \3258 , \3257 , \341 );
and \U$2944 ( \3259 , \3145 , \323 );
and \U$2945 ( \3260 , \3007 , \321 );
nor \U$2946 ( \3261 , \3259 , \3260 );
xnor \U$2947 ( \3262 , \3261 , \328 );
and \U$2948 ( \3263 , \3258 , \3262 );
buf \U$2949 ( \3264 , RIc0c69d8_99);
and \U$2950 ( \3265 , \3264 , \317 );
and \U$2951 ( \3266 , \3262 , \3265 );
and \U$2952 ( \3267 , \3258 , \3265 );
or \U$2953 ( \3268 , \3263 , \3266 , \3267 );
and \U$2954 ( \3269 , \2042 , \579 );
and \U$2955 ( \3270 , \1799 , \577 );
nor \U$2956 ( \3271 , \3269 , \3270 );
xnor \U$2957 ( \3272 , \3271 , \530 );
and \U$2958 ( \3273 , \2233 , \478 );
and \U$2959 ( \3274 , \2047 , \476 );
nor \U$2960 ( \3275 , \3273 , \3274 );
xnor \U$2961 ( \3276 , \3275 , \437 );
and \U$2962 ( \3277 , \3272 , \3276 );
and \U$2963 ( \3278 , \2641 , \408 );
and \U$2964 ( \3279 , \2377 , \406 );
nor \U$2965 ( \3280 , \3278 , \3279 );
xnor \U$2966 ( \3281 , \3280 , \378 );
and \U$2967 ( \3282 , \3276 , \3281 );
and \U$2968 ( \3283 , \3272 , \3281 );
or \U$2969 ( \3284 , \3277 , \3282 , \3283 );
and \U$2970 ( \3285 , \3268 , \3284 );
and \U$2971 ( \3286 , \1379 , \996 );
and \U$2972 ( \3287 , \1274 , \994 );
nor \U$2973 ( \3288 , \3286 , \3287 );
xnor \U$2974 ( \3289 , \3288 , \902 );
and \U$2975 ( \3290 , \1500 , \826 );
and \U$2976 ( \3291 , \1384 , \824 );
nor \U$2977 ( \3292 , \3290 , \3291 );
xnor \U$2978 ( \3293 , \3292 , \754 );
and \U$2979 ( \3294 , \3289 , \3293 );
and \U$2980 ( \3295 , \1791 , \692 );
and \U$2981 ( \3296 , \1615 , \690 );
nor \U$2982 ( \3297 , \3295 , \3296 );
xnor \U$2983 ( \3298 , \3297 , \649 );
and \U$2984 ( \3299 , \3293 , \3298 );
and \U$2985 ( \3300 , \3289 , \3298 );
or \U$2986 ( \3301 , \3294 , \3299 , \3300 );
and \U$2987 ( \3302 , \3284 , \3301 );
and \U$2988 ( \3303 , \3268 , \3301 );
or \U$2989 ( \3304 , \3285 , \3302 , \3303 );
and \U$2990 ( \3305 , \494 , \2300 );
and \U$2991 ( \3306 , \425 , \2298 );
nor \U$2992 ( \3307 , \3305 , \3306 );
xnor \U$2993 ( \3308 , \3307 , \2163 );
and \U$2994 ( \3309 , \553 , \2094 );
and \U$2995 ( \3310 , \499 , \2092 );
nor \U$2996 ( \3311 , \3309 , \3310 );
xnor \U$2997 ( \3312 , \3311 , \1942 );
and \U$2998 ( \3313 , \3308 , \3312 );
and \U$2999 ( \3314 , \681 , \1826 );
and \U$3000 ( \3315 , \604 , \1824 );
nor \U$3001 ( \3316 , \3314 , \3315 );
xnor \U$3002 ( \3317 , \3316 , \1670 );
and \U$3003 ( \3318 , \3312 , \3317 );
and \U$3004 ( \3319 , \3308 , \3317 );
or \U$3005 ( \3320 , \3313 , \3318 , \3319 );
xor \U$3006 ( \3321 , \2766 , \3115 );
xor \U$3007 ( \3322 , \3115 , \3116 );
not \U$3008 ( \3323 , \3322 );
and \U$3009 ( \3324 , \3321 , \3323 );
and \U$3010 ( \3325 , \316 , \3324 );
not \U$3011 ( \3326 , \3325 );
xnor \U$3012 ( \3327 , \3326 , \3119 );
and \U$3013 ( \3328 , \348 , \2918 );
and \U$3014 ( \3329 , \330 , \2916 );
nor \U$3015 ( \3330 , \3328 , \3329 );
xnor \U$3016 ( \3331 , \3330 , \2769 );
and \U$3017 ( \3332 , \3327 , \3331 );
and \U$3018 ( \3333 , \417 , \2596 );
and \U$3019 ( \3334 , \369 , \2594 );
nor \U$3020 ( \3335 , \3333 , \3334 );
xnor \U$3021 ( \3336 , \3335 , \2454 );
and \U$3022 ( \3337 , \3331 , \3336 );
and \U$3023 ( \3338 , \3327 , \3336 );
or \U$3024 ( \3339 , \3332 , \3337 , \3338 );
and \U$3025 ( \3340 , \3320 , \3339 );
and \U$3026 ( \3341 , \789 , \1554 );
and \U$3027 ( \3342 , \709 , \1552 );
nor \U$3028 ( \3343 , \3341 , \3342 );
xnor \U$3029 ( \3344 , \3343 , \1441 );
and \U$3030 ( \3345 , \925 , \1360 );
and \U$3031 ( \3346 , \863 , \1358 );
nor \U$3032 ( \3347 , \3345 , \3346 );
xnor \U$3033 ( \3348 , \3347 , \1224 );
and \U$3034 ( \3349 , \3344 , \3348 );
and \U$3035 ( \3350 , \1186 , \1160 );
and \U$3036 ( \3351 , \988 , \1158 );
nor \U$3037 ( \3352 , \3350 , \3351 );
xnor \U$3038 ( \3353 , \3352 , \1082 );
and \U$3039 ( \3354 , \3348 , \3353 );
and \U$3040 ( \3355 , \3344 , \3353 );
or \U$3041 ( \3356 , \3349 , \3354 , \3355 );
and \U$3042 ( \3357 , \3339 , \3356 );
and \U$3043 ( \3358 , \3320 , \3356 );
or \U$3044 ( \3359 , \3340 , \3357 , \3358 );
and \U$3045 ( \3360 , \3304 , \3359 );
xor \U$3046 ( \3361 , \3139 , \3143 );
xor \U$3047 ( \3362 , \3361 , \3146 );
xor \U$3048 ( \3363 , \3153 , \3157 );
xor \U$3049 ( \3364 , \3363 , \3162 );
and \U$3050 ( \3365 , \3362 , \3364 );
xor \U$3051 ( \3366 , \3170 , \3174 );
xor \U$3052 ( \3367 , \3366 , \3179 );
and \U$3053 ( \3368 , \3364 , \3367 );
and \U$3054 ( \3369 , \3362 , \3367 );
or \U$3055 ( \3370 , \3365 , \3368 , \3369 );
and \U$3056 ( \3371 , \3359 , \3370 );
and \U$3057 ( \3372 , \3304 , \3370 );
or \U$3058 ( \3373 , \3360 , \3371 , \3372 );
xor \U$3059 ( \3374 , \3085 , \3089 );
xor \U$3060 ( \3375 , \3374 , \3094 );
xor \U$3061 ( \3376 , \3101 , \3105 );
xor \U$3062 ( \3377 , \3376 , \3110 );
and \U$3063 ( \3378 , \3375 , \3377 );
xor \U$3064 ( \3379 , \3120 , \3124 );
xor \U$3065 ( \3380 , \3379 , \3129 );
and \U$3066 ( \3381 , \3377 , \3380 );
and \U$3067 ( \3382 , \3375 , \3380 );
or \U$3068 ( \3383 , \3378 , \3381 , \3382 );
xor \U$3069 ( \3384 , \3200 , \3202 );
xor \U$3070 ( \3385 , \3384 , \3205 );
and \U$3071 ( \3386 , \3383 , \3385 );
xor \U$3072 ( \3387 , \3188 , \3190 );
xor \U$3073 ( \3388 , \3387 , \3192 );
and \U$3074 ( \3389 , \3385 , \3388 );
and \U$3075 ( \3390 , \3383 , \3388 );
or \U$3076 ( \3391 , \3386 , \3389 , \3390 );
and \U$3077 ( \3392 , \3373 , \3391 );
xor \U$3078 ( \3393 , \3097 , \3113 );
xor \U$3079 ( \3394 , \3393 , \3132 );
xor \U$3080 ( \3395 , \3149 , \3165 );
xor \U$3081 ( \3396 , \3395 , \3182 );
and \U$3082 ( \3397 , \3394 , \3396 );
and \U$3083 ( \3398 , \3391 , \3397 );
and \U$3084 ( \3399 , \3373 , \3397 );
or \U$3085 ( \3400 , \3392 , \3398 , \3399 );
xor \U$3086 ( \3401 , \3135 , \3185 );
xor \U$3087 ( \3402 , \3401 , \3195 );
xor \U$3088 ( \3403 , \3208 , \3210 );
xor \U$3089 ( \3404 , \3403 , \3213 );
and \U$3090 ( \3405 , \3402 , \3404 );
xor \U$3091 ( \3406 , \3219 , \3221 );
and \U$3092 ( \3407 , \3404 , \3406 );
and \U$3093 ( \3408 , \3402 , \3406 );
or \U$3094 ( \3409 , \3405 , \3407 , \3408 );
and \U$3095 ( \3410 , \3400 , \3409 );
xor \U$3096 ( \3411 , \3227 , \3229 );
xor \U$3097 ( \3412 , \3411 , \3231 );
and \U$3098 ( \3413 , \3409 , \3412 );
and \U$3099 ( \3414 , \3400 , \3412 );
or \U$3100 ( \3415 , \3410 , \3413 , \3414 );
xor \U$3101 ( \3416 , \3025 , \3043 );
xor \U$3102 ( \3417 , \3416 , \3049 );
and \U$3103 ( \3418 , \3415 , \3417 );
xor \U$3104 ( \3419 , \3225 , \3234 );
xor \U$3105 ( \3420 , \3419 , \3237 );
and \U$3106 ( \3421 , \3417 , \3420 );
and \U$3107 ( \3422 , \3415 , \3420 );
or \U$3108 ( \3423 , \3418 , \3421 , \3422 );
xor \U$3109 ( \3424 , \3240 , \3242 );
xor \U$3110 ( \3425 , \3424 , \3245 );
and \U$3111 ( \3426 , \3423 , \3425 );
and \U$3112 ( \3427 , \3254 , \3426 );
xor \U$3113 ( \3428 , \3254 , \3426 );
xor \U$3114 ( \3429 , \3423 , \3425 );
and \U$3115 ( \3430 , \709 , \1826 );
and \U$3116 ( \3431 , \681 , \1824 );
nor \U$3117 ( \3432 , \3430 , \3431 );
xnor \U$3118 ( \3433 , \3432 , \1670 );
and \U$3119 ( \3434 , \863 , \1554 );
and \U$3120 ( \3435 , \789 , \1552 );
nor \U$3121 ( \3436 , \3434 , \3435 );
xnor \U$3122 ( \3437 , \3436 , \1441 );
and \U$3123 ( \3438 , \3433 , \3437 );
and \U$3124 ( \3439 , \988 , \1360 );
and \U$3125 ( \3440 , \925 , \1358 );
nor \U$3126 ( \3441 , \3439 , \3440 );
xnor \U$3127 ( \3442 , \3441 , \1224 );
and \U$3128 ( \3443 , \3437 , \3442 );
and \U$3129 ( \3444 , \3433 , \3442 );
or \U$3130 ( \3445 , \3438 , \3443 , \3444 );
buf \U$3131 ( \3446 , RIc0c86e8_37);
buf \U$3132 ( \3447 , RIc0c8670_38);
and \U$3133 ( \3448 , \3446 , \3447 );
not \U$3134 ( \3449 , \3448 );
and \U$3135 ( \3450 , \3116 , \3449 );
not \U$3136 ( \3451 , \3450 );
and \U$3137 ( \3452 , \330 , \3324 );
and \U$3138 ( \3453 , \316 , \3322 );
nor \U$3139 ( \3454 , \3452 , \3453 );
xnor \U$3140 ( \3455 , \3454 , \3119 );
and \U$3141 ( \3456 , \3451 , \3455 );
and \U$3142 ( \3457 , \369 , \2918 );
and \U$3143 ( \3458 , \348 , \2916 );
nor \U$3144 ( \3459 , \3457 , \3458 );
xnor \U$3145 ( \3460 , \3459 , \2769 );
and \U$3146 ( \3461 , \3455 , \3460 );
and \U$3147 ( \3462 , \3451 , \3460 );
or \U$3148 ( \3463 , \3456 , \3461 , \3462 );
and \U$3149 ( \3464 , \3445 , \3463 );
and \U$3150 ( \3465 , \425 , \2596 );
and \U$3151 ( \3466 , \417 , \2594 );
nor \U$3152 ( \3467 , \3465 , \3466 );
xnor \U$3153 ( \3468 , \3467 , \2454 );
and \U$3154 ( \3469 , \499 , \2300 );
and \U$3155 ( \3470 , \494 , \2298 );
nor \U$3156 ( \3471 , \3469 , \3470 );
xnor \U$3157 ( \3472 , \3471 , \2163 );
and \U$3158 ( \3473 , \3468 , \3472 );
and \U$3159 ( \3474 , \604 , \2094 );
and \U$3160 ( \3475 , \553 , \2092 );
nor \U$3161 ( \3476 , \3474 , \3475 );
xnor \U$3162 ( \3477 , \3476 , \1942 );
and \U$3163 ( \3478 , \3472 , \3477 );
and \U$3164 ( \3479 , \3468 , \3477 );
or \U$3165 ( \3480 , \3473 , \3478 , \3479 );
and \U$3166 ( \3481 , \3463 , \3480 );
and \U$3167 ( \3482 , \3445 , \3480 );
or \U$3168 ( \3483 , \3464 , \3481 , \3482 );
and \U$3169 ( \3484 , \2666 , \408 );
and \U$3170 ( \3485 , \2641 , \406 );
nor \U$3171 ( \3486 , \3484 , \3485 );
xnor \U$3172 ( \3487 , \3486 , \378 );
and \U$3173 ( \3488 , \3007 , \360 );
and \U$3174 ( \3489 , \2840 , \358 );
nor \U$3175 ( \3490 , \3488 , \3489 );
xnor \U$3176 ( \3491 , \3490 , \341 );
and \U$3177 ( \3492 , \3487 , \3491 );
and \U$3178 ( \3493 , \3264 , \323 );
and \U$3179 ( \3494 , \3145 , \321 );
nor \U$3180 ( \3495 , \3493 , \3494 );
xnor \U$3181 ( \3496 , \3495 , \328 );
and \U$3182 ( \3497 , \3491 , \3496 );
and \U$3183 ( \3498 , \3487 , \3496 );
or \U$3184 ( \3499 , \3492 , \3497 , \3498 );
and \U$3185 ( \3500 , \1274 , \1160 );
and \U$3186 ( \3501 , \1186 , \1158 );
nor \U$3187 ( \3502 , \3500 , \3501 );
xnor \U$3188 ( \3503 , \3502 , \1082 );
and \U$3189 ( \3504 , \1384 , \996 );
and \U$3190 ( \3505 , \1379 , \994 );
nor \U$3191 ( \3506 , \3504 , \3505 );
xnor \U$3192 ( \3507 , \3506 , \902 );
and \U$3193 ( \3508 , \3503 , \3507 );
and \U$3194 ( \3509 , \1615 , \826 );
and \U$3195 ( \3510 , \1500 , \824 );
nor \U$3196 ( \3511 , \3509 , \3510 );
xnor \U$3197 ( \3512 , \3511 , \754 );
and \U$3198 ( \3513 , \3507 , \3512 );
and \U$3199 ( \3514 , \3503 , \3512 );
or \U$3200 ( \3515 , \3508 , \3513 , \3514 );
and \U$3201 ( \3516 , \3499 , \3515 );
and \U$3202 ( \3517 , \1799 , \692 );
and \U$3203 ( \3518 , \1791 , \690 );
nor \U$3204 ( \3519 , \3517 , \3518 );
xnor \U$3205 ( \3520 , \3519 , \649 );
and \U$3206 ( \3521 , \2047 , \579 );
and \U$3207 ( \3522 , \2042 , \577 );
nor \U$3208 ( \3523 , \3521 , \3522 );
xnor \U$3209 ( \3524 , \3523 , \530 );
and \U$3210 ( \3525 , \3520 , \3524 );
and \U$3211 ( \3526 , \2377 , \478 );
and \U$3212 ( \3527 , \2233 , \476 );
nor \U$3213 ( \3528 , \3526 , \3527 );
xnor \U$3214 ( \3529 , \3528 , \437 );
and \U$3215 ( \3530 , \3524 , \3529 );
and \U$3216 ( \3531 , \3520 , \3529 );
or \U$3217 ( \3532 , \3525 , \3530 , \3531 );
and \U$3218 ( \3533 , \3515 , \3532 );
and \U$3219 ( \3534 , \3499 , \3532 );
or \U$3220 ( \3535 , \3516 , \3533 , \3534 );
and \U$3221 ( \3536 , \3483 , \3535 );
xor \U$3222 ( \3537 , \3258 , \3262 );
xor \U$3223 ( \3538 , \3537 , \3265 );
xor \U$3224 ( \3539 , \3272 , \3276 );
xor \U$3225 ( \3540 , \3539 , \3281 );
or \U$3226 ( \3541 , \3538 , \3540 );
and \U$3227 ( \3542 , \3535 , \3541 );
and \U$3228 ( \3543 , \3483 , \3541 );
or \U$3229 ( \3544 , \3536 , \3542 , \3543 );
xor \U$3230 ( \3545 , \3308 , \3312 );
xor \U$3231 ( \3546 , \3545 , \3317 );
xor \U$3232 ( \3547 , \3344 , \3348 );
xor \U$3233 ( \3548 , \3547 , \3353 );
and \U$3234 ( \3549 , \3546 , \3548 );
xor \U$3235 ( \3550 , \3289 , \3293 );
xor \U$3236 ( \3551 , \3550 , \3298 );
and \U$3237 ( \3552 , \3548 , \3551 );
and \U$3238 ( \3553 , \3546 , \3551 );
or \U$3239 ( \3554 , \3549 , \3552 , \3553 );
xor \U$3240 ( \3555 , \3362 , \3364 );
xor \U$3241 ( \3556 , \3555 , \3367 );
and \U$3242 ( \3557 , \3554 , \3556 );
xor \U$3243 ( \3558 , \3375 , \3377 );
xor \U$3244 ( \3559 , \3558 , \3380 );
and \U$3245 ( \3560 , \3556 , \3559 );
and \U$3246 ( \3561 , \3554 , \3559 );
or \U$3247 ( \3562 , \3557 , \3560 , \3561 );
and \U$3248 ( \3563 , \3544 , \3562 );
xor \U$3249 ( \3564 , \3268 , \3284 );
xor \U$3250 ( \3565 , \3564 , \3301 );
xor \U$3251 ( \3566 , \3320 , \3339 );
xor \U$3252 ( \3567 , \3566 , \3356 );
and \U$3253 ( \3568 , \3565 , \3567 );
and \U$3254 ( \3569 , \3562 , \3568 );
and \U$3255 ( \3570 , \3544 , \3568 );
or \U$3256 ( \3571 , \3563 , \3569 , \3570 );
xor \U$3257 ( \3572 , \3304 , \3359 );
xor \U$3258 ( \3573 , \3572 , \3370 );
xor \U$3259 ( \3574 , \3383 , \3385 );
xor \U$3260 ( \3575 , \3574 , \3388 );
and \U$3261 ( \3576 , \3573 , \3575 );
xor \U$3262 ( \3577 , \3394 , \3396 );
and \U$3263 ( \3578 , \3575 , \3577 );
and \U$3264 ( \3579 , \3573 , \3577 );
or \U$3265 ( \3580 , \3576 , \3578 , \3579 );
and \U$3266 ( \3581 , \3571 , \3580 );
xor \U$3267 ( \3582 , \3402 , \3404 );
xor \U$3268 ( \3583 , \3582 , \3406 );
and \U$3269 ( \3584 , \3580 , \3583 );
and \U$3270 ( \3585 , \3571 , \3583 );
or \U$3271 ( \3586 , \3581 , \3584 , \3585 );
xor \U$3272 ( \3587 , \3198 , \3216 );
xor \U$3273 ( \3588 , \3587 , \3222 );
and \U$3274 ( \3589 , \3586 , \3588 );
xor \U$3275 ( \3590 , \3400 , \3409 );
xor \U$3276 ( \3591 , \3590 , \3412 );
and \U$3277 ( \3592 , \3588 , \3591 );
and \U$3278 ( \3593 , \3586 , \3591 );
or \U$3279 ( \3594 , \3589 , \3592 , \3593 );
xor \U$3280 ( \3595 , \3415 , \3417 );
xor \U$3281 ( \3596 , \3595 , \3420 );
and \U$3282 ( \3597 , \3594 , \3596 );
and \U$3283 ( \3598 , \3429 , \3597 );
xor \U$3284 ( \3599 , \3429 , \3597 );
xor \U$3285 ( \3600 , \3594 , \3596 );
and \U$3286 ( \3601 , \789 , \1826 );
and \U$3287 ( \3602 , \709 , \1824 );
nor \U$3288 ( \3603 , \3601 , \3602 );
xnor \U$3289 ( \3604 , \3603 , \1670 );
and \U$3290 ( \3605 , \925 , \1554 );
and \U$3291 ( \3606 , \863 , \1552 );
nor \U$3292 ( \3607 , \3605 , \3606 );
xnor \U$3293 ( \3608 , \3607 , \1441 );
and \U$3294 ( \3609 , \3604 , \3608 );
and \U$3295 ( \3610 , \1186 , \1360 );
and \U$3296 ( \3611 , \988 , \1358 );
nor \U$3297 ( \3612 , \3610 , \3611 );
xnor \U$3298 ( \3613 , \3612 , \1224 );
and \U$3299 ( \3614 , \3608 , \3613 );
and \U$3300 ( \3615 , \3604 , \3613 );
or \U$3301 ( \3616 , \3609 , \3614 , \3615 );
and \U$3302 ( \3617 , \494 , \2596 );
and \U$3303 ( \3618 , \425 , \2594 );
nor \U$3304 ( \3619 , \3617 , \3618 );
xnor \U$3305 ( \3620 , \3619 , \2454 );
and \U$3306 ( \3621 , \553 , \2300 );
and \U$3307 ( \3622 , \499 , \2298 );
nor \U$3308 ( \3623 , \3621 , \3622 );
xnor \U$3309 ( \3624 , \3623 , \2163 );
and \U$3310 ( \3625 , \3620 , \3624 );
and \U$3311 ( \3626 , \681 , \2094 );
and \U$3312 ( \3627 , \604 , \2092 );
nor \U$3313 ( \3628 , \3626 , \3627 );
xnor \U$3314 ( \3629 , \3628 , \1942 );
and \U$3315 ( \3630 , \3624 , \3629 );
and \U$3316 ( \3631 , \3620 , \3629 );
or \U$3317 ( \3632 , \3625 , \3630 , \3631 );
and \U$3318 ( \3633 , \3616 , \3632 );
xor \U$3319 ( \3634 , \3116 , \3446 );
xor \U$3320 ( \3635 , \3446 , \3447 );
not \U$3321 ( \3636 , \3635 );
and \U$3322 ( \3637 , \3634 , \3636 );
and \U$3323 ( \3638 , \316 , \3637 );
not \U$3324 ( \3639 , \3638 );
xnor \U$3325 ( \3640 , \3639 , \3450 );
and \U$3326 ( \3641 , \348 , \3324 );
and \U$3327 ( \3642 , \330 , \3322 );
nor \U$3328 ( \3643 , \3641 , \3642 );
xnor \U$3329 ( \3644 , \3643 , \3119 );
and \U$3330 ( \3645 , \3640 , \3644 );
and \U$3331 ( \3646 , \417 , \2918 );
and \U$3332 ( \3647 , \369 , \2916 );
nor \U$3333 ( \3648 , \3646 , \3647 );
xnor \U$3334 ( \3649 , \3648 , \2769 );
and \U$3335 ( \3650 , \3644 , \3649 );
and \U$3336 ( \3651 , \3640 , \3649 );
or \U$3337 ( \3652 , \3645 , \3650 , \3651 );
and \U$3338 ( \3653 , \3632 , \3652 );
and \U$3339 ( \3654 , \3616 , \3652 );
or \U$3340 ( \3655 , \3633 , \3653 , \3654 );
and \U$3341 ( \3656 , \1379 , \1160 );
and \U$3342 ( \3657 , \1274 , \1158 );
nor \U$3343 ( \3658 , \3656 , \3657 );
xnor \U$3344 ( \3659 , \3658 , \1082 );
and \U$3345 ( \3660 , \1500 , \996 );
and \U$3346 ( \3661 , \1384 , \994 );
nor \U$3347 ( \3662 , \3660 , \3661 );
xnor \U$3348 ( \3663 , \3662 , \902 );
and \U$3349 ( \3664 , \3659 , \3663 );
and \U$3350 ( \3665 , \1791 , \826 );
and \U$3351 ( \3666 , \1615 , \824 );
nor \U$3352 ( \3667 , \3665 , \3666 );
xnor \U$3353 ( \3668 , \3667 , \754 );
and \U$3354 ( \3669 , \3663 , \3668 );
and \U$3355 ( \3670 , \3659 , \3668 );
or \U$3356 ( \3671 , \3664 , \3669 , \3670 );
and \U$3357 ( \3672 , \2840 , \408 );
and \U$3358 ( \3673 , \2666 , \406 );
nor \U$3359 ( \3674 , \3672 , \3673 );
xnor \U$3360 ( \3675 , \3674 , \378 );
and \U$3361 ( \3676 , \3145 , \360 );
and \U$3362 ( \3677 , \3007 , \358 );
nor \U$3363 ( \3678 , \3676 , \3677 );
xnor \U$3364 ( \3679 , \3678 , \341 );
and \U$3365 ( \3680 , \3675 , \3679 );
buf \U$3366 ( \3681 , RIc0c6960_100);
and \U$3367 ( \3682 , \3681 , \323 );
and \U$3368 ( \3683 , \3264 , \321 );
nor \U$3369 ( \3684 , \3682 , \3683 );
xnor \U$3370 ( \3685 , \3684 , \328 );
and \U$3371 ( \3686 , \3679 , \3685 );
and \U$3372 ( \3687 , \3675 , \3685 );
or \U$3373 ( \3688 , \3680 , \3686 , \3687 );
and \U$3374 ( \3689 , \3671 , \3688 );
and \U$3375 ( \3690 , \2042 , \692 );
and \U$3376 ( \3691 , \1799 , \690 );
nor \U$3377 ( \3692 , \3690 , \3691 );
xnor \U$3378 ( \3693 , \3692 , \649 );
and \U$3379 ( \3694 , \2233 , \579 );
and \U$3380 ( \3695 , \2047 , \577 );
nor \U$3381 ( \3696 , \3694 , \3695 );
xnor \U$3382 ( \3697 , \3696 , \530 );
and \U$3383 ( \3698 , \3693 , \3697 );
and \U$3384 ( \3699 , \2641 , \478 );
and \U$3385 ( \3700 , \2377 , \476 );
nor \U$3386 ( \3701 , \3699 , \3700 );
xnor \U$3387 ( \3702 , \3701 , \437 );
and \U$3388 ( \3703 , \3697 , \3702 );
and \U$3389 ( \3704 , \3693 , \3702 );
or \U$3390 ( \3705 , \3698 , \3703 , \3704 );
and \U$3391 ( \3706 , \3688 , \3705 );
and \U$3392 ( \3707 , \3671 , \3705 );
or \U$3393 ( \3708 , \3689 , \3706 , \3707 );
and \U$3394 ( \3709 , \3655 , \3708 );
and \U$3395 ( \3710 , \3681 , \317 );
xor \U$3396 ( \3711 , \3487 , \3491 );
xor \U$3397 ( \3712 , \3711 , \3496 );
and \U$3398 ( \3713 , \3710 , \3712 );
xor \U$3399 ( \3714 , \3520 , \3524 );
xor \U$3400 ( \3715 , \3714 , \3529 );
and \U$3401 ( \3716 , \3712 , \3715 );
and \U$3402 ( \3717 , \3710 , \3715 );
or \U$3403 ( \3718 , \3713 , \3716 , \3717 );
and \U$3404 ( \3719 , \3708 , \3718 );
and \U$3405 ( \3720 , \3655 , \3718 );
or \U$3406 ( \3721 , \3709 , \3719 , \3720 );
xor \U$3407 ( \3722 , \3433 , \3437 );
xor \U$3408 ( \3723 , \3722 , \3442 );
xor \U$3409 ( \3724 , \3503 , \3507 );
xor \U$3410 ( \3725 , \3724 , \3512 );
and \U$3411 ( \3726 , \3723 , \3725 );
xor \U$3412 ( \3727 , \3468 , \3472 );
xor \U$3413 ( \3728 , \3727 , \3477 );
and \U$3414 ( \3729 , \3725 , \3728 );
and \U$3415 ( \3730 , \3723 , \3728 );
or \U$3416 ( \3731 , \3726 , \3729 , \3730 );
xor \U$3417 ( \3732 , \3327 , \3331 );
xor \U$3418 ( \3733 , \3732 , \3336 );
and \U$3419 ( \3734 , \3731 , \3733 );
xor \U$3420 ( \3735 , \3546 , \3548 );
xor \U$3421 ( \3736 , \3735 , \3551 );
and \U$3422 ( \3737 , \3733 , \3736 );
and \U$3423 ( \3738 , \3731 , \3736 );
or \U$3424 ( \3739 , \3734 , \3737 , \3738 );
and \U$3425 ( \3740 , \3721 , \3739 );
xor \U$3426 ( \3741 , \3445 , \3463 );
xor \U$3427 ( \3742 , \3741 , \3480 );
xor \U$3428 ( \3743 , \3499 , \3515 );
xor \U$3429 ( \3744 , \3743 , \3532 );
and \U$3430 ( \3745 , \3742 , \3744 );
xnor \U$3431 ( \3746 , \3538 , \3540 );
and \U$3432 ( \3747 , \3744 , \3746 );
and \U$3433 ( \3748 , \3742 , \3746 );
or \U$3434 ( \3749 , \3745 , \3747 , \3748 );
and \U$3435 ( \3750 , \3739 , \3749 );
and \U$3436 ( \3751 , \3721 , \3749 );
or \U$3437 ( \3752 , \3740 , \3750 , \3751 );
xor \U$3438 ( \3753 , \3483 , \3535 );
xor \U$3439 ( \3754 , \3753 , \3541 );
xor \U$3440 ( \3755 , \3554 , \3556 );
xor \U$3441 ( \3756 , \3755 , \3559 );
and \U$3442 ( \3757 , \3754 , \3756 );
xor \U$3443 ( \3758 , \3565 , \3567 );
and \U$3444 ( \3759 , \3756 , \3758 );
and \U$3445 ( \3760 , \3754 , \3758 );
or \U$3446 ( \3761 , \3757 , \3759 , \3760 );
and \U$3447 ( \3762 , \3752 , \3761 );
xor \U$3448 ( \3763 , \3573 , \3575 );
xor \U$3449 ( \3764 , \3763 , \3577 );
and \U$3450 ( \3765 , \3761 , \3764 );
and \U$3451 ( \3766 , \3752 , \3764 );
or \U$3452 ( \3767 , \3762 , \3765 , \3766 );
xor \U$3453 ( \3768 , \3373 , \3391 );
xor \U$3454 ( \3769 , \3768 , \3397 );
and \U$3455 ( \3770 , \3767 , \3769 );
xor \U$3456 ( \3771 , \3571 , \3580 );
xor \U$3457 ( \3772 , \3771 , \3583 );
and \U$3458 ( \3773 , \3769 , \3772 );
and \U$3459 ( \3774 , \3767 , \3772 );
or \U$3460 ( \3775 , \3770 , \3773 , \3774 );
xor \U$3461 ( \3776 , \3586 , \3588 );
xor \U$3462 ( \3777 , \3776 , \3591 );
and \U$3463 ( \3778 , \3775 , \3777 );
and \U$3464 ( \3779 , \3600 , \3778 );
xor \U$3465 ( \3780 , \3600 , \3778 );
xor \U$3466 ( \3781 , \3775 , \3777 );
buf \U$3467 ( \3782 , RIc0c85f8_39);
buf \U$3468 ( \3783 , RIc0c8580_40);
and \U$3469 ( \3784 , \3782 , \3783 );
not \U$3470 ( \3785 , \3784 );
and \U$3471 ( \3786 , \3447 , \3785 );
not \U$3472 ( \3787 , \3786 );
and \U$3473 ( \3788 , \330 , \3637 );
and \U$3474 ( \3789 , \316 , \3635 );
nor \U$3475 ( \3790 , \3788 , \3789 );
xnor \U$3476 ( \3791 , \3790 , \3450 );
and \U$3477 ( \3792 , \3787 , \3791 );
and \U$3478 ( \3793 , \369 , \3324 );
and \U$3479 ( \3794 , \348 , \3322 );
nor \U$3480 ( \3795 , \3793 , \3794 );
xnor \U$3481 ( \3796 , \3795 , \3119 );
and \U$3482 ( \3797 , \3791 , \3796 );
and \U$3483 ( \3798 , \3787 , \3796 );
or \U$3484 ( \3799 , \3792 , \3797 , \3798 );
and \U$3485 ( \3800 , \425 , \2918 );
and \U$3486 ( \3801 , \417 , \2916 );
nor \U$3487 ( \3802 , \3800 , \3801 );
xnor \U$3488 ( \3803 , \3802 , \2769 );
and \U$3489 ( \3804 , \499 , \2596 );
and \U$3490 ( \3805 , \494 , \2594 );
nor \U$3491 ( \3806 , \3804 , \3805 );
xnor \U$3492 ( \3807 , \3806 , \2454 );
and \U$3493 ( \3808 , \3803 , \3807 );
and \U$3494 ( \3809 , \604 , \2300 );
and \U$3495 ( \3810 , \553 , \2298 );
nor \U$3496 ( \3811 , \3809 , \3810 );
xnor \U$3497 ( \3812 , \3811 , \2163 );
and \U$3498 ( \3813 , \3807 , \3812 );
and \U$3499 ( \3814 , \3803 , \3812 );
or \U$3500 ( \3815 , \3808 , \3813 , \3814 );
and \U$3501 ( \3816 , \3799 , \3815 );
and \U$3502 ( \3817 , \709 , \2094 );
and \U$3503 ( \3818 , \681 , \2092 );
nor \U$3504 ( \3819 , \3817 , \3818 );
xnor \U$3505 ( \3820 , \3819 , \1942 );
and \U$3506 ( \3821 , \863 , \1826 );
and \U$3507 ( \3822 , \789 , \1824 );
nor \U$3508 ( \3823 , \3821 , \3822 );
xnor \U$3509 ( \3824 , \3823 , \1670 );
and \U$3510 ( \3825 , \3820 , \3824 );
and \U$3511 ( \3826 , \988 , \1554 );
and \U$3512 ( \3827 , \925 , \1552 );
nor \U$3513 ( \3828 , \3826 , \3827 );
xnor \U$3514 ( \3829 , \3828 , \1441 );
and \U$3515 ( \3830 , \3824 , \3829 );
and \U$3516 ( \3831 , \3820 , \3829 );
or \U$3517 ( \3832 , \3825 , \3830 , \3831 );
and \U$3518 ( \3833 , \3815 , \3832 );
and \U$3519 ( \3834 , \3799 , \3832 );
or \U$3520 ( \3835 , \3816 , \3833 , \3834 );
and \U$3521 ( \3836 , \1799 , \826 );
and \U$3522 ( \3837 , \1791 , \824 );
nor \U$3523 ( \3838 , \3836 , \3837 );
xnor \U$3524 ( \3839 , \3838 , \754 );
and \U$3525 ( \3840 , \2047 , \692 );
and \U$3526 ( \3841 , \2042 , \690 );
nor \U$3527 ( \3842 , \3840 , \3841 );
xnor \U$3528 ( \3843 , \3842 , \649 );
and \U$3529 ( \3844 , \3839 , \3843 );
and \U$3530 ( \3845 , \2377 , \579 );
and \U$3531 ( \3846 , \2233 , \577 );
nor \U$3532 ( \3847 , \3845 , \3846 );
xnor \U$3533 ( \3848 , \3847 , \530 );
and \U$3534 ( \3849 , \3843 , \3848 );
and \U$3535 ( \3850 , \3839 , \3848 );
or \U$3536 ( \3851 , \3844 , \3849 , \3850 );
and \U$3537 ( \3852 , \1274 , \1360 );
and \U$3538 ( \3853 , \1186 , \1358 );
nor \U$3539 ( \3854 , \3852 , \3853 );
xnor \U$3540 ( \3855 , \3854 , \1224 );
and \U$3541 ( \3856 , \1384 , \1160 );
and \U$3542 ( \3857 , \1379 , \1158 );
nor \U$3543 ( \3858 , \3856 , \3857 );
xnor \U$3544 ( \3859 , \3858 , \1082 );
and \U$3545 ( \3860 , \3855 , \3859 );
and \U$3546 ( \3861 , \1615 , \996 );
and \U$3547 ( \3862 , \1500 , \994 );
nor \U$3548 ( \3863 , \3861 , \3862 );
xnor \U$3549 ( \3864 , \3863 , \902 );
and \U$3550 ( \3865 , \3859 , \3864 );
and \U$3551 ( \3866 , \3855 , \3864 );
or \U$3552 ( \3867 , \3860 , \3865 , \3866 );
and \U$3553 ( \3868 , \3851 , \3867 );
and \U$3554 ( \3869 , \2666 , \478 );
and \U$3555 ( \3870 , \2641 , \476 );
nor \U$3556 ( \3871 , \3869 , \3870 );
xnor \U$3557 ( \3872 , \3871 , \437 );
and \U$3558 ( \3873 , \3007 , \408 );
and \U$3559 ( \3874 , \2840 , \406 );
nor \U$3560 ( \3875 , \3873 , \3874 );
xnor \U$3561 ( \3876 , \3875 , \378 );
and \U$3562 ( \3877 , \3872 , \3876 );
and \U$3563 ( \3878 , \3264 , \360 );
and \U$3564 ( \3879 , \3145 , \358 );
nor \U$3565 ( \3880 , \3878 , \3879 );
xnor \U$3566 ( \3881 , \3880 , \341 );
and \U$3567 ( \3882 , \3876 , \3881 );
and \U$3568 ( \3883 , \3872 , \3881 );
or \U$3569 ( \3884 , \3877 , \3882 , \3883 );
and \U$3570 ( \3885 , \3867 , \3884 );
and \U$3571 ( \3886 , \3851 , \3884 );
or \U$3572 ( \3887 , \3868 , \3885 , \3886 );
and \U$3573 ( \3888 , \3835 , \3887 );
buf \U$3574 ( \3889 , RIc0c68e8_101);
and \U$3575 ( \3890 , \3889 , \317 );
xor \U$3576 ( \3891 , \3675 , \3679 );
xor \U$3577 ( \3892 , \3891 , \3685 );
or \U$3578 ( \3893 , \3890 , \3892 );
and \U$3579 ( \3894 , \3887 , \3893 );
and \U$3580 ( \3895 , \3835 , \3893 );
or \U$3581 ( \3896 , \3888 , \3894 , \3895 );
xor \U$3582 ( \3897 , \3604 , \3608 );
xor \U$3583 ( \3898 , \3897 , \3613 );
xor \U$3584 ( \3899 , \3659 , \3663 );
xor \U$3585 ( \3900 , \3899 , \3668 );
and \U$3586 ( \3901 , \3898 , \3900 );
xor \U$3587 ( \3902 , \3693 , \3697 );
xor \U$3588 ( \3903 , \3902 , \3702 );
and \U$3589 ( \3904 , \3900 , \3903 );
and \U$3590 ( \3905 , \3898 , \3903 );
or \U$3591 ( \3906 , \3901 , \3904 , \3905 );
xor \U$3592 ( \3907 , \3451 , \3455 );
xor \U$3593 ( \3908 , \3907 , \3460 );
and \U$3594 ( \3909 , \3906 , \3908 );
xor \U$3595 ( \3910 , \3723 , \3725 );
xor \U$3596 ( \3911 , \3910 , \3728 );
and \U$3597 ( \3912 , \3908 , \3911 );
and \U$3598 ( \3913 , \3906 , \3911 );
or \U$3599 ( \3914 , \3909 , \3912 , \3913 );
and \U$3600 ( \3915 , \3896 , \3914 );
xor \U$3601 ( \3916 , \3616 , \3632 );
xor \U$3602 ( \3917 , \3916 , \3652 );
xor \U$3603 ( \3918 , \3671 , \3688 );
xor \U$3604 ( \3919 , \3918 , \3705 );
and \U$3605 ( \3920 , \3917 , \3919 );
xor \U$3606 ( \3921 , \3710 , \3712 );
xor \U$3607 ( \3922 , \3921 , \3715 );
and \U$3608 ( \3923 , \3919 , \3922 );
and \U$3609 ( \3924 , \3917 , \3922 );
or \U$3610 ( \3925 , \3920 , \3923 , \3924 );
and \U$3611 ( \3926 , \3914 , \3925 );
and \U$3612 ( \3927 , \3896 , \3925 );
or \U$3613 ( \3928 , \3915 , \3926 , \3927 );
xor \U$3614 ( \3929 , \3655 , \3708 );
xor \U$3615 ( \3930 , \3929 , \3718 );
xor \U$3616 ( \3931 , \3731 , \3733 );
xor \U$3617 ( \3932 , \3931 , \3736 );
and \U$3618 ( \3933 , \3930 , \3932 );
xor \U$3619 ( \3934 , \3742 , \3744 );
xor \U$3620 ( \3935 , \3934 , \3746 );
and \U$3621 ( \3936 , \3932 , \3935 );
and \U$3622 ( \3937 , \3930 , \3935 );
or \U$3623 ( \3938 , \3933 , \3936 , \3937 );
and \U$3624 ( \3939 , \3928 , \3938 );
xor \U$3625 ( \3940 , \3754 , \3756 );
xor \U$3626 ( \3941 , \3940 , \3758 );
and \U$3627 ( \3942 , \3938 , \3941 );
and \U$3628 ( \3943 , \3928 , \3941 );
or \U$3629 ( \3944 , \3939 , \3942 , \3943 );
xor \U$3630 ( \3945 , \3544 , \3562 );
xor \U$3631 ( \3946 , \3945 , \3568 );
and \U$3632 ( \3947 , \3944 , \3946 );
xor \U$3633 ( \3948 , \3752 , \3761 );
xor \U$3634 ( \3949 , \3948 , \3764 );
and \U$3635 ( \3950 , \3946 , \3949 );
and \U$3636 ( \3951 , \3944 , \3949 );
or \U$3637 ( \3952 , \3947 , \3950 , \3951 );
xor \U$3638 ( \3953 , \3767 , \3769 );
xor \U$3639 ( \3954 , \3953 , \3772 );
and \U$3640 ( \3955 , \3952 , \3954 );
and \U$3641 ( \3956 , \3781 , \3955 );
xor \U$3642 ( \3957 , \3781 , \3955 );
xor \U$3643 ( \3958 , \3952 , \3954 );
and \U$3644 ( \3959 , \1379 , \1360 );
and \U$3645 ( \3960 , \1274 , \1358 );
nor \U$3646 ( \3961 , \3959 , \3960 );
xnor \U$3647 ( \3962 , \3961 , \1224 );
and \U$3648 ( \3963 , \1500 , \1160 );
and \U$3649 ( \3964 , \1384 , \1158 );
nor \U$3650 ( \3965 , \3963 , \3964 );
xnor \U$3651 ( \3966 , \3965 , \1082 );
and \U$3652 ( \3967 , \3962 , \3966 );
and \U$3653 ( \3968 , \1791 , \996 );
and \U$3654 ( \3969 , \1615 , \994 );
nor \U$3655 ( \3970 , \3968 , \3969 );
xnor \U$3656 ( \3971 , \3970 , \902 );
and \U$3657 ( \3972 , \3966 , \3971 );
and \U$3658 ( \3973 , \3962 , \3971 );
or \U$3659 ( \3974 , \3967 , \3972 , \3973 );
and \U$3660 ( \3975 , \2042 , \826 );
and \U$3661 ( \3976 , \1799 , \824 );
nor \U$3662 ( \3977 , \3975 , \3976 );
xnor \U$3663 ( \3978 , \3977 , \754 );
and \U$3664 ( \3979 , \2233 , \692 );
and \U$3665 ( \3980 , \2047 , \690 );
nor \U$3666 ( \3981 , \3979 , \3980 );
xnor \U$3667 ( \3982 , \3981 , \649 );
and \U$3668 ( \3983 , \3978 , \3982 );
and \U$3669 ( \3984 , \2641 , \579 );
and \U$3670 ( \3985 , \2377 , \577 );
nor \U$3671 ( \3986 , \3984 , \3985 );
xnor \U$3672 ( \3987 , \3986 , \530 );
and \U$3673 ( \3988 , \3982 , \3987 );
and \U$3674 ( \3989 , \3978 , \3987 );
or \U$3675 ( \3990 , \3983 , \3988 , \3989 );
and \U$3676 ( \3991 , \3974 , \3990 );
and \U$3677 ( \3992 , \2840 , \478 );
and \U$3678 ( \3993 , \2666 , \476 );
nor \U$3679 ( \3994 , \3992 , \3993 );
xnor \U$3680 ( \3995 , \3994 , \437 );
and \U$3681 ( \3996 , \3145 , \408 );
and \U$3682 ( \3997 , \3007 , \406 );
nor \U$3683 ( \3998 , \3996 , \3997 );
xnor \U$3684 ( \3999 , \3998 , \378 );
and \U$3685 ( \4000 , \3995 , \3999 );
and \U$3686 ( \4001 , \3681 , \360 );
and \U$3687 ( \4002 , \3264 , \358 );
nor \U$3688 ( \4003 , \4001 , \4002 );
xnor \U$3689 ( \4004 , \4003 , \341 );
and \U$3690 ( \4005 , \3999 , \4004 );
and \U$3691 ( \4006 , \3995 , \4004 );
or \U$3692 ( \4007 , \4000 , \4005 , \4006 );
and \U$3693 ( \4008 , \3990 , \4007 );
and \U$3694 ( \4009 , \3974 , \4007 );
or \U$3695 ( \4010 , \3991 , \4008 , \4009 );
buf \U$3696 ( \4011 , RIc0c6870_102);
and \U$3697 ( \4012 , \4011 , \323 );
and \U$3698 ( \4013 , \3889 , \321 );
nor \U$3699 ( \4014 , \4012 , \4013 );
xnor \U$3700 ( \4015 , \4014 , \328 );
buf \U$3701 ( \4016 , RIc0c67f8_103);
and \U$3702 ( \4017 , \4016 , \317 );
or \U$3703 ( \4018 , \4015 , \4017 );
and \U$3704 ( \4019 , \3889 , \323 );
and \U$3705 ( \4020 , \3681 , \321 );
nor \U$3706 ( \4021 , \4019 , \4020 );
xnor \U$3707 ( \4022 , \4021 , \328 );
and \U$3708 ( \4023 , \4018 , \4022 );
and \U$3709 ( \4024 , \4011 , \317 );
and \U$3710 ( \4025 , \4022 , \4024 );
and \U$3711 ( \4026 , \4018 , \4024 );
or \U$3712 ( \4027 , \4023 , \4025 , \4026 );
and \U$3713 ( \4028 , \4010 , \4027 );
xor \U$3714 ( \4029 , \3447 , \3782 );
xor \U$3715 ( \4030 , \3782 , \3783 );
not \U$3716 ( \4031 , \4030 );
and \U$3717 ( \4032 , \4029 , \4031 );
and \U$3718 ( \4033 , \316 , \4032 );
not \U$3719 ( \4034 , \4033 );
xnor \U$3720 ( \4035 , \4034 , \3786 );
and \U$3721 ( \4036 , \348 , \3637 );
and \U$3722 ( \4037 , \330 , \3635 );
nor \U$3723 ( \4038 , \4036 , \4037 );
xnor \U$3724 ( \4039 , \4038 , \3450 );
and \U$3725 ( \4040 , \4035 , \4039 );
and \U$3726 ( \4041 , \417 , \3324 );
and \U$3727 ( \4042 , \369 , \3322 );
nor \U$3728 ( \4043 , \4041 , \4042 );
xnor \U$3729 ( \4044 , \4043 , \3119 );
and \U$3730 ( \4045 , \4039 , \4044 );
and \U$3731 ( \4046 , \4035 , \4044 );
or \U$3732 ( \4047 , \4040 , \4045 , \4046 );
and \U$3733 ( \4048 , \494 , \2918 );
and \U$3734 ( \4049 , \425 , \2916 );
nor \U$3735 ( \4050 , \4048 , \4049 );
xnor \U$3736 ( \4051 , \4050 , \2769 );
and \U$3737 ( \4052 , \553 , \2596 );
and \U$3738 ( \4053 , \499 , \2594 );
nor \U$3739 ( \4054 , \4052 , \4053 );
xnor \U$3740 ( \4055 , \4054 , \2454 );
and \U$3741 ( \4056 , \4051 , \4055 );
and \U$3742 ( \4057 , \681 , \2300 );
and \U$3743 ( \4058 , \604 , \2298 );
nor \U$3744 ( \4059 , \4057 , \4058 );
xnor \U$3745 ( \4060 , \4059 , \2163 );
and \U$3746 ( \4061 , \4055 , \4060 );
and \U$3747 ( \4062 , \4051 , \4060 );
or \U$3748 ( \4063 , \4056 , \4061 , \4062 );
and \U$3749 ( \4064 , \4047 , \4063 );
and \U$3750 ( \4065 , \789 , \2094 );
and \U$3751 ( \4066 , \709 , \2092 );
nor \U$3752 ( \4067 , \4065 , \4066 );
xnor \U$3753 ( \4068 , \4067 , \1942 );
and \U$3754 ( \4069 , \925 , \1826 );
and \U$3755 ( \4070 , \863 , \1824 );
nor \U$3756 ( \4071 , \4069 , \4070 );
xnor \U$3757 ( \4072 , \4071 , \1670 );
and \U$3758 ( \4073 , \4068 , \4072 );
and \U$3759 ( \4074 , \1186 , \1554 );
and \U$3760 ( \4075 , \988 , \1552 );
nor \U$3761 ( \4076 , \4074 , \4075 );
xnor \U$3762 ( \4077 , \4076 , \1441 );
and \U$3763 ( \4078 , \4072 , \4077 );
and \U$3764 ( \4079 , \4068 , \4077 );
or \U$3765 ( \4080 , \4073 , \4078 , \4079 );
and \U$3766 ( \4081 , \4063 , \4080 );
and \U$3767 ( \4082 , \4047 , \4080 );
or \U$3768 ( \4083 , \4064 , \4081 , \4082 );
and \U$3769 ( \4084 , \4027 , \4083 );
and \U$3770 ( \4085 , \4010 , \4083 );
or \U$3771 ( \4086 , \4028 , \4084 , \4085 );
xor \U$3772 ( \4087 , \3839 , \3843 );
xor \U$3773 ( \4088 , \4087 , \3848 );
xor \U$3774 ( \4089 , \3855 , \3859 );
xor \U$3775 ( \4090 , \4089 , \3864 );
and \U$3776 ( \4091 , \4088 , \4090 );
xor \U$3777 ( \4092 , \3872 , \3876 );
xor \U$3778 ( \4093 , \4092 , \3881 );
and \U$3779 ( \4094 , \4090 , \4093 );
and \U$3780 ( \4095 , \4088 , \4093 );
or \U$3781 ( \4096 , \4091 , \4094 , \4095 );
xor \U$3782 ( \4097 , \3787 , \3791 );
xor \U$3783 ( \4098 , \4097 , \3796 );
xor \U$3784 ( \4099 , \3803 , \3807 );
xor \U$3785 ( \4100 , \4099 , \3812 );
and \U$3786 ( \4101 , \4098 , \4100 );
xor \U$3787 ( \4102 , \3820 , \3824 );
xor \U$3788 ( \4103 , \4102 , \3829 );
and \U$3789 ( \4104 , \4100 , \4103 );
and \U$3790 ( \4105 , \4098 , \4103 );
or \U$3791 ( \4106 , \4101 , \4104 , \4105 );
and \U$3792 ( \4107 , \4096 , \4106 );
xor \U$3793 ( \4108 , \3620 , \3624 );
xor \U$3794 ( \4109 , \4108 , \3629 );
and \U$3795 ( \4110 , \4106 , \4109 );
and \U$3796 ( \4111 , \4096 , \4109 );
or \U$3797 ( \4112 , \4107 , \4110 , \4111 );
and \U$3798 ( \4113 , \4086 , \4112 );
xor \U$3799 ( \4114 , \3640 , \3644 );
xor \U$3800 ( \4115 , \4114 , \3649 );
xor \U$3801 ( \4116 , \3898 , \3900 );
xor \U$3802 ( \4117 , \4116 , \3903 );
and \U$3803 ( \4118 , \4115 , \4117 );
xnor \U$3804 ( \4119 , \3890 , \3892 );
and \U$3805 ( \4120 , \4117 , \4119 );
and \U$3806 ( \4121 , \4115 , \4119 );
or \U$3807 ( \4122 , \4118 , \4120 , \4121 );
and \U$3808 ( \4123 , \4112 , \4122 );
and \U$3809 ( \4124 , \4086 , \4122 );
or \U$3810 ( \4125 , \4113 , \4123 , \4124 );
xor \U$3811 ( \4126 , \3835 , \3887 );
xor \U$3812 ( \4127 , \4126 , \3893 );
xor \U$3813 ( \4128 , \3906 , \3908 );
xor \U$3814 ( \4129 , \4128 , \3911 );
and \U$3815 ( \4130 , \4127 , \4129 );
xor \U$3816 ( \4131 , \3917 , \3919 );
xor \U$3817 ( \4132 , \4131 , \3922 );
and \U$3818 ( \4133 , \4129 , \4132 );
and \U$3819 ( \4134 , \4127 , \4132 );
or \U$3820 ( \4135 , \4130 , \4133 , \4134 );
and \U$3821 ( \4136 , \4125 , \4135 );
xor \U$3822 ( \4137 , \3930 , \3932 );
xor \U$3823 ( \4138 , \4137 , \3935 );
and \U$3824 ( \4139 , \4135 , \4138 );
and \U$3825 ( \4140 , \4125 , \4138 );
or \U$3826 ( \4141 , \4136 , \4139 , \4140 );
xor \U$3827 ( \4142 , \3721 , \3739 );
xor \U$3828 ( \4143 , \4142 , \3749 );
and \U$3829 ( \4144 , \4141 , \4143 );
xor \U$3830 ( \4145 , \3928 , \3938 );
xor \U$3831 ( \4146 , \4145 , \3941 );
and \U$3832 ( \4147 , \4143 , \4146 );
and \U$3833 ( \4148 , \4141 , \4146 );
or \U$3834 ( \4149 , \4144 , \4147 , \4148 );
xor \U$3835 ( \4150 , \3944 , \3946 );
xor \U$3836 ( \4151 , \4150 , \3949 );
and \U$3837 ( \4152 , \4149 , \4151 );
and \U$3838 ( \4153 , \3958 , \4152 );
xor \U$3839 ( \4154 , \3958 , \4152 );
xor \U$3840 ( \4155 , \4149 , \4151 );
and \U$3841 ( \4156 , \1799 , \996 );
and \U$3842 ( \4157 , \1791 , \994 );
nor \U$3843 ( \4158 , \4156 , \4157 );
xnor \U$3844 ( \4159 , \4158 , \902 );
and \U$3845 ( \4160 , \2047 , \826 );
and \U$3846 ( \4161 , \2042 , \824 );
nor \U$3847 ( \4162 , \4160 , \4161 );
xnor \U$3848 ( \4163 , \4162 , \754 );
and \U$3849 ( \4164 , \4159 , \4163 );
and \U$3850 ( \4165 , \2377 , \692 );
and \U$3851 ( \4166 , \2233 , \690 );
nor \U$3852 ( \4167 , \4165 , \4166 );
xnor \U$3853 ( \4168 , \4167 , \649 );
and \U$3854 ( \4169 , \4163 , \4168 );
and \U$3855 ( \4170 , \4159 , \4168 );
or \U$3856 ( \4171 , \4164 , \4169 , \4170 );
and \U$3857 ( \4172 , \1274 , \1554 );
and \U$3858 ( \4173 , \1186 , \1552 );
nor \U$3859 ( \4174 , \4172 , \4173 );
xnor \U$3860 ( \4175 , \4174 , \1441 );
and \U$3861 ( \4176 , \1384 , \1360 );
and \U$3862 ( \4177 , \1379 , \1358 );
nor \U$3863 ( \4178 , \4176 , \4177 );
xnor \U$3864 ( \4179 , \4178 , \1224 );
and \U$3865 ( \4180 , \4175 , \4179 );
and \U$3866 ( \4181 , \1615 , \1160 );
and \U$3867 ( \4182 , \1500 , \1158 );
nor \U$3868 ( \4183 , \4181 , \4182 );
xnor \U$3869 ( \4184 , \4183 , \1082 );
and \U$3870 ( \4185 , \4179 , \4184 );
and \U$3871 ( \4186 , \4175 , \4184 );
or \U$3872 ( \4187 , \4180 , \4185 , \4186 );
and \U$3873 ( \4188 , \4171 , \4187 );
and \U$3874 ( \4189 , \2666 , \579 );
and \U$3875 ( \4190 , \2641 , \577 );
nor \U$3876 ( \4191 , \4189 , \4190 );
xnor \U$3877 ( \4192 , \4191 , \530 );
and \U$3878 ( \4193 , \3007 , \478 );
and \U$3879 ( \4194 , \2840 , \476 );
nor \U$3880 ( \4195 , \4193 , \4194 );
xnor \U$3881 ( \4196 , \4195 , \437 );
and \U$3882 ( \4197 , \4192 , \4196 );
and \U$3883 ( \4198 , \3264 , \408 );
and \U$3884 ( \4199 , \3145 , \406 );
nor \U$3885 ( \4200 , \4198 , \4199 );
xnor \U$3886 ( \4201 , \4200 , \378 );
and \U$3887 ( \4202 , \4196 , \4201 );
and \U$3888 ( \4203 , \4192 , \4201 );
or \U$3889 ( \4204 , \4197 , \4202 , \4203 );
and \U$3890 ( \4205 , \4187 , \4204 );
and \U$3891 ( \4206 , \4171 , \4204 );
or \U$3892 ( \4207 , \4188 , \4205 , \4206 );
buf \U$3893 ( \4208 , RIc0c8508_41);
buf \U$3894 ( \4209 , RIc0c8490_42);
and \U$3895 ( \4210 , \4208 , \4209 );
not \U$3896 ( \4211 , \4210 );
and \U$3897 ( \4212 , \3783 , \4211 );
not \U$3898 ( \4213 , \4212 );
and \U$3899 ( \4214 , \330 , \4032 );
and \U$3900 ( \4215 , \316 , \4030 );
nor \U$3901 ( \4216 , \4214 , \4215 );
xnor \U$3902 ( \4217 , \4216 , \3786 );
and \U$3903 ( \4218 , \4213 , \4217 );
and \U$3904 ( \4219 , \369 , \3637 );
and \U$3905 ( \4220 , \348 , \3635 );
nor \U$3906 ( \4221 , \4219 , \4220 );
xnor \U$3907 ( \4222 , \4221 , \3450 );
and \U$3908 ( \4223 , \4217 , \4222 );
and \U$3909 ( \4224 , \4213 , \4222 );
or \U$3910 ( \4225 , \4218 , \4223 , \4224 );
and \U$3911 ( \4226 , \425 , \3324 );
and \U$3912 ( \4227 , \417 , \3322 );
nor \U$3913 ( \4228 , \4226 , \4227 );
xnor \U$3914 ( \4229 , \4228 , \3119 );
and \U$3915 ( \4230 , \499 , \2918 );
and \U$3916 ( \4231 , \494 , \2916 );
nor \U$3917 ( \4232 , \4230 , \4231 );
xnor \U$3918 ( \4233 , \4232 , \2769 );
and \U$3919 ( \4234 , \4229 , \4233 );
and \U$3920 ( \4235 , \604 , \2596 );
and \U$3921 ( \4236 , \553 , \2594 );
nor \U$3922 ( \4237 , \4235 , \4236 );
xnor \U$3923 ( \4238 , \4237 , \2454 );
and \U$3924 ( \4239 , \4233 , \4238 );
and \U$3925 ( \4240 , \4229 , \4238 );
or \U$3926 ( \4241 , \4234 , \4239 , \4240 );
and \U$3927 ( \4242 , \4225 , \4241 );
and \U$3928 ( \4243 , \709 , \2300 );
and \U$3929 ( \4244 , \681 , \2298 );
nor \U$3930 ( \4245 , \4243 , \4244 );
xnor \U$3931 ( \4246 , \4245 , \2163 );
and \U$3932 ( \4247 , \863 , \2094 );
and \U$3933 ( \4248 , \789 , \2092 );
nor \U$3934 ( \4249 , \4247 , \4248 );
xnor \U$3935 ( \4250 , \4249 , \1942 );
and \U$3936 ( \4251 , \4246 , \4250 );
and \U$3937 ( \4252 , \988 , \1826 );
and \U$3938 ( \4253 , \925 , \1824 );
nor \U$3939 ( \4254 , \4252 , \4253 );
xnor \U$3940 ( \4255 , \4254 , \1670 );
and \U$3941 ( \4256 , \4250 , \4255 );
and \U$3942 ( \4257 , \4246 , \4255 );
or \U$3943 ( \4258 , \4251 , \4256 , \4257 );
and \U$3944 ( \4259 , \4241 , \4258 );
and \U$3945 ( \4260 , \4225 , \4258 );
or \U$3946 ( \4261 , \4242 , \4259 , \4260 );
and \U$3947 ( \4262 , \4207 , \4261 );
and \U$3948 ( \4263 , \3889 , \360 );
and \U$3949 ( \4264 , \3681 , \358 );
nor \U$3950 ( \4265 , \4263 , \4264 );
xnor \U$3951 ( \4266 , \4265 , \341 );
and \U$3952 ( \4267 , \4016 , \323 );
and \U$3953 ( \4268 , \4011 , \321 );
nor \U$3954 ( \4269 , \4267 , \4268 );
xnor \U$3955 ( \4270 , \4269 , \328 );
and \U$3956 ( \4271 , \4266 , \4270 );
buf \U$3957 ( \4272 , RIc0c6780_104);
and \U$3958 ( \4273 , \4272 , \317 );
and \U$3959 ( \4274 , \4270 , \4273 );
and \U$3960 ( \4275 , \4266 , \4273 );
or \U$3961 ( \4276 , \4271 , \4274 , \4275 );
xor \U$3962 ( \4277 , \3995 , \3999 );
xor \U$3963 ( \4278 , \4277 , \4004 );
and \U$3964 ( \4279 , \4276 , \4278 );
xnor \U$3965 ( \4280 , \4015 , \4017 );
and \U$3966 ( \4281 , \4278 , \4280 );
and \U$3967 ( \4282 , \4276 , \4280 );
or \U$3968 ( \4283 , \4279 , \4281 , \4282 );
and \U$3969 ( \4284 , \4261 , \4283 );
and \U$3970 ( \4285 , \4207 , \4283 );
or \U$3971 ( \4286 , \4262 , \4284 , \4285 );
xor \U$3972 ( \4287 , \3962 , \3966 );
xor \U$3973 ( \4288 , \4287 , \3971 );
xor \U$3974 ( \4289 , \3978 , \3982 );
xor \U$3975 ( \4290 , \4289 , \3987 );
and \U$3976 ( \4291 , \4288 , \4290 );
xor \U$3977 ( \4292 , \4068 , \4072 );
xor \U$3978 ( \4293 , \4292 , \4077 );
and \U$3979 ( \4294 , \4290 , \4293 );
and \U$3980 ( \4295 , \4288 , \4293 );
or \U$3981 ( \4296 , \4291 , \4294 , \4295 );
xor \U$3982 ( \4297 , \4035 , \4039 );
xor \U$3983 ( \4298 , \4297 , \4044 );
xor \U$3984 ( \4299 , \4051 , \4055 );
xor \U$3985 ( \4300 , \4299 , \4060 );
and \U$3986 ( \4301 , \4298 , \4300 );
and \U$3987 ( \4302 , \4296 , \4301 );
xor \U$3988 ( \4303 , \4098 , \4100 );
xor \U$3989 ( \4304 , \4303 , \4103 );
and \U$3990 ( \4305 , \4301 , \4304 );
and \U$3991 ( \4306 , \4296 , \4304 );
or \U$3992 ( \4307 , \4302 , \4305 , \4306 );
and \U$3993 ( \4308 , \4286 , \4307 );
xor \U$3994 ( \4309 , \3974 , \3990 );
xor \U$3995 ( \4310 , \4309 , \4007 );
xor \U$3996 ( \4311 , \4018 , \4022 );
xor \U$3997 ( \4312 , \4311 , \4024 );
and \U$3998 ( \4313 , \4310 , \4312 );
xor \U$3999 ( \4314 , \4088 , \4090 );
xor \U$4000 ( \4315 , \4314 , \4093 );
and \U$4001 ( \4316 , \4312 , \4315 );
and \U$4002 ( \4317 , \4310 , \4315 );
or \U$4003 ( \4318 , \4313 , \4316 , \4317 );
and \U$4004 ( \4319 , \4307 , \4318 );
and \U$4005 ( \4320 , \4286 , \4318 );
or \U$4006 ( \4321 , \4308 , \4319 , \4320 );
xor \U$4007 ( \4322 , \3799 , \3815 );
xor \U$4008 ( \4323 , \4322 , \3832 );
xor \U$4009 ( \4324 , \3851 , \3867 );
xor \U$4010 ( \4325 , \4324 , \3884 );
and \U$4011 ( \4326 , \4323 , \4325 );
xor \U$4012 ( \4327 , \4115 , \4117 );
xor \U$4013 ( \4328 , \4327 , \4119 );
and \U$4014 ( \4329 , \4325 , \4328 );
and \U$4015 ( \4330 , \4323 , \4328 );
or \U$4016 ( \4331 , \4326 , \4329 , \4330 );
and \U$4017 ( \4332 , \4321 , \4331 );
xor \U$4018 ( \4333 , \4127 , \4129 );
xor \U$4019 ( \4334 , \4333 , \4132 );
and \U$4020 ( \4335 , \4331 , \4334 );
and \U$4021 ( \4336 , \4321 , \4334 );
or \U$4022 ( \4337 , \4332 , \4335 , \4336 );
xor \U$4023 ( \4338 , \3896 , \3914 );
xor \U$4024 ( \4339 , \4338 , \3925 );
and \U$4025 ( \4340 , \4337 , \4339 );
xor \U$4026 ( \4341 , \4125 , \4135 );
xor \U$4027 ( \4342 , \4341 , \4138 );
and \U$4028 ( \4343 , \4339 , \4342 );
and \U$4029 ( \4344 , \4337 , \4342 );
or \U$4030 ( \4345 , \4340 , \4343 , \4344 );
xor \U$4031 ( \4346 , \4141 , \4143 );
xor \U$4032 ( \4347 , \4346 , \4146 );
and \U$4033 ( \4348 , \4345 , \4347 );
and \U$4034 ( \4349 , \4155 , \4348 );
xor \U$4035 ( \4350 , \4155 , \4348 );
xor \U$4036 ( \4351 , \4345 , \4347 );
xor \U$4037 ( \4352 , \3783 , \4208 );
xor \U$4038 ( \4353 , \4208 , \4209 );
not \U$4039 ( \4354 , \4353 );
and \U$4040 ( \4355 , \4352 , \4354 );
and \U$4041 ( \4356 , \316 , \4355 );
not \U$4042 ( \4357 , \4356 );
xnor \U$4043 ( \4358 , \4357 , \4212 );
and \U$4044 ( \4359 , \348 , \4032 );
and \U$4045 ( \4360 , \330 , \4030 );
nor \U$4046 ( \4361 , \4359 , \4360 );
xnor \U$4047 ( \4362 , \4361 , \3786 );
and \U$4048 ( \4363 , \4358 , \4362 );
and \U$4049 ( \4364 , \417 , \3637 );
and \U$4050 ( \4365 , \369 , \3635 );
nor \U$4051 ( \4366 , \4364 , \4365 );
xnor \U$4052 ( \4367 , \4366 , \3450 );
and \U$4053 ( \4368 , \4362 , \4367 );
and \U$4054 ( \4369 , \4358 , \4367 );
or \U$4055 ( \4370 , \4363 , \4368 , \4369 );
and \U$4056 ( \4371 , \494 , \3324 );
and \U$4057 ( \4372 , \425 , \3322 );
nor \U$4058 ( \4373 , \4371 , \4372 );
xnor \U$4059 ( \4374 , \4373 , \3119 );
and \U$4060 ( \4375 , \553 , \2918 );
and \U$4061 ( \4376 , \499 , \2916 );
nor \U$4062 ( \4377 , \4375 , \4376 );
xnor \U$4063 ( \4378 , \4377 , \2769 );
and \U$4064 ( \4379 , \4374 , \4378 );
and \U$4065 ( \4380 , \681 , \2596 );
and \U$4066 ( \4381 , \604 , \2594 );
nor \U$4067 ( \4382 , \4380 , \4381 );
xnor \U$4068 ( \4383 , \4382 , \2454 );
and \U$4069 ( \4384 , \4378 , \4383 );
and \U$4070 ( \4385 , \4374 , \4383 );
or \U$4071 ( \4386 , \4379 , \4384 , \4385 );
and \U$4072 ( \4387 , \4370 , \4386 );
and \U$4073 ( \4388 , \789 , \2300 );
and \U$4074 ( \4389 , \709 , \2298 );
nor \U$4075 ( \4390 , \4388 , \4389 );
xnor \U$4076 ( \4391 , \4390 , \2163 );
and \U$4077 ( \4392 , \925 , \2094 );
and \U$4078 ( \4393 , \863 , \2092 );
nor \U$4079 ( \4394 , \4392 , \4393 );
xnor \U$4080 ( \4395 , \4394 , \1942 );
and \U$4081 ( \4396 , \4391 , \4395 );
and \U$4082 ( \4397 , \1186 , \1826 );
and \U$4083 ( \4398 , \988 , \1824 );
nor \U$4084 ( \4399 , \4397 , \4398 );
xnor \U$4085 ( \4400 , \4399 , \1670 );
and \U$4086 ( \4401 , \4395 , \4400 );
and \U$4087 ( \4402 , \4391 , \4400 );
or \U$4088 ( \4403 , \4396 , \4401 , \4402 );
and \U$4089 ( \4404 , \4386 , \4403 );
and \U$4090 ( \4405 , \4370 , \4403 );
or \U$4091 ( \4406 , \4387 , \4404 , \4405 );
and \U$4092 ( \4407 , \2840 , \579 );
and \U$4093 ( \4408 , \2666 , \577 );
nor \U$4094 ( \4409 , \4407 , \4408 );
xnor \U$4095 ( \4410 , \4409 , \530 );
and \U$4096 ( \4411 , \3145 , \478 );
and \U$4097 ( \4412 , \3007 , \476 );
nor \U$4098 ( \4413 , \4411 , \4412 );
xnor \U$4099 ( \4414 , \4413 , \437 );
and \U$4100 ( \4415 , \4410 , \4414 );
and \U$4101 ( \4416 , \3681 , \408 );
and \U$4102 ( \4417 , \3264 , \406 );
nor \U$4103 ( \4418 , \4416 , \4417 );
xnor \U$4104 ( \4419 , \4418 , \378 );
and \U$4105 ( \4420 , \4414 , \4419 );
and \U$4106 ( \4421 , \4410 , \4419 );
or \U$4107 ( \4422 , \4415 , \4420 , \4421 );
and \U$4108 ( \4423 , \1379 , \1554 );
and \U$4109 ( \4424 , \1274 , \1552 );
nor \U$4110 ( \4425 , \4423 , \4424 );
xnor \U$4111 ( \4426 , \4425 , \1441 );
and \U$4112 ( \4427 , \1500 , \1360 );
and \U$4113 ( \4428 , \1384 , \1358 );
nor \U$4114 ( \4429 , \4427 , \4428 );
xnor \U$4115 ( \4430 , \4429 , \1224 );
and \U$4116 ( \4431 , \4426 , \4430 );
and \U$4117 ( \4432 , \1791 , \1160 );
and \U$4118 ( \4433 , \1615 , \1158 );
nor \U$4119 ( \4434 , \4432 , \4433 );
xnor \U$4120 ( \4435 , \4434 , \1082 );
and \U$4121 ( \4436 , \4430 , \4435 );
and \U$4122 ( \4437 , \4426 , \4435 );
or \U$4123 ( \4438 , \4431 , \4436 , \4437 );
and \U$4124 ( \4439 , \4422 , \4438 );
and \U$4125 ( \4440 , \2042 , \996 );
and \U$4126 ( \4441 , \1799 , \994 );
nor \U$4127 ( \4442 , \4440 , \4441 );
xnor \U$4128 ( \4443 , \4442 , \902 );
and \U$4129 ( \4444 , \2233 , \826 );
and \U$4130 ( \4445 , \2047 , \824 );
nor \U$4131 ( \4446 , \4444 , \4445 );
xnor \U$4132 ( \4447 , \4446 , \754 );
and \U$4133 ( \4448 , \4443 , \4447 );
and \U$4134 ( \4449 , \2641 , \692 );
and \U$4135 ( \4450 , \2377 , \690 );
nor \U$4136 ( \4451 , \4449 , \4450 );
xnor \U$4137 ( \4452 , \4451 , \649 );
and \U$4138 ( \4453 , \4447 , \4452 );
and \U$4139 ( \4454 , \4443 , \4452 );
or \U$4140 ( \4455 , \4448 , \4453 , \4454 );
and \U$4141 ( \4456 , \4438 , \4455 );
and \U$4142 ( \4457 , \4422 , \4455 );
or \U$4143 ( \4458 , \4439 , \4456 , \4457 );
and \U$4144 ( \4459 , \4406 , \4458 );
and \U$4145 ( \4460 , \4011 , \360 );
and \U$4146 ( \4461 , \3889 , \358 );
nor \U$4147 ( \4462 , \4460 , \4461 );
xnor \U$4148 ( \4463 , \4462 , \341 );
and \U$4149 ( \4464 , \4272 , \323 );
and \U$4150 ( \4465 , \4016 , \321 );
nor \U$4151 ( \4466 , \4464 , \4465 );
xnor \U$4152 ( \4467 , \4466 , \328 );
and \U$4153 ( \4468 , \4463 , \4467 );
buf \U$4154 ( \4469 , RIc0c6708_105);
and \U$4155 ( \4470 , \4469 , \317 );
and \U$4156 ( \4471 , \4467 , \4470 );
and \U$4157 ( \4472 , \4463 , \4470 );
or \U$4158 ( \4473 , \4468 , \4471 , \4472 );
xor \U$4159 ( \4474 , \4266 , \4270 );
xor \U$4160 ( \4475 , \4474 , \4273 );
and \U$4161 ( \4476 , \4473 , \4475 );
xor \U$4162 ( \4477 , \4192 , \4196 );
xor \U$4163 ( \4478 , \4477 , \4201 );
and \U$4164 ( \4479 , \4475 , \4478 );
and \U$4165 ( \4480 , \4473 , \4478 );
or \U$4166 ( \4481 , \4476 , \4479 , \4480 );
and \U$4167 ( \4482 , \4458 , \4481 );
and \U$4168 ( \4483 , \4406 , \4481 );
or \U$4169 ( \4484 , \4459 , \4482 , \4483 );
xor \U$4170 ( \4485 , \4171 , \4187 );
xor \U$4171 ( \4486 , \4485 , \4204 );
xor \U$4172 ( \4487 , \4225 , \4241 );
xor \U$4173 ( \4488 , \4487 , \4258 );
and \U$4174 ( \4489 , \4486 , \4488 );
xor \U$4175 ( \4490 , \4276 , \4278 );
xor \U$4176 ( \4491 , \4490 , \4280 );
and \U$4177 ( \4492 , \4488 , \4491 );
and \U$4178 ( \4493 , \4486 , \4491 );
or \U$4179 ( \4494 , \4489 , \4492 , \4493 );
and \U$4180 ( \4495 , \4484 , \4494 );
xor \U$4181 ( \4496 , \4159 , \4163 );
xor \U$4182 ( \4497 , \4496 , \4168 );
xor \U$4183 ( \4498 , \4175 , \4179 );
xor \U$4184 ( \4499 , \4498 , \4184 );
and \U$4185 ( \4500 , \4497 , \4499 );
xor \U$4186 ( \4501 , \4246 , \4250 );
xor \U$4187 ( \4502 , \4501 , \4255 );
and \U$4188 ( \4503 , \4499 , \4502 );
and \U$4189 ( \4504 , \4497 , \4502 );
or \U$4190 ( \4505 , \4500 , \4503 , \4504 );
xor \U$4191 ( \4506 , \4288 , \4290 );
xor \U$4192 ( \4507 , \4506 , \4293 );
and \U$4193 ( \4508 , \4505 , \4507 );
xor \U$4194 ( \4509 , \4298 , \4300 );
and \U$4195 ( \4510 , \4507 , \4509 );
and \U$4196 ( \4511 , \4505 , \4509 );
or \U$4197 ( \4512 , \4508 , \4510 , \4511 );
and \U$4198 ( \4513 , \4494 , \4512 );
and \U$4199 ( \4514 , \4484 , \4512 );
or \U$4200 ( \4515 , \4495 , \4513 , \4514 );
xor \U$4201 ( \4516 , \4047 , \4063 );
xor \U$4202 ( \4517 , \4516 , \4080 );
xor \U$4203 ( \4518 , \4296 , \4301 );
xor \U$4204 ( \4519 , \4518 , \4304 );
and \U$4205 ( \4520 , \4517 , \4519 );
xor \U$4206 ( \4521 , \4310 , \4312 );
xor \U$4207 ( \4522 , \4521 , \4315 );
and \U$4208 ( \4523 , \4519 , \4522 );
and \U$4209 ( \4524 , \4517 , \4522 );
or \U$4210 ( \4525 , \4520 , \4523 , \4524 );
and \U$4211 ( \4526 , \4515 , \4525 );
xor \U$4212 ( \4527 , \4096 , \4106 );
xor \U$4213 ( \4528 , \4527 , \4109 );
and \U$4214 ( \4529 , \4525 , \4528 );
and \U$4215 ( \4530 , \4515 , \4528 );
or \U$4216 ( \4531 , \4526 , \4529 , \4530 );
xor \U$4217 ( \4532 , \4010 , \4027 );
xor \U$4218 ( \4533 , \4532 , \4083 );
xor \U$4219 ( \4534 , \4286 , \4307 );
xor \U$4220 ( \4535 , \4534 , \4318 );
and \U$4221 ( \4536 , \4533 , \4535 );
xor \U$4222 ( \4537 , \4323 , \4325 );
xor \U$4223 ( \4538 , \4537 , \4328 );
and \U$4224 ( \4539 , \4535 , \4538 );
and \U$4225 ( \4540 , \4533 , \4538 );
or \U$4226 ( \4541 , \4536 , \4539 , \4540 );
and \U$4227 ( \4542 , \4531 , \4541 );
xor \U$4228 ( \4543 , \4086 , \4112 );
xor \U$4229 ( \4544 , \4543 , \4122 );
and \U$4230 ( \4545 , \4541 , \4544 );
and \U$4231 ( \4546 , \4531 , \4544 );
or \U$4232 ( \4547 , \4542 , \4545 , \4546 );
xor \U$4233 ( \4548 , \4337 , \4339 );
xor \U$4234 ( \4549 , \4548 , \4342 );
and \U$4235 ( \4550 , \4547 , \4549 );
and \U$4236 ( \4551 , \4351 , \4550 );
xor \U$4237 ( \4552 , \4351 , \4550 );
xor \U$4238 ( \4553 , \4547 , \4549 );
and \U$4239 ( \4554 , \709 , \2596 );
and \U$4240 ( \4555 , \681 , \2594 );
nor \U$4241 ( \4556 , \4554 , \4555 );
xnor \U$4242 ( \4557 , \4556 , \2454 );
and \U$4243 ( \4558 , \863 , \2300 );
and \U$4244 ( \4559 , \789 , \2298 );
nor \U$4245 ( \4560 , \4558 , \4559 );
xnor \U$4246 ( \4561 , \4560 , \2163 );
and \U$4247 ( \4562 , \4557 , \4561 );
and \U$4248 ( \4563 , \988 , \2094 );
and \U$4249 ( \4564 , \925 , \2092 );
nor \U$4250 ( \4565 , \4563 , \4564 );
xnor \U$4251 ( \4566 , \4565 , \1942 );
and \U$4252 ( \4567 , \4561 , \4566 );
and \U$4253 ( \4568 , \4557 , \4566 );
or \U$4254 ( \4569 , \4562 , \4567 , \4568 );
buf \U$4255 ( \4570 , RIc0c8418_43);
buf \U$4256 ( \4571 , RIc0c83a0_44);
and \U$4257 ( \4572 , \4570 , \4571 );
not \U$4258 ( \4573 , \4572 );
and \U$4259 ( \4574 , \4209 , \4573 );
not \U$4260 ( \4575 , \4574 );
and \U$4261 ( \4576 , \330 , \4355 );
and \U$4262 ( \4577 , \316 , \4353 );
nor \U$4263 ( \4578 , \4576 , \4577 );
xnor \U$4264 ( \4579 , \4578 , \4212 );
and \U$4265 ( \4580 , \4575 , \4579 );
and \U$4266 ( \4581 , \369 , \4032 );
and \U$4267 ( \4582 , \348 , \4030 );
nor \U$4268 ( \4583 , \4581 , \4582 );
xnor \U$4269 ( \4584 , \4583 , \3786 );
and \U$4270 ( \4585 , \4579 , \4584 );
and \U$4271 ( \4586 , \4575 , \4584 );
or \U$4272 ( \4587 , \4580 , \4585 , \4586 );
and \U$4273 ( \4588 , \4569 , \4587 );
and \U$4274 ( \4589 , \425 , \3637 );
and \U$4275 ( \4590 , \417 , \3635 );
nor \U$4276 ( \4591 , \4589 , \4590 );
xnor \U$4277 ( \4592 , \4591 , \3450 );
and \U$4278 ( \4593 , \499 , \3324 );
and \U$4279 ( \4594 , \494 , \3322 );
nor \U$4280 ( \4595 , \4593 , \4594 );
xnor \U$4281 ( \4596 , \4595 , \3119 );
and \U$4282 ( \4597 , \4592 , \4596 );
and \U$4283 ( \4598 , \604 , \2918 );
and \U$4284 ( \4599 , \553 , \2916 );
nor \U$4285 ( \4600 , \4598 , \4599 );
xnor \U$4286 ( \4601 , \4600 , \2769 );
and \U$4287 ( \4602 , \4596 , \4601 );
and \U$4288 ( \4603 , \4592 , \4601 );
or \U$4289 ( \4604 , \4597 , \4602 , \4603 );
and \U$4290 ( \4605 , \4587 , \4604 );
and \U$4291 ( \4606 , \4569 , \4604 );
or \U$4292 ( \4607 , \4588 , \4605 , \4606 );
and \U$4293 ( \4608 , \2666 , \692 );
and \U$4294 ( \4609 , \2641 , \690 );
nor \U$4295 ( \4610 , \4608 , \4609 );
xnor \U$4296 ( \4611 , \4610 , \649 );
and \U$4297 ( \4612 , \3007 , \579 );
and \U$4298 ( \4613 , \2840 , \577 );
nor \U$4299 ( \4614 , \4612 , \4613 );
xnor \U$4300 ( \4615 , \4614 , \530 );
and \U$4301 ( \4616 , \4611 , \4615 );
and \U$4302 ( \4617 , \3264 , \478 );
and \U$4303 ( \4618 , \3145 , \476 );
nor \U$4304 ( \4619 , \4617 , \4618 );
xnor \U$4305 ( \4620 , \4619 , \437 );
and \U$4306 ( \4621 , \4615 , \4620 );
and \U$4307 ( \4622 , \4611 , \4620 );
or \U$4308 ( \4623 , \4616 , \4621 , \4622 );
and \U$4309 ( \4624 , \1274 , \1826 );
and \U$4310 ( \4625 , \1186 , \1824 );
nor \U$4311 ( \4626 , \4624 , \4625 );
xnor \U$4312 ( \4627 , \4626 , \1670 );
and \U$4313 ( \4628 , \1384 , \1554 );
and \U$4314 ( \4629 , \1379 , \1552 );
nor \U$4315 ( \4630 , \4628 , \4629 );
xnor \U$4316 ( \4631 , \4630 , \1441 );
and \U$4317 ( \4632 , \4627 , \4631 );
and \U$4318 ( \4633 , \1615 , \1360 );
and \U$4319 ( \4634 , \1500 , \1358 );
nor \U$4320 ( \4635 , \4633 , \4634 );
xnor \U$4321 ( \4636 , \4635 , \1224 );
and \U$4322 ( \4637 , \4631 , \4636 );
and \U$4323 ( \4638 , \4627 , \4636 );
or \U$4324 ( \4639 , \4632 , \4637 , \4638 );
and \U$4325 ( \4640 , \4623 , \4639 );
and \U$4326 ( \4641 , \1799 , \1160 );
and \U$4327 ( \4642 , \1791 , \1158 );
nor \U$4328 ( \4643 , \4641 , \4642 );
xnor \U$4329 ( \4644 , \4643 , \1082 );
and \U$4330 ( \4645 , \2047 , \996 );
and \U$4331 ( \4646 , \2042 , \994 );
nor \U$4332 ( \4647 , \4645 , \4646 );
xnor \U$4333 ( \4648 , \4647 , \902 );
and \U$4334 ( \4649 , \4644 , \4648 );
and \U$4335 ( \4650 , \2377 , \826 );
and \U$4336 ( \4651 , \2233 , \824 );
nor \U$4337 ( \4652 , \4650 , \4651 );
xnor \U$4338 ( \4653 , \4652 , \754 );
and \U$4339 ( \4654 , \4648 , \4653 );
and \U$4340 ( \4655 , \4644 , \4653 );
or \U$4341 ( \4656 , \4649 , \4654 , \4655 );
and \U$4342 ( \4657 , \4639 , \4656 );
and \U$4343 ( \4658 , \4623 , \4656 );
or \U$4344 ( \4659 , \4640 , \4657 , \4658 );
and \U$4345 ( \4660 , \4607 , \4659 );
and \U$4346 ( \4661 , \3889 , \408 );
and \U$4347 ( \4662 , \3681 , \406 );
nor \U$4348 ( \4663 , \4661 , \4662 );
xnor \U$4349 ( \4664 , \4663 , \378 );
and \U$4350 ( \4665 , \4016 , \360 );
and \U$4351 ( \4666 , \4011 , \358 );
nor \U$4352 ( \4667 , \4665 , \4666 );
xnor \U$4353 ( \4668 , \4667 , \341 );
and \U$4354 ( \4669 , \4664 , \4668 );
and \U$4355 ( \4670 , \4469 , \323 );
and \U$4356 ( \4671 , \4272 , \321 );
nor \U$4357 ( \4672 , \4670 , \4671 );
xnor \U$4358 ( \4673 , \4672 , \328 );
and \U$4359 ( \4674 , \4668 , \4673 );
and \U$4360 ( \4675 , \4664 , \4673 );
or \U$4361 ( \4676 , \4669 , \4674 , \4675 );
xor \U$4362 ( \4677 , \4463 , \4467 );
xor \U$4363 ( \4678 , \4677 , \4470 );
or \U$4364 ( \4679 , \4676 , \4678 );
and \U$4365 ( \4680 , \4659 , \4679 );
and \U$4366 ( \4681 , \4607 , \4679 );
or \U$4367 ( \4682 , \4660 , \4680 , \4681 );
xor \U$4368 ( \4683 , \4410 , \4414 );
xor \U$4369 ( \4684 , \4683 , \4419 );
xor \U$4370 ( \4685 , \4426 , \4430 );
xor \U$4371 ( \4686 , \4685 , \4435 );
and \U$4372 ( \4687 , \4684 , \4686 );
xor \U$4373 ( \4688 , \4443 , \4447 );
xor \U$4374 ( \4689 , \4688 , \4452 );
and \U$4375 ( \4690 , \4686 , \4689 );
and \U$4376 ( \4691 , \4684 , \4689 );
or \U$4377 ( \4692 , \4687 , \4690 , \4691 );
xor \U$4378 ( \4693 , \4358 , \4362 );
xor \U$4379 ( \4694 , \4693 , \4367 );
xor \U$4380 ( \4695 , \4374 , \4378 );
xor \U$4381 ( \4696 , \4695 , \4383 );
and \U$4382 ( \4697 , \4694 , \4696 );
xor \U$4383 ( \4698 , \4391 , \4395 );
xor \U$4384 ( \4699 , \4698 , \4400 );
and \U$4385 ( \4700 , \4696 , \4699 );
and \U$4386 ( \4701 , \4694 , \4699 );
or \U$4387 ( \4702 , \4697 , \4700 , \4701 );
and \U$4388 ( \4703 , \4692 , \4702 );
xor \U$4389 ( \4704 , \4229 , \4233 );
xor \U$4390 ( \4705 , \4704 , \4238 );
and \U$4391 ( \4706 , \4702 , \4705 );
and \U$4392 ( \4707 , \4692 , \4705 );
or \U$4393 ( \4708 , \4703 , \4706 , \4707 );
and \U$4394 ( \4709 , \4682 , \4708 );
xor \U$4395 ( \4710 , \4213 , \4217 );
xor \U$4396 ( \4711 , \4710 , \4222 );
xor \U$4397 ( \4712 , \4497 , \4499 );
xor \U$4398 ( \4713 , \4712 , \4502 );
and \U$4399 ( \4714 , \4711 , \4713 );
xor \U$4400 ( \4715 , \4473 , \4475 );
xor \U$4401 ( \4716 , \4715 , \4478 );
and \U$4402 ( \4717 , \4713 , \4716 );
and \U$4403 ( \4718 , \4711 , \4716 );
or \U$4404 ( \4719 , \4714 , \4717 , \4718 );
and \U$4405 ( \4720 , \4708 , \4719 );
and \U$4406 ( \4721 , \4682 , \4719 );
or \U$4407 ( \4722 , \4709 , \4720 , \4721 );
xor \U$4408 ( \4723 , \4406 , \4458 );
xor \U$4409 ( \4724 , \4723 , \4481 );
xor \U$4410 ( \4725 , \4486 , \4488 );
xor \U$4411 ( \4726 , \4725 , \4491 );
and \U$4412 ( \4727 , \4724 , \4726 );
xor \U$4413 ( \4728 , \4505 , \4507 );
xor \U$4414 ( \4729 , \4728 , \4509 );
and \U$4415 ( \4730 , \4726 , \4729 );
and \U$4416 ( \4731 , \4724 , \4729 );
or \U$4417 ( \4732 , \4727 , \4730 , \4731 );
and \U$4418 ( \4733 , \4722 , \4732 );
xor \U$4419 ( \4734 , \4207 , \4261 );
xor \U$4420 ( \4735 , \4734 , \4283 );
and \U$4421 ( \4736 , \4732 , \4735 );
and \U$4422 ( \4737 , \4722 , \4735 );
or \U$4423 ( \4738 , \4733 , \4736 , \4737 );
xor \U$4424 ( \4739 , \4484 , \4494 );
xor \U$4425 ( \4740 , \4739 , \4512 );
xor \U$4426 ( \4741 , \4517 , \4519 );
xor \U$4427 ( \4742 , \4741 , \4522 );
and \U$4428 ( \4743 , \4740 , \4742 );
and \U$4429 ( \4744 , \4738 , \4743 );
xor \U$4430 ( \4745 , \4533 , \4535 );
xor \U$4431 ( \4746 , \4745 , \4538 );
and \U$4432 ( \4747 , \4743 , \4746 );
and \U$4433 ( \4748 , \4738 , \4746 );
or \U$4434 ( \4749 , \4744 , \4747 , \4748 );
xor \U$4435 ( \4750 , \4531 , \4541 );
xor \U$4436 ( \4751 , \4750 , \4544 );
and \U$4437 ( \4752 , \4749 , \4751 );
xor \U$4438 ( \4753 , \4321 , \4331 );
xor \U$4439 ( \4754 , \4753 , \4334 );
and \U$4440 ( \4755 , \4751 , \4754 );
and \U$4441 ( \4756 , \4749 , \4754 );
or \U$4442 ( \4757 , \4752 , \4755 , \4756 );
and \U$4443 ( \4758 , \4553 , \4757 );
xor \U$4444 ( \4759 , \4553 , \4757 );
xor \U$4445 ( \4760 , \4749 , \4751 );
xor \U$4446 ( \4761 , \4760 , \4754 );
and \U$4447 ( \4762 , \4011 , \408 );
and \U$4448 ( \4763 , \3889 , \406 );
nor \U$4449 ( \4764 , \4762 , \4763 );
xnor \U$4450 ( \4765 , \4764 , \378 );
and \U$4451 ( \4766 , \4272 , \360 );
and \U$4452 ( \4767 , \4016 , \358 );
nor \U$4453 ( \4768 , \4766 , \4767 );
xnor \U$4454 ( \4769 , \4768 , \341 );
and \U$4455 ( \4770 , \4765 , \4769 );
buf \U$4456 ( \4771 , RIc0c6690_106);
and \U$4457 ( \4772 , \4771 , \323 );
and \U$4458 ( \4773 , \4469 , \321 );
nor \U$4459 ( \4774 , \4772 , \4773 );
xnor \U$4460 ( \4775 , \4774 , \328 );
and \U$4461 ( \4776 , \4769 , \4775 );
and \U$4462 ( \4777 , \4765 , \4775 );
or \U$4463 ( \4778 , \4770 , \4776 , \4777 );
buf \U$4464 ( \4779 , RIc0c6618_107);
and \U$4465 ( \4780 , \4779 , \317 );
buf \U$4466 ( \4781 , \4780 );
and \U$4467 ( \4782 , \4778 , \4781 );
and \U$4468 ( \4783 , \4771 , \317 );
and \U$4469 ( \4784 , \4781 , \4783 );
and \U$4470 ( \4785 , \4778 , \4783 );
or \U$4471 ( \4786 , \4782 , \4784 , \4785 );
and \U$4472 ( \4787 , \789 , \2596 );
and \U$4473 ( \4788 , \709 , \2594 );
nor \U$4474 ( \4789 , \4787 , \4788 );
xnor \U$4475 ( \4790 , \4789 , \2454 );
and \U$4476 ( \4791 , \925 , \2300 );
and \U$4477 ( \4792 , \863 , \2298 );
nor \U$4478 ( \4793 , \4791 , \4792 );
xnor \U$4479 ( \4794 , \4793 , \2163 );
and \U$4480 ( \4795 , \4790 , \4794 );
and \U$4481 ( \4796 , \1186 , \2094 );
and \U$4482 ( \4797 , \988 , \2092 );
nor \U$4483 ( \4798 , \4796 , \4797 );
xnor \U$4484 ( \4799 , \4798 , \1942 );
and \U$4485 ( \4800 , \4794 , \4799 );
and \U$4486 ( \4801 , \4790 , \4799 );
or \U$4487 ( \4802 , \4795 , \4800 , \4801 );
xor \U$4488 ( \4803 , \4209 , \4570 );
xor \U$4489 ( \4804 , \4570 , \4571 );
not \U$4490 ( \4805 , \4804 );
and \U$4491 ( \4806 , \4803 , \4805 );
and \U$4492 ( \4807 , \316 , \4806 );
not \U$4493 ( \4808 , \4807 );
xnor \U$4494 ( \4809 , \4808 , \4574 );
and \U$4495 ( \4810 , \348 , \4355 );
and \U$4496 ( \4811 , \330 , \4353 );
nor \U$4497 ( \4812 , \4810 , \4811 );
xnor \U$4498 ( \4813 , \4812 , \4212 );
and \U$4499 ( \4814 , \4809 , \4813 );
and \U$4500 ( \4815 , \417 , \4032 );
and \U$4501 ( \4816 , \369 , \4030 );
nor \U$4502 ( \4817 , \4815 , \4816 );
xnor \U$4503 ( \4818 , \4817 , \3786 );
and \U$4504 ( \4819 , \4813 , \4818 );
and \U$4505 ( \4820 , \4809 , \4818 );
or \U$4506 ( \4821 , \4814 , \4819 , \4820 );
and \U$4507 ( \4822 , \4802 , \4821 );
and \U$4508 ( \4823 , \494 , \3637 );
and \U$4509 ( \4824 , \425 , \3635 );
nor \U$4510 ( \4825 , \4823 , \4824 );
xnor \U$4511 ( \4826 , \4825 , \3450 );
and \U$4512 ( \4827 , \553 , \3324 );
and \U$4513 ( \4828 , \499 , \3322 );
nor \U$4514 ( \4829 , \4827 , \4828 );
xnor \U$4515 ( \4830 , \4829 , \3119 );
and \U$4516 ( \4831 , \4826 , \4830 );
and \U$4517 ( \4832 , \681 , \2918 );
and \U$4518 ( \4833 , \604 , \2916 );
nor \U$4519 ( \4834 , \4832 , \4833 );
xnor \U$4520 ( \4835 , \4834 , \2769 );
and \U$4521 ( \4836 , \4830 , \4835 );
and \U$4522 ( \4837 , \4826 , \4835 );
or \U$4523 ( \4838 , \4831 , \4836 , \4837 );
and \U$4524 ( \4839 , \4821 , \4838 );
and \U$4525 ( \4840 , \4802 , \4838 );
or \U$4526 ( \4841 , \4822 , \4839 , \4840 );
and \U$4527 ( \4842 , \4786 , \4841 );
and \U$4528 ( \4843 , \2840 , \692 );
and \U$4529 ( \4844 , \2666 , \690 );
nor \U$4530 ( \4845 , \4843 , \4844 );
xnor \U$4531 ( \4846 , \4845 , \649 );
and \U$4532 ( \4847 , \3145 , \579 );
and \U$4533 ( \4848 , \3007 , \577 );
nor \U$4534 ( \4849 , \4847 , \4848 );
xnor \U$4535 ( \4850 , \4849 , \530 );
and \U$4536 ( \4851 , \4846 , \4850 );
and \U$4537 ( \4852 , \3681 , \478 );
and \U$4538 ( \4853 , \3264 , \476 );
nor \U$4539 ( \4854 , \4852 , \4853 );
xnor \U$4540 ( \4855 , \4854 , \437 );
and \U$4541 ( \4856 , \4850 , \4855 );
and \U$4542 ( \4857 , \4846 , \4855 );
or \U$4543 ( \4858 , \4851 , \4856 , \4857 );
and \U$4544 ( \4859 , \2042 , \1160 );
and \U$4545 ( \4860 , \1799 , \1158 );
nor \U$4546 ( \4861 , \4859 , \4860 );
xnor \U$4547 ( \4862 , \4861 , \1082 );
and \U$4548 ( \4863 , \2233 , \996 );
and \U$4549 ( \4864 , \2047 , \994 );
nor \U$4550 ( \4865 , \4863 , \4864 );
xnor \U$4551 ( \4866 , \4865 , \902 );
and \U$4552 ( \4867 , \4862 , \4866 );
and \U$4553 ( \4868 , \2641 , \826 );
and \U$4554 ( \4869 , \2377 , \824 );
nor \U$4555 ( \4870 , \4868 , \4869 );
xnor \U$4556 ( \4871 , \4870 , \754 );
and \U$4557 ( \4872 , \4866 , \4871 );
and \U$4558 ( \4873 , \4862 , \4871 );
or \U$4559 ( \4874 , \4867 , \4872 , \4873 );
and \U$4560 ( \4875 , \4858 , \4874 );
and \U$4561 ( \4876 , \1379 , \1826 );
and \U$4562 ( \4877 , \1274 , \1824 );
nor \U$4563 ( \4878 , \4876 , \4877 );
xnor \U$4564 ( \4879 , \4878 , \1670 );
and \U$4565 ( \4880 , \1500 , \1554 );
and \U$4566 ( \4881 , \1384 , \1552 );
nor \U$4567 ( \4882 , \4880 , \4881 );
xnor \U$4568 ( \4883 , \4882 , \1441 );
and \U$4569 ( \4884 , \4879 , \4883 );
and \U$4570 ( \4885 , \1791 , \1360 );
and \U$4571 ( \4886 , \1615 , \1358 );
nor \U$4572 ( \4887 , \4885 , \4886 );
xnor \U$4573 ( \4888 , \4887 , \1224 );
and \U$4574 ( \4889 , \4883 , \4888 );
and \U$4575 ( \4890 , \4879 , \4888 );
or \U$4576 ( \4891 , \4884 , \4889 , \4890 );
and \U$4577 ( \4892 , \4874 , \4891 );
and \U$4578 ( \4893 , \4858 , \4891 );
or \U$4579 ( \4894 , \4875 , \4892 , \4893 );
and \U$4580 ( \4895 , \4841 , \4894 );
and \U$4581 ( \4896 , \4786 , \4894 );
or \U$4582 ( \4897 , \4842 , \4895 , \4896 );
xor \U$4583 ( \4898 , \4611 , \4615 );
xor \U$4584 ( \4899 , \4898 , \4620 );
xor \U$4585 ( \4900 , \4644 , \4648 );
xor \U$4586 ( \4901 , \4900 , \4653 );
and \U$4587 ( \4902 , \4899 , \4901 );
xor \U$4588 ( \4903 , \4664 , \4668 );
xor \U$4589 ( \4904 , \4903 , \4673 );
and \U$4590 ( \4905 , \4901 , \4904 );
and \U$4591 ( \4906 , \4899 , \4904 );
or \U$4592 ( \4907 , \4902 , \4905 , \4906 );
xor \U$4593 ( \4908 , \4557 , \4561 );
xor \U$4594 ( \4909 , \4908 , \4566 );
xor \U$4595 ( \4910 , \4627 , \4631 );
xor \U$4596 ( \4911 , \4910 , \4636 );
and \U$4597 ( \4912 , \4909 , \4911 );
xor \U$4598 ( \4913 , \4592 , \4596 );
xor \U$4599 ( \4914 , \4913 , \4601 );
and \U$4600 ( \4915 , \4911 , \4914 );
and \U$4601 ( \4916 , \4909 , \4914 );
or \U$4602 ( \4917 , \4912 , \4915 , \4916 );
and \U$4603 ( \4918 , \4907 , \4917 );
xor \U$4604 ( \4919 , \4694 , \4696 );
xor \U$4605 ( \4920 , \4919 , \4699 );
and \U$4606 ( \4921 , \4917 , \4920 );
and \U$4607 ( \4922 , \4907 , \4920 );
or \U$4608 ( \4923 , \4918 , \4921 , \4922 );
and \U$4609 ( \4924 , \4897 , \4923 );
xor \U$4610 ( \4925 , \4623 , \4639 );
xor \U$4611 ( \4926 , \4925 , \4656 );
xor \U$4612 ( \4927 , \4684 , \4686 );
xor \U$4613 ( \4928 , \4927 , \4689 );
and \U$4614 ( \4929 , \4926 , \4928 );
xnor \U$4615 ( \4930 , \4676 , \4678 );
and \U$4616 ( \4931 , \4928 , \4930 );
and \U$4617 ( \4932 , \4926 , \4930 );
or \U$4618 ( \4933 , \4929 , \4931 , \4932 );
and \U$4619 ( \4934 , \4923 , \4933 );
and \U$4620 ( \4935 , \4897 , \4933 );
or \U$4621 ( \4936 , \4924 , \4934 , \4935 );
xor \U$4622 ( \4937 , \4370 , \4386 );
xor \U$4623 ( \4938 , \4937 , \4403 );
xor \U$4624 ( \4939 , \4422 , \4438 );
xor \U$4625 ( \4940 , \4939 , \4455 );
and \U$4626 ( \4941 , \4938 , \4940 );
xor \U$4627 ( \4942 , \4711 , \4713 );
xor \U$4628 ( \4943 , \4942 , \4716 );
and \U$4629 ( \4944 , \4940 , \4943 );
and \U$4630 ( \4945 , \4938 , \4943 );
or \U$4631 ( \4946 , \4941 , \4944 , \4945 );
and \U$4632 ( \4947 , \4936 , \4946 );
xor \U$4633 ( \4948 , \4724 , \4726 );
xor \U$4634 ( \4949 , \4948 , \4729 );
and \U$4635 ( \4950 , \4946 , \4949 );
and \U$4636 ( \4951 , \4936 , \4949 );
or \U$4637 ( \4952 , \4947 , \4950 , \4951 );
xor \U$4638 ( \4953 , \4722 , \4732 );
xor \U$4639 ( \4954 , \4953 , \4735 );
and \U$4640 ( \4955 , \4952 , \4954 );
xor \U$4641 ( \4956 , \4740 , \4742 );
and \U$4642 ( \4957 , \4954 , \4956 );
and \U$4643 ( \4958 , \4952 , \4956 );
or \U$4644 ( \4959 , \4955 , \4957 , \4958 );
xor \U$4645 ( \4960 , \4515 , \4525 );
xor \U$4646 ( \4961 , \4960 , \4528 );
and \U$4647 ( \4962 , \4959 , \4961 );
xor \U$4648 ( \4963 , \4738 , \4743 );
xor \U$4649 ( \4964 , \4963 , \4746 );
and \U$4650 ( \4965 , \4961 , \4964 );
and \U$4651 ( \4966 , \4959 , \4964 );
or \U$4652 ( \4967 , \4962 , \4965 , \4966 );
and \U$4653 ( \4968 , \4761 , \4967 );
xor \U$4654 ( \4969 , \4761 , \4967 );
xor \U$4655 ( \4970 , \4959 , \4961 );
xor \U$4656 ( \4971 , \4970 , \4964 );
and \U$4657 ( \4972 , \709 , \2918 );
and \U$4658 ( \4973 , \681 , \2916 );
nor \U$4659 ( \4974 , \4972 , \4973 );
xnor \U$4660 ( \4975 , \4974 , \2769 );
and \U$4661 ( \4976 , \863 , \2596 );
and \U$4662 ( \4977 , \789 , \2594 );
nor \U$4663 ( \4978 , \4976 , \4977 );
xnor \U$4664 ( \4979 , \4978 , \2454 );
and \U$4665 ( \4980 , \4975 , \4979 );
and \U$4666 ( \4981 , \988 , \2300 );
and \U$4667 ( \4982 , \925 , \2298 );
nor \U$4668 ( \4983 , \4981 , \4982 );
xnor \U$4669 ( \4984 , \4983 , \2163 );
and \U$4670 ( \4985 , \4979 , \4984 );
and \U$4671 ( \4986 , \4975 , \4984 );
or \U$4672 ( \4987 , \4980 , \4985 , \4986 );
buf \U$4673 ( \4988 , RIc0c8328_45);
buf \U$4674 ( \4989 , RIc0c82b0_46);
and \U$4675 ( \4990 , \4988 , \4989 );
not \U$4676 ( \4991 , \4990 );
and \U$4677 ( \4992 , \4571 , \4991 );
not \U$4678 ( \4993 , \4992 );
and \U$4679 ( \4994 , \330 , \4806 );
and \U$4680 ( \4995 , \316 , \4804 );
nor \U$4681 ( \4996 , \4994 , \4995 );
xnor \U$4682 ( \4997 , \4996 , \4574 );
and \U$4683 ( \4998 , \4993 , \4997 );
and \U$4684 ( \4999 , \369 , \4355 );
and \U$4685 ( \5000 , \348 , \4353 );
nor \U$4686 ( \5001 , \4999 , \5000 );
xnor \U$4687 ( \5002 , \5001 , \4212 );
and \U$4688 ( \5003 , \4997 , \5002 );
and \U$4689 ( \5004 , \4993 , \5002 );
or \U$4690 ( \5005 , \4998 , \5003 , \5004 );
and \U$4691 ( \5006 , \4987 , \5005 );
and \U$4692 ( \5007 , \425 , \4032 );
and \U$4693 ( \5008 , \417 , \4030 );
nor \U$4694 ( \5009 , \5007 , \5008 );
xnor \U$4695 ( \5010 , \5009 , \3786 );
and \U$4696 ( \5011 , \499 , \3637 );
and \U$4697 ( \5012 , \494 , \3635 );
nor \U$4698 ( \5013 , \5011 , \5012 );
xnor \U$4699 ( \5014 , \5013 , \3450 );
and \U$4700 ( \5015 , \5010 , \5014 );
and \U$4701 ( \5016 , \604 , \3324 );
and \U$4702 ( \5017 , \553 , \3322 );
nor \U$4703 ( \5018 , \5016 , \5017 );
xnor \U$4704 ( \5019 , \5018 , \3119 );
and \U$4705 ( \5020 , \5014 , \5019 );
and \U$4706 ( \5021 , \5010 , \5019 );
or \U$4707 ( \5022 , \5015 , \5020 , \5021 );
and \U$4708 ( \5023 , \5005 , \5022 );
and \U$4709 ( \5024 , \4987 , \5022 );
or \U$4710 ( \5025 , \5006 , \5023 , \5024 );
and \U$4711 ( \5026 , \1274 , \2094 );
and \U$4712 ( \5027 , \1186 , \2092 );
nor \U$4713 ( \5028 , \5026 , \5027 );
xnor \U$4714 ( \5029 , \5028 , \1942 );
and \U$4715 ( \5030 , \1384 , \1826 );
and \U$4716 ( \5031 , \1379 , \1824 );
nor \U$4717 ( \5032 , \5030 , \5031 );
xnor \U$4718 ( \5033 , \5032 , \1670 );
and \U$4719 ( \5034 , \5029 , \5033 );
and \U$4720 ( \5035 , \1615 , \1554 );
and \U$4721 ( \5036 , \1500 , \1552 );
nor \U$4722 ( \5037 , \5035 , \5036 );
xnor \U$4723 ( \5038 , \5037 , \1441 );
and \U$4724 ( \5039 , \5033 , \5038 );
and \U$4725 ( \5040 , \5029 , \5038 );
or \U$4726 ( \5041 , \5034 , \5039 , \5040 );
and \U$4727 ( \5042 , \2666 , \826 );
and \U$4728 ( \5043 , \2641 , \824 );
nor \U$4729 ( \5044 , \5042 , \5043 );
xnor \U$4730 ( \5045 , \5044 , \754 );
and \U$4731 ( \5046 , \3007 , \692 );
and \U$4732 ( \5047 , \2840 , \690 );
nor \U$4733 ( \5048 , \5046 , \5047 );
xnor \U$4734 ( \5049 , \5048 , \649 );
and \U$4735 ( \5050 , \5045 , \5049 );
and \U$4736 ( \5051 , \3264 , \579 );
and \U$4737 ( \5052 , \3145 , \577 );
nor \U$4738 ( \5053 , \5051 , \5052 );
xnor \U$4739 ( \5054 , \5053 , \530 );
and \U$4740 ( \5055 , \5049 , \5054 );
and \U$4741 ( \5056 , \5045 , \5054 );
or \U$4742 ( \5057 , \5050 , \5055 , \5056 );
and \U$4743 ( \5058 , \5041 , \5057 );
and \U$4744 ( \5059 , \1799 , \1360 );
and \U$4745 ( \5060 , \1791 , \1358 );
nor \U$4746 ( \5061 , \5059 , \5060 );
xnor \U$4747 ( \5062 , \5061 , \1224 );
and \U$4748 ( \5063 , \2047 , \1160 );
and \U$4749 ( \5064 , \2042 , \1158 );
nor \U$4750 ( \5065 , \5063 , \5064 );
xnor \U$4751 ( \5066 , \5065 , \1082 );
and \U$4752 ( \5067 , \5062 , \5066 );
and \U$4753 ( \5068 , \2377 , \996 );
and \U$4754 ( \5069 , \2233 , \994 );
nor \U$4755 ( \5070 , \5068 , \5069 );
xnor \U$4756 ( \5071 , \5070 , \902 );
and \U$4757 ( \5072 , \5066 , \5071 );
and \U$4758 ( \5073 , \5062 , \5071 );
or \U$4759 ( \5074 , \5067 , \5072 , \5073 );
and \U$4760 ( \5075 , \5057 , \5074 );
and \U$4761 ( \5076 , \5041 , \5074 );
or \U$4762 ( \5077 , \5058 , \5075 , \5076 );
and \U$4763 ( \5078 , \5025 , \5077 );
and \U$4764 ( \5079 , \3889 , \478 );
and \U$4765 ( \5080 , \3681 , \476 );
nor \U$4766 ( \5081 , \5079 , \5080 );
xnor \U$4767 ( \5082 , \5081 , \437 );
and \U$4768 ( \5083 , \4016 , \408 );
and \U$4769 ( \5084 , \4011 , \406 );
nor \U$4770 ( \5085 , \5083 , \5084 );
xnor \U$4771 ( \5086 , \5085 , \378 );
and \U$4772 ( \5087 , \5082 , \5086 );
and \U$4773 ( \5088 , \4469 , \360 );
and \U$4774 ( \5089 , \4272 , \358 );
nor \U$4775 ( \5090 , \5088 , \5089 );
xnor \U$4776 ( \5091 , \5090 , \341 );
and \U$4777 ( \5092 , \5086 , \5091 );
and \U$4778 ( \5093 , \5082 , \5091 );
or \U$4779 ( \5094 , \5087 , \5092 , \5093 );
xor \U$4780 ( \5095 , \4765 , \4769 );
xor \U$4781 ( \5096 , \5095 , \4775 );
and \U$4782 ( \5097 , \5094 , \5096 );
not \U$4783 ( \5098 , \4780 );
and \U$4784 ( \5099 , \5096 , \5098 );
and \U$4785 ( \5100 , \5094 , \5098 );
or \U$4786 ( \5101 , \5097 , \5099 , \5100 );
and \U$4787 ( \5102 , \5077 , \5101 );
and \U$4788 ( \5103 , \5025 , \5101 );
or \U$4789 ( \5104 , \5078 , \5102 , \5103 );
xor \U$4790 ( \5105 , \4846 , \4850 );
xor \U$4791 ( \5106 , \5105 , \4855 );
xor \U$4792 ( \5107 , \4862 , \4866 );
xor \U$4793 ( \5108 , \5107 , \4871 );
and \U$4794 ( \5109 , \5106 , \5108 );
xor \U$4795 ( \5110 , \4879 , \4883 );
xor \U$4796 ( \5111 , \5110 , \4888 );
and \U$4797 ( \5112 , \5108 , \5111 );
and \U$4798 ( \5113 , \5106 , \5111 );
or \U$4799 ( \5114 , \5109 , \5112 , \5113 );
xor \U$4800 ( \5115 , \4790 , \4794 );
xor \U$4801 ( \5116 , \5115 , \4799 );
xor \U$4802 ( \5117 , \4809 , \4813 );
xor \U$4803 ( \5118 , \5117 , \4818 );
and \U$4804 ( \5119 , \5116 , \5118 );
xor \U$4805 ( \5120 , \4826 , \4830 );
xor \U$4806 ( \5121 , \5120 , \4835 );
and \U$4807 ( \5122 , \5118 , \5121 );
and \U$4808 ( \5123 , \5116 , \5121 );
or \U$4809 ( \5124 , \5119 , \5122 , \5123 );
and \U$4810 ( \5125 , \5114 , \5124 );
xor \U$4811 ( \5126 , \4575 , \4579 );
xor \U$4812 ( \5127 , \5126 , \4584 );
and \U$4813 ( \5128 , \5124 , \5127 );
and \U$4814 ( \5129 , \5114 , \5127 );
or \U$4815 ( \5130 , \5125 , \5128 , \5129 );
and \U$4816 ( \5131 , \5104 , \5130 );
xor \U$4817 ( \5132 , \4778 , \4781 );
xor \U$4818 ( \5133 , \5132 , \4783 );
xor \U$4819 ( \5134 , \4899 , \4901 );
xor \U$4820 ( \5135 , \5134 , \4904 );
and \U$4821 ( \5136 , \5133 , \5135 );
xor \U$4822 ( \5137 , \4909 , \4911 );
xor \U$4823 ( \5138 , \5137 , \4914 );
and \U$4824 ( \5139 , \5135 , \5138 );
and \U$4825 ( \5140 , \5133 , \5138 );
or \U$4826 ( \5141 , \5136 , \5139 , \5140 );
and \U$4827 ( \5142 , \5130 , \5141 );
and \U$4828 ( \5143 , \5104 , \5141 );
or \U$4829 ( \5144 , \5131 , \5142 , \5143 );
xor \U$4830 ( \5145 , \4569 , \4587 );
xor \U$4831 ( \5146 , \5145 , \4604 );
xor \U$4832 ( \5147 , \4907 , \4917 );
xor \U$4833 ( \5148 , \5147 , \4920 );
and \U$4834 ( \5149 , \5146 , \5148 );
xor \U$4835 ( \5150 , \4926 , \4928 );
xor \U$4836 ( \5151 , \5150 , \4930 );
and \U$4837 ( \5152 , \5148 , \5151 );
and \U$4838 ( \5153 , \5146 , \5151 );
or \U$4839 ( \5154 , \5149 , \5152 , \5153 );
and \U$4840 ( \5155 , \5144 , \5154 );
xor \U$4841 ( \5156 , \4692 , \4702 );
xor \U$4842 ( \5157 , \5156 , \4705 );
and \U$4843 ( \5158 , \5154 , \5157 );
and \U$4844 ( \5159 , \5144 , \5157 );
or \U$4845 ( \5160 , \5155 , \5158 , \5159 );
xor \U$4846 ( \5161 , \4607 , \4659 );
xor \U$4847 ( \5162 , \5161 , \4679 );
xor \U$4848 ( \5163 , \4897 , \4923 );
xor \U$4849 ( \5164 , \5163 , \4933 );
and \U$4850 ( \5165 , \5162 , \5164 );
xor \U$4851 ( \5166 , \4938 , \4940 );
xor \U$4852 ( \5167 , \5166 , \4943 );
and \U$4853 ( \5168 , \5164 , \5167 );
and \U$4854 ( \5169 , \5162 , \5167 );
or \U$4855 ( \5170 , \5165 , \5168 , \5169 );
and \U$4856 ( \5171 , \5160 , \5170 );
xor \U$4857 ( \5172 , \4682 , \4708 );
xor \U$4858 ( \5173 , \5172 , \4719 );
and \U$4859 ( \5174 , \5170 , \5173 );
and \U$4860 ( \5175 , \5160 , \5173 );
or \U$4861 ( \5176 , \5171 , \5174 , \5175 );
xor \U$4862 ( \5177 , \4571 , \4988 );
xor \U$4863 ( \5178 , \4988 , \4989 );
not \U$4864 ( \5179 , \5178 );
and \U$4865 ( \5180 , \5177 , \5179 );
and \U$4866 ( \5181 , \316 , \5180 );
not \U$4867 ( \5182 , \5181 );
xnor \U$4868 ( \5183 , \5182 , \4992 );
and \U$4869 ( \5184 , \348 , \4806 );
and \U$4870 ( \5185 , \330 , \4804 );
nor \U$4871 ( \5186 , \5184 , \5185 );
xnor \U$4872 ( \5187 , \5186 , \4574 );
and \U$4873 ( \5188 , \5183 , \5187 );
and \U$4874 ( \5189 , \417 , \4355 );
and \U$4875 ( \5190 , \369 , \4353 );
nor \U$4876 ( \5191 , \5189 , \5190 );
xnor \U$4877 ( \5192 , \5191 , \4212 );
and \U$4878 ( \5193 , \5187 , \5192 );
and \U$4879 ( \5194 , \5183 , \5192 );
or \U$4880 ( \5195 , \5188 , \5193 , \5194 );
and \U$4881 ( \5196 , \789 , \2918 );
and \U$4882 ( \5197 , \709 , \2916 );
nor \U$4883 ( \5198 , \5196 , \5197 );
xnor \U$4884 ( \5199 , \5198 , \2769 );
and \U$4885 ( \5200 , \925 , \2596 );
and \U$4886 ( \5201 , \863 , \2594 );
nor \U$4887 ( \5202 , \5200 , \5201 );
xnor \U$4888 ( \5203 , \5202 , \2454 );
and \U$4889 ( \5204 , \5199 , \5203 );
and \U$4890 ( \5205 , \1186 , \2300 );
and \U$4891 ( \5206 , \988 , \2298 );
nor \U$4892 ( \5207 , \5205 , \5206 );
xnor \U$4893 ( \5208 , \5207 , \2163 );
and \U$4894 ( \5209 , \5203 , \5208 );
and \U$4895 ( \5210 , \5199 , \5208 );
or \U$4896 ( \5211 , \5204 , \5209 , \5210 );
and \U$4897 ( \5212 , \5195 , \5211 );
and \U$4898 ( \5213 , \494 , \4032 );
and \U$4899 ( \5214 , \425 , \4030 );
nor \U$4900 ( \5215 , \5213 , \5214 );
xnor \U$4901 ( \5216 , \5215 , \3786 );
and \U$4902 ( \5217 , \553 , \3637 );
and \U$4903 ( \5218 , \499 , \3635 );
nor \U$4904 ( \5219 , \5217 , \5218 );
xnor \U$4905 ( \5220 , \5219 , \3450 );
and \U$4906 ( \5221 , \5216 , \5220 );
and \U$4907 ( \5222 , \681 , \3324 );
and \U$4908 ( \5223 , \604 , \3322 );
nor \U$4909 ( \5224 , \5222 , \5223 );
xnor \U$4910 ( \5225 , \5224 , \3119 );
and \U$4911 ( \5226 , \5220 , \5225 );
and \U$4912 ( \5227 , \5216 , \5225 );
or \U$4913 ( \5228 , \5221 , \5226 , \5227 );
and \U$4914 ( \5229 , \5211 , \5228 );
and \U$4915 ( \5230 , \5195 , \5228 );
or \U$4916 ( \5231 , \5212 , \5229 , \5230 );
and \U$4917 ( \5232 , \4011 , \478 );
and \U$4918 ( \5233 , \3889 , \476 );
nor \U$4919 ( \5234 , \5232 , \5233 );
xnor \U$4920 ( \5235 , \5234 , \437 );
and \U$4921 ( \5236 , \4272 , \408 );
and \U$4922 ( \5237 , \4016 , \406 );
nor \U$4923 ( \5238 , \5236 , \5237 );
xnor \U$4924 ( \5239 , \5238 , \378 );
and \U$4925 ( \5240 , \5235 , \5239 );
and \U$4926 ( \5241 , \4771 , \360 );
and \U$4927 ( \5242 , \4469 , \358 );
nor \U$4928 ( \5243 , \5241 , \5242 );
xnor \U$4929 ( \5244 , \5243 , \341 );
and \U$4930 ( \5245 , \5239 , \5244 );
and \U$4931 ( \5246 , \5235 , \5244 );
or \U$4932 ( \5247 , \5240 , \5245 , \5246 );
buf \U$4933 ( \5248 , RIc0c65a0_108);
and \U$4934 ( \5249 , \5248 , \323 );
and \U$4935 ( \5250 , \4779 , \321 );
nor \U$4936 ( \5251 , \5249 , \5250 );
xnor \U$4937 ( \5252 , \5251 , \328 );
buf \U$4938 ( \5253 , RIc0c6528_109);
and \U$4939 ( \5254 , \5253 , \317 );
or \U$4940 ( \5255 , \5252 , \5254 );
and \U$4941 ( \5256 , \5247 , \5255 );
and \U$4942 ( \5257 , \4779 , \323 );
and \U$4943 ( \5258 , \4771 , \321 );
nor \U$4944 ( \5259 , \5257 , \5258 );
xnor \U$4945 ( \5260 , \5259 , \328 );
and \U$4946 ( \5261 , \5255 , \5260 );
and \U$4947 ( \5262 , \5247 , \5260 );
or \U$4948 ( \5263 , \5256 , \5261 , \5262 );
and \U$4949 ( \5264 , \5231 , \5263 );
and \U$4950 ( \5265 , \1379 , \2094 );
and \U$4951 ( \5266 , \1274 , \2092 );
nor \U$4952 ( \5267 , \5265 , \5266 );
xnor \U$4953 ( \5268 , \5267 , \1942 );
and \U$4954 ( \5269 , \1500 , \1826 );
and \U$4955 ( \5270 , \1384 , \1824 );
nor \U$4956 ( \5271 , \5269 , \5270 );
xnor \U$4957 ( \5272 , \5271 , \1670 );
and \U$4958 ( \5273 , \5268 , \5272 );
and \U$4959 ( \5274 , \1791 , \1554 );
and \U$4960 ( \5275 , \1615 , \1552 );
nor \U$4961 ( \5276 , \5274 , \5275 );
xnor \U$4962 ( \5277 , \5276 , \1441 );
and \U$4963 ( \5278 , \5272 , \5277 );
and \U$4964 ( \5279 , \5268 , \5277 );
or \U$4965 ( \5280 , \5273 , \5278 , \5279 );
and \U$4966 ( \5281 , \2042 , \1360 );
and \U$4967 ( \5282 , \1799 , \1358 );
nor \U$4968 ( \5283 , \5281 , \5282 );
xnor \U$4969 ( \5284 , \5283 , \1224 );
and \U$4970 ( \5285 , \2233 , \1160 );
and \U$4971 ( \5286 , \2047 , \1158 );
nor \U$4972 ( \5287 , \5285 , \5286 );
xnor \U$4973 ( \5288 , \5287 , \1082 );
and \U$4974 ( \5289 , \5284 , \5288 );
and \U$4975 ( \5290 , \2641 , \996 );
and \U$4976 ( \5291 , \2377 , \994 );
nor \U$4977 ( \5292 , \5290 , \5291 );
xnor \U$4978 ( \5293 , \5292 , \902 );
and \U$4979 ( \5294 , \5288 , \5293 );
and \U$4980 ( \5295 , \5284 , \5293 );
or \U$4981 ( \5296 , \5289 , \5294 , \5295 );
and \U$4982 ( \5297 , \5280 , \5296 );
and \U$4983 ( \5298 , \2840 , \826 );
and \U$4984 ( \5299 , \2666 , \824 );
nor \U$4985 ( \5300 , \5298 , \5299 );
xnor \U$4986 ( \5301 , \5300 , \754 );
and \U$4987 ( \5302 , \3145 , \692 );
and \U$4988 ( \5303 , \3007 , \690 );
nor \U$4989 ( \5304 , \5302 , \5303 );
xnor \U$4990 ( \5305 , \5304 , \649 );
and \U$4991 ( \5306 , \5301 , \5305 );
and \U$4992 ( \5307 , \3681 , \579 );
and \U$4993 ( \5308 , \3264 , \577 );
nor \U$4994 ( \5309 , \5307 , \5308 );
xnor \U$4995 ( \5310 , \5309 , \530 );
and \U$4996 ( \5311 , \5305 , \5310 );
and \U$4997 ( \5312 , \5301 , \5310 );
or \U$4998 ( \5313 , \5306 , \5311 , \5312 );
and \U$4999 ( \5314 , \5296 , \5313 );
and \U$5000 ( \5315 , \5280 , \5313 );
or \U$5001 ( \5316 , \5297 , \5314 , \5315 );
and \U$5002 ( \5317 , \5263 , \5316 );
and \U$5003 ( \5318 , \5231 , \5316 );
or \U$5004 ( \5319 , \5264 , \5317 , \5318 );
and \U$5005 ( \5320 , \5248 , \317 );
xor \U$5006 ( \5321 , \5082 , \5086 );
xor \U$5007 ( \5322 , \5321 , \5091 );
and \U$5008 ( \5323 , \5320 , \5322 );
xor \U$5009 ( \5324 , \5045 , \5049 );
xor \U$5010 ( \5325 , \5324 , \5054 );
and \U$5011 ( \5326 , \5322 , \5325 );
and \U$5012 ( \5327 , \5320 , \5325 );
or \U$5013 ( \5328 , \5323 , \5326 , \5327 );
xor \U$5014 ( \5329 , \5029 , \5033 );
xor \U$5015 ( \5330 , \5329 , \5038 );
xor \U$5016 ( \5331 , \4975 , \4979 );
xor \U$5017 ( \5332 , \5331 , \4984 );
and \U$5018 ( \5333 , \5330 , \5332 );
xor \U$5019 ( \5334 , \5062 , \5066 );
xor \U$5020 ( \5335 , \5334 , \5071 );
and \U$5021 ( \5336 , \5332 , \5335 );
and \U$5022 ( \5337 , \5330 , \5335 );
or \U$5023 ( \5338 , \5333 , \5336 , \5337 );
and \U$5024 ( \5339 , \5328 , \5338 );
xor \U$5025 ( \5340 , \5116 , \5118 );
xor \U$5026 ( \5341 , \5340 , \5121 );
and \U$5027 ( \5342 , \5338 , \5341 );
and \U$5028 ( \5343 , \5328 , \5341 );
or \U$5029 ( \5344 , \5339 , \5342 , \5343 );
and \U$5030 ( \5345 , \5319 , \5344 );
xor \U$5031 ( \5346 , \5041 , \5057 );
xor \U$5032 ( \5347 , \5346 , \5074 );
xor \U$5033 ( \5348 , \5106 , \5108 );
xor \U$5034 ( \5349 , \5348 , \5111 );
and \U$5035 ( \5350 , \5347 , \5349 );
xor \U$5036 ( \5351 , \5094 , \5096 );
xor \U$5037 ( \5352 , \5351 , \5098 );
and \U$5038 ( \5353 , \5349 , \5352 );
and \U$5039 ( \5354 , \5347 , \5352 );
or \U$5040 ( \5355 , \5350 , \5353 , \5354 );
and \U$5041 ( \5356 , \5344 , \5355 );
and \U$5042 ( \5357 , \5319 , \5355 );
or \U$5043 ( \5358 , \5345 , \5356 , \5357 );
xor \U$5044 ( \5359 , \4802 , \4821 );
xor \U$5045 ( \5360 , \5359 , \4838 );
xor \U$5046 ( \5361 , \4858 , \4874 );
xor \U$5047 ( \5362 , \5361 , \4891 );
and \U$5048 ( \5363 , \5360 , \5362 );
xor \U$5049 ( \5364 , \5133 , \5135 );
xor \U$5050 ( \5365 , \5364 , \5138 );
and \U$5051 ( \5366 , \5362 , \5365 );
and \U$5052 ( \5367 , \5360 , \5365 );
or \U$5053 ( \5368 , \5363 , \5366 , \5367 );
and \U$5054 ( \5369 , \5358 , \5368 );
xor \U$5055 ( \5370 , \4786 , \4841 );
xor \U$5056 ( \5371 , \5370 , \4894 );
and \U$5057 ( \5372 , \5368 , \5371 );
and \U$5058 ( \5373 , \5358 , \5371 );
or \U$5059 ( \5374 , \5369 , \5372 , \5373 );
xor \U$5060 ( \5375 , \5144 , \5154 );
xor \U$5061 ( \5376 , \5375 , \5157 );
and \U$5062 ( \5377 , \5374 , \5376 );
xor \U$5063 ( \5378 , \5162 , \5164 );
xor \U$5064 ( \5379 , \5378 , \5167 );
and \U$5065 ( \5380 , \5376 , \5379 );
and \U$5066 ( \5381 , \5374 , \5379 );
or \U$5067 ( \5382 , \5377 , \5380 , \5381 );
xor \U$5068 ( \5383 , \5160 , \5170 );
xor \U$5069 ( \5384 , \5383 , \5173 );
and \U$5070 ( \5385 , \5382 , \5384 );
xor \U$5071 ( \5386 , \4936 , \4946 );
xor \U$5072 ( \5387 , \5386 , \4949 );
and \U$5073 ( \5388 , \5384 , \5387 );
and \U$5074 ( \5389 , \5382 , \5387 );
or \U$5075 ( \5390 , \5385 , \5388 , \5389 );
and \U$5076 ( \5391 , \5176 , \5390 );
xor \U$5077 ( \5392 , \4952 , \4954 );
xor \U$5078 ( \5393 , \5392 , \4956 );
and \U$5079 ( \5394 , \5390 , \5393 );
and \U$5080 ( \5395 , \5176 , \5393 );
or \U$5081 ( \5396 , \5391 , \5394 , \5395 );
and \U$5082 ( \5397 , \4971 , \5396 );
xor \U$5083 ( \5398 , \4971 , \5396 );
xor \U$5084 ( \5399 , \5176 , \5390 );
xor \U$5085 ( \5400 , \5399 , \5393 );
buf \U$5086 ( \5401 , RIc0c8238_47);
buf \U$5087 ( \5402 , RIc0c81c0_48);
and \U$5088 ( \5403 , \5401 , \5402 );
not \U$5089 ( \5404 , \5403 );
and \U$5090 ( \5405 , \4989 , \5404 );
not \U$5091 ( \5406 , \5405 );
and \U$5092 ( \5407 , \330 , \5180 );
and \U$5093 ( \5408 , \316 , \5178 );
nor \U$5094 ( \5409 , \5407 , \5408 );
xnor \U$5095 ( \5410 , \5409 , \4992 );
and \U$5096 ( \5411 , \5406 , \5410 );
and \U$5097 ( \5412 , \369 , \4806 );
and \U$5098 ( \5413 , \348 , \4804 );
nor \U$5099 ( \5414 , \5412 , \5413 );
xnor \U$5100 ( \5415 , \5414 , \4574 );
and \U$5101 ( \5416 , \5410 , \5415 );
and \U$5102 ( \5417 , \5406 , \5415 );
or \U$5103 ( \5418 , \5411 , \5416 , \5417 );
and \U$5104 ( \5419 , \425 , \4355 );
and \U$5105 ( \5420 , \417 , \4353 );
nor \U$5106 ( \5421 , \5419 , \5420 );
xnor \U$5107 ( \5422 , \5421 , \4212 );
and \U$5108 ( \5423 , \499 , \4032 );
and \U$5109 ( \5424 , \494 , \4030 );
nor \U$5110 ( \5425 , \5423 , \5424 );
xnor \U$5111 ( \5426 , \5425 , \3786 );
and \U$5112 ( \5427 , \5422 , \5426 );
and \U$5113 ( \5428 , \604 , \3637 );
and \U$5114 ( \5429 , \553 , \3635 );
nor \U$5115 ( \5430 , \5428 , \5429 );
xnor \U$5116 ( \5431 , \5430 , \3450 );
and \U$5117 ( \5432 , \5426 , \5431 );
and \U$5118 ( \5433 , \5422 , \5431 );
or \U$5119 ( \5434 , \5427 , \5432 , \5433 );
and \U$5120 ( \5435 , \5418 , \5434 );
and \U$5121 ( \5436 , \709 , \3324 );
and \U$5122 ( \5437 , \681 , \3322 );
nor \U$5123 ( \5438 , \5436 , \5437 );
xnor \U$5124 ( \5439 , \5438 , \3119 );
and \U$5125 ( \5440 , \863 , \2918 );
and \U$5126 ( \5441 , \789 , \2916 );
nor \U$5127 ( \5442 , \5440 , \5441 );
xnor \U$5128 ( \5443 , \5442 , \2769 );
and \U$5129 ( \5444 , \5439 , \5443 );
and \U$5130 ( \5445 , \988 , \2596 );
and \U$5131 ( \5446 , \925 , \2594 );
nor \U$5132 ( \5447 , \5445 , \5446 );
xnor \U$5133 ( \5448 , \5447 , \2454 );
and \U$5134 ( \5449 , \5443 , \5448 );
and \U$5135 ( \5450 , \5439 , \5448 );
or \U$5136 ( \5451 , \5444 , \5449 , \5450 );
and \U$5137 ( \5452 , \5434 , \5451 );
and \U$5138 ( \5453 , \5418 , \5451 );
or \U$5139 ( \5454 , \5435 , \5452 , \5453 );
and \U$5140 ( \5455 , \1274 , \2300 );
and \U$5141 ( \5456 , \1186 , \2298 );
nor \U$5142 ( \5457 , \5455 , \5456 );
xnor \U$5143 ( \5458 , \5457 , \2163 );
and \U$5144 ( \5459 , \1384 , \2094 );
and \U$5145 ( \5460 , \1379 , \2092 );
nor \U$5146 ( \5461 , \5459 , \5460 );
xnor \U$5147 ( \5462 , \5461 , \1942 );
and \U$5148 ( \5463 , \5458 , \5462 );
and \U$5149 ( \5464 , \1615 , \1826 );
and \U$5150 ( \5465 , \1500 , \1824 );
nor \U$5151 ( \5466 , \5464 , \5465 );
xnor \U$5152 ( \5467 , \5466 , \1670 );
and \U$5153 ( \5468 , \5462 , \5467 );
and \U$5154 ( \5469 , \5458 , \5467 );
or \U$5155 ( \5470 , \5463 , \5468 , \5469 );
and \U$5156 ( \5471 , \1799 , \1554 );
and \U$5157 ( \5472 , \1791 , \1552 );
nor \U$5158 ( \5473 , \5471 , \5472 );
xnor \U$5159 ( \5474 , \5473 , \1441 );
and \U$5160 ( \5475 , \2047 , \1360 );
and \U$5161 ( \5476 , \2042 , \1358 );
nor \U$5162 ( \5477 , \5475 , \5476 );
xnor \U$5163 ( \5478 , \5477 , \1224 );
and \U$5164 ( \5479 , \5474 , \5478 );
and \U$5165 ( \5480 , \2377 , \1160 );
and \U$5166 ( \5481 , \2233 , \1158 );
nor \U$5167 ( \5482 , \5480 , \5481 );
xnor \U$5168 ( \5483 , \5482 , \1082 );
and \U$5169 ( \5484 , \5478 , \5483 );
and \U$5170 ( \5485 , \5474 , \5483 );
or \U$5171 ( \5486 , \5479 , \5484 , \5485 );
and \U$5172 ( \5487 , \5470 , \5486 );
and \U$5173 ( \5488 , \2666 , \996 );
and \U$5174 ( \5489 , \2641 , \994 );
nor \U$5175 ( \5490 , \5488 , \5489 );
xnor \U$5176 ( \5491 , \5490 , \902 );
and \U$5177 ( \5492 , \3007 , \826 );
and \U$5178 ( \5493 , \2840 , \824 );
nor \U$5179 ( \5494 , \5492 , \5493 );
xnor \U$5180 ( \5495 , \5494 , \754 );
and \U$5181 ( \5496 , \5491 , \5495 );
and \U$5182 ( \5497 , \3264 , \692 );
and \U$5183 ( \5498 , \3145 , \690 );
nor \U$5184 ( \5499 , \5497 , \5498 );
xnor \U$5185 ( \5500 , \5499 , \649 );
and \U$5186 ( \5501 , \5495 , \5500 );
and \U$5187 ( \5502 , \5491 , \5500 );
or \U$5188 ( \5503 , \5496 , \5501 , \5502 );
and \U$5189 ( \5504 , \5486 , \5503 );
and \U$5190 ( \5505 , \5470 , \5503 );
or \U$5191 ( \5506 , \5487 , \5504 , \5505 );
and \U$5192 ( \5507 , \5454 , \5506 );
and \U$5193 ( \5508 , \4779 , \360 );
and \U$5194 ( \5509 , \4771 , \358 );
nor \U$5195 ( \5510 , \5508 , \5509 );
xnor \U$5196 ( \5511 , \5510 , \341 );
and \U$5197 ( \5512 , \5253 , \323 );
and \U$5198 ( \5513 , \5248 , \321 );
nor \U$5199 ( \5514 , \5512 , \5513 );
xnor \U$5200 ( \5515 , \5514 , \328 );
and \U$5201 ( \5516 , \5511 , \5515 );
buf \U$5202 ( \5517 , RIc0c64b0_110);
and \U$5203 ( \5518 , \5517 , \317 );
and \U$5204 ( \5519 , \5515 , \5518 );
and \U$5205 ( \5520 , \5511 , \5518 );
or \U$5206 ( \5521 , \5516 , \5519 , \5520 );
and \U$5207 ( \5522 , \3889 , \579 );
and \U$5208 ( \5523 , \3681 , \577 );
nor \U$5209 ( \5524 , \5522 , \5523 );
xnor \U$5210 ( \5525 , \5524 , \530 );
and \U$5211 ( \5526 , \4016 , \478 );
and \U$5212 ( \5527 , \4011 , \476 );
nor \U$5213 ( \5528 , \5526 , \5527 );
xnor \U$5214 ( \5529 , \5528 , \437 );
and \U$5215 ( \5530 , \5525 , \5529 );
and \U$5216 ( \5531 , \4469 , \408 );
and \U$5217 ( \5532 , \4272 , \406 );
nor \U$5218 ( \5533 , \5531 , \5532 );
xnor \U$5219 ( \5534 , \5533 , \378 );
and \U$5220 ( \5535 , \5529 , \5534 );
and \U$5221 ( \5536 , \5525 , \5534 );
or \U$5222 ( \5537 , \5530 , \5535 , \5536 );
and \U$5223 ( \5538 , \5521 , \5537 );
xnor \U$5224 ( \5539 , \5252 , \5254 );
and \U$5225 ( \5540 , \5537 , \5539 );
and \U$5226 ( \5541 , \5521 , \5539 );
or \U$5227 ( \5542 , \5538 , \5540 , \5541 );
and \U$5228 ( \5543 , \5506 , \5542 );
and \U$5229 ( \5544 , \5454 , \5542 );
or \U$5230 ( \5545 , \5507 , \5543 , \5544 );
xor \U$5231 ( \5546 , \5235 , \5239 );
xor \U$5232 ( \5547 , \5546 , \5244 );
xor \U$5233 ( \5548 , \5284 , \5288 );
xor \U$5234 ( \5549 , \5548 , \5293 );
and \U$5235 ( \5550 , \5547 , \5549 );
xor \U$5236 ( \5551 , \5301 , \5305 );
xor \U$5237 ( \5552 , \5551 , \5310 );
and \U$5238 ( \5553 , \5549 , \5552 );
and \U$5239 ( \5554 , \5547 , \5552 );
or \U$5240 ( \5555 , \5550 , \5553 , \5554 );
xor \U$5241 ( \5556 , \5268 , \5272 );
xor \U$5242 ( \5557 , \5556 , \5277 );
xor \U$5243 ( \5558 , \5199 , \5203 );
xor \U$5244 ( \5559 , \5558 , \5208 );
and \U$5245 ( \5560 , \5557 , \5559 );
xor \U$5246 ( \5561 , \5216 , \5220 );
xor \U$5247 ( \5562 , \5561 , \5225 );
and \U$5248 ( \5563 , \5559 , \5562 );
and \U$5249 ( \5564 , \5557 , \5562 );
or \U$5250 ( \5565 , \5560 , \5563 , \5564 );
and \U$5251 ( \5566 , \5555 , \5565 );
xor \U$5252 ( \5567 , \5010 , \5014 );
xor \U$5253 ( \5568 , \5567 , \5019 );
and \U$5254 ( \5569 , \5565 , \5568 );
and \U$5255 ( \5570 , \5555 , \5568 );
or \U$5256 ( \5571 , \5566 , \5569 , \5570 );
and \U$5257 ( \5572 , \5545 , \5571 );
xor \U$5258 ( \5573 , \4993 , \4997 );
xor \U$5259 ( \5574 , \5573 , \5002 );
xor \U$5260 ( \5575 , \5320 , \5322 );
xor \U$5261 ( \5576 , \5575 , \5325 );
and \U$5262 ( \5577 , \5574 , \5576 );
xor \U$5263 ( \5578 , \5330 , \5332 );
xor \U$5264 ( \5579 , \5578 , \5335 );
and \U$5265 ( \5580 , \5576 , \5579 );
and \U$5266 ( \5581 , \5574 , \5579 );
or \U$5267 ( \5582 , \5577 , \5580 , \5581 );
and \U$5268 ( \5583 , \5571 , \5582 );
and \U$5269 ( \5584 , \5545 , \5582 );
or \U$5270 ( \5585 , \5572 , \5583 , \5584 );
xor \U$5271 ( \5586 , \5195 , \5211 );
xor \U$5272 ( \5587 , \5586 , \5228 );
xor \U$5273 ( \5588 , \5247 , \5255 );
xor \U$5274 ( \5589 , \5588 , \5260 );
and \U$5275 ( \5590 , \5587 , \5589 );
xor \U$5276 ( \5591 , \5280 , \5296 );
xor \U$5277 ( \5592 , \5591 , \5313 );
and \U$5278 ( \5593 , \5589 , \5592 );
and \U$5279 ( \5594 , \5587 , \5592 );
or \U$5280 ( \5595 , \5590 , \5593 , \5594 );
xor \U$5281 ( \5596 , \4987 , \5005 );
xor \U$5282 ( \5597 , \5596 , \5022 );
and \U$5283 ( \5598 , \5595 , \5597 );
xor \U$5284 ( \5599 , \5347 , \5349 );
xor \U$5285 ( \5600 , \5599 , \5352 );
and \U$5286 ( \5601 , \5597 , \5600 );
and \U$5287 ( \5602 , \5595 , \5600 );
or \U$5288 ( \5603 , \5598 , \5601 , \5602 );
and \U$5289 ( \5604 , \5585 , \5603 );
xor \U$5290 ( \5605 , \5114 , \5124 );
xor \U$5291 ( \5606 , \5605 , \5127 );
and \U$5292 ( \5607 , \5603 , \5606 );
and \U$5293 ( \5608 , \5585 , \5606 );
or \U$5294 ( \5609 , \5604 , \5607 , \5608 );
xor \U$5295 ( \5610 , \5025 , \5077 );
xor \U$5296 ( \5611 , \5610 , \5101 );
xor \U$5297 ( \5612 , \5319 , \5344 );
xor \U$5298 ( \5613 , \5612 , \5355 );
and \U$5299 ( \5614 , \5611 , \5613 );
xor \U$5300 ( \5615 , \5360 , \5362 );
xor \U$5301 ( \5616 , \5615 , \5365 );
and \U$5302 ( \5617 , \5613 , \5616 );
and \U$5303 ( \5618 , \5611 , \5616 );
or \U$5304 ( \5619 , \5614 , \5617 , \5618 );
and \U$5305 ( \5620 , \5609 , \5619 );
xor \U$5306 ( \5621 , \5146 , \5148 );
xor \U$5307 ( \5622 , \5621 , \5151 );
and \U$5308 ( \5623 , \5619 , \5622 );
and \U$5309 ( \5624 , \5609 , \5622 );
or \U$5310 ( \5625 , \5620 , \5623 , \5624 );
xor \U$5311 ( \5626 , \5104 , \5130 );
xor \U$5312 ( \5627 , \5626 , \5141 );
xor \U$5313 ( \5628 , \5358 , \5368 );
xor \U$5314 ( \5629 , \5628 , \5371 );
and \U$5315 ( \5630 , \5627 , \5629 );
and \U$5316 ( \5631 , \5625 , \5630 );
xor \U$5317 ( \5632 , \5374 , \5376 );
xor \U$5318 ( \5633 , \5632 , \5379 );
and \U$5319 ( \5634 , \5630 , \5633 );
and \U$5320 ( \5635 , \5625 , \5633 );
or \U$5321 ( \5636 , \5631 , \5634 , \5635 );
xor \U$5322 ( \5637 , \5382 , \5384 );
xor \U$5323 ( \5638 , \5637 , \5387 );
and \U$5324 ( \5639 , \5636 , \5638 );
and \U$5325 ( \5640 , \5400 , \5639 );
xor \U$5326 ( \5641 , \5400 , \5639 );
xor \U$5327 ( \5642 , \5636 , \5638 );
xor \U$5328 ( \5643 , \4989 , \5401 );
xor \U$5329 ( \5644 , \5401 , \5402 );
not \U$5330 ( \5645 , \5644 );
and \U$5331 ( \5646 , \5643 , \5645 );
and \U$5332 ( \5647 , \316 , \5646 );
not \U$5333 ( \5648 , \5647 );
xnor \U$5334 ( \5649 , \5648 , \5405 );
and \U$5335 ( \5650 , \348 , \5180 );
and \U$5336 ( \5651 , \330 , \5178 );
nor \U$5337 ( \5652 , \5650 , \5651 );
xnor \U$5338 ( \5653 , \5652 , \4992 );
and \U$5339 ( \5654 , \5649 , \5653 );
and \U$5340 ( \5655 , \417 , \4806 );
and \U$5341 ( \5656 , \369 , \4804 );
nor \U$5342 ( \5657 , \5655 , \5656 );
xnor \U$5343 ( \5658 , \5657 , \4574 );
and \U$5344 ( \5659 , \5653 , \5658 );
and \U$5345 ( \5660 , \5649 , \5658 );
or \U$5346 ( \5661 , \5654 , \5659 , \5660 );
and \U$5347 ( \5662 , \494 , \4355 );
and \U$5348 ( \5663 , \425 , \4353 );
nor \U$5349 ( \5664 , \5662 , \5663 );
xnor \U$5350 ( \5665 , \5664 , \4212 );
and \U$5351 ( \5666 , \553 , \4032 );
and \U$5352 ( \5667 , \499 , \4030 );
nor \U$5353 ( \5668 , \5666 , \5667 );
xnor \U$5354 ( \5669 , \5668 , \3786 );
and \U$5355 ( \5670 , \5665 , \5669 );
and \U$5356 ( \5671 , \681 , \3637 );
and \U$5357 ( \5672 , \604 , \3635 );
nor \U$5358 ( \5673 , \5671 , \5672 );
xnor \U$5359 ( \5674 , \5673 , \3450 );
and \U$5360 ( \5675 , \5669 , \5674 );
and \U$5361 ( \5676 , \5665 , \5674 );
or \U$5362 ( \5677 , \5670 , \5675 , \5676 );
and \U$5363 ( \5678 , \5661 , \5677 );
and \U$5364 ( \5679 , \789 , \3324 );
and \U$5365 ( \5680 , \709 , \3322 );
nor \U$5366 ( \5681 , \5679 , \5680 );
xnor \U$5367 ( \5682 , \5681 , \3119 );
and \U$5368 ( \5683 , \925 , \2918 );
and \U$5369 ( \5684 , \863 , \2916 );
nor \U$5370 ( \5685 , \5683 , \5684 );
xnor \U$5371 ( \5686 , \5685 , \2769 );
and \U$5372 ( \5687 , \5682 , \5686 );
and \U$5373 ( \5688 , \1186 , \2596 );
and \U$5374 ( \5689 , \988 , \2594 );
nor \U$5375 ( \5690 , \5688 , \5689 );
xnor \U$5376 ( \5691 , \5690 , \2454 );
and \U$5377 ( \5692 , \5686 , \5691 );
and \U$5378 ( \5693 , \5682 , \5691 );
or \U$5379 ( \5694 , \5687 , \5692 , \5693 );
and \U$5380 ( \5695 , \5677 , \5694 );
and \U$5381 ( \5696 , \5661 , \5694 );
or \U$5382 ( \5697 , \5678 , \5695 , \5696 );
and \U$5383 ( \5698 , \1379 , \2300 );
and \U$5384 ( \5699 , \1274 , \2298 );
nor \U$5385 ( \5700 , \5698 , \5699 );
xnor \U$5386 ( \5701 , \5700 , \2163 );
and \U$5387 ( \5702 , \1500 , \2094 );
and \U$5388 ( \5703 , \1384 , \2092 );
nor \U$5389 ( \5704 , \5702 , \5703 );
xnor \U$5390 ( \5705 , \5704 , \1942 );
and \U$5391 ( \5706 , \5701 , \5705 );
and \U$5392 ( \5707 , \1791 , \1826 );
and \U$5393 ( \5708 , \1615 , \1824 );
nor \U$5394 ( \5709 , \5707 , \5708 );
xnor \U$5395 ( \5710 , \5709 , \1670 );
and \U$5396 ( \5711 , \5705 , \5710 );
and \U$5397 ( \5712 , \5701 , \5710 );
or \U$5398 ( \5713 , \5706 , \5711 , \5712 );
and \U$5399 ( \5714 , \2042 , \1554 );
and \U$5400 ( \5715 , \1799 , \1552 );
nor \U$5401 ( \5716 , \5714 , \5715 );
xnor \U$5402 ( \5717 , \5716 , \1441 );
and \U$5403 ( \5718 , \2233 , \1360 );
and \U$5404 ( \5719 , \2047 , \1358 );
nor \U$5405 ( \5720 , \5718 , \5719 );
xnor \U$5406 ( \5721 , \5720 , \1224 );
and \U$5407 ( \5722 , \5717 , \5721 );
and \U$5408 ( \5723 , \2641 , \1160 );
and \U$5409 ( \5724 , \2377 , \1158 );
nor \U$5410 ( \5725 , \5723 , \5724 );
xnor \U$5411 ( \5726 , \5725 , \1082 );
and \U$5412 ( \5727 , \5721 , \5726 );
and \U$5413 ( \5728 , \5717 , \5726 );
or \U$5414 ( \5729 , \5722 , \5727 , \5728 );
and \U$5415 ( \5730 , \5713 , \5729 );
and \U$5416 ( \5731 , \2840 , \996 );
and \U$5417 ( \5732 , \2666 , \994 );
nor \U$5418 ( \5733 , \5731 , \5732 );
xnor \U$5419 ( \5734 , \5733 , \902 );
and \U$5420 ( \5735 , \3145 , \826 );
and \U$5421 ( \5736 , \3007 , \824 );
nor \U$5422 ( \5737 , \5735 , \5736 );
xnor \U$5423 ( \5738 , \5737 , \754 );
and \U$5424 ( \5739 , \5734 , \5738 );
and \U$5425 ( \5740 , \3681 , \692 );
and \U$5426 ( \5741 , \3264 , \690 );
nor \U$5427 ( \5742 , \5740 , \5741 );
xnor \U$5428 ( \5743 , \5742 , \649 );
and \U$5429 ( \5744 , \5738 , \5743 );
and \U$5430 ( \5745 , \5734 , \5743 );
or \U$5431 ( \5746 , \5739 , \5744 , \5745 );
and \U$5432 ( \5747 , \5729 , \5746 );
and \U$5433 ( \5748 , \5713 , \5746 );
or \U$5434 ( \5749 , \5730 , \5747 , \5748 );
and \U$5435 ( \5750 , \5697 , \5749 );
and \U$5436 ( \5751 , \4011 , \579 );
and \U$5437 ( \5752 , \3889 , \577 );
nor \U$5438 ( \5753 , \5751 , \5752 );
xnor \U$5439 ( \5754 , \5753 , \530 );
and \U$5440 ( \5755 , \4272 , \478 );
and \U$5441 ( \5756 , \4016 , \476 );
nor \U$5442 ( \5757 , \5755 , \5756 );
xnor \U$5443 ( \5758 , \5757 , \437 );
and \U$5444 ( \5759 , \5754 , \5758 );
and \U$5445 ( \5760 , \4771 , \408 );
and \U$5446 ( \5761 , \4469 , \406 );
nor \U$5447 ( \5762 , \5760 , \5761 );
xnor \U$5448 ( \5763 , \5762 , \378 );
and \U$5449 ( \5764 , \5758 , \5763 );
and \U$5450 ( \5765 , \5754 , \5763 );
or \U$5451 ( \5766 , \5759 , \5764 , \5765 );
and \U$5452 ( \5767 , \5248 , \360 );
and \U$5453 ( \5768 , \4779 , \358 );
nor \U$5454 ( \5769 , \5767 , \5768 );
xnor \U$5455 ( \5770 , \5769 , \341 );
and \U$5456 ( \5771 , \5517 , \323 );
and \U$5457 ( \5772 , \5253 , \321 );
nor \U$5458 ( \5773 , \5771 , \5772 );
xnor \U$5459 ( \5774 , \5773 , \328 );
and \U$5460 ( \5775 , \5770 , \5774 );
buf \U$5461 ( \5776 , RIc0c6438_111);
and \U$5462 ( \5777 , \5776 , \317 );
and \U$5463 ( \5778 , \5774 , \5777 );
and \U$5464 ( \5779 , \5770 , \5777 );
or \U$5465 ( \5780 , \5775 , \5778 , \5779 );
and \U$5466 ( \5781 , \5766 , \5780 );
xor \U$5467 ( \5782 , \5511 , \5515 );
xor \U$5468 ( \5783 , \5782 , \5518 );
and \U$5469 ( \5784 , \5780 , \5783 );
and \U$5470 ( \5785 , \5766 , \5783 );
or \U$5471 ( \5786 , \5781 , \5784 , \5785 );
and \U$5472 ( \5787 , \5749 , \5786 );
and \U$5473 ( \5788 , \5697 , \5786 );
or \U$5474 ( \5789 , \5750 , \5787 , \5788 );
xor \U$5475 ( \5790 , \5458 , \5462 );
xor \U$5476 ( \5791 , \5790 , \5467 );
xor \U$5477 ( \5792 , \5422 , \5426 );
xor \U$5478 ( \5793 , \5792 , \5431 );
and \U$5479 ( \5794 , \5791 , \5793 );
xor \U$5480 ( \5795 , \5439 , \5443 );
xor \U$5481 ( \5796 , \5795 , \5448 );
and \U$5482 ( \5797 , \5793 , \5796 );
and \U$5483 ( \5798 , \5791 , \5796 );
or \U$5484 ( \5799 , \5794 , \5797 , \5798 );
xor \U$5485 ( \5800 , \5474 , \5478 );
xor \U$5486 ( \5801 , \5800 , \5483 );
xor \U$5487 ( \5802 , \5491 , \5495 );
xor \U$5488 ( \5803 , \5802 , \5500 );
and \U$5489 ( \5804 , \5801 , \5803 );
xor \U$5490 ( \5805 , \5525 , \5529 );
xor \U$5491 ( \5806 , \5805 , \5534 );
and \U$5492 ( \5807 , \5803 , \5806 );
and \U$5493 ( \5808 , \5801 , \5806 );
or \U$5494 ( \5809 , \5804 , \5807 , \5808 );
and \U$5495 ( \5810 , \5799 , \5809 );
xor \U$5496 ( \5811 , \5183 , \5187 );
xor \U$5497 ( \5812 , \5811 , \5192 );
and \U$5498 ( \5813 , \5809 , \5812 );
and \U$5499 ( \5814 , \5799 , \5812 );
or \U$5500 ( \5815 , \5810 , \5813 , \5814 );
and \U$5501 ( \5816 , \5789 , \5815 );
xor \U$5502 ( \5817 , \5547 , \5549 );
xor \U$5503 ( \5818 , \5817 , \5552 );
xor \U$5504 ( \5819 , \5557 , \5559 );
xor \U$5505 ( \5820 , \5819 , \5562 );
and \U$5506 ( \5821 , \5818 , \5820 );
xor \U$5507 ( \5822 , \5521 , \5537 );
xor \U$5508 ( \5823 , \5822 , \5539 );
and \U$5509 ( \5824 , \5820 , \5823 );
and \U$5510 ( \5825 , \5818 , \5823 );
or \U$5511 ( \5826 , \5821 , \5824 , \5825 );
and \U$5512 ( \5827 , \5815 , \5826 );
and \U$5513 ( \5828 , \5789 , \5826 );
or \U$5514 ( \5829 , \5816 , \5827 , \5828 );
xor \U$5515 ( \5830 , \5555 , \5565 );
xor \U$5516 ( \5831 , \5830 , \5568 );
xor \U$5517 ( \5832 , \5587 , \5589 );
xor \U$5518 ( \5833 , \5832 , \5592 );
and \U$5519 ( \5834 , \5831 , \5833 );
xor \U$5520 ( \5835 , \5574 , \5576 );
xor \U$5521 ( \5836 , \5835 , \5579 );
and \U$5522 ( \5837 , \5833 , \5836 );
and \U$5523 ( \5838 , \5831 , \5836 );
or \U$5524 ( \5839 , \5834 , \5837 , \5838 );
and \U$5525 ( \5840 , \5829 , \5839 );
xor \U$5526 ( \5841 , \5328 , \5338 );
xor \U$5527 ( \5842 , \5841 , \5341 );
and \U$5528 ( \5843 , \5839 , \5842 );
and \U$5529 ( \5844 , \5829 , \5842 );
or \U$5530 ( \5845 , \5840 , \5843 , \5844 );
xor \U$5531 ( \5846 , \5231 , \5263 );
xor \U$5532 ( \5847 , \5846 , \5316 );
xor \U$5533 ( \5848 , \5545 , \5571 );
xor \U$5534 ( \5849 , \5848 , \5582 );
and \U$5535 ( \5850 , \5847 , \5849 );
xor \U$5536 ( \5851 , \5595 , \5597 );
xor \U$5537 ( \5852 , \5851 , \5600 );
and \U$5538 ( \5853 , \5849 , \5852 );
and \U$5539 ( \5854 , \5847 , \5852 );
or \U$5540 ( \5855 , \5850 , \5853 , \5854 );
and \U$5541 ( \5856 , \5845 , \5855 );
xor \U$5542 ( \5857 , \5611 , \5613 );
xor \U$5543 ( \5858 , \5857 , \5616 );
and \U$5544 ( \5859 , \5855 , \5858 );
and \U$5545 ( \5860 , \5845 , \5858 );
or \U$5546 ( \5861 , \5856 , \5859 , \5860 );
xor \U$5547 ( \5862 , \5609 , \5619 );
xor \U$5548 ( \5863 , \5862 , \5622 );
and \U$5549 ( \5864 , \5861 , \5863 );
xor \U$5550 ( \5865 , \5627 , \5629 );
and \U$5551 ( \5866 , \5863 , \5865 );
and \U$5552 ( \5867 , \5861 , \5865 );
or \U$5553 ( \5868 , \5864 , \5866 , \5867 );
xor \U$5554 ( \5869 , \5625 , \5630 );
xor \U$5555 ( \5870 , \5869 , \5633 );
and \U$5556 ( \5871 , \5868 , \5870 );
and \U$5557 ( \5872 , \5642 , \5871 );
xor \U$5558 ( \5873 , \5642 , \5871 );
xor \U$5559 ( \5874 , \5868 , \5870 );
and \U$5560 ( \5875 , \425 , \4806 );
and \U$5561 ( \5876 , \417 , \4804 );
nor \U$5562 ( \5877 , \5875 , \5876 );
xnor \U$5563 ( \5878 , \5877 , \4574 );
and \U$5564 ( \5879 , \499 , \4355 );
and \U$5565 ( \5880 , \494 , \4353 );
nor \U$5566 ( \5881 , \5879 , \5880 );
xnor \U$5567 ( \5882 , \5881 , \4212 );
and \U$5568 ( \5883 , \5878 , \5882 );
and \U$5569 ( \5884 , \604 , \4032 );
and \U$5570 ( \5885 , \553 , \4030 );
nor \U$5571 ( \5886 , \5884 , \5885 );
xnor \U$5572 ( \5887 , \5886 , \3786 );
and \U$5573 ( \5888 , \5882 , \5887 );
and \U$5574 ( \5889 , \5878 , \5887 );
or \U$5575 ( \5890 , \5883 , \5888 , \5889 );
buf \U$5576 ( \5891 , RIc0c8148_49);
buf \U$5577 ( \5892 , RIc0c80d0_50);
and \U$5578 ( \5893 , \5891 , \5892 );
not \U$5579 ( \5894 , \5893 );
and \U$5580 ( \5895 , \5402 , \5894 );
not \U$5581 ( \5896 , \5895 );
and \U$5582 ( \5897 , \330 , \5646 );
and \U$5583 ( \5898 , \316 , \5644 );
nor \U$5584 ( \5899 , \5897 , \5898 );
xnor \U$5585 ( \5900 , \5899 , \5405 );
and \U$5586 ( \5901 , \5896 , \5900 );
and \U$5587 ( \5902 , \369 , \5180 );
and \U$5588 ( \5903 , \348 , \5178 );
nor \U$5589 ( \5904 , \5902 , \5903 );
xnor \U$5590 ( \5905 , \5904 , \4992 );
and \U$5591 ( \5906 , \5900 , \5905 );
and \U$5592 ( \5907 , \5896 , \5905 );
or \U$5593 ( \5908 , \5901 , \5906 , \5907 );
and \U$5594 ( \5909 , \5890 , \5908 );
and \U$5595 ( \5910 , \709 , \3637 );
and \U$5596 ( \5911 , \681 , \3635 );
nor \U$5597 ( \5912 , \5910 , \5911 );
xnor \U$5598 ( \5913 , \5912 , \3450 );
and \U$5599 ( \5914 , \863 , \3324 );
and \U$5600 ( \5915 , \789 , \3322 );
nor \U$5601 ( \5916 , \5914 , \5915 );
xnor \U$5602 ( \5917 , \5916 , \3119 );
and \U$5603 ( \5918 , \5913 , \5917 );
and \U$5604 ( \5919 , \988 , \2918 );
and \U$5605 ( \5920 , \925 , \2916 );
nor \U$5606 ( \5921 , \5919 , \5920 );
xnor \U$5607 ( \5922 , \5921 , \2769 );
and \U$5608 ( \5923 , \5917 , \5922 );
and \U$5609 ( \5924 , \5913 , \5922 );
or \U$5610 ( \5925 , \5918 , \5923 , \5924 );
and \U$5611 ( \5926 , \5908 , \5925 );
and \U$5612 ( \5927 , \5890 , \5925 );
or \U$5613 ( \5928 , \5909 , \5926 , \5927 );
and \U$5614 ( \5929 , \2666 , \1160 );
and \U$5615 ( \5930 , \2641 , \1158 );
nor \U$5616 ( \5931 , \5929 , \5930 );
xnor \U$5617 ( \5932 , \5931 , \1082 );
and \U$5618 ( \5933 , \3007 , \996 );
and \U$5619 ( \5934 , \2840 , \994 );
nor \U$5620 ( \5935 , \5933 , \5934 );
xnor \U$5621 ( \5936 , \5935 , \902 );
and \U$5622 ( \5937 , \5932 , \5936 );
and \U$5623 ( \5938 , \3264 , \826 );
and \U$5624 ( \5939 , \3145 , \824 );
nor \U$5625 ( \5940 , \5938 , \5939 );
xnor \U$5626 ( \5941 , \5940 , \754 );
and \U$5627 ( \5942 , \5936 , \5941 );
and \U$5628 ( \5943 , \5932 , \5941 );
or \U$5629 ( \5944 , \5937 , \5942 , \5943 );
and \U$5630 ( \5945 , \1799 , \1826 );
and \U$5631 ( \5946 , \1791 , \1824 );
nor \U$5632 ( \5947 , \5945 , \5946 );
xnor \U$5633 ( \5948 , \5947 , \1670 );
and \U$5634 ( \5949 , \2047 , \1554 );
and \U$5635 ( \5950 , \2042 , \1552 );
nor \U$5636 ( \5951 , \5949 , \5950 );
xnor \U$5637 ( \5952 , \5951 , \1441 );
and \U$5638 ( \5953 , \5948 , \5952 );
and \U$5639 ( \5954 , \2377 , \1360 );
and \U$5640 ( \5955 , \2233 , \1358 );
nor \U$5641 ( \5956 , \5954 , \5955 );
xnor \U$5642 ( \5957 , \5956 , \1224 );
and \U$5643 ( \5958 , \5952 , \5957 );
and \U$5644 ( \5959 , \5948 , \5957 );
or \U$5645 ( \5960 , \5953 , \5958 , \5959 );
and \U$5646 ( \5961 , \5944 , \5960 );
and \U$5647 ( \5962 , \1274 , \2596 );
and \U$5648 ( \5963 , \1186 , \2594 );
nor \U$5649 ( \5964 , \5962 , \5963 );
xnor \U$5650 ( \5965 , \5964 , \2454 );
and \U$5651 ( \5966 , \1384 , \2300 );
and \U$5652 ( \5967 , \1379 , \2298 );
nor \U$5653 ( \5968 , \5966 , \5967 );
xnor \U$5654 ( \5969 , \5968 , \2163 );
and \U$5655 ( \5970 , \5965 , \5969 );
and \U$5656 ( \5971 , \1615 , \2094 );
and \U$5657 ( \5972 , \1500 , \2092 );
nor \U$5658 ( \5973 , \5971 , \5972 );
xnor \U$5659 ( \5974 , \5973 , \1942 );
and \U$5660 ( \5975 , \5969 , \5974 );
and \U$5661 ( \5976 , \5965 , \5974 );
or \U$5662 ( \5977 , \5970 , \5975 , \5976 );
and \U$5663 ( \5978 , \5960 , \5977 );
and \U$5664 ( \5979 , \5944 , \5977 );
or \U$5665 ( \5980 , \5961 , \5978 , \5979 );
and \U$5666 ( \5981 , \5928 , \5980 );
and \U$5667 ( \5982 , \3889 , \692 );
and \U$5668 ( \5983 , \3681 , \690 );
nor \U$5669 ( \5984 , \5982 , \5983 );
xnor \U$5670 ( \5985 , \5984 , \649 );
and \U$5671 ( \5986 , \4016 , \579 );
and \U$5672 ( \5987 , \4011 , \577 );
nor \U$5673 ( \5988 , \5986 , \5987 );
xnor \U$5674 ( \5989 , \5988 , \530 );
and \U$5675 ( \5990 , \5985 , \5989 );
and \U$5676 ( \5991 , \4469 , \478 );
and \U$5677 ( \5992 , \4272 , \476 );
nor \U$5678 ( \5993 , \5991 , \5992 );
xnor \U$5679 ( \5994 , \5993 , \437 );
and \U$5680 ( \5995 , \5989 , \5994 );
and \U$5681 ( \5996 , \5985 , \5994 );
or \U$5682 ( \5997 , \5990 , \5995 , \5996 );
and \U$5683 ( \5998 , \4779 , \408 );
and \U$5684 ( \5999 , \4771 , \406 );
nor \U$5685 ( \6000 , \5998 , \5999 );
xnor \U$5686 ( \6001 , \6000 , \378 );
and \U$5687 ( \6002 , \5253 , \360 );
and \U$5688 ( \6003 , \5248 , \358 );
nor \U$5689 ( \6004 , \6002 , \6003 );
xnor \U$5690 ( \6005 , \6004 , \341 );
and \U$5691 ( \6006 , \6001 , \6005 );
and \U$5692 ( \6007 , \5776 , \323 );
and \U$5693 ( \6008 , \5517 , \321 );
nor \U$5694 ( \6009 , \6007 , \6008 );
xnor \U$5695 ( \6010 , \6009 , \328 );
and \U$5696 ( \6011 , \6005 , \6010 );
and \U$5697 ( \6012 , \6001 , \6010 );
or \U$5698 ( \6013 , \6006 , \6011 , \6012 );
or \U$5699 ( \6014 , \5997 , \6013 );
and \U$5700 ( \6015 , \5980 , \6014 );
and \U$5701 ( \6016 , \5928 , \6014 );
or \U$5702 ( \6017 , \5981 , \6015 , \6016 );
xor \U$5703 ( \6018 , \5701 , \5705 );
xor \U$5704 ( \6019 , \6018 , \5710 );
xor \U$5705 ( \6020 , \5717 , \5721 );
xor \U$5706 ( \6021 , \6020 , \5726 );
and \U$5707 ( \6022 , \6019 , \6021 );
xor \U$5708 ( \6023 , \5682 , \5686 );
xor \U$5709 ( \6024 , \6023 , \5691 );
and \U$5710 ( \6025 , \6021 , \6024 );
and \U$5711 ( \6026 , \6019 , \6024 );
or \U$5712 ( \6027 , \6022 , \6025 , \6026 );
xor \U$5713 ( \6028 , \5734 , \5738 );
xor \U$5714 ( \6029 , \6028 , \5743 );
xor \U$5715 ( \6030 , \5754 , \5758 );
xor \U$5716 ( \6031 , \6030 , \5763 );
and \U$5717 ( \6032 , \6029 , \6031 );
xor \U$5718 ( \6033 , \5770 , \5774 );
xor \U$5719 ( \6034 , \6033 , \5777 );
and \U$5720 ( \6035 , \6031 , \6034 );
and \U$5721 ( \6036 , \6029 , \6034 );
or \U$5722 ( \6037 , \6032 , \6035 , \6036 );
and \U$5723 ( \6038 , \6027 , \6037 );
xor \U$5724 ( \6039 , \5649 , \5653 );
xor \U$5725 ( \6040 , \6039 , \5658 );
xor \U$5726 ( \6041 , \5665 , \5669 );
xor \U$5727 ( \6042 , \6041 , \5674 );
and \U$5728 ( \6043 , \6040 , \6042 );
and \U$5729 ( \6044 , \6037 , \6043 );
and \U$5730 ( \6045 , \6027 , \6043 );
or \U$5731 ( \6046 , \6038 , \6044 , \6045 );
and \U$5732 ( \6047 , \6017 , \6046 );
xor \U$5733 ( \6048 , \5406 , \5410 );
xor \U$5734 ( \6049 , \6048 , \5415 );
xor \U$5735 ( \6050 , \5791 , \5793 );
xor \U$5736 ( \6051 , \6050 , \5796 );
and \U$5737 ( \6052 , \6049 , \6051 );
xor \U$5738 ( \6053 , \5801 , \5803 );
xor \U$5739 ( \6054 , \6053 , \5806 );
and \U$5740 ( \6055 , \6051 , \6054 );
and \U$5741 ( \6056 , \6049 , \6054 );
or \U$5742 ( \6057 , \6052 , \6055 , \6056 );
and \U$5743 ( \6058 , \6046 , \6057 );
and \U$5744 ( \6059 , \6017 , \6057 );
or \U$5745 ( \6060 , \6047 , \6058 , \6059 );
xor \U$5746 ( \6061 , \5661 , \5677 );
xor \U$5747 ( \6062 , \6061 , \5694 );
xor \U$5748 ( \6063 , \5713 , \5729 );
xor \U$5749 ( \6064 , \6063 , \5746 );
and \U$5750 ( \6065 , \6062 , \6064 );
xor \U$5751 ( \6066 , \5766 , \5780 );
xor \U$5752 ( \6067 , \6066 , \5783 );
and \U$5753 ( \6068 , \6064 , \6067 );
and \U$5754 ( \6069 , \6062 , \6067 );
or \U$5755 ( \6070 , \6065 , \6068 , \6069 );
xor \U$5756 ( \6071 , \5418 , \5434 );
xor \U$5757 ( \6072 , \6071 , \5451 );
and \U$5758 ( \6073 , \6070 , \6072 );
xor \U$5759 ( \6074 , \5470 , \5486 );
xor \U$5760 ( \6075 , \6074 , \5503 );
and \U$5761 ( \6076 , \6072 , \6075 );
and \U$5762 ( \6077 , \6070 , \6075 );
or \U$5763 ( \6078 , \6073 , \6076 , \6077 );
and \U$5764 ( \6079 , \6060 , \6078 );
xor \U$5765 ( \6080 , \5697 , \5749 );
xor \U$5766 ( \6081 , \6080 , \5786 );
xor \U$5767 ( \6082 , \5799 , \5809 );
xor \U$5768 ( \6083 , \6082 , \5812 );
and \U$5769 ( \6084 , \6081 , \6083 );
xor \U$5770 ( \6085 , \5818 , \5820 );
xor \U$5771 ( \6086 , \6085 , \5823 );
and \U$5772 ( \6087 , \6083 , \6086 );
and \U$5773 ( \6088 , \6081 , \6086 );
or \U$5774 ( \6089 , \6084 , \6087 , \6088 );
and \U$5775 ( \6090 , \6078 , \6089 );
and \U$5776 ( \6091 , \6060 , \6089 );
or \U$5777 ( \6092 , \6079 , \6090 , \6091 );
xor \U$5778 ( \6093 , \5454 , \5506 );
xor \U$5779 ( \6094 , \6093 , \5542 );
xor \U$5780 ( \6095 , \5789 , \5815 );
xor \U$5781 ( \6096 , \6095 , \5826 );
and \U$5782 ( \6097 , \6094 , \6096 );
xor \U$5783 ( \6098 , \5831 , \5833 );
xor \U$5784 ( \6099 , \6098 , \5836 );
and \U$5785 ( \6100 , \6096 , \6099 );
and \U$5786 ( \6101 , \6094 , \6099 );
or \U$5787 ( \6102 , \6097 , \6100 , \6101 );
and \U$5788 ( \6103 , \6092 , \6102 );
xor \U$5789 ( \6104 , \5847 , \5849 );
xor \U$5790 ( \6105 , \6104 , \5852 );
and \U$5791 ( \6106 , \6102 , \6105 );
and \U$5792 ( \6107 , \6092 , \6105 );
or \U$5793 ( \6108 , \6103 , \6106 , \6107 );
xor \U$5794 ( \6109 , \5585 , \5603 );
xor \U$5795 ( \6110 , \6109 , \5606 );
and \U$5796 ( \6111 , \6108 , \6110 );
xor \U$5797 ( \6112 , \5845 , \5855 );
xor \U$5798 ( \6113 , \6112 , \5858 );
and \U$5799 ( \6114 , \6110 , \6113 );
and \U$5800 ( \6115 , \6108 , \6113 );
or \U$5801 ( \6116 , \6111 , \6114 , \6115 );
xor \U$5802 ( \6117 , \5861 , \5863 );
xor \U$5803 ( \6118 , \6117 , \5865 );
and \U$5804 ( \6119 , \6116 , \6118 );
and \U$5805 ( \6120 , \5874 , \6119 );
xor \U$5806 ( \6121 , \5874 , \6119 );
xor \U$5807 ( \6122 , \6116 , \6118 );
and \U$5808 ( \6123 , \4011 , \692 );
and \U$5809 ( \6124 , \3889 , \690 );
nor \U$5810 ( \6125 , \6123 , \6124 );
xnor \U$5811 ( \6126 , \6125 , \649 );
and \U$5812 ( \6127 , \4272 , \579 );
and \U$5813 ( \6128 , \4016 , \577 );
nor \U$5814 ( \6129 , \6127 , \6128 );
xnor \U$5815 ( \6130 , \6129 , \530 );
and \U$5816 ( \6131 , \6126 , \6130 );
and \U$5817 ( \6132 , \4771 , \478 );
and \U$5818 ( \6133 , \4469 , \476 );
nor \U$5819 ( \6134 , \6132 , \6133 );
xnor \U$5820 ( \6135 , \6134 , \437 );
and \U$5821 ( \6136 , \6130 , \6135 );
and \U$5822 ( \6137 , \6126 , \6135 );
or \U$5823 ( \6138 , \6131 , \6136 , \6137 );
and \U$5824 ( \6139 , \5248 , \408 );
and \U$5825 ( \6140 , \4779 , \406 );
nor \U$5826 ( \6141 , \6139 , \6140 );
xnor \U$5827 ( \6142 , \6141 , \378 );
and \U$5828 ( \6143 , \5517 , \360 );
and \U$5829 ( \6144 , \5253 , \358 );
nor \U$5830 ( \6145 , \6143 , \6144 );
xnor \U$5831 ( \6146 , \6145 , \341 );
and \U$5832 ( \6147 , \6142 , \6146 );
buf \U$5833 ( \6148 , RIc0c63c0_112);
and \U$5834 ( \6149 , \6148 , \323 );
and \U$5835 ( \6150 , \5776 , \321 );
nor \U$5836 ( \6151 , \6149 , \6150 );
xnor \U$5837 ( \6152 , \6151 , \328 );
and \U$5838 ( \6153 , \6146 , \6152 );
and \U$5839 ( \6154 , \6142 , \6152 );
or \U$5840 ( \6155 , \6147 , \6153 , \6154 );
and \U$5841 ( \6156 , \6138 , \6155 );
buf \U$5842 ( \6157 , RIc0c6348_113);
and \U$5843 ( \6158 , \6157 , \317 );
buf \U$5844 ( \6159 , \6158 );
and \U$5845 ( \6160 , \6155 , \6159 );
and \U$5846 ( \6161 , \6138 , \6159 );
or \U$5847 ( \6162 , \6156 , \6160 , \6161 );
and \U$5848 ( \6163 , \2042 , \1826 );
and \U$5849 ( \6164 , \1799 , \1824 );
nor \U$5850 ( \6165 , \6163 , \6164 );
xnor \U$5851 ( \6166 , \6165 , \1670 );
and \U$5852 ( \6167 , \2233 , \1554 );
and \U$5853 ( \6168 , \2047 , \1552 );
nor \U$5854 ( \6169 , \6167 , \6168 );
xnor \U$5855 ( \6170 , \6169 , \1441 );
and \U$5856 ( \6171 , \6166 , \6170 );
and \U$5857 ( \6172 , \2641 , \1360 );
and \U$5858 ( \6173 , \2377 , \1358 );
nor \U$5859 ( \6174 , \6172 , \6173 );
xnor \U$5860 ( \6175 , \6174 , \1224 );
and \U$5861 ( \6176 , \6170 , \6175 );
and \U$5862 ( \6177 , \6166 , \6175 );
or \U$5863 ( \6178 , \6171 , \6176 , \6177 );
and \U$5864 ( \6179 , \1379 , \2596 );
and \U$5865 ( \6180 , \1274 , \2594 );
nor \U$5866 ( \6181 , \6179 , \6180 );
xnor \U$5867 ( \6182 , \6181 , \2454 );
and \U$5868 ( \6183 , \1500 , \2300 );
and \U$5869 ( \6184 , \1384 , \2298 );
nor \U$5870 ( \6185 , \6183 , \6184 );
xnor \U$5871 ( \6186 , \6185 , \2163 );
and \U$5872 ( \6187 , \6182 , \6186 );
and \U$5873 ( \6188 , \1791 , \2094 );
and \U$5874 ( \6189 , \1615 , \2092 );
nor \U$5875 ( \6190 , \6188 , \6189 );
xnor \U$5876 ( \6191 , \6190 , \1942 );
and \U$5877 ( \6192 , \6186 , \6191 );
and \U$5878 ( \6193 , \6182 , \6191 );
or \U$5879 ( \6194 , \6187 , \6192 , \6193 );
and \U$5880 ( \6195 , \6178 , \6194 );
and \U$5881 ( \6196 , \2840 , \1160 );
and \U$5882 ( \6197 , \2666 , \1158 );
nor \U$5883 ( \6198 , \6196 , \6197 );
xnor \U$5884 ( \6199 , \6198 , \1082 );
and \U$5885 ( \6200 , \3145 , \996 );
and \U$5886 ( \6201 , \3007 , \994 );
nor \U$5887 ( \6202 , \6200 , \6201 );
xnor \U$5888 ( \6203 , \6202 , \902 );
and \U$5889 ( \6204 , \6199 , \6203 );
and \U$5890 ( \6205 , \3681 , \826 );
and \U$5891 ( \6206 , \3264 , \824 );
nor \U$5892 ( \6207 , \6205 , \6206 );
xnor \U$5893 ( \6208 , \6207 , \754 );
and \U$5894 ( \6209 , \6203 , \6208 );
and \U$5895 ( \6210 , \6199 , \6208 );
or \U$5896 ( \6211 , \6204 , \6209 , \6210 );
and \U$5897 ( \6212 , \6194 , \6211 );
and \U$5898 ( \6213 , \6178 , \6211 );
or \U$5899 ( \6214 , \6195 , \6212 , \6213 );
and \U$5900 ( \6215 , \6162 , \6214 );
and \U$5901 ( \6216 , \494 , \4806 );
and \U$5902 ( \6217 , \425 , \4804 );
nor \U$5903 ( \6218 , \6216 , \6217 );
xnor \U$5904 ( \6219 , \6218 , \4574 );
and \U$5905 ( \6220 , \553 , \4355 );
and \U$5906 ( \6221 , \499 , \4353 );
nor \U$5907 ( \6222 , \6220 , \6221 );
xnor \U$5908 ( \6223 , \6222 , \4212 );
and \U$5909 ( \6224 , \6219 , \6223 );
and \U$5910 ( \6225 , \681 , \4032 );
and \U$5911 ( \6226 , \604 , \4030 );
nor \U$5912 ( \6227 , \6225 , \6226 );
xnor \U$5913 ( \6228 , \6227 , \3786 );
and \U$5914 ( \6229 , \6223 , \6228 );
and \U$5915 ( \6230 , \6219 , \6228 );
or \U$5916 ( \6231 , \6224 , \6229 , \6230 );
xor \U$5917 ( \6232 , \5402 , \5891 );
xor \U$5918 ( \6233 , \5891 , \5892 );
not \U$5919 ( \6234 , \6233 );
and \U$5920 ( \6235 , \6232 , \6234 );
and \U$5921 ( \6236 , \316 , \6235 );
not \U$5922 ( \6237 , \6236 );
xnor \U$5923 ( \6238 , \6237 , \5895 );
and \U$5924 ( \6239 , \348 , \5646 );
and \U$5925 ( \6240 , \330 , \5644 );
nor \U$5926 ( \6241 , \6239 , \6240 );
xnor \U$5927 ( \6242 , \6241 , \5405 );
and \U$5928 ( \6243 , \6238 , \6242 );
and \U$5929 ( \6244 , \417 , \5180 );
and \U$5930 ( \6245 , \369 , \5178 );
nor \U$5931 ( \6246 , \6244 , \6245 );
xnor \U$5932 ( \6247 , \6246 , \4992 );
and \U$5933 ( \6248 , \6242 , \6247 );
and \U$5934 ( \6249 , \6238 , \6247 );
or \U$5935 ( \6250 , \6243 , \6248 , \6249 );
and \U$5936 ( \6251 , \6231 , \6250 );
and \U$5937 ( \6252 , \789 , \3637 );
and \U$5938 ( \6253 , \709 , \3635 );
nor \U$5939 ( \6254 , \6252 , \6253 );
xnor \U$5940 ( \6255 , \6254 , \3450 );
and \U$5941 ( \6256 , \925 , \3324 );
and \U$5942 ( \6257 , \863 , \3322 );
nor \U$5943 ( \6258 , \6256 , \6257 );
xnor \U$5944 ( \6259 , \6258 , \3119 );
and \U$5945 ( \6260 , \6255 , \6259 );
and \U$5946 ( \6261 , \1186 , \2918 );
and \U$5947 ( \6262 , \988 , \2916 );
nor \U$5948 ( \6263 , \6261 , \6262 );
xnor \U$5949 ( \6264 , \6263 , \2769 );
and \U$5950 ( \6265 , \6259 , \6264 );
and \U$5951 ( \6266 , \6255 , \6264 );
or \U$5952 ( \6267 , \6260 , \6265 , \6266 );
and \U$5953 ( \6268 , \6250 , \6267 );
and \U$5954 ( \6269 , \6231 , \6267 );
or \U$5955 ( \6270 , \6251 , \6268 , \6269 );
and \U$5956 ( \6271 , \6214 , \6270 );
and \U$5957 ( \6272 , \6162 , \6270 );
or \U$5958 ( \6273 , \6215 , \6271 , \6272 );
xor \U$5959 ( \6274 , \5878 , \5882 );
xor \U$5960 ( \6275 , \6274 , \5887 );
xor \U$5961 ( \6276 , \5896 , \5900 );
xor \U$5962 ( \6277 , \6276 , \5905 );
and \U$5963 ( \6278 , \6275 , \6277 );
xor \U$5964 ( \6279 , \5913 , \5917 );
xor \U$5965 ( \6280 , \6279 , \5922 );
and \U$5966 ( \6281 , \6277 , \6280 );
and \U$5967 ( \6282 , \6275 , \6280 );
or \U$5968 ( \6283 , \6278 , \6281 , \6282 );
xor \U$5969 ( \6284 , \5932 , \5936 );
xor \U$5970 ( \6285 , \6284 , \5941 );
xor \U$5971 ( \6286 , \5948 , \5952 );
xor \U$5972 ( \6287 , \6286 , \5957 );
and \U$5973 ( \6288 , \6285 , \6287 );
xor \U$5974 ( \6289 , \5965 , \5969 );
xor \U$5975 ( \6290 , \6289 , \5974 );
and \U$5976 ( \6291 , \6287 , \6290 );
and \U$5977 ( \6292 , \6285 , \6290 );
or \U$5978 ( \6293 , \6288 , \6291 , \6292 );
and \U$5979 ( \6294 , \6283 , \6293 );
and \U$5980 ( \6295 , \6148 , \317 );
xor \U$5981 ( \6296 , \5985 , \5989 );
xor \U$5982 ( \6297 , \6296 , \5994 );
and \U$5983 ( \6298 , \6295 , \6297 );
xor \U$5984 ( \6299 , \6001 , \6005 );
xor \U$5985 ( \6300 , \6299 , \6010 );
and \U$5986 ( \6301 , \6297 , \6300 );
and \U$5987 ( \6302 , \6295 , \6300 );
or \U$5988 ( \6303 , \6298 , \6301 , \6302 );
and \U$5989 ( \6304 , \6293 , \6303 );
and \U$5990 ( \6305 , \6283 , \6303 );
or \U$5991 ( \6306 , \6294 , \6304 , \6305 );
and \U$5992 ( \6307 , \6273 , \6306 );
xor \U$5993 ( \6308 , \6019 , \6021 );
xor \U$5994 ( \6309 , \6308 , \6024 );
xor \U$5995 ( \6310 , \6029 , \6031 );
xor \U$5996 ( \6311 , \6310 , \6034 );
and \U$5997 ( \6312 , \6309 , \6311 );
xor \U$5998 ( \6313 , \6040 , \6042 );
and \U$5999 ( \6314 , \6311 , \6313 );
and \U$6000 ( \6315 , \6309 , \6313 );
or \U$6001 ( \6316 , \6312 , \6314 , \6315 );
and \U$6002 ( \6317 , \6306 , \6316 );
and \U$6003 ( \6318 , \6273 , \6316 );
or \U$6004 ( \6319 , \6307 , \6317 , \6318 );
xor \U$6005 ( \6320 , \5890 , \5908 );
xor \U$6006 ( \6321 , \6320 , \5925 );
xor \U$6007 ( \6322 , \5944 , \5960 );
xor \U$6008 ( \6323 , \6322 , \5977 );
and \U$6009 ( \6324 , \6321 , \6323 );
xnor \U$6010 ( \6325 , \5997 , \6013 );
and \U$6011 ( \6326 , \6323 , \6325 );
and \U$6012 ( \6327 , \6321 , \6325 );
or \U$6013 ( \6328 , \6324 , \6326 , \6327 );
xor \U$6014 ( \6329 , \6049 , \6051 );
xor \U$6015 ( \6330 , \6329 , \6054 );
and \U$6016 ( \6331 , \6328 , \6330 );
xor \U$6017 ( \6332 , \6062 , \6064 );
xor \U$6018 ( \6333 , \6332 , \6067 );
and \U$6019 ( \6334 , \6330 , \6333 );
and \U$6020 ( \6335 , \6328 , \6333 );
or \U$6021 ( \6336 , \6331 , \6334 , \6335 );
and \U$6022 ( \6337 , \6319 , \6336 );
xor \U$6023 ( \6338 , \5928 , \5980 );
xor \U$6024 ( \6339 , \6338 , \6014 );
xor \U$6025 ( \6340 , \6027 , \6037 );
xor \U$6026 ( \6341 , \6340 , \6043 );
and \U$6027 ( \6342 , \6339 , \6341 );
and \U$6028 ( \6343 , \6336 , \6342 );
and \U$6029 ( \6344 , \6319 , \6342 );
or \U$6030 ( \6345 , \6337 , \6343 , \6344 );
xor \U$6031 ( \6346 , \6017 , \6046 );
xor \U$6032 ( \6347 , \6346 , \6057 );
xor \U$6033 ( \6348 , \6070 , \6072 );
xor \U$6034 ( \6349 , \6348 , \6075 );
and \U$6035 ( \6350 , \6347 , \6349 );
xor \U$6036 ( \6351 , \6081 , \6083 );
xor \U$6037 ( \6352 , \6351 , \6086 );
and \U$6038 ( \6353 , \6349 , \6352 );
and \U$6039 ( \6354 , \6347 , \6352 );
or \U$6040 ( \6355 , \6350 , \6353 , \6354 );
and \U$6041 ( \6356 , \6345 , \6355 );
xor \U$6042 ( \6357 , \6094 , \6096 );
xor \U$6043 ( \6358 , \6357 , \6099 );
and \U$6044 ( \6359 , \6355 , \6358 );
and \U$6045 ( \6360 , \6345 , \6358 );
or \U$6046 ( \6361 , \6356 , \6359 , \6360 );
xor \U$6047 ( \6362 , \5829 , \5839 );
xor \U$6048 ( \6363 , \6362 , \5842 );
and \U$6049 ( \6364 , \6361 , \6363 );
xor \U$6050 ( \6365 , \6092 , \6102 );
xor \U$6051 ( \6366 , \6365 , \6105 );
and \U$6052 ( \6367 , \6363 , \6366 );
and \U$6053 ( \6368 , \6361 , \6366 );
or \U$6054 ( \6369 , \6364 , \6367 , \6368 );
xor \U$6055 ( \6370 , \6108 , \6110 );
xor \U$6056 ( \6371 , \6370 , \6113 );
and \U$6057 ( \6372 , \6369 , \6371 );
and \U$6058 ( \6373 , \6122 , \6372 );
xor \U$6059 ( \6374 , \6122 , \6372 );
xor \U$6060 ( \6375 , \6369 , \6371 );
xor \U$6061 ( \6376 , \6166 , \6170 );
xor \U$6062 ( \6377 , \6376 , \6175 );
xor \U$6063 ( \6378 , \6182 , \6186 );
xor \U$6064 ( \6379 , \6378 , \6191 );
and \U$6065 ( \6380 , \6377 , \6379 );
xor \U$6066 ( \6381 , \6199 , \6203 );
xor \U$6067 ( \6382 , \6381 , \6208 );
and \U$6068 ( \6383 , \6379 , \6382 );
and \U$6069 ( \6384 , \6377 , \6382 );
or \U$6070 ( \6385 , \6380 , \6383 , \6384 );
xor \U$6071 ( \6386 , \6219 , \6223 );
xor \U$6072 ( \6387 , \6386 , \6228 );
xor \U$6073 ( \6388 , \6238 , \6242 );
xor \U$6074 ( \6389 , \6388 , \6247 );
and \U$6075 ( \6390 , \6387 , \6389 );
xor \U$6076 ( \6391 , \6255 , \6259 );
xor \U$6077 ( \6392 , \6391 , \6264 );
and \U$6078 ( \6393 , \6389 , \6392 );
and \U$6079 ( \6394 , \6387 , \6392 );
or \U$6080 ( \6395 , \6390 , \6393 , \6394 );
and \U$6081 ( \6396 , \6385 , \6395 );
xor \U$6082 ( \6397 , \6126 , \6130 );
xor \U$6083 ( \6398 , \6397 , \6135 );
xor \U$6084 ( \6399 , \6142 , \6146 );
xor \U$6085 ( \6400 , \6399 , \6152 );
and \U$6086 ( \6401 , \6398 , \6400 );
not \U$6087 ( \6402 , \6158 );
and \U$6088 ( \6403 , \6400 , \6402 );
and \U$6089 ( \6404 , \6398 , \6402 );
or \U$6090 ( \6405 , \6401 , \6403 , \6404 );
and \U$6091 ( \6406 , \6395 , \6405 );
and \U$6092 ( \6407 , \6385 , \6405 );
or \U$6093 ( \6408 , \6396 , \6406 , \6407 );
and \U$6094 ( \6409 , \425 , \5180 );
and \U$6095 ( \6410 , \417 , \5178 );
nor \U$6096 ( \6411 , \6409 , \6410 );
xnor \U$6097 ( \6412 , \6411 , \4992 );
and \U$6098 ( \6413 , \499 , \4806 );
and \U$6099 ( \6414 , \494 , \4804 );
nor \U$6100 ( \6415 , \6413 , \6414 );
xnor \U$6101 ( \6416 , \6415 , \4574 );
and \U$6102 ( \6417 , \6412 , \6416 );
and \U$6103 ( \6418 , \604 , \4355 );
and \U$6104 ( \6419 , \553 , \4353 );
nor \U$6105 ( \6420 , \6418 , \6419 );
xnor \U$6106 ( \6421 , \6420 , \4212 );
and \U$6107 ( \6422 , \6416 , \6421 );
and \U$6108 ( \6423 , \6412 , \6421 );
or \U$6109 ( \6424 , \6417 , \6422 , \6423 );
buf \U$6110 ( \6425 , RIc0c8058_51);
buf \U$6111 ( \6426 , RIc0c7fe0_52);
and \U$6112 ( \6427 , \6425 , \6426 );
not \U$6113 ( \6428 , \6427 );
and \U$6114 ( \6429 , \5892 , \6428 );
not \U$6115 ( \6430 , \6429 );
and \U$6116 ( \6431 , \330 , \6235 );
and \U$6117 ( \6432 , \316 , \6233 );
nor \U$6118 ( \6433 , \6431 , \6432 );
xnor \U$6119 ( \6434 , \6433 , \5895 );
and \U$6120 ( \6435 , \6430 , \6434 );
and \U$6121 ( \6436 , \369 , \5646 );
and \U$6122 ( \6437 , \348 , \5644 );
nor \U$6123 ( \6438 , \6436 , \6437 );
xnor \U$6124 ( \6439 , \6438 , \5405 );
and \U$6125 ( \6440 , \6434 , \6439 );
and \U$6126 ( \6441 , \6430 , \6439 );
or \U$6127 ( \6442 , \6435 , \6440 , \6441 );
and \U$6128 ( \6443 , \6424 , \6442 );
and \U$6129 ( \6444 , \709 , \4032 );
and \U$6130 ( \6445 , \681 , \4030 );
nor \U$6131 ( \6446 , \6444 , \6445 );
xnor \U$6132 ( \6447 , \6446 , \3786 );
and \U$6133 ( \6448 , \863 , \3637 );
and \U$6134 ( \6449 , \789 , \3635 );
nor \U$6135 ( \6450 , \6448 , \6449 );
xnor \U$6136 ( \6451 , \6450 , \3450 );
and \U$6137 ( \6452 , \6447 , \6451 );
and \U$6138 ( \6453 , \988 , \3324 );
and \U$6139 ( \6454 , \925 , \3322 );
nor \U$6140 ( \6455 , \6453 , \6454 );
xnor \U$6141 ( \6456 , \6455 , \3119 );
and \U$6142 ( \6457 , \6451 , \6456 );
and \U$6143 ( \6458 , \6447 , \6456 );
or \U$6144 ( \6459 , \6452 , \6457 , \6458 );
and \U$6145 ( \6460 , \6442 , \6459 );
and \U$6146 ( \6461 , \6424 , \6459 );
or \U$6147 ( \6462 , \6443 , \6460 , \6461 );
and \U$6148 ( \6463 , \3889 , \826 );
and \U$6149 ( \6464 , \3681 , \824 );
nor \U$6150 ( \6465 , \6463 , \6464 );
xnor \U$6151 ( \6466 , \6465 , \754 );
and \U$6152 ( \6467 , \4016 , \692 );
and \U$6153 ( \6468 , \4011 , \690 );
nor \U$6154 ( \6469 , \6467 , \6468 );
xnor \U$6155 ( \6470 , \6469 , \649 );
and \U$6156 ( \6471 , \6466 , \6470 );
and \U$6157 ( \6472 , \4469 , \579 );
and \U$6158 ( \6473 , \4272 , \577 );
nor \U$6159 ( \6474 , \6472 , \6473 );
xnor \U$6160 ( \6475 , \6474 , \530 );
and \U$6161 ( \6476 , \6470 , \6475 );
and \U$6162 ( \6477 , \6466 , \6475 );
or \U$6163 ( \6478 , \6471 , \6476 , \6477 );
and \U$6164 ( \6479 , \4779 , \478 );
and \U$6165 ( \6480 , \4771 , \476 );
nor \U$6166 ( \6481 , \6479 , \6480 );
xnor \U$6167 ( \6482 , \6481 , \437 );
and \U$6168 ( \6483 , \5253 , \408 );
and \U$6169 ( \6484 , \5248 , \406 );
nor \U$6170 ( \6485 , \6483 , \6484 );
xnor \U$6171 ( \6486 , \6485 , \378 );
and \U$6172 ( \6487 , \6482 , \6486 );
and \U$6173 ( \6488 , \5776 , \360 );
and \U$6174 ( \6489 , \5517 , \358 );
nor \U$6175 ( \6490 , \6488 , \6489 );
xnor \U$6176 ( \6491 , \6490 , \341 );
and \U$6177 ( \6492 , \6486 , \6491 );
and \U$6178 ( \6493 , \6482 , \6491 );
or \U$6179 ( \6494 , \6487 , \6492 , \6493 );
and \U$6180 ( \6495 , \6478 , \6494 );
and \U$6181 ( \6496 , \6157 , \323 );
and \U$6182 ( \6497 , \6148 , \321 );
nor \U$6183 ( \6498 , \6496 , \6497 );
xnor \U$6184 ( \6499 , \6498 , \328 );
buf \U$6185 ( \6500 , RIc0c62d0_114);
and \U$6186 ( \6501 , \6500 , \317 );
and \U$6187 ( \6502 , \6499 , \6501 );
and \U$6188 ( \6503 , \6494 , \6502 );
and \U$6189 ( \6504 , \6478 , \6502 );
or \U$6190 ( \6505 , \6495 , \6503 , \6504 );
and \U$6191 ( \6506 , \6462 , \6505 );
and \U$6192 ( \6507 , \1274 , \2918 );
and \U$6193 ( \6508 , \1186 , \2916 );
nor \U$6194 ( \6509 , \6507 , \6508 );
xnor \U$6195 ( \6510 , \6509 , \2769 );
and \U$6196 ( \6511 , \1384 , \2596 );
and \U$6197 ( \6512 , \1379 , \2594 );
nor \U$6198 ( \6513 , \6511 , \6512 );
xnor \U$6199 ( \6514 , \6513 , \2454 );
and \U$6200 ( \6515 , \6510 , \6514 );
and \U$6201 ( \6516 , \1615 , \2300 );
and \U$6202 ( \6517 , \1500 , \2298 );
nor \U$6203 ( \6518 , \6516 , \6517 );
xnor \U$6204 ( \6519 , \6518 , \2163 );
and \U$6205 ( \6520 , \6514 , \6519 );
and \U$6206 ( \6521 , \6510 , \6519 );
or \U$6207 ( \6522 , \6515 , \6520 , \6521 );
and \U$6208 ( \6523 , \1799 , \2094 );
and \U$6209 ( \6524 , \1791 , \2092 );
nor \U$6210 ( \6525 , \6523 , \6524 );
xnor \U$6211 ( \6526 , \6525 , \1942 );
and \U$6212 ( \6527 , \2047 , \1826 );
and \U$6213 ( \6528 , \2042 , \1824 );
nor \U$6214 ( \6529 , \6527 , \6528 );
xnor \U$6215 ( \6530 , \6529 , \1670 );
and \U$6216 ( \6531 , \6526 , \6530 );
and \U$6217 ( \6532 , \2377 , \1554 );
and \U$6218 ( \6533 , \2233 , \1552 );
nor \U$6219 ( \6534 , \6532 , \6533 );
xnor \U$6220 ( \6535 , \6534 , \1441 );
and \U$6221 ( \6536 , \6530 , \6535 );
and \U$6222 ( \6537 , \6526 , \6535 );
or \U$6223 ( \6538 , \6531 , \6536 , \6537 );
and \U$6224 ( \6539 , \6522 , \6538 );
and \U$6225 ( \6540 , \2666 , \1360 );
and \U$6226 ( \6541 , \2641 , \1358 );
nor \U$6227 ( \6542 , \6540 , \6541 );
xnor \U$6228 ( \6543 , \6542 , \1224 );
and \U$6229 ( \6544 , \3007 , \1160 );
and \U$6230 ( \6545 , \2840 , \1158 );
nor \U$6231 ( \6546 , \6544 , \6545 );
xnor \U$6232 ( \6547 , \6546 , \1082 );
and \U$6233 ( \6548 , \6543 , \6547 );
and \U$6234 ( \6549 , \3264 , \996 );
and \U$6235 ( \6550 , \3145 , \994 );
nor \U$6236 ( \6551 , \6549 , \6550 );
xnor \U$6237 ( \6552 , \6551 , \902 );
and \U$6238 ( \6553 , \6547 , \6552 );
and \U$6239 ( \6554 , \6543 , \6552 );
or \U$6240 ( \6555 , \6548 , \6553 , \6554 );
and \U$6241 ( \6556 , \6538 , \6555 );
and \U$6242 ( \6557 , \6522 , \6555 );
or \U$6243 ( \6558 , \6539 , \6556 , \6557 );
and \U$6244 ( \6559 , \6505 , \6558 );
and \U$6245 ( \6560 , \6462 , \6558 );
or \U$6246 ( \6561 , \6506 , \6559 , \6560 );
and \U$6247 ( \6562 , \6408 , \6561 );
xor \U$6248 ( \6563 , \6275 , \6277 );
xor \U$6249 ( \6564 , \6563 , \6280 );
xor \U$6250 ( \6565 , \6285 , \6287 );
xor \U$6251 ( \6566 , \6565 , \6290 );
and \U$6252 ( \6567 , \6564 , \6566 );
xor \U$6253 ( \6568 , \6295 , \6297 );
xor \U$6254 ( \6569 , \6568 , \6300 );
and \U$6255 ( \6570 , \6566 , \6569 );
and \U$6256 ( \6571 , \6564 , \6569 );
or \U$6257 ( \6572 , \6567 , \6570 , \6571 );
and \U$6258 ( \6573 , \6561 , \6572 );
and \U$6259 ( \6574 , \6408 , \6572 );
or \U$6260 ( \6575 , \6562 , \6573 , \6574 );
xor \U$6261 ( \6576 , \6138 , \6155 );
xor \U$6262 ( \6577 , \6576 , \6159 );
xor \U$6263 ( \6578 , \6178 , \6194 );
xor \U$6264 ( \6579 , \6578 , \6211 );
and \U$6265 ( \6580 , \6577 , \6579 );
xor \U$6266 ( \6581 , \6231 , \6250 );
xor \U$6267 ( \6582 , \6581 , \6267 );
and \U$6268 ( \6583 , \6579 , \6582 );
and \U$6269 ( \6584 , \6577 , \6582 );
or \U$6270 ( \6585 , \6580 , \6583 , \6584 );
xor \U$6271 ( \6586 , \6321 , \6323 );
xor \U$6272 ( \6587 , \6586 , \6325 );
and \U$6273 ( \6588 , \6585 , \6587 );
xor \U$6274 ( \6589 , \6309 , \6311 );
xor \U$6275 ( \6590 , \6589 , \6313 );
and \U$6276 ( \6591 , \6587 , \6590 );
and \U$6277 ( \6592 , \6585 , \6590 );
or \U$6278 ( \6593 , \6588 , \6591 , \6592 );
and \U$6279 ( \6594 , \6575 , \6593 );
xor \U$6280 ( \6595 , \6162 , \6214 );
xor \U$6281 ( \6596 , \6595 , \6270 );
xor \U$6282 ( \6597 , \6283 , \6293 );
xor \U$6283 ( \6598 , \6597 , \6303 );
and \U$6284 ( \6599 , \6596 , \6598 );
and \U$6285 ( \6600 , \6593 , \6599 );
and \U$6286 ( \6601 , \6575 , \6599 );
or \U$6287 ( \6602 , \6594 , \6600 , \6601 );
xor \U$6288 ( \6603 , \6273 , \6306 );
xor \U$6289 ( \6604 , \6603 , \6316 );
xor \U$6290 ( \6605 , \6328 , \6330 );
xor \U$6291 ( \6606 , \6605 , \6333 );
and \U$6292 ( \6607 , \6604 , \6606 );
xor \U$6293 ( \6608 , \6339 , \6341 );
and \U$6294 ( \6609 , \6606 , \6608 );
and \U$6295 ( \6610 , \6604 , \6608 );
or \U$6296 ( \6611 , \6607 , \6609 , \6610 );
and \U$6297 ( \6612 , \6602 , \6611 );
xor \U$6298 ( \6613 , \6347 , \6349 );
xor \U$6299 ( \6614 , \6613 , \6352 );
and \U$6300 ( \6615 , \6611 , \6614 );
and \U$6301 ( \6616 , \6602 , \6614 );
or \U$6302 ( \6617 , \6612 , \6615 , \6616 );
xor \U$6303 ( \6618 , \6060 , \6078 );
xor \U$6304 ( \6619 , \6618 , \6089 );
and \U$6305 ( \6620 , \6617 , \6619 );
xor \U$6306 ( \6621 , \6345 , \6355 );
xor \U$6307 ( \6622 , \6621 , \6358 );
and \U$6308 ( \6623 , \6619 , \6622 );
and \U$6309 ( \6624 , \6617 , \6622 );
or \U$6310 ( \6625 , \6620 , \6623 , \6624 );
xor \U$6311 ( \6626 , \6361 , \6363 );
xor \U$6312 ( \6627 , \6626 , \6366 );
and \U$6313 ( \6628 , \6625 , \6627 );
and \U$6314 ( \6629 , \6375 , \6628 );
xor \U$6315 ( \6630 , \6375 , \6628 );
xor \U$6316 ( \6631 , \6625 , \6627 );
xor \U$6317 ( \6632 , \6510 , \6514 );
xor \U$6318 ( \6633 , \6632 , \6519 );
xor \U$6319 ( \6634 , \6526 , \6530 );
xor \U$6320 ( \6635 , \6634 , \6535 );
and \U$6321 ( \6636 , \6633 , \6635 );
xor \U$6322 ( \6637 , \6543 , \6547 );
xor \U$6323 ( \6638 , \6637 , \6552 );
and \U$6324 ( \6639 , \6635 , \6638 );
and \U$6325 ( \6640 , \6633 , \6638 );
or \U$6326 ( \6641 , \6636 , \6639 , \6640 );
xor \U$6327 ( \6642 , \6412 , \6416 );
xor \U$6328 ( \6643 , \6642 , \6421 );
xor \U$6329 ( \6644 , \6430 , \6434 );
xor \U$6330 ( \6645 , \6644 , \6439 );
and \U$6331 ( \6646 , \6643 , \6645 );
xor \U$6332 ( \6647 , \6447 , \6451 );
xor \U$6333 ( \6648 , \6647 , \6456 );
and \U$6334 ( \6649 , \6645 , \6648 );
and \U$6335 ( \6650 , \6643 , \6648 );
or \U$6336 ( \6651 , \6646 , \6649 , \6650 );
and \U$6337 ( \6652 , \6641 , \6651 );
xor \U$6338 ( \6653 , \6466 , \6470 );
xor \U$6339 ( \6654 , \6653 , \6475 );
xor \U$6340 ( \6655 , \6482 , \6486 );
xor \U$6341 ( \6656 , \6655 , \6491 );
and \U$6342 ( \6657 , \6654 , \6656 );
xor \U$6343 ( \6658 , \6499 , \6501 );
and \U$6344 ( \6659 , \6656 , \6658 );
and \U$6345 ( \6660 , \6654 , \6658 );
or \U$6346 ( \6661 , \6657 , \6659 , \6660 );
and \U$6347 ( \6662 , \6651 , \6661 );
and \U$6348 ( \6663 , \6641 , \6661 );
or \U$6349 ( \6664 , \6652 , \6662 , \6663 );
and \U$6350 ( \6665 , \4011 , \826 );
and \U$6351 ( \6666 , \3889 , \824 );
nor \U$6352 ( \6667 , \6665 , \6666 );
xnor \U$6353 ( \6668 , \6667 , \754 );
and \U$6354 ( \6669 , \4272 , \692 );
and \U$6355 ( \6670 , \4016 , \690 );
nor \U$6356 ( \6671 , \6669 , \6670 );
xnor \U$6357 ( \6672 , \6671 , \649 );
and \U$6358 ( \6673 , \6668 , \6672 );
and \U$6359 ( \6674 , \4771 , \579 );
and \U$6360 ( \6675 , \4469 , \577 );
nor \U$6361 ( \6676 , \6674 , \6675 );
xnor \U$6362 ( \6677 , \6676 , \530 );
and \U$6363 ( \6678 , \6672 , \6677 );
and \U$6364 ( \6679 , \6668 , \6677 );
or \U$6365 ( \6680 , \6673 , \6678 , \6679 );
and \U$6366 ( \6681 , \5248 , \478 );
and \U$6367 ( \6682 , \4779 , \476 );
nor \U$6368 ( \6683 , \6681 , \6682 );
xnor \U$6369 ( \6684 , \6683 , \437 );
and \U$6370 ( \6685 , \5517 , \408 );
and \U$6371 ( \6686 , \5253 , \406 );
nor \U$6372 ( \6687 , \6685 , \6686 );
xnor \U$6373 ( \6688 , \6687 , \378 );
and \U$6374 ( \6689 , \6684 , \6688 );
and \U$6375 ( \6690 , \6148 , \360 );
and \U$6376 ( \6691 , \5776 , \358 );
nor \U$6377 ( \6692 , \6690 , \6691 );
xnor \U$6378 ( \6693 , \6692 , \341 );
and \U$6379 ( \6694 , \6688 , \6693 );
and \U$6380 ( \6695 , \6684 , \6693 );
or \U$6381 ( \6696 , \6689 , \6694 , \6695 );
and \U$6382 ( \6697 , \6680 , \6696 );
and \U$6383 ( \6698 , \6500 , \323 );
and \U$6384 ( \6699 , \6157 , \321 );
nor \U$6385 ( \6700 , \6698 , \6699 );
xnor \U$6386 ( \6701 , \6700 , \328 );
buf \U$6387 ( \6702 , RIc0c6258_115);
and \U$6388 ( \6703 , \6702 , \317 );
or \U$6389 ( \6704 , \6701 , \6703 );
and \U$6390 ( \6705 , \6696 , \6704 );
and \U$6391 ( \6706 , \6680 , \6704 );
or \U$6392 ( \6707 , \6697 , \6705 , \6706 );
and \U$6393 ( \6708 , \789 , \4032 );
and \U$6394 ( \6709 , \709 , \4030 );
nor \U$6395 ( \6710 , \6708 , \6709 );
xnor \U$6396 ( \6711 , \6710 , \3786 );
and \U$6397 ( \6712 , \925 , \3637 );
and \U$6398 ( \6713 , \863 , \3635 );
nor \U$6399 ( \6714 , \6712 , \6713 );
xnor \U$6400 ( \6715 , \6714 , \3450 );
and \U$6401 ( \6716 , \6711 , \6715 );
and \U$6402 ( \6717 , \1186 , \3324 );
and \U$6403 ( \6718 , \988 , \3322 );
nor \U$6404 ( \6719 , \6717 , \6718 );
xnor \U$6405 ( \6720 , \6719 , \3119 );
and \U$6406 ( \6721 , \6715 , \6720 );
and \U$6407 ( \6722 , \6711 , \6720 );
or \U$6408 ( \6723 , \6716 , \6721 , \6722 );
and \U$6409 ( \6724 , \494 , \5180 );
and \U$6410 ( \6725 , \425 , \5178 );
nor \U$6411 ( \6726 , \6724 , \6725 );
xnor \U$6412 ( \6727 , \6726 , \4992 );
and \U$6413 ( \6728 , \553 , \4806 );
and \U$6414 ( \6729 , \499 , \4804 );
nor \U$6415 ( \6730 , \6728 , \6729 );
xnor \U$6416 ( \6731 , \6730 , \4574 );
and \U$6417 ( \6732 , \6727 , \6731 );
and \U$6418 ( \6733 , \681 , \4355 );
and \U$6419 ( \6734 , \604 , \4353 );
nor \U$6420 ( \6735 , \6733 , \6734 );
xnor \U$6421 ( \6736 , \6735 , \4212 );
and \U$6422 ( \6737 , \6731 , \6736 );
and \U$6423 ( \6738 , \6727 , \6736 );
or \U$6424 ( \6739 , \6732 , \6737 , \6738 );
and \U$6425 ( \6740 , \6723 , \6739 );
xor \U$6426 ( \6741 , \5892 , \6425 );
xor \U$6427 ( \6742 , \6425 , \6426 );
not \U$6428 ( \6743 , \6742 );
and \U$6429 ( \6744 , \6741 , \6743 );
and \U$6430 ( \6745 , \316 , \6744 );
not \U$6431 ( \6746 , \6745 );
xnor \U$6432 ( \6747 , \6746 , \6429 );
and \U$6433 ( \6748 , \348 , \6235 );
and \U$6434 ( \6749 , \330 , \6233 );
nor \U$6435 ( \6750 , \6748 , \6749 );
xnor \U$6436 ( \6751 , \6750 , \5895 );
and \U$6437 ( \6752 , \6747 , \6751 );
and \U$6438 ( \6753 , \417 , \5646 );
and \U$6439 ( \6754 , \369 , \5644 );
nor \U$6440 ( \6755 , \6753 , \6754 );
xnor \U$6441 ( \6756 , \6755 , \5405 );
and \U$6442 ( \6757 , \6751 , \6756 );
and \U$6443 ( \6758 , \6747 , \6756 );
or \U$6444 ( \6759 , \6752 , \6757 , \6758 );
and \U$6445 ( \6760 , \6739 , \6759 );
and \U$6446 ( \6761 , \6723 , \6759 );
or \U$6447 ( \6762 , \6740 , \6760 , \6761 );
and \U$6448 ( \6763 , \6707 , \6762 );
and \U$6449 ( \6764 , \2042 , \2094 );
and \U$6450 ( \6765 , \1799 , \2092 );
nor \U$6451 ( \6766 , \6764 , \6765 );
xnor \U$6452 ( \6767 , \6766 , \1942 );
and \U$6453 ( \6768 , \2233 , \1826 );
and \U$6454 ( \6769 , \2047 , \1824 );
nor \U$6455 ( \6770 , \6768 , \6769 );
xnor \U$6456 ( \6771 , \6770 , \1670 );
and \U$6457 ( \6772 , \6767 , \6771 );
and \U$6458 ( \6773 , \2641 , \1554 );
and \U$6459 ( \6774 , \2377 , \1552 );
nor \U$6460 ( \6775 , \6773 , \6774 );
xnor \U$6461 ( \6776 , \6775 , \1441 );
and \U$6462 ( \6777 , \6771 , \6776 );
and \U$6463 ( \6778 , \6767 , \6776 );
or \U$6464 ( \6779 , \6772 , \6777 , \6778 );
and \U$6465 ( \6780 , \2840 , \1360 );
and \U$6466 ( \6781 , \2666 , \1358 );
nor \U$6467 ( \6782 , \6780 , \6781 );
xnor \U$6468 ( \6783 , \6782 , \1224 );
and \U$6469 ( \6784 , \3145 , \1160 );
and \U$6470 ( \6785 , \3007 , \1158 );
nor \U$6471 ( \6786 , \6784 , \6785 );
xnor \U$6472 ( \6787 , \6786 , \1082 );
and \U$6473 ( \6788 , \6783 , \6787 );
and \U$6474 ( \6789 , \3681 , \996 );
and \U$6475 ( \6790 , \3264 , \994 );
nor \U$6476 ( \6791 , \6789 , \6790 );
xnor \U$6477 ( \6792 , \6791 , \902 );
and \U$6478 ( \6793 , \6787 , \6792 );
and \U$6479 ( \6794 , \6783 , \6792 );
or \U$6480 ( \6795 , \6788 , \6793 , \6794 );
and \U$6481 ( \6796 , \6779 , \6795 );
and \U$6482 ( \6797 , \1379 , \2918 );
and \U$6483 ( \6798 , \1274 , \2916 );
nor \U$6484 ( \6799 , \6797 , \6798 );
xnor \U$6485 ( \6800 , \6799 , \2769 );
and \U$6486 ( \6801 , \1500 , \2596 );
and \U$6487 ( \6802 , \1384 , \2594 );
nor \U$6488 ( \6803 , \6801 , \6802 );
xnor \U$6489 ( \6804 , \6803 , \2454 );
and \U$6490 ( \6805 , \6800 , \6804 );
and \U$6491 ( \6806 , \1791 , \2300 );
and \U$6492 ( \6807 , \1615 , \2298 );
nor \U$6493 ( \6808 , \6806 , \6807 );
xnor \U$6494 ( \6809 , \6808 , \2163 );
and \U$6495 ( \6810 , \6804 , \6809 );
and \U$6496 ( \6811 , \6800 , \6809 );
or \U$6497 ( \6812 , \6805 , \6810 , \6811 );
and \U$6498 ( \6813 , \6795 , \6812 );
and \U$6499 ( \6814 , \6779 , \6812 );
or \U$6500 ( \6815 , \6796 , \6813 , \6814 );
and \U$6501 ( \6816 , \6762 , \6815 );
and \U$6502 ( \6817 , \6707 , \6815 );
or \U$6503 ( \6818 , \6763 , \6816 , \6817 );
and \U$6504 ( \6819 , \6664 , \6818 );
xor \U$6505 ( \6820 , \6377 , \6379 );
xor \U$6506 ( \6821 , \6820 , \6382 );
xor \U$6507 ( \6822 , \6387 , \6389 );
xor \U$6508 ( \6823 , \6822 , \6392 );
and \U$6509 ( \6824 , \6821 , \6823 );
xor \U$6510 ( \6825 , \6398 , \6400 );
xor \U$6511 ( \6826 , \6825 , \6402 );
and \U$6512 ( \6827 , \6823 , \6826 );
and \U$6513 ( \6828 , \6821 , \6826 );
or \U$6514 ( \6829 , \6824 , \6827 , \6828 );
and \U$6515 ( \6830 , \6818 , \6829 );
and \U$6516 ( \6831 , \6664 , \6829 );
or \U$6517 ( \6832 , \6819 , \6830 , \6831 );
xor \U$6518 ( \6833 , \6424 , \6442 );
xor \U$6519 ( \6834 , \6833 , \6459 );
xor \U$6520 ( \6835 , \6478 , \6494 );
xor \U$6521 ( \6836 , \6835 , \6502 );
and \U$6522 ( \6837 , \6834 , \6836 );
xor \U$6523 ( \6838 , \6522 , \6538 );
xor \U$6524 ( \6839 , \6838 , \6555 );
and \U$6525 ( \6840 , \6836 , \6839 );
and \U$6526 ( \6841 , \6834 , \6839 );
or \U$6527 ( \6842 , \6837 , \6840 , \6841 );
xor \U$6528 ( \6843 , \6577 , \6579 );
xor \U$6529 ( \6844 , \6843 , \6582 );
and \U$6530 ( \6845 , \6842 , \6844 );
xor \U$6531 ( \6846 , \6564 , \6566 );
xor \U$6532 ( \6847 , \6846 , \6569 );
and \U$6533 ( \6848 , \6844 , \6847 );
and \U$6534 ( \6849 , \6842 , \6847 );
or \U$6535 ( \6850 , \6845 , \6848 , \6849 );
and \U$6536 ( \6851 , \6832 , \6850 );
xor \U$6537 ( \6852 , \6385 , \6395 );
xor \U$6538 ( \6853 , \6852 , \6405 );
xor \U$6539 ( \6854 , \6462 , \6505 );
xor \U$6540 ( \6855 , \6854 , \6558 );
and \U$6541 ( \6856 , \6853 , \6855 );
and \U$6542 ( \6857 , \6850 , \6856 );
and \U$6543 ( \6858 , \6832 , \6856 );
or \U$6544 ( \6859 , \6851 , \6857 , \6858 );
xor \U$6545 ( \6860 , \6408 , \6561 );
xor \U$6546 ( \6861 , \6860 , \6572 );
xor \U$6547 ( \6862 , \6585 , \6587 );
xor \U$6548 ( \6863 , \6862 , \6590 );
and \U$6549 ( \6864 , \6861 , \6863 );
xor \U$6550 ( \6865 , \6596 , \6598 );
and \U$6551 ( \6866 , \6863 , \6865 );
and \U$6552 ( \6867 , \6861 , \6865 );
or \U$6553 ( \6868 , \6864 , \6866 , \6867 );
and \U$6554 ( \6869 , \6859 , \6868 );
xor \U$6555 ( \6870 , \6604 , \6606 );
xor \U$6556 ( \6871 , \6870 , \6608 );
and \U$6557 ( \6872 , \6868 , \6871 );
and \U$6558 ( \6873 , \6859 , \6871 );
or \U$6559 ( \6874 , \6869 , \6872 , \6873 );
xor \U$6560 ( \6875 , \6319 , \6336 );
xor \U$6561 ( \6876 , \6875 , \6342 );
and \U$6562 ( \6877 , \6874 , \6876 );
xor \U$6563 ( \6878 , \6602 , \6611 );
xor \U$6564 ( \6879 , \6878 , \6614 );
and \U$6565 ( \6880 , \6876 , \6879 );
and \U$6566 ( \6881 , \6874 , \6879 );
or \U$6567 ( \6882 , \6877 , \6880 , \6881 );
xor \U$6568 ( \6883 , \6617 , \6619 );
xor \U$6569 ( \6884 , \6883 , \6622 );
and \U$6570 ( \6885 , \6882 , \6884 );
and \U$6571 ( \6886 , \6631 , \6885 );
xor \U$6572 ( \6887 , \6631 , \6885 );
xor \U$6573 ( \6888 , \6882 , \6884 );
and \U$6574 ( \6889 , \1274 , \3324 );
and \U$6575 ( \6890 , \1186 , \3322 );
nor \U$6576 ( \6891 , \6889 , \6890 );
xnor \U$6577 ( \6892 , \6891 , \3119 );
and \U$6578 ( \6893 , \1384 , \2918 );
and \U$6579 ( \6894 , \1379 , \2916 );
nor \U$6580 ( \6895 , \6893 , \6894 );
xnor \U$6581 ( \6896 , \6895 , \2769 );
and \U$6582 ( \6897 , \6892 , \6896 );
and \U$6583 ( \6898 , \1615 , \2596 );
and \U$6584 ( \6899 , \1500 , \2594 );
nor \U$6585 ( \6900 , \6898 , \6899 );
xnor \U$6586 ( \6901 , \6900 , \2454 );
and \U$6587 ( \6902 , \6896 , \6901 );
and \U$6588 ( \6903 , \6892 , \6901 );
or \U$6589 ( \6904 , \6897 , \6902 , \6903 );
and \U$6590 ( \6905 , \1799 , \2300 );
and \U$6591 ( \6906 , \1791 , \2298 );
nor \U$6592 ( \6907 , \6905 , \6906 );
xnor \U$6593 ( \6908 , \6907 , \2163 );
and \U$6594 ( \6909 , \2047 , \2094 );
and \U$6595 ( \6910 , \2042 , \2092 );
nor \U$6596 ( \6911 , \6909 , \6910 );
xnor \U$6597 ( \6912 , \6911 , \1942 );
and \U$6598 ( \6913 , \6908 , \6912 );
and \U$6599 ( \6914 , \2377 , \1826 );
and \U$6600 ( \6915 , \2233 , \1824 );
nor \U$6601 ( \6916 , \6914 , \6915 );
xnor \U$6602 ( \6917 , \6916 , \1670 );
and \U$6603 ( \6918 , \6912 , \6917 );
and \U$6604 ( \6919 , \6908 , \6917 );
or \U$6605 ( \6920 , \6913 , \6918 , \6919 );
and \U$6606 ( \6921 , \6904 , \6920 );
and \U$6607 ( \6922 , \2666 , \1554 );
and \U$6608 ( \6923 , \2641 , \1552 );
nor \U$6609 ( \6924 , \6922 , \6923 );
xnor \U$6610 ( \6925 , \6924 , \1441 );
and \U$6611 ( \6926 , \3007 , \1360 );
and \U$6612 ( \6927 , \2840 , \1358 );
nor \U$6613 ( \6928 , \6926 , \6927 );
xnor \U$6614 ( \6929 , \6928 , \1224 );
and \U$6615 ( \6930 , \6925 , \6929 );
and \U$6616 ( \6931 , \3264 , \1160 );
and \U$6617 ( \6932 , \3145 , \1158 );
nor \U$6618 ( \6933 , \6931 , \6932 );
xnor \U$6619 ( \6934 , \6933 , \1082 );
and \U$6620 ( \6935 , \6929 , \6934 );
and \U$6621 ( \6936 , \6925 , \6934 );
or \U$6622 ( \6937 , \6930 , \6935 , \6936 );
and \U$6623 ( \6938 , \6920 , \6937 );
and \U$6624 ( \6939 , \6904 , \6937 );
or \U$6625 ( \6940 , \6921 , \6938 , \6939 );
and \U$6626 ( \6941 , \425 , \5646 );
and \U$6627 ( \6942 , \417 , \5644 );
nor \U$6628 ( \6943 , \6941 , \6942 );
xnor \U$6629 ( \6944 , \6943 , \5405 );
and \U$6630 ( \6945 , \499 , \5180 );
and \U$6631 ( \6946 , \494 , \5178 );
nor \U$6632 ( \6947 , \6945 , \6946 );
xnor \U$6633 ( \6948 , \6947 , \4992 );
and \U$6634 ( \6949 , \6944 , \6948 );
and \U$6635 ( \6950 , \604 , \4806 );
and \U$6636 ( \6951 , \553 , \4804 );
nor \U$6637 ( \6952 , \6950 , \6951 );
xnor \U$6638 ( \6953 , \6952 , \4574 );
and \U$6639 ( \6954 , \6948 , \6953 );
and \U$6640 ( \6955 , \6944 , \6953 );
or \U$6641 ( \6956 , \6949 , \6954 , \6955 );
and \U$6642 ( \6957 , \709 , \4355 );
and \U$6643 ( \6958 , \681 , \4353 );
nor \U$6644 ( \6959 , \6957 , \6958 );
xnor \U$6645 ( \6960 , \6959 , \4212 );
and \U$6646 ( \6961 , \863 , \4032 );
and \U$6647 ( \6962 , \789 , \4030 );
nor \U$6648 ( \6963 , \6961 , \6962 );
xnor \U$6649 ( \6964 , \6963 , \3786 );
and \U$6650 ( \6965 , \6960 , \6964 );
and \U$6651 ( \6966 , \988 , \3637 );
and \U$6652 ( \6967 , \925 , \3635 );
nor \U$6653 ( \6968 , \6966 , \6967 );
xnor \U$6654 ( \6969 , \6968 , \3450 );
and \U$6655 ( \6970 , \6964 , \6969 );
and \U$6656 ( \6971 , \6960 , \6969 );
or \U$6657 ( \6972 , \6965 , \6970 , \6971 );
and \U$6658 ( \6973 , \6956 , \6972 );
buf \U$6659 ( \6974 , RIc0c7f68_53);
buf \U$6660 ( \6975 , RIc0c7ef0_54);
and \U$6661 ( \6976 , \6974 , \6975 );
not \U$6662 ( \6977 , \6976 );
and \U$6663 ( \6978 , \6426 , \6977 );
not \U$6664 ( \6979 , \6978 );
and \U$6665 ( \6980 , \330 , \6744 );
and \U$6666 ( \6981 , \316 , \6742 );
nor \U$6667 ( \6982 , \6980 , \6981 );
xnor \U$6668 ( \6983 , \6982 , \6429 );
and \U$6669 ( \6984 , \6979 , \6983 );
and \U$6670 ( \6985 , \369 , \6235 );
and \U$6671 ( \6986 , \348 , \6233 );
nor \U$6672 ( \6987 , \6985 , \6986 );
xnor \U$6673 ( \6988 , \6987 , \5895 );
and \U$6674 ( \6989 , \6983 , \6988 );
and \U$6675 ( \6990 , \6979 , \6988 );
or \U$6676 ( \6991 , \6984 , \6989 , \6990 );
and \U$6677 ( \6992 , \6972 , \6991 );
and \U$6678 ( \6993 , \6956 , \6991 );
or \U$6679 ( \6994 , \6973 , \6992 , \6993 );
and \U$6680 ( \6995 , \6940 , \6994 );
and \U$6681 ( \6996 , \6157 , \360 );
and \U$6682 ( \6997 , \6148 , \358 );
nor \U$6683 ( \6998 , \6996 , \6997 );
xnor \U$6684 ( \6999 , \6998 , \341 );
and \U$6685 ( \7000 , \6702 , \323 );
and \U$6686 ( \7001 , \6500 , \321 );
nor \U$6687 ( \7002 , \7000 , \7001 );
xnor \U$6688 ( \7003 , \7002 , \328 );
and \U$6689 ( \7004 , \6999 , \7003 );
buf \U$6690 ( \7005 , RIc0c61e0_116);
and \U$6691 ( \7006 , \7005 , \317 );
and \U$6692 ( \7007 , \7003 , \7006 );
and \U$6693 ( \7008 , \6999 , \7006 );
or \U$6694 ( \7009 , \7004 , \7007 , \7008 );
and \U$6695 ( \7010 , \3889 , \996 );
and \U$6696 ( \7011 , \3681 , \994 );
nor \U$6697 ( \7012 , \7010 , \7011 );
xnor \U$6698 ( \7013 , \7012 , \902 );
and \U$6699 ( \7014 , \4016 , \826 );
and \U$6700 ( \7015 , \4011 , \824 );
nor \U$6701 ( \7016 , \7014 , \7015 );
xnor \U$6702 ( \7017 , \7016 , \754 );
and \U$6703 ( \7018 , \7013 , \7017 );
and \U$6704 ( \7019 , \4469 , \692 );
and \U$6705 ( \7020 , \4272 , \690 );
nor \U$6706 ( \7021 , \7019 , \7020 );
xnor \U$6707 ( \7022 , \7021 , \649 );
and \U$6708 ( \7023 , \7017 , \7022 );
and \U$6709 ( \7024 , \7013 , \7022 );
or \U$6710 ( \7025 , \7018 , \7023 , \7024 );
and \U$6711 ( \7026 , \7009 , \7025 );
and \U$6712 ( \7027 , \4779 , \579 );
and \U$6713 ( \7028 , \4771 , \577 );
nor \U$6714 ( \7029 , \7027 , \7028 );
xnor \U$6715 ( \7030 , \7029 , \530 );
and \U$6716 ( \7031 , \5253 , \478 );
and \U$6717 ( \7032 , \5248 , \476 );
nor \U$6718 ( \7033 , \7031 , \7032 );
xnor \U$6719 ( \7034 , \7033 , \437 );
and \U$6720 ( \7035 , \7030 , \7034 );
and \U$6721 ( \7036 , \5776 , \408 );
and \U$6722 ( \7037 , \5517 , \406 );
nor \U$6723 ( \7038 , \7036 , \7037 );
xnor \U$6724 ( \7039 , \7038 , \378 );
and \U$6725 ( \7040 , \7034 , \7039 );
and \U$6726 ( \7041 , \7030 , \7039 );
or \U$6727 ( \7042 , \7035 , \7040 , \7041 );
and \U$6728 ( \7043 , \7025 , \7042 );
and \U$6729 ( \7044 , \7009 , \7042 );
or \U$6730 ( \7045 , \7026 , \7043 , \7044 );
and \U$6731 ( \7046 , \6994 , \7045 );
and \U$6732 ( \7047 , \6940 , \7045 );
or \U$6733 ( \7048 , \6995 , \7046 , \7047 );
xor \U$6734 ( \7049 , \6767 , \6771 );
xor \U$6735 ( \7050 , \7049 , \6776 );
xor \U$6736 ( \7051 , \6783 , \6787 );
xor \U$6737 ( \7052 , \7051 , \6792 );
and \U$6738 ( \7053 , \7050 , \7052 );
xor \U$6739 ( \7054 , \6800 , \6804 );
xor \U$6740 ( \7055 , \7054 , \6809 );
and \U$6741 ( \7056 , \7052 , \7055 );
and \U$6742 ( \7057 , \7050 , \7055 );
or \U$6743 ( \7058 , \7053 , \7056 , \7057 );
xor \U$6744 ( \7059 , \6711 , \6715 );
xor \U$6745 ( \7060 , \7059 , \6720 );
xor \U$6746 ( \7061 , \6727 , \6731 );
xor \U$6747 ( \7062 , \7061 , \6736 );
and \U$6748 ( \7063 , \7060 , \7062 );
xor \U$6749 ( \7064 , \6747 , \6751 );
xor \U$6750 ( \7065 , \7064 , \6756 );
and \U$6751 ( \7066 , \7062 , \7065 );
and \U$6752 ( \7067 , \7060 , \7065 );
or \U$6753 ( \7068 , \7063 , \7066 , \7067 );
and \U$6754 ( \7069 , \7058 , \7068 );
xor \U$6755 ( \7070 , \6668 , \6672 );
xor \U$6756 ( \7071 , \7070 , \6677 );
xor \U$6757 ( \7072 , \6684 , \6688 );
xor \U$6758 ( \7073 , \7072 , \6693 );
and \U$6759 ( \7074 , \7071 , \7073 );
xnor \U$6760 ( \7075 , \6701 , \6703 );
and \U$6761 ( \7076 , \7073 , \7075 );
and \U$6762 ( \7077 , \7071 , \7075 );
or \U$6763 ( \7078 , \7074 , \7076 , \7077 );
and \U$6764 ( \7079 , \7068 , \7078 );
and \U$6765 ( \7080 , \7058 , \7078 );
or \U$6766 ( \7081 , \7069 , \7079 , \7080 );
and \U$6767 ( \7082 , \7048 , \7081 );
xor \U$6768 ( \7083 , \6633 , \6635 );
xor \U$6769 ( \7084 , \7083 , \6638 );
xor \U$6770 ( \7085 , \6643 , \6645 );
xor \U$6771 ( \7086 , \7085 , \6648 );
and \U$6772 ( \7087 , \7084 , \7086 );
xor \U$6773 ( \7088 , \6654 , \6656 );
xor \U$6774 ( \7089 , \7088 , \6658 );
and \U$6775 ( \7090 , \7086 , \7089 );
and \U$6776 ( \7091 , \7084 , \7089 );
or \U$6777 ( \7092 , \7087 , \7090 , \7091 );
and \U$6778 ( \7093 , \7081 , \7092 );
and \U$6779 ( \7094 , \7048 , \7092 );
or \U$6780 ( \7095 , \7082 , \7093 , \7094 );
xor \U$6781 ( \7096 , \6680 , \6696 );
xor \U$6782 ( \7097 , \7096 , \6704 );
xor \U$6783 ( \7098 , \6723 , \6739 );
xor \U$6784 ( \7099 , \7098 , \6759 );
and \U$6785 ( \7100 , \7097 , \7099 );
xor \U$6786 ( \7101 , \6779 , \6795 );
xor \U$6787 ( \7102 , \7101 , \6812 );
and \U$6788 ( \7103 , \7099 , \7102 );
and \U$6789 ( \7104 , \7097 , \7102 );
or \U$6790 ( \7105 , \7100 , \7103 , \7104 );
xor \U$6791 ( \7106 , \6834 , \6836 );
xor \U$6792 ( \7107 , \7106 , \6839 );
and \U$6793 ( \7108 , \7105 , \7107 );
xor \U$6794 ( \7109 , \6821 , \6823 );
xor \U$6795 ( \7110 , \7109 , \6826 );
and \U$6796 ( \7111 , \7107 , \7110 );
and \U$6797 ( \7112 , \7105 , \7110 );
or \U$6798 ( \7113 , \7108 , \7111 , \7112 );
and \U$6799 ( \7114 , \7095 , \7113 );
xor \U$6800 ( \7115 , \6641 , \6651 );
xor \U$6801 ( \7116 , \7115 , \6661 );
xor \U$6802 ( \7117 , \6707 , \6762 );
xor \U$6803 ( \7118 , \7117 , \6815 );
and \U$6804 ( \7119 , \7116 , \7118 );
and \U$6805 ( \7120 , \7113 , \7119 );
and \U$6806 ( \7121 , \7095 , \7119 );
or \U$6807 ( \7122 , \7114 , \7120 , \7121 );
xor \U$6808 ( \7123 , \6664 , \6818 );
xor \U$6809 ( \7124 , \7123 , \6829 );
xor \U$6810 ( \7125 , \6842 , \6844 );
xor \U$6811 ( \7126 , \7125 , \6847 );
and \U$6812 ( \7127 , \7124 , \7126 );
xor \U$6813 ( \7128 , \6853 , \6855 );
and \U$6814 ( \7129 , \7126 , \7128 );
and \U$6815 ( \7130 , \7124 , \7128 );
or \U$6816 ( \7131 , \7127 , \7129 , \7130 );
and \U$6817 ( \7132 , \7122 , \7131 );
xor \U$6818 ( \7133 , \6861 , \6863 );
xor \U$6819 ( \7134 , \7133 , \6865 );
and \U$6820 ( \7135 , \7131 , \7134 );
and \U$6821 ( \7136 , \7122 , \7134 );
or \U$6822 ( \7137 , \7132 , \7135 , \7136 );
xor \U$6823 ( \7138 , \6575 , \6593 );
xor \U$6824 ( \7139 , \7138 , \6599 );
and \U$6825 ( \7140 , \7137 , \7139 );
xor \U$6826 ( \7141 , \6859 , \6868 );
xor \U$6827 ( \7142 , \7141 , \6871 );
and \U$6828 ( \7143 , \7139 , \7142 );
and \U$6829 ( \7144 , \7137 , \7142 );
or \U$6830 ( \7145 , \7140 , \7143 , \7144 );
xor \U$6831 ( \7146 , \6874 , \6876 );
xor \U$6832 ( \7147 , \7146 , \6879 );
and \U$6833 ( \7148 , \7145 , \7147 );
and \U$6834 ( \7149 , \6888 , \7148 );
xor \U$6835 ( \7150 , \6888 , \7148 );
xor \U$6836 ( \7151 , \7145 , \7147 );
and \U$6837 ( \7152 , \4011 , \996 );
and \U$6838 ( \7153 , \3889 , \994 );
nor \U$6839 ( \7154 , \7152 , \7153 );
xnor \U$6840 ( \7155 , \7154 , \902 );
and \U$6841 ( \7156 , \4272 , \826 );
and \U$6842 ( \7157 , \4016 , \824 );
nor \U$6843 ( \7158 , \7156 , \7157 );
xnor \U$6844 ( \7159 , \7158 , \754 );
and \U$6845 ( \7160 , \7155 , \7159 );
and \U$6846 ( \7161 , \4771 , \692 );
and \U$6847 ( \7162 , \4469 , \690 );
nor \U$6848 ( \7163 , \7161 , \7162 );
xnor \U$6849 ( \7164 , \7163 , \649 );
and \U$6850 ( \7165 , \7159 , \7164 );
and \U$6851 ( \7166 , \7155 , \7164 );
or \U$6852 ( \7167 , \7160 , \7165 , \7166 );
and \U$6853 ( \7168 , \6500 , \360 );
and \U$6854 ( \7169 , \6157 , \358 );
nor \U$6855 ( \7170 , \7168 , \7169 );
xnor \U$6856 ( \7171 , \7170 , \341 );
and \U$6857 ( \7172 , \7005 , \323 );
and \U$6858 ( \7173 , \6702 , \321 );
nor \U$6859 ( \7174 , \7172 , \7173 );
xnor \U$6860 ( \7175 , \7174 , \328 );
and \U$6861 ( \7176 , \7171 , \7175 );
buf \U$6862 ( \7177 , RIc0c6168_117);
and \U$6863 ( \7178 , \7177 , \317 );
and \U$6864 ( \7179 , \7175 , \7178 );
and \U$6865 ( \7180 , \7171 , \7178 );
or \U$6866 ( \7181 , \7176 , \7179 , \7180 );
and \U$6867 ( \7182 , \7167 , \7181 );
and \U$6868 ( \7183 , \5248 , \579 );
and \U$6869 ( \7184 , \4779 , \577 );
nor \U$6870 ( \7185 , \7183 , \7184 );
xnor \U$6871 ( \7186 , \7185 , \530 );
and \U$6872 ( \7187 , \5517 , \478 );
and \U$6873 ( \7188 , \5253 , \476 );
nor \U$6874 ( \7189 , \7187 , \7188 );
xnor \U$6875 ( \7190 , \7189 , \437 );
and \U$6876 ( \7191 , \7186 , \7190 );
and \U$6877 ( \7192 , \6148 , \408 );
and \U$6878 ( \7193 , \5776 , \406 );
nor \U$6879 ( \7194 , \7192 , \7193 );
xnor \U$6880 ( \7195 , \7194 , \378 );
and \U$6881 ( \7196 , \7190 , \7195 );
and \U$6882 ( \7197 , \7186 , \7195 );
or \U$6883 ( \7198 , \7191 , \7196 , \7197 );
and \U$6884 ( \7199 , \7181 , \7198 );
and \U$6885 ( \7200 , \7167 , \7198 );
or \U$6886 ( \7201 , \7182 , \7199 , \7200 );
and \U$6887 ( \7202 , \494 , \5646 );
and \U$6888 ( \7203 , \425 , \5644 );
nor \U$6889 ( \7204 , \7202 , \7203 );
xnor \U$6890 ( \7205 , \7204 , \5405 );
and \U$6891 ( \7206 , \553 , \5180 );
and \U$6892 ( \7207 , \499 , \5178 );
nor \U$6893 ( \7208 , \7206 , \7207 );
xnor \U$6894 ( \7209 , \7208 , \4992 );
and \U$6895 ( \7210 , \7205 , \7209 );
and \U$6896 ( \7211 , \681 , \4806 );
and \U$6897 ( \7212 , \604 , \4804 );
nor \U$6898 ( \7213 , \7211 , \7212 );
xnor \U$6899 ( \7214 , \7213 , \4574 );
and \U$6900 ( \7215 , \7209 , \7214 );
and \U$6901 ( \7216 , \7205 , \7214 );
or \U$6902 ( \7217 , \7210 , \7215 , \7216 );
and \U$6903 ( \7218 , \789 , \4355 );
and \U$6904 ( \7219 , \709 , \4353 );
nor \U$6905 ( \7220 , \7218 , \7219 );
xnor \U$6906 ( \7221 , \7220 , \4212 );
and \U$6907 ( \7222 , \925 , \4032 );
and \U$6908 ( \7223 , \863 , \4030 );
nor \U$6909 ( \7224 , \7222 , \7223 );
xnor \U$6910 ( \7225 , \7224 , \3786 );
and \U$6911 ( \7226 , \7221 , \7225 );
and \U$6912 ( \7227 , \1186 , \3637 );
and \U$6913 ( \7228 , \988 , \3635 );
nor \U$6914 ( \7229 , \7227 , \7228 );
xnor \U$6915 ( \7230 , \7229 , \3450 );
and \U$6916 ( \7231 , \7225 , \7230 );
and \U$6917 ( \7232 , \7221 , \7230 );
or \U$6918 ( \7233 , \7226 , \7231 , \7232 );
and \U$6919 ( \7234 , \7217 , \7233 );
xor \U$6920 ( \7235 , \6426 , \6974 );
xor \U$6921 ( \7236 , \6974 , \6975 );
not \U$6922 ( \7237 , \7236 );
and \U$6923 ( \7238 , \7235 , \7237 );
and \U$6924 ( \7239 , \316 , \7238 );
not \U$6925 ( \7240 , \7239 );
xnor \U$6926 ( \7241 , \7240 , \6978 );
and \U$6927 ( \7242 , \348 , \6744 );
and \U$6928 ( \7243 , \330 , \6742 );
nor \U$6929 ( \7244 , \7242 , \7243 );
xnor \U$6930 ( \7245 , \7244 , \6429 );
and \U$6931 ( \7246 , \7241 , \7245 );
and \U$6932 ( \7247 , \417 , \6235 );
and \U$6933 ( \7248 , \369 , \6233 );
nor \U$6934 ( \7249 , \7247 , \7248 );
xnor \U$6935 ( \7250 , \7249 , \5895 );
and \U$6936 ( \7251 , \7245 , \7250 );
and \U$6937 ( \7252 , \7241 , \7250 );
or \U$6938 ( \7253 , \7246 , \7251 , \7252 );
and \U$6939 ( \7254 , \7233 , \7253 );
and \U$6940 ( \7255 , \7217 , \7253 );
or \U$6941 ( \7256 , \7234 , \7254 , \7255 );
and \U$6942 ( \7257 , \7201 , \7256 );
and \U$6943 ( \7258 , \1379 , \3324 );
and \U$6944 ( \7259 , \1274 , \3322 );
nor \U$6945 ( \7260 , \7258 , \7259 );
xnor \U$6946 ( \7261 , \7260 , \3119 );
and \U$6947 ( \7262 , \1500 , \2918 );
and \U$6948 ( \7263 , \1384 , \2916 );
nor \U$6949 ( \7264 , \7262 , \7263 );
xnor \U$6950 ( \7265 , \7264 , \2769 );
and \U$6951 ( \7266 , \7261 , \7265 );
and \U$6952 ( \7267 , \1791 , \2596 );
and \U$6953 ( \7268 , \1615 , \2594 );
nor \U$6954 ( \7269 , \7267 , \7268 );
xnor \U$6955 ( \7270 , \7269 , \2454 );
and \U$6956 ( \7271 , \7265 , \7270 );
and \U$6957 ( \7272 , \7261 , \7270 );
or \U$6958 ( \7273 , \7266 , \7271 , \7272 );
and \U$6959 ( \7274 , \2042 , \2300 );
and \U$6960 ( \7275 , \1799 , \2298 );
nor \U$6961 ( \7276 , \7274 , \7275 );
xnor \U$6962 ( \7277 , \7276 , \2163 );
and \U$6963 ( \7278 , \2233 , \2094 );
and \U$6964 ( \7279 , \2047 , \2092 );
nor \U$6965 ( \7280 , \7278 , \7279 );
xnor \U$6966 ( \7281 , \7280 , \1942 );
and \U$6967 ( \7282 , \7277 , \7281 );
and \U$6968 ( \7283 , \2641 , \1826 );
and \U$6969 ( \7284 , \2377 , \1824 );
nor \U$6970 ( \7285 , \7283 , \7284 );
xnor \U$6971 ( \7286 , \7285 , \1670 );
and \U$6972 ( \7287 , \7281 , \7286 );
and \U$6973 ( \7288 , \7277 , \7286 );
or \U$6974 ( \7289 , \7282 , \7287 , \7288 );
and \U$6975 ( \7290 , \7273 , \7289 );
and \U$6976 ( \7291 , \2840 , \1554 );
and \U$6977 ( \7292 , \2666 , \1552 );
nor \U$6978 ( \7293 , \7291 , \7292 );
xnor \U$6979 ( \7294 , \7293 , \1441 );
and \U$6980 ( \7295 , \3145 , \1360 );
and \U$6981 ( \7296 , \3007 , \1358 );
nor \U$6982 ( \7297 , \7295 , \7296 );
xnor \U$6983 ( \7298 , \7297 , \1224 );
and \U$6984 ( \7299 , \7294 , \7298 );
and \U$6985 ( \7300 , \3681 , \1160 );
and \U$6986 ( \7301 , \3264 , \1158 );
nor \U$6987 ( \7302 , \7300 , \7301 );
xnor \U$6988 ( \7303 , \7302 , \1082 );
and \U$6989 ( \7304 , \7298 , \7303 );
and \U$6990 ( \7305 , \7294 , \7303 );
or \U$6991 ( \7306 , \7299 , \7304 , \7305 );
and \U$6992 ( \7307 , \7289 , \7306 );
and \U$6993 ( \7308 , \7273 , \7306 );
or \U$6994 ( \7309 , \7290 , \7307 , \7308 );
and \U$6995 ( \7310 , \7256 , \7309 );
and \U$6996 ( \7311 , \7201 , \7309 );
or \U$6997 ( \7312 , \7257 , \7310 , \7311 );
xor \U$6998 ( \7313 , \6999 , \7003 );
xor \U$6999 ( \7314 , \7313 , \7006 );
xor \U$7000 ( \7315 , \7013 , \7017 );
xor \U$7001 ( \7316 , \7315 , \7022 );
and \U$7002 ( \7317 , \7314 , \7316 );
xor \U$7003 ( \7318 , \7030 , \7034 );
xor \U$7004 ( \7319 , \7318 , \7039 );
and \U$7005 ( \7320 , \7316 , \7319 );
and \U$7006 ( \7321 , \7314 , \7319 );
or \U$7007 ( \7322 , \7317 , \7320 , \7321 );
xor \U$7008 ( \7323 , \6892 , \6896 );
xor \U$7009 ( \7324 , \7323 , \6901 );
xor \U$7010 ( \7325 , \6908 , \6912 );
xor \U$7011 ( \7326 , \7325 , \6917 );
and \U$7012 ( \7327 , \7324 , \7326 );
xor \U$7013 ( \7328 , \6925 , \6929 );
xor \U$7014 ( \7329 , \7328 , \6934 );
and \U$7015 ( \7330 , \7326 , \7329 );
and \U$7016 ( \7331 , \7324 , \7329 );
or \U$7017 ( \7332 , \7327 , \7330 , \7331 );
and \U$7018 ( \7333 , \7322 , \7332 );
xor \U$7019 ( \7334 , \6944 , \6948 );
xor \U$7020 ( \7335 , \7334 , \6953 );
xor \U$7021 ( \7336 , \6960 , \6964 );
xor \U$7022 ( \7337 , \7336 , \6969 );
and \U$7023 ( \7338 , \7335 , \7337 );
xor \U$7024 ( \7339 , \6979 , \6983 );
xor \U$7025 ( \7340 , \7339 , \6988 );
and \U$7026 ( \7341 , \7337 , \7340 );
and \U$7027 ( \7342 , \7335 , \7340 );
or \U$7028 ( \7343 , \7338 , \7341 , \7342 );
and \U$7029 ( \7344 , \7332 , \7343 );
and \U$7030 ( \7345 , \7322 , \7343 );
or \U$7031 ( \7346 , \7333 , \7344 , \7345 );
and \U$7032 ( \7347 , \7312 , \7346 );
xor \U$7033 ( \7348 , \7050 , \7052 );
xor \U$7034 ( \7349 , \7348 , \7055 );
xor \U$7035 ( \7350 , \7060 , \7062 );
xor \U$7036 ( \7351 , \7350 , \7065 );
and \U$7037 ( \7352 , \7349 , \7351 );
xor \U$7038 ( \7353 , \7071 , \7073 );
xor \U$7039 ( \7354 , \7353 , \7075 );
and \U$7040 ( \7355 , \7351 , \7354 );
and \U$7041 ( \7356 , \7349 , \7354 );
or \U$7042 ( \7357 , \7352 , \7355 , \7356 );
and \U$7043 ( \7358 , \7346 , \7357 );
and \U$7044 ( \7359 , \7312 , \7357 );
or \U$7045 ( \7360 , \7347 , \7358 , \7359 );
xor \U$7046 ( \7361 , \6904 , \6920 );
xor \U$7047 ( \7362 , \7361 , \6937 );
xor \U$7048 ( \7363 , \6956 , \6972 );
xor \U$7049 ( \7364 , \7363 , \6991 );
and \U$7050 ( \7365 , \7362 , \7364 );
xor \U$7051 ( \7366 , \7009 , \7025 );
xor \U$7052 ( \7367 , \7366 , \7042 );
and \U$7053 ( \7368 , \7364 , \7367 );
and \U$7054 ( \7369 , \7362 , \7367 );
or \U$7055 ( \7370 , \7365 , \7368 , \7369 );
xor \U$7056 ( \7371 , \7097 , \7099 );
xor \U$7057 ( \7372 , \7371 , \7102 );
and \U$7058 ( \7373 , \7370 , \7372 );
xor \U$7059 ( \7374 , \7084 , \7086 );
xor \U$7060 ( \7375 , \7374 , \7089 );
and \U$7061 ( \7376 , \7372 , \7375 );
and \U$7062 ( \7377 , \7370 , \7375 );
or \U$7063 ( \7378 , \7373 , \7376 , \7377 );
and \U$7064 ( \7379 , \7360 , \7378 );
xor \U$7065 ( \7380 , \6940 , \6994 );
xor \U$7066 ( \7381 , \7380 , \7045 );
xor \U$7067 ( \7382 , \7058 , \7068 );
xor \U$7068 ( \7383 , \7382 , \7078 );
and \U$7069 ( \7384 , \7381 , \7383 );
and \U$7070 ( \7385 , \7378 , \7384 );
and \U$7071 ( \7386 , \7360 , \7384 );
or \U$7072 ( \7387 , \7379 , \7385 , \7386 );
xor \U$7073 ( \7388 , \7048 , \7081 );
xor \U$7074 ( \7389 , \7388 , \7092 );
xor \U$7075 ( \7390 , \7105 , \7107 );
xor \U$7076 ( \7391 , \7390 , \7110 );
and \U$7077 ( \7392 , \7389 , \7391 );
xor \U$7078 ( \7393 , \7116 , \7118 );
and \U$7079 ( \7394 , \7391 , \7393 );
and \U$7080 ( \7395 , \7389 , \7393 );
or \U$7081 ( \7396 , \7392 , \7394 , \7395 );
and \U$7082 ( \7397 , \7387 , \7396 );
xor \U$7083 ( \7398 , \7124 , \7126 );
xor \U$7084 ( \7399 , \7398 , \7128 );
and \U$7085 ( \7400 , \7396 , \7399 );
and \U$7086 ( \7401 , \7387 , \7399 );
or \U$7087 ( \7402 , \7397 , \7400 , \7401 );
xor \U$7088 ( \7403 , \6832 , \6850 );
xor \U$7089 ( \7404 , \7403 , \6856 );
and \U$7090 ( \7405 , \7402 , \7404 );
xor \U$7091 ( \7406 , \7122 , \7131 );
xor \U$7092 ( \7407 , \7406 , \7134 );
and \U$7093 ( \7408 , \7404 , \7407 );
and \U$7094 ( \7409 , \7402 , \7407 );
or \U$7095 ( \7410 , \7405 , \7408 , \7409 );
xor \U$7096 ( \7411 , \7137 , \7139 );
xor \U$7097 ( \7412 , \7411 , \7142 );
and \U$7098 ( \7413 , \7410 , \7412 );
and \U$7099 ( \7414 , \7151 , \7413 );
xor \U$7100 ( \7415 , \7151 , \7413 );
xor \U$7101 ( \7416 , \7410 , \7412 );
xor \U$7102 ( \7417 , \7205 , \7209 );
xor \U$7103 ( \7418 , \7417 , \7214 );
xor \U$7104 ( \7419 , \7261 , \7265 );
xor \U$7105 ( \7420 , \7419 , \7270 );
and \U$7106 ( \7421 , \7418 , \7420 );
xor \U$7107 ( \7422 , \7221 , \7225 );
xor \U$7108 ( \7423 , \7422 , \7230 );
and \U$7109 ( \7424 , \7420 , \7423 );
and \U$7110 ( \7425 , \7418 , \7423 );
or \U$7111 ( \7426 , \7421 , \7424 , \7425 );
xor \U$7112 ( \7427 , \7277 , \7281 );
xor \U$7113 ( \7428 , \7427 , \7286 );
xor \U$7114 ( \7429 , \7155 , \7159 );
xor \U$7115 ( \7430 , \7429 , \7164 );
and \U$7116 ( \7431 , \7428 , \7430 );
xor \U$7117 ( \7432 , \7294 , \7298 );
xor \U$7118 ( \7433 , \7432 , \7303 );
and \U$7119 ( \7434 , \7430 , \7433 );
and \U$7120 ( \7435 , \7428 , \7433 );
or \U$7121 ( \7436 , \7431 , \7434 , \7435 );
and \U$7122 ( \7437 , \7426 , \7436 );
xor \U$7123 ( \7438 , \7171 , \7175 );
xor \U$7124 ( \7439 , \7438 , \7178 );
xor \U$7125 ( \7440 , \7186 , \7190 );
xor \U$7126 ( \7441 , \7440 , \7195 );
or \U$7127 ( \7442 , \7439 , \7441 );
and \U$7128 ( \7443 , \7436 , \7442 );
and \U$7129 ( \7444 , \7426 , \7442 );
or \U$7130 ( \7445 , \7437 , \7443 , \7444 );
and \U$7131 ( \7446 , \1799 , \2596 );
and \U$7132 ( \7447 , \1791 , \2594 );
nor \U$7133 ( \7448 , \7446 , \7447 );
xnor \U$7134 ( \7449 , \7448 , \2454 );
and \U$7135 ( \7450 , \2047 , \2300 );
and \U$7136 ( \7451 , \2042 , \2298 );
nor \U$7137 ( \7452 , \7450 , \7451 );
xnor \U$7138 ( \7453 , \7452 , \2163 );
and \U$7139 ( \7454 , \7449 , \7453 );
and \U$7140 ( \7455 , \2377 , \2094 );
and \U$7141 ( \7456 , \2233 , \2092 );
nor \U$7142 ( \7457 , \7455 , \7456 );
xnor \U$7143 ( \7458 , \7457 , \1942 );
and \U$7144 ( \7459 , \7453 , \7458 );
and \U$7145 ( \7460 , \7449 , \7458 );
or \U$7146 ( \7461 , \7454 , \7459 , \7460 );
and \U$7147 ( \7462 , \1274 , \3637 );
and \U$7148 ( \7463 , \1186 , \3635 );
nor \U$7149 ( \7464 , \7462 , \7463 );
xnor \U$7150 ( \7465 , \7464 , \3450 );
and \U$7151 ( \7466 , \1384 , \3324 );
and \U$7152 ( \7467 , \1379 , \3322 );
nor \U$7153 ( \7468 , \7466 , \7467 );
xnor \U$7154 ( \7469 , \7468 , \3119 );
and \U$7155 ( \7470 , \7465 , \7469 );
and \U$7156 ( \7471 , \1615 , \2918 );
and \U$7157 ( \7472 , \1500 , \2916 );
nor \U$7158 ( \7473 , \7471 , \7472 );
xnor \U$7159 ( \7474 , \7473 , \2769 );
and \U$7160 ( \7475 , \7469 , \7474 );
and \U$7161 ( \7476 , \7465 , \7474 );
or \U$7162 ( \7477 , \7470 , \7475 , \7476 );
and \U$7163 ( \7478 , \7461 , \7477 );
and \U$7164 ( \7479 , \2666 , \1826 );
and \U$7165 ( \7480 , \2641 , \1824 );
nor \U$7166 ( \7481 , \7479 , \7480 );
xnor \U$7167 ( \7482 , \7481 , \1670 );
and \U$7168 ( \7483 , \3007 , \1554 );
and \U$7169 ( \7484 , \2840 , \1552 );
nor \U$7170 ( \7485 , \7483 , \7484 );
xnor \U$7171 ( \7486 , \7485 , \1441 );
and \U$7172 ( \7487 , \7482 , \7486 );
and \U$7173 ( \7488 , \3264 , \1360 );
and \U$7174 ( \7489 , \3145 , \1358 );
nor \U$7175 ( \7490 , \7488 , \7489 );
xnor \U$7176 ( \7491 , \7490 , \1224 );
and \U$7177 ( \7492 , \7486 , \7491 );
and \U$7178 ( \7493 , \7482 , \7491 );
or \U$7179 ( \7494 , \7487 , \7492 , \7493 );
and \U$7180 ( \7495 , \7477 , \7494 );
and \U$7181 ( \7496 , \7461 , \7494 );
or \U$7182 ( \7497 , \7478 , \7495 , \7496 );
and \U$7183 ( \7498 , \425 , \6235 );
and \U$7184 ( \7499 , \417 , \6233 );
nor \U$7185 ( \7500 , \7498 , \7499 );
xnor \U$7186 ( \7501 , \7500 , \5895 );
and \U$7187 ( \7502 , \499 , \5646 );
and \U$7188 ( \7503 , \494 , \5644 );
nor \U$7189 ( \7504 , \7502 , \7503 );
xnor \U$7190 ( \7505 , \7504 , \5405 );
and \U$7191 ( \7506 , \7501 , \7505 );
and \U$7192 ( \7507 , \604 , \5180 );
and \U$7193 ( \7508 , \553 , \5178 );
nor \U$7194 ( \7509 , \7507 , \7508 );
xnor \U$7195 ( \7510 , \7509 , \4992 );
and \U$7196 ( \7511 , \7505 , \7510 );
and \U$7197 ( \7512 , \7501 , \7510 );
or \U$7198 ( \7513 , \7506 , \7511 , \7512 );
buf \U$7199 ( \7514 , RIc0c7e78_55);
buf \U$7200 ( \7515 , RIc0c7e00_56);
and \U$7201 ( \7516 , \7514 , \7515 );
not \U$7202 ( \7517 , \7516 );
and \U$7203 ( \7518 , \6975 , \7517 );
not \U$7204 ( \7519 , \7518 );
and \U$7205 ( \7520 , \330 , \7238 );
and \U$7206 ( \7521 , \316 , \7236 );
nor \U$7207 ( \7522 , \7520 , \7521 );
xnor \U$7208 ( \7523 , \7522 , \6978 );
and \U$7209 ( \7524 , \7519 , \7523 );
and \U$7210 ( \7525 , \369 , \6744 );
and \U$7211 ( \7526 , \348 , \6742 );
nor \U$7212 ( \7527 , \7525 , \7526 );
xnor \U$7213 ( \7528 , \7527 , \6429 );
and \U$7214 ( \7529 , \7523 , \7528 );
and \U$7215 ( \7530 , \7519 , \7528 );
or \U$7216 ( \7531 , \7524 , \7529 , \7530 );
and \U$7217 ( \7532 , \7513 , \7531 );
and \U$7218 ( \7533 , \709 , \4806 );
and \U$7219 ( \7534 , \681 , \4804 );
nor \U$7220 ( \7535 , \7533 , \7534 );
xnor \U$7221 ( \7536 , \7535 , \4574 );
and \U$7222 ( \7537 , \863 , \4355 );
and \U$7223 ( \7538 , \789 , \4353 );
nor \U$7224 ( \7539 , \7537 , \7538 );
xnor \U$7225 ( \7540 , \7539 , \4212 );
and \U$7226 ( \7541 , \7536 , \7540 );
and \U$7227 ( \7542 , \988 , \4032 );
and \U$7228 ( \7543 , \925 , \4030 );
nor \U$7229 ( \7544 , \7542 , \7543 );
xnor \U$7230 ( \7545 , \7544 , \3786 );
and \U$7231 ( \7546 , \7540 , \7545 );
and \U$7232 ( \7547 , \7536 , \7545 );
or \U$7233 ( \7548 , \7541 , \7546 , \7547 );
and \U$7234 ( \7549 , \7531 , \7548 );
and \U$7235 ( \7550 , \7513 , \7548 );
or \U$7236 ( \7551 , \7532 , \7549 , \7550 );
and \U$7237 ( \7552 , \7497 , \7551 );
and \U$7238 ( \7553 , \3889 , \1160 );
and \U$7239 ( \7554 , \3681 , \1158 );
nor \U$7240 ( \7555 , \7553 , \7554 );
xnor \U$7241 ( \7556 , \7555 , \1082 );
and \U$7242 ( \7557 , \4016 , \996 );
and \U$7243 ( \7558 , \4011 , \994 );
nor \U$7244 ( \7559 , \7557 , \7558 );
xnor \U$7245 ( \7560 , \7559 , \902 );
and \U$7246 ( \7561 , \7556 , \7560 );
and \U$7247 ( \7562 , \4469 , \826 );
and \U$7248 ( \7563 , \4272 , \824 );
nor \U$7249 ( \7564 , \7562 , \7563 );
xnor \U$7250 ( \7565 , \7564 , \754 );
and \U$7251 ( \7566 , \7560 , \7565 );
and \U$7252 ( \7567 , \7556 , \7565 );
or \U$7253 ( \7568 , \7561 , \7566 , \7567 );
and \U$7254 ( \7569 , \4779 , \692 );
and \U$7255 ( \7570 , \4771 , \690 );
nor \U$7256 ( \7571 , \7569 , \7570 );
xnor \U$7257 ( \7572 , \7571 , \649 );
and \U$7258 ( \7573 , \5253 , \579 );
and \U$7259 ( \7574 , \5248 , \577 );
nor \U$7260 ( \7575 , \7573 , \7574 );
xnor \U$7261 ( \7576 , \7575 , \530 );
and \U$7262 ( \7577 , \7572 , \7576 );
and \U$7263 ( \7578 , \5776 , \478 );
and \U$7264 ( \7579 , \5517 , \476 );
nor \U$7265 ( \7580 , \7578 , \7579 );
xnor \U$7266 ( \7581 , \7580 , \437 );
and \U$7267 ( \7582 , \7576 , \7581 );
and \U$7268 ( \7583 , \7572 , \7581 );
or \U$7269 ( \7584 , \7577 , \7582 , \7583 );
and \U$7270 ( \7585 , \7568 , \7584 );
and \U$7271 ( \7586 , \6157 , \408 );
and \U$7272 ( \7587 , \6148 , \406 );
nor \U$7273 ( \7588 , \7586 , \7587 );
xnor \U$7274 ( \7589 , \7588 , \378 );
and \U$7275 ( \7590 , \6702 , \360 );
and \U$7276 ( \7591 , \6500 , \358 );
nor \U$7277 ( \7592 , \7590 , \7591 );
xnor \U$7278 ( \7593 , \7592 , \341 );
and \U$7279 ( \7594 , \7589 , \7593 );
and \U$7280 ( \7595 , \7177 , \323 );
and \U$7281 ( \7596 , \7005 , \321 );
nor \U$7282 ( \7597 , \7595 , \7596 );
xnor \U$7283 ( \7598 , \7597 , \328 );
and \U$7284 ( \7599 , \7593 , \7598 );
and \U$7285 ( \7600 , \7589 , \7598 );
or \U$7286 ( \7601 , \7594 , \7599 , \7600 );
and \U$7287 ( \7602 , \7584 , \7601 );
and \U$7288 ( \7603 , \7568 , \7601 );
or \U$7289 ( \7604 , \7585 , \7602 , \7603 );
and \U$7290 ( \7605 , \7551 , \7604 );
and \U$7291 ( \7606 , \7497 , \7604 );
or \U$7292 ( \7607 , \7552 , \7605 , \7606 );
and \U$7293 ( \7608 , \7445 , \7607 );
xor \U$7294 ( \7609 , \7314 , \7316 );
xor \U$7295 ( \7610 , \7609 , \7319 );
xor \U$7296 ( \7611 , \7324 , \7326 );
xor \U$7297 ( \7612 , \7611 , \7329 );
and \U$7298 ( \7613 , \7610 , \7612 );
xor \U$7299 ( \7614 , \7335 , \7337 );
xor \U$7300 ( \7615 , \7614 , \7340 );
and \U$7301 ( \7616 , \7612 , \7615 );
and \U$7302 ( \7617 , \7610 , \7615 );
or \U$7303 ( \7618 , \7613 , \7616 , \7617 );
and \U$7304 ( \7619 , \7607 , \7618 );
and \U$7305 ( \7620 , \7445 , \7618 );
or \U$7306 ( \7621 , \7608 , \7619 , \7620 );
xor \U$7307 ( \7622 , \7167 , \7181 );
xor \U$7308 ( \7623 , \7622 , \7198 );
xor \U$7309 ( \7624 , \7217 , \7233 );
xor \U$7310 ( \7625 , \7624 , \7253 );
and \U$7311 ( \7626 , \7623 , \7625 );
xor \U$7312 ( \7627 , \7273 , \7289 );
xor \U$7313 ( \7628 , \7627 , \7306 );
and \U$7314 ( \7629 , \7625 , \7628 );
and \U$7315 ( \7630 , \7623 , \7628 );
or \U$7316 ( \7631 , \7626 , \7629 , \7630 );
xor \U$7317 ( \7632 , \7362 , \7364 );
xor \U$7318 ( \7633 , \7632 , \7367 );
and \U$7319 ( \7634 , \7631 , \7633 );
xor \U$7320 ( \7635 , \7349 , \7351 );
xor \U$7321 ( \7636 , \7635 , \7354 );
and \U$7322 ( \7637 , \7633 , \7636 );
and \U$7323 ( \7638 , \7631 , \7636 );
or \U$7324 ( \7639 , \7634 , \7637 , \7638 );
and \U$7325 ( \7640 , \7621 , \7639 );
xor \U$7326 ( \7641 , \7201 , \7256 );
xor \U$7327 ( \7642 , \7641 , \7309 );
xor \U$7328 ( \7643 , \7322 , \7332 );
xor \U$7329 ( \7644 , \7643 , \7343 );
and \U$7330 ( \7645 , \7642 , \7644 );
and \U$7331 ( \7646 , \7639 , \7645 );
and \U$7332 ( \7647 , \7621 , \7645 );
or \U$7333 ( \7648 , \7640 , \7646 , \7647 );
xor \U$7334 ( \7649 , \7312 , \7346 );
xor \U$7335 ( \7650 , \7649 , \7357 );
xor \U$7336 ( \7651 , \7370 , \7372 );
xor \U$7337 ( \7652 , \7651 , \7375 );
and \U$7338 ( \7653 , \7650 , \7652 );
xor \U$7339 ( \7654 , \7381 , \7383 );
and \U$7340 ( \7655 , \7652 , \7654 );
and \U$7341 ( \7656 , \7650 , \7654 );
or \U$7342 ( \7657 , \7653 , \7655 , \7656 );
and \U$7343 ( \7658 , \7648 , \7657 );
xor \U$7344 ( \7659 , \7389 , \7391 );
xor \U$7345 ( \7660 , \7659 , \7393 );
and \U$7346 ( \7661 , \7657 , \7660 );
and \U$7347 ( \7662 , \7648 , \7660 );
or \U$7348 ( \7663 , \7658 , \7661 , \7662 );
xor \U$7349 ( \7664 , \7095 , \7113 );
xor \U$7350 ( \7665 , \7664 , \7119 );
and \U$7351 ( \7666 , \7663 , \7665 );
xor \U$7352 ( \7667 , \7387 , \7396 );
xor \U$7353 ( \7668 , \7667 , \7399 );
and \U$7354 ( \7669 , \7665 , \7668 );
and \U$7355 ( \7670 , \7663 , \7668 );
or \U$7356 ( \7671 , \7666 , \7669 , \7670 );
xor \U$7357 ( \7672 , \7402 , \7404 );
xor \U$7358 ( \7673 , \7672 , \7407 );
and \U$7359 ( \7674 , \7671 , \7673 );
and \U$7360 ( \7675 , \7416 , \7674 );
xor \U$7361 ( \7676 , \7416 , \7674 );
xor \U$7362 ( \7677 , \7671 , \7673 );
and \U$7363 ( \7678 , \4011 , \1160 );
and \U$7364 ( \7679 , \3889 , \1158 );
nor \U$7365 ( \7680 , \7678 , \7679 );
xnor \U$7366 ( \7681 , \7680 , \1082 );
and \U$7367 ( \7682 , \4272 , \996 );
and \U$7368 ( \7683 , \4016 , \994 );
nor \U$7369 ( \7684 , \7682 , \7683 );
xnor \U$7370 ( \7685 , \7684 , \902 );
and \U$7371 ( \7686 , \7681 , \7685 );
and \U$7372 ( \7687 , \4771 , \826 );
and \U$7373 ( \7688 , \4469 , \824 );
nor \U$7374 ( \7689 , \7687 , \7688 );
xnor \U$7375 ( \7690 , \7689 , \754 );
and \U$7376 ( \7691 , \7685 , \7690 );
and \U$7377 ( \7692 , \7681 , \7690 );
or \U$7378 ( \7693 , \7686 , \7691 , \7692 );
and \U$7379 ( \7694 , \6500 , \408 );
and \U$7380 ( \7695 , \6157 , \406 );
nor \U$7381 ( \7696 , \7694 , \7695 );
xnor \U$7382 ( \7697 , \7696 , \378 );
and \U$7383 ( \7698 , \7005 , \360 );
and \U$7384 ( \7699 , \6702 , \358 );
nor \U$7385 ( \7700 , \7698 , \7699 );
xnor \U$7386 ( \7701 , \7700 , \341 );
and \U$7387 ( \7702 , \7697 , \7701 );
buf \U$7388 ( \7703 , RIc0c60f0_118);
and \U$7389 ( \7704 , \7703 , \323 );
and \U$7390 ( \7705 , \7177 , \321 );
nor \U$7391 ( \7706 , \7704 , \7705 );
xnor \U$7392 ( \7707 , \7706 , \328 );
and \U$7393 ( \7708 , \7701 , \7707 );
and \U$7394 ( \7709 , \7697 , \7707 );
or \U$7395 ( \7710 , \7702 , \7708 , \7709 );
and \U$7396 ( \7711 , \7693 , \7710 );
and \U$7397 ( \7712 , \5248 , \692 );
and \U$7398 ( \7713 , \4779 , \690 );
nor \U$7399 ( \7714 , \7712 , \7713 );
xnor \U$7400 ( \7715 , \7714 , \649 );
and \U$7401 ( \7716 , \5517 , \579 );
and \U$7402 ( \7717 , \5253 , \577 );
nor \U$7403 ( \7718 , \7716 , \7717 );
xnor \U$7404 ( \7719 , \7718 , \530 );
and \U$7405 ( \7720 , \7715 , \7719 );
and \U$7406 ( \7721 , \6148 , \478 );
and \U$7407 ( \7722 , \5776 , \476 );
nor \U$7408 ( \7723 , \7721 , \7722 );
xnor \U$7409 ( \7724 , \7723 , \437 );
and \U$7410 ( \7725 , \7719 , \7724 );
and \U$7411 ( \7726 , \7715 , \7724 );
or \U$7412 ( \7727 , \7720 , \7725 , \7726 );
and \U$7413 ( \7728 , \7710 , \7727 );
and \U$7414 ( \7729 , \7693 , \7727 );
or \U$7415 ( \7730 , \7711 , \7728 , \7729 );
and \U$7416 ( \7731 , \494 , \6235 );
and \U$7417 ( \7732 , \425 , \6233 );
nor \U$7418 ( \7733 , \7731 , \7732 );
xnor \U$7419 ( \7734 , \7733 , \5895 );
and \U$7420 ( \7735 , \553 , \5646 );
and \U$7421 ( \7736 , \499 , \5644 );
nor \U$7422 ( \7737 , \7735 , \7736 );
xnor \U$7423 ( \7738 , \7737 , \5405 );
and \U$7424 ( \7739 , \7734 , \7738 );
and \U$7425 ( \7740 , \681 , \5180 );
and \U$7426 ( \7741 , \604 , \5178 );
nor \U$7427 ( \7742 , \7740 , \7741 );
xnor \U$7428 ( \7743 , \7742 , \4992 );
and \U$7429 ( \7744 , \7738 , \7743 );
and \U$7430 ( \7745 , \7734 , \7743 );
or \U$7431 ( \7746 , \7739 , \7744 , \7745 );
and \U$7432 ( \7747 , \789 , \4806 );
and \U$7433 ( \7748 , \709 , \4804 );
nor \U$7434 ( \7749 , \7747 , \7748 );
xnor \U$7435 ( \7750 , \7749 , \4574 );
and \U$7436 ( \7751 , \925 , \4355 );
and \U$7437 ( \7752 , \863 , \4353 );
nor \U$7438 ( \7753 , \7751 , \7752 );
xnor \U$7439 ( \7754 , \7753 , \4212 );
and \U$7440 ( \7755 , \7750 , \7754 );
and \U$7441 ( \7756 , \1186 , \4032 );
and \U$7442 ( \7757 , \988 , \4030 );
nor \U$7443 ( \7758 , \7756 , \7757 );
xnor \U$7444 ( \7759 , \7758 , \3786 );
and \U$7445 ( \7760 , \7754 , \7759 );
and \U$7446 ( \7761 , \7750 , \7759 );
or \U$7447 ( \7762 , \7755 , \7760 , \7761 );
and \U$7448 ( \7763 , \7746 , \7762 );
xor \U$7449 ( \7764 , \6975 , \7514 );
xor \U$7450 ( \7765 , \7514 , \7515 );
not \U$7451 ( \7766 , \7765 );
and \U$7452 ( \7767 , \7764 , \7766 );
and \U$7453 ( \7768 , \316 , \7767 );
not \U$7454 ( \7769 , \7768 );
xnor \U$7455 ( \7770 , \7769 , \7518 );
and \U$7456 ( \7771 , \348 , \7238 );
and \U$7457 ( \7772 , \330 , \7236 );
nor \U$7458 ( \7773 , \7771 , \7772 );
xnor \U$7459 ( \7774 , \7773 , \6978 );
and \U$7460 ( \7775 , \7770 , \7774 );
and \U$7461 ( \7776 , \417 , \6744 );
and \U$7462 ( \7777 , \369 , \6742 );
nor \U$7463 ( \7778 , \7776 , \7777 );
xnor \U$7464 ( \7779 , \7778 , \6429 );
and \U$7465 ( \7780 , \7774 , \7779 );
and \U$7466 ( \7781 , \7770 , \7779 );
or \U$7467 ( \7782 , \7775 , \7780 , \7781 );
and \U$7468 ( \7783 , \7762 , \7782 );
and \U$7469 ( \7784 , \7746 , \7782 );
or \U$7470 ( \7785 , \7763 , \7783 , \7784 );
and \U$7471 ( \7786 , \7730 , \7785 );
and \U$7472 ( \7787 , \2840 , \1826 );
and \U$7473 ( \7788 , \2666 , \1824 );
nor \U$7474 ( \7789 , \7787 , \7788 );
xnor \U$7475 ( \7790 , \7789 , \1670 );
and \U$7476 ( \7791 , \3145 , \1554 );
and \U$7477 ( \7792 , \3007 , \1552 );
nor \U$7478 ( \7793 , \7791 , \7792 );
xnor \U$7479 ( \7794 , \7793 , \1441 );
and \U$7480 ( \7795 , \7790 , \7794 );
and \U$7481 ( \7796 , \3681 , \1360 );
and \U$7482 ( \7797 , \3264 , \1358 );
nor \U$7483 ( \7798 , \7796 , \7797 );
xnor \U$7484 ( \7799 , \7798 , \1224 );
and \U$7485 ( \7800 , \7794 , \7799 );
and \U$7486 ( \7801 , \7790 , \7799 );
or \U$7487 ( \7802 , \7795 , \7800 , \7801 );
and \U$7488 ( \7803 , \1379 , \3637 );
and \U$7489 ( \7804 , \1274 , \3635 );
nor \U$7490 ( \7805 , \7803 , \7804 );
xnor \U$7491 ( \7806 , \7805 , \3450 );
and \U$7492 ( \7807 , \1500 , \3324 );
and \U$7493 ( \7808 , \1384 , \3322 );
nor \U$7494 ( \7809 , \7807 , \7808 );
xnor \U$7495 ( \7810 , \7809 , \3119 );
and \U$7496 ( \7811 , \7806 , \7810 );
and \U$7497 ( \7812 , \1791 , \2918 );
and \U$7498 ( \7813 , \1615 , \2916 );
nor \U$7499 ( \7814 , \7812 , \7813 );
xnor \U$7500 ( \7815 , \7814 , \2769 );
and \U$7501 ( \7816 , \7810 , \7815 );
and \U$7502 ( \7817 , \7806 , \7815 );
or \U$7503 ( \7818 , \7811 , \7816 , \7817 );
and \U$7504 ( \7819 , \7802 , \7818 );
and \U$7505 ( \7820 , \2042 , \2596 );
and \U$7506 ( \7821 , \1799 , \2594 );
nor \U$7507 ( \7822 , \7820 , \7821 );
xnor \U$7508 ( \7823 , \7822 , \2454 );
and \U$7509 ( \7824 , \2233 , \2300 );
and \U$7510 ( \7825 , \2047 , \2298 );
nor \U$7511 ( \7826 , \7824 , \7825 );
xnor \U$7512 ( \7827 , \7826 , \2163 );
and \U$7513 ( \7828 , \7823 , \7827 );
and \U$7514 ( \7829 , \2641 , \2094 );
and \U$7515 ( \7830 , \2377 , \2092 );
nor \U$7516 ( \7831 , \7829 , \7830 );
xnor \U$7517 ( \7832 , \7831 , \1942 );
and \U$7518 ( \7833 , \7827 , \7832 );
and \U$7519 ( \7834 , \7823 , \7832 );
or \U$7520 ( \7835 , \7828 , \7833 , \7834 );
and \U$7521 ( \7836 , \7818 , \7835 );
and \U$7522 ( \7837 , \7802 , \7835 );
or \U$7523 ( \7838 , \7819 , \7836 , \7837 );
and \U$7524 ( \7839 , \7785 , \7838 );
and \U$7525 ( \7840 , \7730 , \7838 );
or \U$7526 ( \7841 , \7786 , \7839 , \7840 );
xor \U$7527 ( \7842 , \7501 , \7505 );
xor \U$7528 ( \7843 , \7842 , \7510 );
xor \U$7529 ( \7844 , \7465 , \7469 );
xor \U$7530 ( \7845 , \7844 , \7474 );
and \U$7531 ( \7846 , \7843 , \7845 );
xor \U$7532 ( \7847 , \7536 , \7540 );
xor \U$7533 ( \7848 , \7847 , \7545 );
and \U$7534 ( \7849 , \7845 , \7848 );
and \U$7535 ( \7850 , \7843 , \7848 );
or \U$7536 ( \7851 , \7846 , \7849 , \7850 );
and \U$7537 ( \7852 , \7703 , \317 );
xor \U$7538 ( \7853 , \7572 , \7576 );
xor \U$7539 ( \7854 , \7853 , \7581 );
and \U$7540 ( \7855 , \7852 , \7854 );
xor \U$7541 ( \7856 , \7589 , \7593 );
xor \U$7542 ( \7857 , \7856 , \7598 );
and \U$7543 ( \7858 , \7854 , \7857 );
and \U$7544 ( \7859 , \7852 , \7857 );
or \U$7545 ( \7860 , \7855 , \7858 , \7859 );
and \U$7546 ( \7861 , \7851 , \7860 );
xor \U$7547 ( \7862 , \7556 , \7560 );
xor \U$7548 ( \7863 , \7862 , \7565 );
xor \U$7549 ( \7864 , \7449 , \7453 );
xor \U$7550 ( \7865 , \7864 , \7458 );
and \U$7551 ( \7866 , \7863 , \7865 );
xor \U$7552 ( \7867 , \7482 , \7486 );
xor \U$7553 ( \7868 , \7867 , \7491 );
and \U$7554 ( \7869 , \7865 , \7868 );
and \U$7555 ( \7870 , \7863 , \7868 );
or \U$7556 ( \7871 , \7866 , \7869 , \7870 );
and \U$7557 ( \7872 , \7860 , \7871 );
and \U$7558 ( \7873 , \7851 , \7871 );
or \U$7559 ( \7874 , \7861 , \7872 , \7873 );
and \U$7560 ( \7875 , \7841 , \7874 );
xor \U$7561 ( \7876 , \7241 , \7245 );
xor \U$7562 ( \7877 , \7876 , \7250 );
xor \U$7563 ( \7878 , \7418 , \7420 );
xor \U$7564 ( \7879 , \7878 , \7423 );
and \U$7565 ( \7880 , \7877 , \7879 );
xor \U$7566 ( \7881 , \7428 , \7430 );
xor \U$7567 ( \7882 , \7881 , \7433 );
and \U$7568 ( \7883 , \7879 , \7882 );
and \U$7569 ( \7884 , \7877 , \7882 );
or \U$7570 ( \7885 , \7880 , \7883 , \7884 );
and \U$7571 ( \7886 , \7874 , \7885 );
and \U$7572 ( \7887 , \7841 , \7885 );
or \U$7573 ( \7888 , \7875 , \7886 , \7887 );
xor \U$7574 ( \7889 , \7461 , \7477 );
xor \U$7575 ( \7890 , \7889 , \7494 );
xor \U$7576 ( \7891 , \7568 , \7584 );
xor \U$7577 ( \7892 , \7891 , \7601 );
and \U$7578 ( \7893 , \7890 , \7892 );
xnor \U$7579 ( \7894 , \7439 , \7441 );
and \U$7580 ( \7895 , \7892 , \7894 );
and \U$7581 ( \7896 , \7890 , \7894 );
or \U$7582 ( \7897 , \7893 , \7895 , \7896 );
xor \U$7583 ( \7898 , \7623 , \7625 );
xor \U$7584 ( \7899 , \7898 , \7628 );
and \U$7585 ( \7900 , \7897 , \7899 );
xor \U$7586 ( \7901 , \7610 , \7612 );
xor \U$7587 ( \7902 , \7901 , \7615 );
and \U$7588 ( \7903 , \7899 , \7902 );
and \U$7589 ( \7904 , \7897 , \7902 );
or \U$7590 ( \7905 , \7900 , \7903 , \7904 );
and \U$7591 ( \7906 , \7888 , \7905 );
xor \U$7592 ( \7907 , \7426 , \7436 );
xor \U$7593 ( \7908 , \7907 , \7442 );
xor \U$7594 ( \7909 , \7497 , \7551 );
xor \U$7595 ( \7910 , \7909 , \7604 );
and \U$7596 ( \7911 , \7908 , \7910 );
and \U$7597 ( \7912 , \7905 , \7911 );
and \U$7598 ( \7913 , \7888 , \7911 );
or \U$7599 ( \7914 , \7906 , \7912 , \7913 );
xor \U$7600 ( \7915 , \7445 , \7607 );
xor \U$7601 ( \7916 , \7915 , \7618 );
xor \U$7602 ( \7917 , \7631 , \7633 );
xor \U$7603 ( \7918 , \7917 , \7636 );
and \U$7604 ( \7919 , \7916 , \7918 );
xor \U$7605 ( \7920 , \7642 , \7644 );
and \U$7606 ( \7921 , \7918 , \7920 );
and \U$7607 ( \7922 , \7916 , \7920 );
or \U$7608 ( \7923 , \7919 , \7921 , \7922 );
and \U$7609 ( \7924 , \7914 , \7923 );
xor \U$7610 ( \7925 , \7650 , \7652 );
xor \U$7611 ( \7926 , \7925 , \7654 );
and \U$7612 ( \7927 , \7923 , \7926 );
and \U$7613 ( \7928 , \7914 , \7926 );
or \U$7614 ( \7929 , \7924 , \7927 , \7928 );
xor \U$7615 ( \7930 , \7360 , \7378 );
xor \U$7616 ( \7931 , \7930 , \7384 );
and \U$7617 ( \7932 , \7929 , \7931 );
xor \U$7618 ( \7933 , \7648 , \7657 );
xor \U$7619 ( \7934 , \7933 , \7660 );
and \U$7620 ( \7935 , \7931 , \7934 );
and \U$7621 ( \7936 , \7929 , \7934 );
or \U$7622 ( \7937 , \7932 , \7935 , \7936 );
xor \U$7623 ( \7938 , \7663 , \7665 );
xor \U$7624 ( \7939 , \7938 , \7668 );
and \U$7625 ( \7940 , \7937 , \7939 );
and \U$7626 ( \7941 , \7677 , \7940 );
xor \U$7627 ( \7942 , \7677 , \7940 );
xor \U$7628 ( \7943 , \7937 , \7939 );
and \U$7629 ( \7944 , \2666 , \2094 );
and \U$7630 ( \7945 , \2641 , \2092 );
nor \U$7631 ( \7946 , \7944 , \7945 );
xnor \U$7632 ( \7947 , \7946 , \1942 );
and \U$7633 ( \7948 , \3007 , \1826 );
and \U$7634 ( \7949 , \2840 , \1824 );
nor \U$7635 ( \7950 , \7948 , \7949 );
xnor \U$7636 ( \7951 , \7950 , \1670 );
and \U$7637 ( \7952 , \7947 , \7951 );
and \U$7638 ( \7953 , \3264 , \1554 );
and \U$7639 ( \7954 , \3145 , \1552 );
nor \U$7640 ( \7955 , \7953 , \7954 );
xnor \U$7641 ( \7956 , \7955 , \1441 );
and \U$7642 ( \7957 , \7951 , \7956 );
and \U$7643 ( \7958 , \7947 , \7956 );
or \U$7644 ( \7959 , \7952 , \7957 , \7958 );
and \U$7645 ( \7960 , \1274 , \4032 );
and \U$7646 ( \7961 , \1186 , \4030 );
nor \U$7647 ( \7962 , \7960 , \7961 );
xnor \U$7648 ( \7963 , \7962 , \3786 );
and \U$7649 ( \7964 , \1384 , \3637 );
and \U$7650 ( \7965 , \1379 , \3635 );
nor \U$7651 ( \7966 , \7964 , \7965 );
xnor \U$7652 ( \7967 , \7966 , \3450 );
and \U$7653 ( \7968 , \7963 , \7967 );
and \U$7654 ( \7969 , \1615 , \3324 );
and \U$7655 ( \7970 , \1500 , \3322 );
nor \U$7656 ( \7971 , \7969 , \7970 );
xnor \U$7657 ( \7972 , \7971 , \3119 );
and \U$7658 ( \7973 , \7967 , \7972 );
and \U$7659 ( \7974 , \7963 , \7972 );
or \U$7660 ( \7975 , \7968 , \7973 , \7974 );
and \U$7661 ( \7976 , \7959 , \7975 );
and \U$7662 ( \7977 , \1799 , \2918 );
and \U$7663 ( \7978 , \1791 , \2916 );
nor \U$7664 ( \7979 , \7977 , \7978 );
xnor \U$7665 ( \7980 , \7979 , \2769 );
and \U$7666 ( \7981 , \2047 , \2596 );
and \U$7667 ( \7982 , \2042 , \2594 );
nor \U$7668 ( \7983 , \7981 , \7982 );
xnor \U$7669 ( \7984 , \7983 , \2454 );
and \U$7670 ( \7985 , \7980 , \7984 );
and \U$7671 ( \7986 , \2377 , \2300 );
and \U$7672 ( \7987 , \2233 , \2298 );
nor \U$7673 ( \7988 , \7986 , \7987 );
xnor \U$7674 ( \7989 , \7988 , \2163 );
and \U$7675 ( \7990 , \7984 , \7989 );
and \U$7676 ( \7991 , \7980 , \7989 );
or \U$7677 ( \7992 , \7985 , \7990 , \7991 );
and \U$7678 ( \7993 , \7975 , \7992 );
and \U$7679 ( \7994 , \7959 , \7992 );
or \U$7680 ( \7995 , \7976 , \7993 , \7994 );
and \U$7681 ( \7996 , \709 , \5180 );
and \U$7682 ( \7997 , \681 , \5178 );
nor \U$7683 ( \7998 , \7996 , \7997 );
xnor \U$7684 ( \7999 , \7998 , \4992 );
and \U$7685 ( \8000 , \863 , \4806 );
and \U$7686 ( \8001 , \789 , \4804 );
nor \U$7687 ( \8002 , \8000 , \8001 );
xnor \U$7688 ( \8003 , \8002 , \4574 );
and \U$7689 ( \8004 , \7999 , \8003 );
and \U$7690 ( \8005 , \988 , \4355 );
and \U$7691 ( \8006 , \925 , \4353 );
nor \U$7692 ( \8007 , \8005 , \8006 );
xnor \U$7693 ( \8008 , \8007 , \4212 );
and \U$7694 ( \8009 , \8003 , \8008 );
and \U$7695 ( \8010 , \7999 , \8008 );
or \U$7696 ( \8011 , \8004 , \8009 , \8010 );
buf \U$7697 ( \8012 , RIc0c7d88_57);
buf \U$7698 ( \8013 , RIc0c7d10_58);
and \U$7699 ( \8014 , \8012 , \8013 );
not \U$7700 ( \8015 , \8014 );
and \U$7701 ( \8016 , \7515 , \8015 );
not \U$7702 ( \8017 , \8016 );
and \U$7703 ( \8018 , \330 , \7767 );
and \U$7704 ( \8019 , \316 , \7765 );
nor \U$7705 ( \8020 , \8018 , \8019 );
xnor \U$7706 ( \8021 , \8020 , \7518 );
and \U$7707 ( \8022 , \8017 , \8021 );
and \U$7708 ( \8023 , \369 , \7238 );
and \U$7709 ( \8024 , \348 , \7236 );
nor \U$7710 ( \8025 , \8023 , \8024 );
xnor \U$7711 ( \8026 , \8025 , \6978 );
and \U$7712 ( \8027 , \8021 , \8026 );
and \U$7713 ( \8028 , \8017 , \8026 );
or \U$7714 ( \8029 , \8022 , \8027 , \8028 );
and \U$7715 ( \8030 , \8011 , \8029 );
and \U$7716 ( \8031 , \425 , \6744 );
and \U$7717 ( \8032 , \417 , \6742 );
nor \U$7718 ( \8033 , \8031 , \8032 );
xnor \U$7719 ( \8034 , \8033 , \6429 );
and \U$7720 ( \8035 , \499 , \6235 );
and \U$7721 ( \8036 , \494 , \6233 );
nor \U$7722 ( \8037 , \8035 , \8036 );
xnor \U$7723 ( \8038 , \8037 , \5895 );
and \U$7724 ( \8039 , \8034 , \8038 );
and \U$7725 ( \8040 , \604 , \5646 );
and \U$7726 ( \8041 , \553 , \5644 );
nor \U$7727 ( \8042 , \8040 , \8041 );
xnor \U$7728 ( \8043 , \8042 , \5405 );
and \U$7729 ( \8044 , \8038 , \8043 );
and \U$7730 ( \8045 , \8034 , \8043 );
or \U$7731 ( \8046 , \8039 , \8044 , \8045 );
and \U$7732 ( \8047 , \8029 , \8046 );
and \U$7733 ( \8048 , \8011 , \8046 );
or \U$7734 ( \8049 , \8030 , \8047 , \8048 );
and \U$7735 ( \8050 , \7995 , \8049 );
and \U$7736 ( \8051 , \4779 , \826 );
and \U$7737 ( \8052 , \4771 , \824 );
nor \U$7738 ( \8053 , \8051 , \8052 );
xnor \U$7739 ( \8054 , \8053 , \754 );
and \U$7740 ( \8055 , \5253 , \692 );
and \U$7741 ( \8056 , \5248 , \690 );
nor \U$7742 ( \8057 , \8055 , \8056 );
xnor \U$7743 ( \8058 , \8057 , \649 );
and \U$7744 ( \8059 , \8054 , \8058 );
and \U$7745 ( \8060 , \5776 , \579 );
and \U$7746 ( \8061 , \5517 , \577 );
nor \U$7747 ( \8062 , \8060 , \8061 );
xnor \U$7748 ( \8063 , \8062 , \530 );
and \U$7749 ( \8064 , \8058 , \8063 );
and \U$7750 ( \8065 , \8054 , \8063 );
or \U$7751 ( \8066 , \8059 , \8064 , \8065 );
and \U$7752 ( \8067 , \6157 , \478 );
and \U$7753 ( \8068 , \6148 , \476 );
nor \U$7754 ( \8069 , \8067 , \8068 );
xnor \U$7755 ( \8070 , \8069 , \437 );
and \U$7756 ( \8071 , \6702 , \408 );
and \U$7757 ( \8072 , \6500 , \406 );
nor \U$7758 ( \8073 , \8071 , \8072 );
xnor \U$7759 ( \8074 , \8073 , \378 );
and \U$7760 ( \8075 , \8070 , \8074 );
and \U$7761 ( \8076 , \7177 , \360 );
and \U$7762 ( \8077 , \7005 , \358 );
nor \U$7763 ( \8078 , \8076 , \8077 );
xnor \U$7764 ( \8079 , \8078 , \341 );
and \U$7765 ( \8080 , \8074 , \8079 );
and \U$7766 ( \8081 , \8070 , \8079 );
or \U$7767 ( \8082 , \8075 , \8080 , \8081 );
and \U$7768 ( \8083 , \8066 , \8082 );
and \U$7769 ( \8084 , \3889 , \1360 );
and \U$7770 ( \8085 , \3681 , \1358 );
nor \U$7771 ( \8086 , \8084 , \8085 );
xnor \U$7772 ( \8087 , \8086 , \1224 );
and \U$7773 ( \8088 , \4016 , \1160 );
and \U$7774 ( \8089 , \4011 , \1158 );
nor \U$7775 ( \8090 , \8088 , \8089 );
xnor \U$7776 ( \8091 , \8090 , \1082 );
and \U$7777 ( \8092 , \8087 , \8091 );
and \U$7778 ( \8093 , \4469 , \996 );
and \U$7779 ( \8094 , \4272 , \994 );
nor \U$7780 ( \8095 , \8093 , \8094 );
xnor \U$7781 ( \8096 , \8095 , \902 );
and \U$7782 ( \8097 , \8091 , \8096 );
and \U$7783 ( \8098 , \8087 , \8096 );
or \U$7784 ( \8099 , \8092 , \8097 , \8098 );
and \U$7785 ( \8100 , \8082 , \8099 );
and \U$7786 ( \8101 , \8066 , \8099 );
or \U$7787 ( \8102 , \8083 , \8100 , \8101 );
and \U$7788 ( \8103 , \8049 , \8102 );
and \U$7789 ( \8104 , \7995 , \8102 );
or \U$7790 ( \8105 , \8050 , \8103 , \8104 );
xor \U$7791 ( \8106 , \7681 , \7685 );
xor \U$7792 ( \8107 , \8106 , \7690 );
xor \U$7793 ( \8108 , \7790 , \7794 );
xor \U$7794 ( \8109 , \8108 , \7799 );
and \U$7795 ( \8110 , \8107 , \8109 );
xor \U$7796 ( \8111 , \7715 , \7719 );
xor \U$7797 ( \8112 , \8111 , \7724 );
and \U$7798 ( \8113 , \8109 , \8112 );
and \U$7799 ( \8114 , \8107 , \8112 );
or \U$7800 ( \8115 , \8110 , \8113 , \8114 );
xor \U$7801 ( \8116 , \7750 , \7754 );
xor \U$7802 ( \8117 , \8116 , \7759 );
xor \U$7803 ( \8118 , \7806 , \7810 );
xor \U$7804 ( \8119 , \8118 , \7815 );
and \U$7805 ( \8120 , \8117 , \8119 );
xor \U$7806 ( \8121 , \7823 , \7827 );
xor \U$7807 ( \8122 , \8121 , \7832 );
and \U$7808 ( \8123 , \8119 , \8122 );
and \U$7809 ( \8124 , \8117 , \8122 );
or \U$7810 ( \8125 , \8120 , \8123 , \8124 );
and \U$7811 ( \8126 , \8115 , \8125 );
buf \U$7812 ( \8127 , RIc0c6078_119);
and \U$7813 ( \8128 , \8127 , \317 );
xor \U$7814 ( \8129 , \7697 , \7701 );
xor \U$7815 ( \8130 , \8129 , \7707 );
or \U$7816 ( \8131 , \8128 , \8130 );
and \U$7817 ( \8132 , \8125 , \8131 );
and \U$7818 ( \8133 , \8115 , \8131 );
or \U$7819 ( \8134 , \8126 , \8132 , \8133 );
and \U$7820 ( \8135 , \8105 , \8134 );
xor \U$7821 ( \8136 , \7519 , \7523 );
xor \U$7822 ( \8137 , \8136 , \7528 );
xor \U$7823 ( \8138 , \7843 , \7845 );
xor \U$7824 ( \8139 , \8138 , \7848 );
and \U$7825 ( \8140 , \8137 , \8139 );
xor \U$7826 ( \8141 , \7863 , \7865 );
xor \U$7827 ( \8142 , \8141 , \7868 );
and \U$7828 ( \8143 , \8139 , \8142 );
and \U$7829 ( \8144 , \8137 , \8142 );
or \U$7830 ( \8145 , \8140 , \8143 , \8144 );
and \U$7831 ( \8146 , \8134 , \8145 );
and \U$7832 ( \8147 , \8105 , \8145 );
or \U$7833 ( \8148 , \8135 , \8146 , \8147 );
xor \U$7834 ( \8149 , \7730 , \7785 );
xor \U$7835 ( \8150 , \8149 , \7838 );
xor \U$7836 ( \8151 , \7851 , \7860 );
xor \U$7837 ( \8152 , \8151 , \7871 );
and \U$7838 ( \8153 , \8150 , \8152 );
xor \U$7839 ( \8154 , \7877 , \7879 );
xor \U$7840 ( \8155 , \8154 , \7882 );
and \U$7841 ( \8156 , \8152 , \8155 );
and \U$7842 ( \8157 , \8150 , \8155 );
or \U$7843 ( \8158 , \8153 , \8156 , \8157 );
and \U$7844 ( \8159 , \8148 , \8158 );
xor \U$7845 ( \8160 , \7693 , \7710 );
xor \U$7846 ( \8161 , \8160 , \7727 );
xor \U$7847 ( \8162 , \7802 , \7818 );
xor \U$7848 ( \8163 , \8162 , \7835 );
and \U$7849 ( \8164 , \8161 , \8163 );
xor \U$7850 ( \8165 , \7852 , \7854 );
xor \U$7851 ( \8166 , \8165 , \7857 );
and \U$7852 ( \8167 , \8163 , \8166 );
and \U$7853 ( \8168 , \8161 , \8166 );
or \U$7854 ( \8169 , \8164 , \8167 , \8168 );
xor \U$7855 ( \8170 , \7513 , \7531 );
xor \U$7856 ( \8171 , \8170 , \7548 );
and \U$7857 ( \8172 , \8169 , \8171 );
xor \U$7858 ( \8173 , \7890 , \7892 );
xor \U$7859 ( \8174 , \8173 , \7894 );
and \U$7860 ( \8175 , \8171 , \8174 );
and \U$7861 ( \8176 , \8169 , \8174 );
or \U$7862 ( \8177 , \8172 , \8175 , \8176 );
and \U$7863 ( \8178 , \8158 , \8177 );
and \U$7864 ( \8179 , \8148 , \8177 );
or \U$7865 ( \8180 , \8159 , \8178 , \8179 );
xor \U$7866 ( \8181 , \7841 , \7874 );
xor \U$7867 ( \8182 , \8181 , \7885 );
xor \U$7868 ( \8183 , \7897 , \7899 );
xor \U$7869 ( \8184 , \8183 , \7902 );
and \U$7870 ( \8185 , \8182 , \8184 );
xor \U$7871 ( \8186 , \7908 , \7910 );
and \U$7872 ( \8187 , \8184 , \8186 );
and \U$7873 ( \8188 , \8182 , \8186 );
or \U$7874 ( \8189 , \8185 , \8187 , \8188 );
and \U$7875 ( \8190 , \8180 , \8189 );
xor \U$7876 ( \8191 , \7916 , \7918 );
xor \U$7877 ( \8192 , \8191 , \7920 );
and \U$7878 ( \8193 , \8189 , \8192 );
and \U$7879 ( \8194 , \8180 , \8192 );
or \U$7880 ( \8195 , \8190 , \8193 , \8194 );
xor \U$7881 ( \8196 , \7621 , \7639 );
xor \U$7882 ( \8197 , \8196 , \7645 );
and \U$7883 ( \8198 , \8195 , \8197 );
xor \U$7884 ( \8199 , \7914 , \7923 );
xor \U$7885 ( \8200 , \8199 , \7926 );
and \U$7886 ( \8201 , \8197 , \8200 );
and \U$7887 ( \8202 , \8195 , \8200 );
or \U$7888 ( \8203 , \8198 , \8201 , \8202 );
xor \U$7889 ( \8204 , \7929 , \7931 );
xor \U$7890 ( \8205 , \8204 , \7934 );
and \U$7891 ( \8206 , \8203 , \8205 );
and \U$7892 ( \8207 , \7943 , \8206 );
xor \U$7893 ( \8208 , \7943 , \8206 );
xor \U$7894 ( \8209 , \8203 , \8205 );
and \U$7895 ( \8210 , \2042 , \2918 );
and \U$7896 ( \8211 , \1799 , \2916 );
nor \U$7897 ( \8212 , \8210 , \8211 );
xnor \U$7898 ( \8213 , \8212 , \2769 );
and \U$7899 ( \8214 , \2233 , \2596 );
and \U$7900 ( \8215 , \2047 , \2594 );
nor \U$7901 ( \8216 , \8214 , \8215 );
xnor \U$7902 ( \8217 , \8216 , \2454 );
and \U$7903 ( \8218 , \8213 , \8217 );
and \U$7904 ( \8219 , \2641 , \2300 );
and \U$7905 ( \8220 , \2377 , \2298 );
nor \U$7906 ( \8221 , \8219 , \8220 );
xnor \U$7907 ( \8222 , \8221 , \2163 );
and \U$7908 ( \8223 , \8217 , \8222 );
and \U$7909 ( \8224 , \8213 , \8222 );
or \U$7910 ( \8225 , \8218 , \8223 , \8224 );
and \U$7911 ( \8226 , \2840 , \2094 );
and \U$7912 ( \8227 , \2666 , \2092 );
nor \U$7913 ( \8228 , \8226 , \8227 );
xnor \U$7914 ( \8229 , \8228 , \1942 );
and \U$7915 ( \8230 , \3145 , \1826 );
and \U$7916 ( \8231 , \3007 , \1824 );
nor \U$7917 ( \8232 , \8230 , \8231 );
xnor \U$7918 ( \8233 , \8232 , \1670 );
and \U$7919 ( \8234 , \8229 , \8233 );
and \U$7920 ( \8235 , \3681 , \1554 );
and \U$7921 ( \8236 , \3264 , \1552 );
nor \U$7922 ( \8237 , \8235 , \8236 );
xnor \U$7923 ( \8238 , \8237 , \1441 );
and \U$7924 ( \8239 , \8233 , \8238 );
and \U$7925 ( \8240 , \8229 , \8238 );
or \U$7926 ( \8241 , \8234 , \8239 , \8240 );
and \U$7927 ( \8242 , \8225 , \8241 );
and \U$7928 ( \8243 , \1379 , \4032 );
and \U$7929 ( \8244 , \1274 , \4030 );
nor \U$7930 ( \8245 , \8243 , \8244 );
xnor \U$7931 ( \8246 , \8245 , \3786 );
and \U$7932 ( \8247 , \1500 , \3637 );
and \U$7933 ( \8248 , \1384 , \3635 );
nor \U$7934 ( \8249 , \8247 , \8248 );
xnor \U$7935 ( \8250 , \8249 , \3450 );
and \U$7936 ( \8251 , \8246 , \8250 );
and \U$7937 ( \8252 , \1791 , \3324 );
and \U$7938 ( \8253 , \1615 , \3322 );
nor \U$7939 ( \8254 , \8252 , \8253 );
xnor \U$7940 ( \8255 , \8254 , \3119 );
and \U$7941 ( \8256 , \8250 , \8255 );
and \U$7942 ( \8257 , \8246 , \8255 );
or \U$7943 ( \8258 , \8251 , \8256 , \8257 );
and \U$7944 ( \8259 , \8241 , \8258 );
and \U$7945 ( \8260 , \8225 , \8258 );
or \U$7946 ( \8261 , \8242 , \8259 , \8260 );
and \U$7947 ( \8262 , \5248 , \826 );
and \U$7948 ( \8263 , \4779 , \824 );
nor \U$7949 ( \8264 , \8262 , \8263 );
xnor \U$7950 ( \8265 , \8264 , \754 );
and \U$7951 ( \8266 , \5517 , \692 );
and \U$7952 ( \8267 , \5253 , \690 );
nor \U$7953 ( \8268 , \8266 , \8267 );
xnor \U$7954 ( \8269 , \8268 , \649 );
and \U$7955 ( \8270 , \8265 , \8269 );
and \U$7956 ( \8271 , \6148 , \579 );
and \U$7957 ( \8272 , \5776 , \577 );
nor \U$7958 ( \8273 , \8271 , \8272 );
xnor \U$7959 ( \8274 , \8273 , \530 );
and \U$7960 ( \8275 , \8269 , \8274 );
and \U$7961 ( \8276 , \8265 , \8274 );
or \U$7962 ( \8277 , \8270 , \8275 , \8276 );
and \U$7963 ( \8278 , \4011 , \1360 );
and \U$7964 ( \8279 , \3889 , \1358 );
nor \U$7965 ( \8280 , \8278 , \8279 );
xnor \U$7966 ( \8281 , \8280 , \1224 );
and \U$7967 ( \8282 , \4272 , \1160 );
and \U$7968 ( \8283 , \4016 , \1158 );
nor \U$7969 ( \8284 , \8282 , \8283 );
xnor \U$7970 ( \8285 , \8284 , \1082 );
and \U$7971 ( \8286 , \8281 , \8285 );
and \U$7972 ( \8287 , \4771 , \996 );
and \U$7973 ( \8288 , \4469 , \994 );
nor \U$7974 ( \8289 , \8287 , \8288 );
xnor \U$7975 ( \8290 , \8289 , \902 );
and \U$7976 ( \8291 , \8285 , \8290 );
and \U$7977 ( \8292 , \8281 , \8290 );
or \U$7978 ( \8293 , \8286 , \8291 , \8292 );
and \U$7979 ( \8294 , \8277 , \8293 );
and \U$7980 ( \8295 , \6500 , \478 );
and \U$7981 ( \8296 , \6157 , \476 );
nor \U$7982 ( \8297 , \8295 , \8296 );
xnor \U$7983 ( \8298 , \8297 , \437 );
and \U$7984 ( \8299 , \7005 , \408 );
and \U$7985 ( \8300 , \6702 , \406 );
nor \U$7986 ( \8301 , \8299 , \8300 );
xnor \U$7987 ( \8302 , \8301 , \378 );
and \U$7988 ( \8303 , \8298 , \8302 );
and \U$7989 ( \8304 , \7703 , \360 );
and \U$7990 ( \8305 , \7177 , \358 );
nor \U$7991 ( \8306 , \8304 , \8305 );
xnor \U$7992 ( \8307 , \8306 , \341 );
and \U$7993 ( \8308 , \8302 , \8307 );
and \U$7994 ( \8309 , \8298 , \8307 );
or \U$7995 ( \8310 , \8303 , \8308 , \8309 );
and \U$7996 ( \8311 , \8293 , \8310 );
and \U$7997 ( \8312 , \8277 , \8310 );
or \U$7998 ( \8313 , \8294 , \8311 , \8312 );
and \U$7999 ( \8314 , \8261 , \8313 );
and \U$8000 ( \8315 , \789 , \5180 );
and \U$8001 ( \8316 , \709 , \5178 );
nor \U$8002 ( \8317 , \8315 , \8316 );
xnor \U$8003 ( \8318 , \8317 , \4992 );
and \U$8004 ( \8319 , \925 , \4806 );
and \U$8005 ( \8320 , \863 , \4804 );
nor \U$8006 ( \8321 , \8319 , \8320 );
xnor \U$8007 ( \8322 , \8321 , \4574 );
and \U$8008 ( \8323 , \8318 , \8322 );
and \U$8009 ( \8324 , \1186 , \4355 );
and \U$8010 ( \8325 , \988 , \4353 );
nor \U$8011 ( \8326 , \8324 , \8325 );
xnor \U$8012 ( \8327 , \8326 , \4212 );
and \U$8013 ( \8328 , \8322 , \8327 );
and \U$8014 ( \8329 , \8318 , \8327 );
or \U$8015 ( \8330 , \8323 , \8328 , \8329 );
xor \U$8016 ( \8331 , \7515 , \8012 );
xor \U$8017 ( \8332 , \8012 , \8013 );
not \U$8018 ( \8333 , \8332 );
and \U$8019 ( \8334 , \8331 , \8333 );
and \U$8020 ( \8335 , \316 , \8334 );
not \U$8021 ( \8336 , \8335 );
xnor \U$8022 ( \8337 , \8336 , \8016 );
and \U$8023 ( \8338 , \348 , \7767 );
and \U$8024 ( \8339 , \330 , \7765 );
nor \U$8025 ( \8340 , \8338 , \8339 );
xnor \U$8026 ( \8341 , \8340 , \7518 );
and \U$8027 ( \8342 , \8337 , \8341 );
and \U$8028 ( \8343 , \417 , \7238 );
and \U$8029 ( \8344 , \369 , \7236 );
nor \U$8030 ( \8345 , \8343 , \8344 );
xnor \U$8031 ( \8346 , \8345 , \6978 );
and \U$8032 ( \8347 , \8341 , \8346 );
and \U$8033 ( \8348 , \8337 , \8346 );
or \U$8034 ( \8349 , \8342 , \8347 , \8348 );
and \U$8035 ( \8350 , \8330 , \8349 );
and \U$8036 ( \8351 , \494 , \6744 );
and \U$8037 ( \8352 , \425 , \6742 );
nor \U$8038 ( \8353 , \8351 , \8352 );
xnor \U$8039 ( \8354 , \8353 , \6429 );
and \U$8040 ( \8355 , \553 , \6235 );
and \U$8041 ( \8356 , \499 , \6233 );
nor \U$8042 ( \8357 , \8355 , \8356 );
xnor \U$8043 ( \8358 , \8357 , \5895 );
and \U$8044 ( \8359 , \8354 , \8358 );
and \U$8045 ( \8360 , \681 , \5646 );
and \U$8046 ( \8361 , \604 , \5644 );
nor \U$8047 ( \8362 , \8360 , \8361 );
xnor \U$8048 ( \8363 , \8362 , \5405 );
and \U$8049 ( \8364 , \8358 , \8363 );
and \U$8050 ( \8365 , \8354 , \8363 );
or \U$8051 ( \8366 , \8359 , \8364 , \8365 );
and \U$8052 ( \8367 , \8349 , \8366 );
and \U$8053 ( \8368 , \8330 , \8366 );
or \U$8054 ( \8369 , \8350 , \8367 , \8368 );
and \U$8055 ( \8370 , \8313 , \8369 );
and \U$8056 ( \8371 , \8261 , \8369 );
or \U$8057 ( \8372 , \8314 , \8370 , \8371 );
buf \U$8058 ( \8373 , RIc0c6000_120);
and \U$8059 ( \8374 , \8373 , \323 );
and \U$8060 ( \8375 , \8127 , \321 );
nor \U$8061 ( \8376 , \8374 , \8375 );
xnor \U$8062 ( \8377 , \8376 , \328 );
buf \U$8063 ( \8378 , RIc0c5f88_121);
and \U$8064 ( \8379 , \8378 , \317 );
or \U$8065 ( \8380 , \8377 , \8379 );
and \U$8066 ( \8381 , \8127 , \323 );
and \U$8067 ( \8382 , \7703 , \321 );
nor \U$8068 ( \8383 , \8381 , \8382 );
xnor \U$8069 ( \8384 , \8383 , \328 );
and \U$8070 ( \8385 , \8380 , \8384 );
and \U$8071 ( \8386 , \8373 , \317 );
and \U$8072 ( \8387 , \8384 , \8386 );
and \U$8073 ( \8388 , \8380 , \8386 );
or \U$8074 ( \8389 , \8385 , \8387 , \8388 );
xor \U$8075 ( \8390 , \8054 , \8058 );
xor \U$8076 ( \8391 , \8390 , \8063 );
xor \U$8077 ( \8392 , \8070 , \8074 );
xor \U$8078 ( \8393 , \8392 , \8079 );
and \U$8079 ( \8394 , \8391 , \8393 );
xor \U$8080 ( \8395 , \8087 , \8091 );
xor \U$8081 ( \8396 , \8395 , \8096 );
and \U$8082 ( \8397 , \8393 , \8396 );
and \U$8083 ( \8398 , \8391 , \8396 );
or \U$8084 ( \8399 , \8394 , \8397 , \8398 );
and \U$8085 ( \8400 , \8389 , \8399 );
xor \U$8086 ( \8401 , \7947 , \7951 );
xor \U$8087 ( \8402 , \8401 , \7956 );
xor \U$8088 ( \8403 , \7963 , \7967 );
xor \U$8089 ( \8404 , \8403 , \7972 );
and \U$8090 ( \8405 , \8402 , \8404 );
xor \U$8091 ( \8406 , \7980 , \7984 );
xor \U$8092 ( \8407 , \8406 , \7989 );
and \U$8093 ( \8408 , \8404 , \8407 );
and \U$8094 ( \8409 , \8402 , \8407 );
or \U$8095 ( \8410 , \8405 , \8408 , \8409 );
and \U$8096 ( \8411 , \8399 , \8410 );
and \U$8097 ( \8412 , \8389 , \8410 );
or \U$8098 ( \8413 , \8400 , \8411 , \8412 );
and \U$8099 ( \8414 , \8372 , \8413 );
xor \U$8100 ( \8415 , \7999 , \8003 );
xor \U$8101 ( \8416 , \8415 , \8008 );
xor \U$8102 ( \8417 , \8017 , \8021 );
xor \U$8103 ( \8418 , \8417 , \8026 );
and \U$8104 ( \8419 , \8416 , \8418 );
xor \U$8105 ( \8420 , \8034 , \8038 );
xor \U$8106 ( \8421 , \8420 , \8043 );
and \U$8107 ( \8422 , \8418 , \8421 );
and \U$8108 ( \8423 , \8416 , \8421 );
or \U$8109 ( \8424 , \8419 , \8422 , \8423 );
xor \U$8110 ( \8425 , \7734 , \7738 );
xor \U$8111 ( \8426 , \8425 , \7743 );
and \U$8112 ( \8427 , \8424 , \8426 );
xor \U$8113 ( \8428 , \7770 , \7774 );
xor \U$8114 ( \8429 , \8428 , \7779 );
and \U$8115 ( \8430 , \8426 , \8429 );
and \U$8116 ( \8431 , \8424 , \8429 );
or \U$8117 ( \8432 , \8427 , \8430 , \8431 );
and \U$8118 ( \8433 , \8413 , \8432 );
and \U$8119 ( \8434 , \8372 , \8432 );
or \U$8120 ( \8435 , \8414 , \8433 , \8434 );
xor \U$8121 ( \8436 , \7959 , \7975 );
xor \U$8122 ( \8437 , \8436 , \7992 );
xor \U$8123 ( \8438 , \8011 , \8029 );
xor \U$8124 ( \8439 , \8438 , \8046 );
and \U$8125 ( \8440 , \8437 , \8439 );
xor \U$8126 ( \8441 , \8066 , \8082 );
xor \U$8127 ( \8442 , \8441 , \8099 );
and \U$8128 ( \8443 , \8439 , \8442 );
and \U$8129 ( \8444 , \8437 , \8442 );
or \U$8130 ( \8445 , \8440 , \8443 , \8444 );
xor \U$8131 ( \8446 , \8107 , \8109 );
xor \U$8132 ( \8447 , \8446 , \8112 );
xor \U$8133 ( \8448 , \8117 , \8119 );
xor \U$8134 ( \8449 , \8448 , \8122 );
and \U$8135 ( \8450 , \8447 , \8449 );
xnor \U$8136 ( \8451 , \8128 , \8130 );
and \U$8137 ( \8452 , \8449 , \8451 );
and \U$8138 ( \8453 , \8447 , \8451 );
or \U$8139 ( \8454 , \8450 , \8452 , \8453 );
and \U$8140 ( \8455 , \8445 , \8454 );
xor \U$8141 ( \8456 , \7746 , \7762 );
xor \U$8142 ( \8457 , \8456 , \7782 );
and \U$8143 ( \8458 , \8454 , \8457 );
and \U$8144 ( \8459 , \8445 , \8457 );
or \U$8145 ( \8460 , \8455 , \8458 , \8459 );
and \U$8146 ( \8461 , \8435 , \8460 );
xor \U$8147 ( \8462 , \8115 , \8125 );
xor \U$8148 ( \8463 , \8462 , \8131 );
xor \U$8149 ( \8464 , \8161 , \8163 );
xor \U$8150 ( \8465 , \8464 , \8166 );
and \U$8151 ( \8466 , \8463 , \8465 );
xor \U$8152 ( \8467 , \8137 , \8139 );
xor \U$8153 ( \8468 , \8467 , \8142 );
and \U$8154 ( \8469 , \8465 , \8468 );
and \U$8155 ( \8470 , \8463 , \8468 );
or \U$8156 ( \8471 , \8466 , \8469 , \8470 );
and \U$8157 ( \8472 , \8460 , \8471 );
and \U$8158 ( \8473 , \8435 , \8471 );
or \U$8159 ( \8474 , \8461 , \8472 , \8473 );
xor \U$8160 ( \8475 , \8105 , \8134 );
xor \U$8161 ( \8476 , \8475 , \8145 );
xor \U$8162 ( \8477 , \8150 , \8152 );
xor \U$8163 ( \8478 , \8477 , \8155 );
and \U$8164 ( \8479 , \8476 , \8478 );
xor \U$8165 ( \8480 , \8169 , \8171 );
xor \U$8166 ( \8481 , \8480 , \8174 );
and \U$8167 ( \8482 , \8478 , \8481 );
and \U$8168 ( \8483 , \8476 , \8481 );
or \U$8169 ( \8484 , \8479 , \8482 , \8483 );
and \U$8170 ( \8485 , \8474 , \8484 );
xor \U$8171 ( \8486 , \8182 , \8184 );
xor \U$8172 ( \8487 , \8486 , \8186 );
and \U$8173 ( \8488 , \8484 , \8487 );
and \U$8174 ( \8489 , \8474 , \8487 );
or \U$8175 ( \8490 , \8485 , \8488 , \8489 );
xor \U$8176 ( \8491 , \7888 , \7905 );
xor \U$8177 ( \8492 , \8491 , \7911 );
and \U$8178 ( \8493 , \8490 , \8492 );
xor \U$8179 ( \8494 , \8180 , \8189 );
xor \U$8180 ( \8495 , \8494 , \8192 );
and \U$8181 ( \8496 , \8492 , \8495 );
and \U$8182 ( \8497 , \8490 , \8495 );
or \U$8183 ( \8498 , \8493 , \8496 , \8497 );
xor \U$8184 ( \8499 , \8195 , \8197 );
xor \U$8185 ( \8500 , \8499 , \8200 );
and \U$8186 ( \8501 , \8498 , \8500 );
and \U$8187 ( \8502 , \8209 , \8501 );
xor \U$8188 ( \8503 , \8209 , \8501 );
xor \U$8189 ( \8504 , \8498 , \8500 );
and \U$8190 ( \8505 , \425 , \7238 );
and \U$8191 ( \8506 , \417 , \7236 );
nor \U$8192 ( \8507 , \8505 , \8506 );
xnor \U$8193 ( \8508 , \8507 , \6978 );
and \U$8194 ( \8509 , \499 , \6744 );
and \U$8195 ( \8510 , \494 , \6742 );
nor \U$8196 ( \8511 , \8509 , \8510 );
xnor \U$8197 ( \8512 , \8511 , \6429 );
and \U$8198 ( \8513 , \8508 , \8512 );
and \U$8199 ( \8514 , \604 , \6235 );
and \U$8200 ( \8515 , \553 , \6233 );
nor \U$8201 ( \8516 , \8514 , \8515 );
xnor \U$8202 ( \8517 , \8516 , \5895 );
and \U$8203 ( \8518 , \8512 , \8517 );
and \U$8204 ( \8519 , \8508 , \8517 );
or \U$8205 ( \8520 , \8513 , \8518 , \8519 );
buf \U$8206 ( \8521 , RIc0c7c98_59);
buf \U$8207 ( \8522 , RIc0c7c20_60);
and \U$8208 ( \8523 , \8521 , \8522 );
not \U$8209 ( \8524 , \8523 );
and \U$8210 ( \8525 , \8013 , \8524 );
not \U$8211 ( \8526 , \8525 );
and \U$8212 ( \8527 , \330 , \8334 );
and \U$8213 ( \8528 , \316 , \8332 );
nor \U$8214 ( \8529 , \8527 , \8528 );
xnor \U$8215 ( \8530 , \8529 , \8016 );
and \U$8216 ( \8531 , \8526 , \8530 );
and \U$8217 ( \8532 , \369 , \7767 );
and \U$8218 ( \8533 , \348 , \7765 );
nor \U$8219 ( \8534 , \8532 , \8533 );
xnor \U$8220 ( \8535 , \8534 , \7518 );
and \U$8221 ( \8536 , \8530 , \8535 );
and \U$8222 ( \8537 , \8526 , \8535 );
or \U$8223 ( \8538 , \8531 , \8536 , \8537 );
and \U$8224 ( \8539 , \8520 , \8538 );
and \U$8225 ( \8540 , \709 , \5646 );
and \U$8226 ( \8541 , \681 , \5644 );
nor \U$8227 ( \8542 , \8540 , \8541 );
xnor \U$8228 ( \8543 , \8542 , \5405 );
and \U$8229 ( \8544 , \863 , \5180 );
and \U$8230 ( \8545 , \789 , \5178 );
nor \U$8231 ( \8546 , \8544 , \8545 );
xnor \U$8232 ( \8547 , \8546 , \4992 );
and \U$8233 ( \8548 , \8543 , \8547 );
and \U$8234 ( \8549 , \988 , \4806 );
and \U$8235 ( \8550 , \925 , \4804 );
nor \U$8236 ( \8551 , \8549 , \8550 );
xnor \U$8237 ( \8552 , \8551 , \4574 );
and \U$8238 ( \8553 , \8547 , \8552 );
and \U$8239 ( \8554 , \8543 , \8552 );
or \U$8240 ( \8555 , \8548 , \8553 , \8554 );
and \U$8241 ( \8556 , \8538 , \8555 );
and \U$8242 ( \8557 , \8520 , \8555 );
or \U$8243 ( \8558 , \8539 , \8556 , \8557 );
and \U$8244 ( \8559 , \2666 , \2300 );
and \U$8245 ( \8560 , \2641 , \2298 );
nor \U$8246 ( \8561 , \8559 , \8560 );
xnor \U$8247 ( \8562 , \8561 , \2163 );
and \U$8248 ( \8563 , \3007 , \2094 );
and \U$8249 ( \8564 , \2840 , \2092 );
nor \U$8250 ( \8565 , \8563 , \8564 );
xnor \U$8251 ( \8566 , \8565 , \1942 );
and \U$8252 ( \8567 , \8562 , \8566 );
and \U$8253 ( \8568 , \3264 , \1826 );
and \U$8254 ( \8569 , \3145 , \1824 );
nor \U$8255 ( \8570 , \8568 , \8569 );
xnor \U$8256 ( \8571 , \8570 , \1670 );
and \U$8257 ( \8572 , \8566 , \8571 );
and \U$8258 ( \8573 , \8562 , \8571 );
or \U$8259 ( \8574 , \8567 , \8572 , \8573 );
and \U$8260 ( \8575 , \1799 , \3324 );
and \U$8261 ( \8576 , \1791 , \3322 );
nor \U$8262 ( \8577 , \8575 , \8576 );
xnor \U$8263 ( \8578 , \8577 , \3119 );
and \U$8264 ( \8579 , \2047 , \2918 );
and \U$8265 ( \8580 , \2042 , \2916 );
nor \U$8266 ( \8581 , \8579 , \8580 );
xnor \U$8267 ( \8582 , \8581 , \2769 );
and \U$8268 ( \8583 , \8578 , \8582 );
and \U$8269 ( \8584 , \2377 , \2596 );
and \U$8270 ( \8585 , \2233 , \2594 );
nor \U$8271 ( \8586 , \8584 , \8585 );
xnor \U$8272 ( \8587 , \8586 , \2454 );
and \U$8273 ( \8588 , \8582 , \8587 );
and \U$8274 ( \8589 , \8578 , \8587 );
or \U$8275 ( \8590 , \8583 , \8588 , \8589 );
and \U$8276 ( \8591 , \8574 , \8590 );
and \U$8277 ( \8592 , \1274 , \4355 );
and \U$8278 ( \8593 , \1186 , \4353 );
nor \U$8279 ( \8594 , \8592 , \8593 );
xnor \U$8280 ( \8595 , \8594 , \4212 );
and \U$8281 ( \8596 , \1384 , \4032 );
and \U$8282 ( \8597 , \1379 , \4030 );
nor \U$8283 ( \8598 , \8596 , \8597 );
xnor \U$8284 ( \8599 , \8598 , \3786 );
and \U$8285 ( \8600 , \8595 , \8599 );
and \U$8286 ( \8601 , \1615 , \3637 );
and \U$8287 ( \8602 , \1500 , \3635 );
nor \U$8288 ( \8603 , \8601 , \8602 );
xnor \U$8289 ( \8604 , \8603 , \3450 );
and \U$8290 ( \8605 , \8599 , \8604 );
and \U$8291 ( \8606 , \8595 , \8604 );
or \U$8292 ( \8607 , \8600 , \8605 , \8606 );
and \U$8293 ( \8608 , \8590 , \8607 );
and \U$8294 ( \8609 , \8574 , \8607 );
or \U$8295 ( \8610 , \8591 , \8608 , \8609 );
and \U$8296 ( \8611 , \8558 , \8610 );
and \U$8297 ( \8612 , \4779 , \996 );
and \U$8298 ( \8613 , \4771 , \994 );
nor \U$8299 ( \8614 , \8612 , \8613 );
xnor \U$8300 ( \8615 , \8614 , \902 );
and \U$8301 ( \8616 , \5253 , \826 );
and \U$8302 ( \8617 , \5248 , \824 );
nor \U$8303 ( \8618 , \8616 , \8617 );
xnor \U$8304 ( \8619 , \8618 , \754 );
and \U$8305 ( \8620 , \8615 , \8619 );
and \U$8306 ( \8621 , \5776 , \692 );
and \U$8307 ( \8622 , \5517 , \690 );
nor \U$8308 ( \8623 , \8621 , \8622 );
xnor \U$8309 ( \8624 , \8623 , \649 );
and \U$8310 ( \8625 , \8619 , \8624 );
and \U$8311 ( \8626 , \8615 , \8624 );
or \U$8312 ( \8627 , \8620 , \8625 , \8626 );
and \U$8313 ( \8628 , \3889 , \1554 );
and \U$8314 ( \8629 , \3681 , \1552 );
nor \U$8315 ( \8630 , \8628 , \8629 );
xnor \U$8316 ( \8631 , \8630 , \1441 );
and \U$8317 ( \8632 , \4016 , \1360 );
and \U$8318 ( \8633 , \4011 , \1358 );
nor \U$8319 ( \8634 , \8632 , \8633 );
xnor \U$8320 ( \8635 , \8634 , \1224 );
and \U$8321 ( \8636 , \8631 , \8635 );
and \U$8322 ( \8637 , \4469 , \1160 );
and \U$8323 ( \8638 , \4272 , \1158 );
nor \U$8324 ( \8639 , \8637 , \8638 );
xnor \U$8325 ( \8640 , \8639 , \1082 );
and \U$8326 ( \8641 , \8635 , \8640 );
and \U$8327 ( \8642 , \8631 , \8640 );
or \U$8328 ( \8643 , \8636 , \8641 , \8642 );
and \U$8329 ( \8644 , \8627 , \8643 );
and \U$8330 ( \8645 , \6157 , \579 );
and \U$8331 ( \8646 , \6148 , \577 );
nor \U$8332 ( \8647 , \8645 , \8646 );
xnor \U$8333 ( \8648 , \8647 , \530 );
and \U$8334 ( \8649 , \6702 , \478 );
and \U$8335 ( \8650 , \6500 , \476 );
nor \U$8336 ( \8651 , \8649 , \8650 );
xnor \U$8337 ( \8652 , \8651 , \437 );
and \U$8338 ( \8653 , \8648 , \8652 );
and \U$8339 ( \8654 , \7177 , \408 );
and \U$8340 ( \8655 , \7005 , \406 );
nor \U$8341 ( \8656 , \8654 , \8655 );
xnor \U$8342 ( \8657 , \8656 , \378 );
and \U$8343 ( \8658 , \8652 , \8657 );
and \U$8344 ( \8659 , \8648 , \8657 );
or \U$8345 ( \8660 , \8653 , \8658 , \8659 );
and \U$8346 ( \8661 , \8643 , \8660 );
and \U$8347 ( \8662 , \8627 , \8660 );
or \U$8348 ( \8663 , \8644 , \8661 , \8662 );
and \U$8349 ( \8664 , \8610 , \8663 );
and \U$8350 ( \8665 , \8558 , \8663 );
or \U$8351 ( \8666 , \8611 , \8664 , \8665 );
xor \U$8352 ( \8667 , \8213 , \8217 );
xor \U$8353 ( \8668 , \8667 , \8222 );
xor \U$8354 ( \8669 , \8318 , \8322 );
xor \U$8355 ( \8670 , \8669 , \8327 );
and \U$8356 ( \8671 , \8668 , \8670 );
xor \U$8357 ( \8672 , \8246 , \8250 );
xor \U$8358 ( \8673 , \8672 , \8255 );
and \U$8359 ( \8674 , \8670 , \8673 );
and \U$8360 ( \8675 , \8668 , \8673 );
or \U$8361 ( \8676 , \8671 , \8674 , \8675 );
xor \U$8362 ( \8677 , \8229 , \8233 );
xor \U$8363 ( \8678 , \8677 , \8238 );
xor \U$8364 ( \8679 , \8265 , \8269 );
xor \U$8365 ( \8680 , \8679 , \8274 );
and \U$8366 ( \8681 , \8678 , \8680 );
xor \U$8367 ( \8682 , \8281 , \8285 );
xor \U$8368 ( \8683 , \8682 , \8290 );
and \U$8369 ( \8684 , \8680 , \8683 );
and \U$8370 ( \8685 , \8678 , \8683 );
or \U$8371 ( \8686 , \8681 , \8684 , \8685 );
and \U$8372 ( \8687 , \8676 , \8686 );
and \U$8373 ( \8688 , \8127 , \360 );
and \U$8374 ( \8689 , \7703 , \358 );
nor \U$8375 ( \8690 , \8688 , \8689 );
xnor \U$8376 ( \8691 , \8690 , \341 );
and \U$8377 ( \8692 , \8378 , \323 );
and \U$8378 ( \8693 , \8373 , \321 );
nor \U$8379 ( \8694 , \8692 , \8693 );
xnor \U$8380 ( \8695 , \8694 , \328 );
and \U$8381 ( \8696 , \8691 , \8695 );
buf \U$8382 ( \8697 , RIc0c5f10_122);
and \U$8383 ( \8698 , \8697 , \317 );
and \U$8384 ( \8699 , \8695 , \8698 );
and \U$8385 ( \8700 , \8691 , \8698 );
or \U$8386 ( \8701 , \8696 , \8699 , \8700 );
xor \U$8387 ( \8702 , \8298 , \8302 );
xor \U$8388 ( \8703 , \8702 , \8307 );
and \U$8389 ( \8704 , \8701 , \8703 );
xnor \U$8390 ( \8705 , \8377 , \8379 );
and \U$8391 ( \8706 , \8703 , \8705 );
and \U$8392 ( \8707 , \8701 , \8705 );
or \U$8393 ( \8708 , \8704 , \8706 , \8707 );
and \U$8394 ( \8709 , \8686 , \8708 );
and \U$8395 ( \8710 , \8676 , \8708 );
or \U$8396 ( \8711 , \8687 , \8709 , \8710 );
and \U$8397 ( \8712 , \8666 , \8711 );
xor \U$8398 ( \8713 , \8391 , \8393 );
xor \U$8399 ( \8714 , \8713 , \8396 );
xor \U$8400 ( \8715 , \8402 , \8404 );
xor \U$8401 ( \8716 , \8715 , \8407 );
and \U$8402 ( \8717 , \8714 , \8716 );
xor \U$8403 ( \8718 , \8416 , \8418 );
xor \U$8404 ( \8719 , \8718 , \8421 );
and \U$8405 ( \8720 , \8716 , \8719 );
and \U$8406 ( \8721 , \8714 , \8719 );
or \U$8407 ( \8722 , \8717 , \8720 , \8721 );
and \U$8408 ( \8723 , \8711 , \8722 );
and \U$8409 ( \8724 , \8666 , \8722 );
or \U$8410 ( \8725 , \8712 , \8723 , \8724 );
xor \U$8411 ( \8726 , \8261 , \8313 );
xor \U$8412 ( \8727 , \8726 , \8369 );
xor \U$8413 ( \8728 , \8389 , \8399 );
xor \U$8414 ( \8729 , \8728 , \8410 );
and \U$8415 ( \8730 , \8727 , \8729 );
xor \U$8416 ( \8731 , \8424 , \8426 );
xor \U$8417 ( \8732 , \8731 , \8429 );
and \U$8418 ( \8733 , \8729 , \8732 );
and \U$8419 ( \8734 , \8727 , \8732 );
or \U$8420 ( \8735 , \8730 , \8733 , \8734 );
and \U$8421 ( \8736 , \8725 , \8735 );
xor \U$8422 ( \8737 , \8225 , \8241 );
xor \U$8423 ( \8738 , \8737 , \8258 );
xor \U$8424 ( \8739 , \8277 , \8293 );
xor \U$8425 ( \8740 , \8739 , \8310 );
and \U$8426 ( \8741 , \8738 , \8740 );
xor \U$8427 ( \8742 , \8380 , \8384 );
xor \U$8428 ( \8743 , \8742 , \8386 );
and \U$8429 ( \8744 , \8740 , \8743 );
and \U$8430 ( \8745 , \8738 , \8743 );
or \U$8431 ( \8746 , \8741 , \8744 , \8745 );
xor \U$8432 ( \8747 , \8437 , \8439 );
xor \U$8433 ( \8748 , \8747 , \8442 );
and \U$8434 ( \8749 , \8746 , \8748 );
xor \U$8435 ( \8750 , \8447 , \8449 );
xor \U$8436 ( \8751 , \8750 , \8451 );
and \U$8437 ( \8752 , \8748 , \8751 );
and \U$8438 ( \8753 , \8746 , \8751 );
or \U$8439 ( \8754 , \8749 , \8752 , \8753 );
and \U$8440 ( \8755 , \8735 , \8754 );
and \U$8441 ( \8756 , \8725 , \8754 );
or \U$8442 ( \8757 , \8736 , \8755 , \8756 );
xor \U$8443 ( \8758 , \7995 , \8049 );
xor \U$8444 ( \8759 , \8758 , \8102 );
xor \U$8445 ( \8760 , \8445 , \8454 );
xor \U$8446 ( \8761 , \8760 , \8457 );
and \U$8447 ( \8762 , \8759 , \8761 );
xor \U$8448 ( \8763 , \8463 , \8465 );
xor \U$8449 ( \8764 , \8763 , \8468 );
and \U$8450 ( \8765 , \8761 , \8764 );
and \U$8451 ( \8766 , \8759 , \8764 );
or \U$8452 ( \8767 , \8762 , \8765 , \8766 );
and \U$8453 ( \8768 , \8757 , \8767 );
xor \U$8454 ( \8769 , \8476 , \8478 );
xor \U$8455 ( \8770 , \8769 , \8481 );
and \U$8456 ( \8771 , \8767 , \8770 );
and \U$8457 ( \8772 , \8757 , \8770 );
or \U$8458 ( \8773 , \8768 , \8771 , \8772 );
xor \U$8459 ( \8774 , \8148 , \8158 );
xor \U$8460 ( \8775 , \8774 , \8177 );
and \U$8461 ( \8776 , \8773 , \8775 );
xor \U$8462 ( \8777 , \8474 , \8484 );
xor \U$8463 ( \8778 , \8777 , \8487 );
and \U$8464 ( \8779 , \8775 , \8778 );
and \U$8465 ( \8780 , \8773 , \8778 );
or \U$8466 ( \8781 , \8776 , \8779 , \8780 );
xor \U$8467 ( \8782 , \8490 , \8492 );
xor \U$8468 ( \8783 , \8782 , \8495 );
and \U$8469 ( \8784 , \8781 , \8783 );
and \U$8470 ( \8785 , \8504 , \8784 );
xor \U$8471 ( \8786 , \8504 , \8784 );
xor \U$8472 ( \8787 , \8781 , \8783 );
and \U$8473 ( \8788 , \2840 , \2300 );
and \U$8474 ( \8789 , \2666 , \2298 );
nor \U$8475 ( \8790 , \8788 , \8789 );
xnor \U$8476 ( \8791 , \8790 , \2163 );
and \U$8477 ( \8792 , \3145 , \2094 );
and \U$8478 ( \8793 , \3007 , \2092 );
nor \U$8479 ( \8794 , \8792 , \8793 );
xnor \U$8480 ( \8795 , \8794 , \1942 );
and \U$8481 ( \8796 , \8791 , \8795 );
and \U$8482 ( \8797 , \3681 , \1826 );
and \U$8483 ( \8798 , \3264 , \1824 );
nor \U$8484 ( \8799 , \8797 , \8798 );
xnor \U$8485 ( \8800 , \8799 , \1670 );
and \U$8486 ( \8801 , \8795 , \8800 );
and \U$8487 ( \8802 , \8791 , \8800 );
or \U$8488 ( \8803 , \8796 , \8801 , \8802 );
and \U$8489 ( \8804 , \1379 , \4355 );
and \U$8490 ( \8805 , \1274 , \4353 );
nor \U$8491 ( \8806 , \8804 , \8805 );
xnor \U$8492 ( \8807 , \8806 , \4212 );
and \U$8493 ( \8808 , \1500 , \4032 );
and \U$8494 ( \8809 , \1384 , \4030 );
nor \U$8495 ( \8810 , \8808 , \8809 );
xnor \U$8496 ( \8811 , \8810 , \3786 );
and \U$8497 ( \8812 , \8807 , \8811 );
and \U$8498 ( \8813 , \1791 , \3637 );
and \U$8499 ( \8814 , \1615 , \3635 );
nor \U$8500 ( \8815 , \8813 , \8814 );
xnor \U$8501 ( \8816 , \8815 , \3450 );
and \U$8502 ( \8817 , \8811 , \8816 );
and \U$8503 ( \8818 , \8807 , \8816 );
or \U$8504 ( \8819 , \8812 , \8817 , \8818 );
and \U$8505 ( \8820 , \8803 , \8819 );
and \U$8506 ( \8821 , \2042 , \3324 );
and \U$8507 ( \8822 , \1799 , \3322 );
nor \U$8508 ( \8823 , \8821 , \8822 );
xnor \U$8509 ( \8824 , \8823 , \3119 );
and \U$8510 ( \8825 , \2233 , \2918 );
and \U$8511 ( \8826 , \2047 , \2916 );
nor \U$8512 ( \8827 , \8825 , \8826 );
xnor \U$8513 ( \8828 , \8827 , \2769 );
and \U$8514 ( \8829 , \8824 , \8828 );
and \U$8515 ( \8830 , \2641 , \2596 );
and \U$8516 ( \8831 , \2377 , \2594 );
nor \U$8517 ( \8832 , \8830 , \8831 );
xnor \U$8518 ( \8833 , \8832 , \2454 );
and \U$8519 ( \8834 , \8828 , \8833 );
and \U$8520 ( \8835 , \8824 , \8833 );
or \U$8521 ( \8836 , \8829 , \8834 , \8835 );
and \U$8522 ( \8837 , \8819 , \8836 );
and \U$8523 ( \8838 , \8803 , \8836 );
or \U$8524 ( \8839 , \8820 , \8837 , \8838 );
and \U$8525 ( \8840 , \6500 , \579 );
and \U$8526 ( \8841 , \6157 , \577 );
nor \U$8527 ( \8842 , \8840 , \8841 );
xnor \U$8528 ( \8843 , \8842 , \530 );
and \U$8529 ( \8844 , \7005 , \478 );
and \U$8530 ( \8845 , \6702 , \476 );
nor \U$8531 ( \8846 , \8844 , \8845 );
xnor \U$8532 ( \8847 , \8846 , \437 );
and \U$8533 ( \8848 , \8843 , \8847 );
and \U$8534 ( \8849 , \7703 , \408 );
and \U$8535 ( \8850 , \7177 , \406 );
nor \U$8536 ( \8851 , \8849 , \8850 );
xnor \U$8537 ( \8852 , \8851 , \378 );
and \U$8538 ( \8853 , \8847 , \8852 );
and \U$8539 ( \8854 , \8843 , \8852 );
or \U$8540 ( \8855 , \8848 , \8853 , \8854 );
and \U$8541 ( \8856 , \5248 , \996 );
and \U$8542 ( \8857 , \4779 , \994 );
nor \U$8543 ( \8858 , \8856 , \8857 );
xnor \U$8544 ( \8859 , \8858 , \902 );
and \U$8545 ( \8860 , \5517 , \826 );
and \U$8546 ( \8861 , \5253 , \824 );
nor \U$8547 ( \8862 , \8860 , \8861 );
xnor \U$8548 ( \8863 , \8862 , \754 );
and \U$8549 ( \8864 , \8859 , \8863 );
and \U$8550 ( \8865 , \6148 , \692 );
and \U$8551 ( \8866 , \5776 , \690 );
nor \U$8552 ( \8867 , \8865 , \8866 );
xnor \U$8553 ( \8868 , \8867 , \649 );
and \U$8554 ( \8869 , \8863 , \8868 );
and \U$8555 ( \8870 , \8859 , \8868 );
or \U$8556 ( \8871 , \8864 , \8869 , \8870 );
and \U$8557 ( \8872 , \8855 , \8871 );
and \U$8558 ( \8873 , \4011 , \1554 );
and \U$8559 ( \8874 , \3889 , \1552 );
nor \U$8560 ( \8875 , \8873 , \8874 );
xnor \U$8561 ( \8876 , \8875 , \1441 );
and \U$8562 ( \8877 , \4272 , \1360 );
and \U$8563 ( \8878 , \4016 , \1358 );
nor \U$8564 ( \8879 , \8877 , \8878 );
xnor \U$8565 ( \8880 , \8879 , \1224 );
and \U$8566 ( \8881 , \8876 , \8880 );
and \U$8567 ( \8882 , \4771 , \1160 );
and \U$8568 ( \8883 , \4469 , \1158 );
nor \U$8569 ( \8884 , \8882 , \8883 );
xnor \U$8570 ( \8885 , \8884 , \1082 );
and \U$8571 ( \8886 , \8880 , \8885 );
and \U$8572 ( \8887 , \8876 , \8885 );
or \U$8573 ( \8888 , \8881 , \8886 , \8887 );
and \U$8574 ( \8889 , \8871 , \8888 );
and \U$8575 ( \8890 , \8855 , \8888 );
or \U$8576 ( \8891 , \8872 , \8889 , \8890 );
and \U$8577 ( \8892 , \8839 , \8891 );
xor \U$8578 ( \8893 , \8013 , \8521 );
xor \U$8579 ( \8894 , \8521 , \8522 );
not \U$8580 ( \8895 , \8894 );
and \U$8581 ( \8896 , \8893 , \8895 );
and \U$8582 ( \8897 , \316 , \8896 );
not \U$8583 ( \8898 , \8897 );
xnor \U$8584 ( \8899 , \8898 , \8525 );
and \U$8585 ( \8900 , \348 , \8334 );
and \U$8586 ( \8901 , \330 , \8332 );
nor \U$8587 ( \8902 , \8900 , \8901 );
xnor \U$8588 ( \8903 , \8902 , \8016 );
and \U$8589 ( \8904 , \8899 , \8903 );
and \U$8590 ( \8905 , \417 , \7767 );
and \U$8591 ( \8906 , \369 , \7765 );
nor \U$8592 ( \8907 , \8905 , \8906 );
xnor \U$8593 ( \8908 , \8907 , \7518 );
and \U$8594 ( \8909 , \8903 , \8908 );
and \U$8595 ( \8910 , \8899 , \8908 );
or \U$8596 ( \8911 , \8904 , \8909 , \8910 );
and \U$8597 ( \8912 , \789 , \5646 );
and \U$8598 ( \8913 , \709 , \5644 );
nor \U$8599 ( \8914 , \8912 , \8913 );
xnor \U$8600 ( \8915 , \8914 , \5405 );
and \U$8601 ( \8916 , \925 , \5180 );
and \U$8602 ( \8917 , \863 , \5178 );
nor \U$8603 ( \8918 , \8916 , \8917 );
xnor \U$8604 ( \8919 , \8918 , \4992 );
and \U$8605 ( \8920 , \8915 , \8919 );
and \U$8606 ( \8921 , \1186 , \4806 );
and \U$8607 ( \8922 , \988 , \4804 );
nor \U$8608 ( \8923 , \8921 , \8922 );
xnor \U$8609 ( \8924 , \8923 , \4574 );
and \U$8610 ( \8925 , \8919 , \8924 );
and \U$8611 ( \8926 , \8915 , \8924 );
or \U$8612 ( \8927 , \8920 , \8925 , \8926 );
and \U$8613 ( \8928 , \8911 , \8927 );
and \U$8614 ( \8929 , \494 , \7238 );
and \U$8615 ( \8930 , \425 , \7236 );
nor \U$8616 ( \8931 , \8929 , \8930 );
xnor \U$8617 ( \8932 , \8931 , \6978 );
and \U$8618 ( \8933 , \553 , \6744 );
and \U$8619 ( \8934 , \499 , \6742 );
nor \U$8620 ( \8935 , \8933 , \8934 );
xnor \U$8621 ( \8936 , \8935 , \6429 );
and \U$8622 ( \8937 , \8932 , \8936 );
and \U$8623 ( \8938 , \681 , \6235 );
and \U$8624 ( \8939 , \604 , \6233 );
nor \U$8625 ( \8940 , \8938 , \8939 );
xnor \U$8626 ( \8941 , \8940 , \5895 );
and \U$8627 ( \8942 , \8936 , \8941 );
and \U$8628 ( \8943 , \8932 , \8941 );
or \U$8629 ( \8944 , \8937 , \8942 , \8943 );
and \U$8630 ( \8945 , \8927 , \8944 );
and \U$8631 ( \8946 , \8911 , \8944 );
or \U$8632 ( \8947 , \8928 , \8945 , \8946 );
and \U$8633 ( \8948 , \8891 , \8947 );
and \U$8634 ( \8949 , \8839 , \8947 );
or \U$8635 ( \8950 , \8892 , \8948 , \8949 );
xor \U$8636 ( \8951 , \8543 , \8547 );
xor \U$8637 ( \8952 , \8951 , \8552 );
xor \U$8638 ( \8953 , \8578 , \8582 );
xor \U$8639 ( \8954 , \8953 , \8587 );
and \U$8640 ( \8955 , \8952 , \8954 );
xor \U$8641 ( \8956 , \8595 , \8599 );
xor \U$8642 ( \8957 , \8956 , \8604 );
and \U$8643 ( \8958 , \8954 , \8957 );
and \U$8644 ( \8959 , \8952 , \8957 );
or \U$8645 ( \8960 , \8955 , \8958 , \8959 );
xor \U$8646 ( \8961 , \8562 , \8566 );
xor \U$8647 ( \8962 , \8961 , \8571 );
xor \U$8648 ( \8963 , \8615 , \8619 );
xor \U$8649 ( \8964 , \8963 , \8624 );
and \U$8650 ( \8965 , \8962 , \8964 );
xor \U$8651 ( \8966 , \8631 , \8635 );
xor \U$8652 ( \8967 , \8966 , \8640 );
and \U$8653 ( \8968 , \8964 , \8967 );
and \U$8654 ( \8969 , \8962 , \8967 );
or \U$8655 ( \8970 , \8965 , \8968 , \8969 );
and \U$8656 ( \8971 , \8960 , \8970 );
and \U$8657 ( \8972 , \8373 , \360 );
and \U$8658 ( \8973 , \8127 , \358 );
nor \U$8659 ( \8974 , \8972 , \8973 );
xnor \U$8660 ( \8975 , \8974 , \341 );
and \U$8661 ( \8976 , \8697 , \323 );
and \U$8662 ( \8977 , \8378 , \321 );
nor \U$8663 ( \8978 , \8976 , \8977 );
xnor \U$8664 ( \8979 , \8978 , \328 );
and \U$8665 ( \8980 , \8975 , \8979 );
buf \U$8666 ( \8981 , RIc0c5e98_123);
and \U$8667 ( \8982 , \8981 , \317 );
and \U$8668 ( \8983 , \8979 , \8982 );
and \U$8669 ( \8984 , \8975 , \8982 );
or \U$8670 ( \8985 , \8980 , \8983 , \8984 );
xor \U$8671 ( \8986 , \8691 , \8695 );
xor \U$8672 ( \8987 , \8986 , \8698 );
and \U$8673 ( \8988 , \8985 , \8987 );
xor \U$8674 ( \8989 , \8648 , \8652 );
xor \U$8675 ( \8990 , \8989 , \8657 );
and \U$8676 ( \8991 , \8987 , \8990 );
and \U$8677 ( \8992 , \8985 , \8990 );
or \U$8678 ( \8993 , \8988 , \8991 , \8992 );
and \U$8679 ( \8994 , \8970 , \8993 );
and \U$8680 ( \8995 , \8960 , \8993 );
or \U$8681 ( \8996 , \8971 , \8994 , \8995 );
and \U$8682 ( \8997 , \8950 , \8996 );
xor \U$8683 ( \8998 , \8337 , \8341 );
xor \U$8684 ( \8999 , \8998 , \8346 );
xor \U$8685 ( \9000 , \8354 , \8358 );
xor \U$8686 ( \9001 , \9000 , \8363 );
and \U$8687 ( \9002 , \8999 , \9001 );
xor \U$8688 ( \9003 , \8668 , \8670 );
xor \U$8689 ( \9004 , \9003 , \8673 );
and \U$8690 ( \9005 , \9001 , \9004 );
and \U$8691 ( \9006 , \8999 , \9004 );
or \U$8692 ( \9007 , \9002 , \9005 , \9006 );
and \U$8693 ( \9008 , \8996 , \9007 );
and \U$8694 ( \9009 , \8950 , \9007 );
or \U$8695 ( \9010 , \8997 , \9008 , \9009 );
xor \U$8696 ( \9011 , \8627 , \8643 );
xor \U$8697 ( \9012 , \9011 , \8660 );
xor \U$8698 ( \9013 , \8678 , \8680 );
xor \U$8699 ( \9014 , \9013 , \8683 );
and \U$8700 ( \9015 , \9012 , \9014 );
xor \U$8701 ( \9016 , \8701 , \8703 );
xor \U$8702 ( \9017 , \9016 , \8705 );
and \U$8703 ( \9018 , \9014 , \9017 );
and \U$8704 ( \9019 , \9012 , \9017 );
or \U$8705 ( \9020 , \9015 , \9018 , \9019 );
xor \U$8706 ( \9021 , \8330 , \8349 );
xor \U$8707 ( \9022 , \9021 , \8366 );
and \U$8708 ( \9023 , \9020 , \9022 );
xor \U$8709 ( \9024 , \8738 , \8740 );
xor \U$8710 ( \9025 , \9024 , \8743 );
and \U$8711 ( \9026 , \9022 , \9025 );
and \U$8712 ( \9027 , \9020 , \9025 );
or \U$8713 ( \9028 , \9023 , \9026 , \9027 );
and \U$8714 ( \9029 , \9010 , \9028 );
xor \U$8715 ( \9030 , \8558 , \8610 );
xor \U$8716 ( \9031 , \9030 , \8663 );
xor \U$8717 ( \9032 , \8676 , \8686 );
xor \U$8718 ( \9033 , \9032 , \8708 );
and \U$8719 ( \9034 , \9031 , \9033 );
xor \U$8720 ( \9035 , \8714 , \8716 );
xor \U$8721 ( \9036 , \9035 , \8719 );
and \U$8722 ( \9037 , \9033 , \9036 );
and \U$8723 ( \9038 , \9031 , \9036 );
or \U$8724 ( \9039 , \9034 , \9037 , \9038 );
and \U$8725 ( \9040 , \9028 , \9039 );
and \U$8726 ( \9041 , \9010 , \9039 );
or \U$8727 ( \9042 , \9029 , \9040 , \9041 );
xor \U$8728 ( \9043 , \8666 , \8711 );
xor \U$8729 ( \9044 , \9043 , \8722 );
xor \U$8730 ( \9045 , \8727 , \8729 );
xor \U$8731 ( \9046 , \9045 , \8732 );
and \U$8732 ( \9047 , \9044 , \9046 );
xor \U$8733 ( \9048 , \8746 , \8748 );
xor \U$8734 ( \9049 , \9048 , \8751 );
and \U$8735 ( \9050 , \9046 , \9049 );
and \U$8736 ( \9051 , \9044 , \9049 );
or \U$8737 ( \9052 , \9047 , \9050 , \9051 );
and \U$8738 ( \9053 , \9042 , \9052 );
xor \U$8739 ( \9054 , \8372 , \8413 );
xor \U$8740 ( \9055 , \9054 , \8432 );
and \U$8741 ( \9056 , \9052 , \9055 );
and \U$8742 ( \9057 , \9042 , \9055 );
or \U$8743 ( \9058 , \9053 , \9056 , \9057 );
xor \U$8744 ( \9059 , \8725 , \8735 );
xor \U$8745 ( \9060 , \9059 , \8754 );
xor \U$8746 ( \9061 , \8759 , \8761 );
xor \U$8747 ( \9062 , \9061 , \8764 );
and \U$8748 ( \9063 , \9060 , \9062 );
and \U$8749 ( \9064 , \9058 , \9063 );
xor \U$8750 ( \9065 , \8435 , \8460 );
xor \U$8751 ( \9066 , \9065 , \8471 );
and \U$8752 ( \9067 , \9063 , \9066 );
and \U$8753 ( \9068 , \9058 , \9066 );
or \U$8754 ( \9069 , \9064 , \9067 , \9068 );
xor \U$8755 ( \9070 , \8773 , \8775 );
xor \U$8756 ( \9071 , \9070 , \8778 );
and \U$8757 ( \9072 , \9069 , \9071 );
and \U$8758 ( \9073 , \8787 , \9072 );
xor \U$8759 ( \9074 , \8787 , \9072 );
xor \U$8760 ( \9075 , \9069 , \9071 );
xor \U$8761 ( \9076 , \8843 , \8847 );
xor \U$8762 ( \9077 , \9076 , \8852 );
xor \U$8763 ( \9078 , \8859 , \8863 );
xor \U$8764 ( \9079 , \9078 , \8868 );
and \U$8765 ( \9080 , \9077 , \9079 );
xor \U$8766 ( \9081 , \8876 , \8880 );
xor \U$8767 ( \9082 , \9081 , \8885 );
and \U$8768 ( \9083 , \9079 , \9082 );
and \U$8769 ( \9084 , \9077 , \9082 );
or \U$8770 ( \9085 , \9080 , \9083 , \9084 );
xor \U$8771 ( \9086 , \8791 , \8795 );
xor \U$8772 ( \9087 , \9086 , \8800 );
xor \U$8773 ( \9088 , \8807 , \8811 );
xor \U$8774 ( \9089 , \9088 , \8816 );
and \U$8775 ( \9090 , \9087 , \9089 );
xor \U$8776 ( \9091 , \8824 , \8828 );
xor \U$8777 ( \9092 , \9091 , \8833 );
and \U$8778 ( \9093 , \9089 , \9092 );
and \U$8779 ( \9094 , \9087 , \9092 );
or \U$8780 ( \9095 , \9090 , \9093 , \9094 );
and \U$8781 ( \9096 , \9085 , \9095 );
and \U$8782 ( \9097 , \8127 , \408 );
and \U$8783 ( \9098 , \7703 , \406 );
nor \U$8784 ( \9099 , \9097 , \9098 );
xnor \U$8785 ( \9100 , \9099 , \378 );
and \U$8786 ( \9101 , \8378 , \360 );
and \U$8787 ( \9102 , \8373 , \358 );
nor \U$8788 ( \9103 , \9101 , \9102 );
xnor \U$8789 ( \9104 , \9103 , \341 );
and \U$8790 ( \9105 , \9100 , \9104 );
and \U$8791 ( \9106 , \8981 , \323 );
and \U$8792 ( \9107 , \8697 , \321 );
nor \U$8793 ( \9108 , \9106 , \9107 );
xnor \U$8794 ( \9109 , \9108 , \328 );
and \U$8795 ( \9110 , \9104 , \9109 );
and \U$8796 ( \9111 , \9100 , \9109 );
or \U$8797 ( \9112 , \9105 , \9110 , \9111 );
xor \U$8798 ( \9113 , \8975 , \8979 );
xor \U$8799 ( \9114 , \9113 , \8982 );
or \U$8800 ( \9115 , \9112 , \9114 );
and \U$8801 ( \9116 , \9095 , \9115 );
and \U$8802 ( \9117 , \9085 , \9115 );
or \U$8803 ( \9118 , \9096 , \9116 , \9117 );
buf \U$8804 ( \9119 , RIc0c7ba8_61);
buf \U$8805 ( \9120 , RIc0c7b30_62);
and \U$8806 ( \9121 , \9119 , \9120 );
not \U$8807 ( \9122 , \9121 );
and \U$8808 ( \9123 , \8522 , \9122 );
not \U$8809 ( \9124 , \9123 );
and \U$8810 ( \9125 , \330 , \8896 );
and \U$8811 ( \9126 , \316 , \8894 );
nor \U$8812 ( \9127 , \9125 , \9126 );
xnor \U$8813 ( \9128 , \9127 , \8525 );
and \U$8814 ( \9129 , \9124 , \9128 );
and \U$8815 ( \9130 , \369 , \8334 );
and \U$8816 ( \9131 , \348 , \8332 );
nor \U$8817 ( \9132 , \9130 , \9131 );
xnor \U$8818 ( \9133 , \9132 , \8016 );
and \U$8819 ( \9134 , \9128 , \9133 );
and \U$8820 ( \9135 , \9124 , \9133 );
or \U$8821 ( \9136 , \9129 , \9134 , \9135 );
and \U$8822 ( \9137 , \709 , \6235 );
and \U$8823 ( \9138 , \681 , \6233 );
nor \U$8824 ( \9139 , \9137 , \9138 );
xnor \U$8825 ( \9140 , \9139 , \5895 );
and \U$8826 ( \9141 , \863 , \5646 );
and \U$8827 ( \9142 , \789 , \5644 );
nor \U$8828 ( \9143 , \9141 , \9142 );
xnor \U$8829 ( \9144 , \9143 , \5405 );
and \U$8830 ( \9145 , \9140 , \9144 );
and \U$8831 ( \9146 , \988 , \5180 );
and \U$8832 ( \9147 , \925 , \5178 );
nor \U$8833 ( \9148 , \9146 , \9147 );
xnor \U$8834 ( \9149 , \9148 , \4992 );
and \U$8835 ( \9150 , \9144 , \9149 );
and \U$8836 ( \9151 , \9140 , \9149 );
or \U$8837 ( \9152 , \9145 , \9150 , \9151 );
and \U$8838 ( \9153 , \9136 , \9152 );
and \U$8839 ( \9154 , \425 , \7767 );
and \U$8840 ( \9155 , \417 , \7765 );
nor \U$8841 ( \9156 , \9154 , \9155 );
xnor \U$8842 ( \9157 , \9156 , \7518 );
and \U$8843 ( \9158 , \499 , \7238 );
and \U$8844 ( \9159 , \494 , \7236 );
nor \U$8845 ( \9160 , \9158 , \9159 );
xnor \U$8846 ( \9161 , \9160 , \6978 );
and \U$8847 ( \9162 , \9157 , \9161 );
and \U$8848 ( \9163 , \604 , \6744 );
and \U$8849 ( \9164 , \553 , \6742 );
nor \U$8850 ( \9165 , \9163 , \9164 );
xnor \U$8851 ( \9166 , \9165 , \6429 );
and \U$8852 ( \9167 , \9161 , \9166 );
and \U$8853 ( \9168 , \9157 , \9166 );
or \U$8854 ( \9169 , \9162 , \9167 , \9168 );
and \U$8855 ( \9170 , \9152 , \9169 );
and \U$8856 ( \9171 , \9136 , \9169 );
or \U$8857 ( \9172 , \9153 , \9170 , \9171 );
and \U$8858 ( \9173 , \1799 , \3637 );
and \U$8859 ( \9174 , \1791 , \3635 );
nor \U$8860 ( \9175 , \9173 , \9174 );
xnor \U$8861 ( \9176 , \9175 , \3450 );
and \U$8862 ( \9177 , \2047 , \3324 );
and \U$8863 ( \9178 , \2042 , \3322 );
nor \U$8864 ( \9179 , \9177 , \9178 );
xnor \U$8865 ( \9180 , \9179 , \3119 );
and \U$8866 ( \9181 , \9176 , \9180 );
and \U$8867 ( \9182 , \2377 , \2918 );
and \U$8868 ( \9183 , \2233 , \2916 );
nor \U$8869 ( \9184 , \9182 , \9183 );
xnor \U$8870 ( \9185 , \9184 , \2769 );
and \U$8871 ( \9186 , \9180 , \9185 );
and \U$8872 ( \9187 , \9176 , \9185 );
or \U$8873 ( \9188 , \9181 , \9186 , \9187 );
and \U$8874 ( \9189 , \2666 , \2596 );
and \U$8875 ( \9190 , \2641 , \2594 );
nor \U$8876 ( \9191 , \9189 , \9190 );
xnor \U$8877 ( \9192 , \9191 , \2454 );
and \U$8878 ( \9193 , \3007 , \2300 );
and \U$8879 ( \9194 , \2840 , \2298 );
nor \U$8880 ( \9195 , \9193 , \9194 );
xnor \U$8881 ( \9196 , \9195 , \2163 );
and \U$8882 ( \9197 , \9192 , \9196 );
and \U$8883 ( \9198 , \3264 , \2094 );
and \U$8884 ( \9199 , \3145 , \2092 );
nor \U$8885 ( \9200 , \9198 , \9199 );
xnor \U$8886 ( \9201 , \9200 , \1942 );
and \U$8887 ( \9202 , \9196 , \9201 );
and \U$8888 ( \9203 , \9192 , \9201 );
or \U$8889 ( \9204 , \9197 , \9202 , \9203 );
and \U$8890 ( \9205 , \9188 , \9204 );
and \U$8891 ( \9206 , \1274 , \4806 );
and \U$8892 ( \9207 , \1186 , \4804 );
nor \U$8893 ( \9208 , \9206 , \9207 );
xnor \U$8894 ( \9209 , \9208 , \4574 );
and \U$8895 ( \9210 , \1384 , \4355 );
and \U$8896 ( \9211 , \1379 , \4353 );
nor \U$8897 ( \9212 , \9210 , \9211 );
xnor \U$8898 ( \9213 , \9212 , \4212 );
and \U$8899 ( \9214 , \9209 , \9213 );
and \U$8900 ( \9215 , \1615 , \4032 );
and \U$8901 ( \9216 , \1500 , \4030 );
nor \U$8902 ( \9217 , \9215 , \9216 );
xnor \U$8903 ( \9218 , \9217 , \3786 );
and \U$8904 ( \9219 , \9213 , \9218 );
and \U$8905 ( \9220 , \9209 , \9218 );
or \U$8906 ( \9221 , \9214 , \9219 , \9220 );
and \U$8907 ( \9222 , \9204 , \9221 );
and \U$8908 ( \9223 , \9188 , \9221 );
or \U$8909 ( \9224 , \9205 , \9222 , \9223 );
and \U$8910 ( \9225 , \9172 , \9224 );
and \U$8911 ( \9226 , \6157 , \692 );
and \U$8912 ( \9227 , \6148 , \690 );
nor \U$8913 ( \9228 , \9226 , \9227 );
xnor \U$8914 ( \9229 , \9228 , \649 );
and \U$8915 ( \9230 , \6702 , \579 );
and \U$8916 ( \9231 , \6500 , \577 );
nor \U$8917 ( \9232 , \9230 , \9231 );
xnor \U$8918 ( \9233 , \9232 , \530 );
and \U$8919 ( \9234 , \9229 , \9233 );
and \U$8920 ( \9235 , \7177 , \478 );
and \U$8921 ( \9236 , \7005 , \476 );
nor \U$8922 ( \9237 , \9235 , \9236 );
xnor \U$8923 ( \9238 , \9237 , \437 );
and \U$8924 ( \9239 , \9233 , \9238 );
and \U$8925 ( \9240 , \9229 , \9238 );
or \U$8926 ( \9241 , \9234 , \9239 , \9240 );
and \U$8927 ( \9242 , \4779 , \1160 );
and \U$8928 ( \9243 , \4771 , \1158 );
nor \U$8929 ( \9244 , \9242 , \9243 );
xnor \U$8930 ( \9245 , \9244 , \1082 );
and \U$8931 ( \9246 , \5253 , \996 );
and \U$8932 ( \9247 , \5248 , \994 );
nor \U$8933 ( \9248 , \9246 , \9247 );
xnor \U$8934 ( \9249 , \9248 , \902 );
and \U$8935 ( \9250 , \9245 , \9249 );
and \U$8936 ( \9251 , \5776 , \826 );
and \U$8937 ( \9252 , \5517 , \824 );
nor \U$8938 ( \9253 , \9251 , \9252 );
xnor \U$8939 ( \9254 , \9253 , \754 );
and \U$8940 ( \9255 , \9249 , \9254 );
and \U$8941 ( \9256 , \9245 , \9254 );
or \U$8942 ( \9257 , \9250 , \9255 , \9256 );
and \U$8943 ( \9258 , \9241 , \9257 );
and \U$8944 ( \9259 , \3889 , \1826 );
and \U$8945 ( \9260 , \3681 , \1824 );
nor \U$8946 ( \9261 , \9259 , \9260 );
xnor \U$8947 ( \9262 , \9261 , \1670 );
and \U$8948 ( \9263 , \4016 , \1554 );
and \U$8949 ( \9264 , \4011 , \1552 );
nor \U$8950 ( \9265 , \9263 , \9264 );
xnor \U$8951 ( \9266 , \9265 , \1441 );
and \U$8952 ( \9267 , \9262 , \9266 );
and \U$8953 ( \9268 , \4469 , \1360 );
and \U$8954 ( \9269 , \4272 , \1358 );
nor \U$8955 ( \9270 , \9268 , \9269 );
xnor \U$8956 ( \9271 , \9270 , \1224 );
and \U$8957 ( \9272 , \9266 , \9271 );
and \U$8958 ( \9273 , \9262 , \9271 );
or \U$8959 ( \9274 , \9267 , \9272 , \9273 );
and \U$8960 ( \9275 , \9257 , \9274 );
and \U$8961 ( \9276 , \9241 , \9274 );
or \U$8962 ( \9277 , \9258 , \9275 , \9276 );
and \U$8963 ( \9278 , \9224 , \9277 );
and \U$8964 ( \9279 , \9172 , \9277 );
or \U$8965 ( \9280 , \9225 , \9278 , \9279 );
and \U$8966 ( \9281 , \9118 , \9280 );
xor \U$8967 ( \9282 , \8899 , \8903 );
xor \U$8968 ( \9283 , \9282 , \8908 );
xor \U$8969 ( \9284 , \8915 , \8919 );
xor \U$8970 ( \9285 , \9284 , \8924 );
and \U$8971 ( \9286 , \9283 , \9285 );
xor \U$8972 ( \9287 , \8932 , \8936 );
xor \U$8973 ( \9288 , \9287 , \8941 );
and \U$8974 ( \9289 , \9285 , \9288 );
and \U$8975 ( \9290 , \9283 , \9288 );
or \U$8976 ( \9291 , \9286 , \9289 , \9290 );
xor \U$8977 ( \9292 , \8508 , \8512 );
xor \U$8978 ( \9293 , \9292 , \8517 );
and \U$8979 ( \9294 , \9291 , \9293 );
xor \U$8980 ( \9295 , \8526 , \8530 );
xor \U$8981 ( \9296 , \9295 , \8535 );
and \U$8982 ( \9297 , \9293 , \9296 );
and \U$8983 ( \9298 , \9291 , \9296 );
or \U$8984 ( \9299 , \9294 , \9297 , \9298 );
and \U$8985 ( \9300 , \9280 , \9299 );
and \U$8986 ( \9301 , \9118 , \9299 );
or \U$8987 ( \9302 , \9281 , \9300 , \9301 );
xor \U$8988 ( \9303 , \8803 , \8819 );
xor \U$8989 ( \9304 , \9303 , \8836 );
xor \U$8990 ( \9305 , \8855 , \8871 );
xor \U$8991 ( \9306 , \9305 , \8888 );
and \U$8992 ( \9307 , \9304 , \9306 );
xor \U$8993 ( \9308 , \8911 , \8927 );
xor \U$8994 ( \9309 , \9308 , \8944 );
and \U$8995 ( \9310 , \9306 , \9309 );
and \U$8996 ( \9311 , \9304 , \9309 );
or \U$8997 ( \9312 , \9307 , \9310 , \9311 );
xor \U$8998 ( \9313 , \8952 , \8954 );
xor \U$8999 ( \9314 , \9313 , \8957 );
xor \U$9000 ( \9315 , \8962 , \8964 );
xor \U$9001 ( \9316 , \9315 , \8967 );
and \U$9002 ( \9317 , \9314 , \9316 );
xor \U$9003 ( \9318 , \8985 , \8987 );
xor \U$9004 ( \9319 , \9318 , \8990 );
and \U$9005 ( \9320 , \9316 , \9319 );
and \U$9006 ( \9321 , \9314 , \9319 );
or \U$9007 ( \9322 , \9317 , \9320 , \9321 );
and \U$9008 ( \9323 , \9312 , \9322 );
xor \U$9009 ( \9324 , \8574 , \8590 );
xor \U$9010 ( \9325 , \9324 , \8607 );
and \U$9011 ( \9326 , \9322 , \9325 );
and \U$9012 ( \9327 , \9312 , \9325 );
or \U$9013 ( \9328 , \9323 , \9326 , \9327 );
and \U$9014 ( \9329 , \9302 , \9328 );
xor \U$9015 ( \9330 , \8520 , \8538 );
xor \U$9016 ( \9331 , \9330 , \8555 );
xor \U$9017 ( \9332 , \8999 , \9001 );
xor \U$9018 ( \9333 , \9332 , \9004 );
and \U$9019 ( \9334 , \9331 , \9333 );
xor \U$9020 ( \9335 , \9012 , \9014 );
xor \U$9021 ( \9336 , \9335 , \9017 );
and \U$9022 ( \9337 , \9333 , \9336 );
and \U$9023 ( \9338 , \9331 , \9336 );
or \U$9024 ( \9339 , \9334 , \9337 , \9338 );
and \U$9025 ( \9340 , \9328 , \9339 );
and \U$9026 ( \9341 , \9302 , \9339 );
or \U$9027 ( \9342 , \9329 , \9340 , \9341 );
xor \U$9028 ( \9343 , \8950 , \8996 );
xor \U$9029 ( \9344 , \9343 , \9007 );
xor \U$9030 ( \9345 , \9020 , \9022 );
xor \U$9031 ( \9346 , \9345 , \9025 );
and \U$9032 ( \9347 , \9344 , \9346 );
xor \U$9033 ( \9348 , \9031 , \9033 );
xor \U$9034 ( \9349 , \9348 , \9036 );
and \U$9035 ( \9350 , \9346 , \9349 );
and \U$9036 ( \9351 , \9344 , \9349 );
or \U$9037 ( \9352 , \9347 , \9350 , \9351 );
and \U$9038 ( \9353 , \9342 , \9352 );
xor \U$9039 ( \9354 , \9044 , \9046 );
xor \U$9040 ( \9355 , \9354 , \9049 );
and \U$9041 ( \9356 , \9352 , \9355 );
and \U$9042 ( \9357 , \9342 , \9355 );
or \U$9043 ( \9358 , \9353 , \9356 , \9357 );
xor \U$9044 ( \9359 , \9042 , \9052 );
xor \U$9045 ( \9360 , \9359 , \9055 );
and \U$9046 ( \9361 , \9358 , \9360 );
xor \U$9047 ( \9362 , \9060 , \9062 );
and \U$9048 ( \9363 , \9360 , \9362 );
and \U$9049 ( \9364 , \9358 , \9362 );
or \U$9050 ( \9365 , \9361 , \9363 , \9364 );
xor \U$9051 ( \9366 , \9058 , \9063 );
xor \U$9052 ( \9367 , \9366 , \9066 );
and \U$9053 ( \9368 , \9365 , \9367 );
xor \U$9054 ( \9369 , \8757 , \8767 );
xor \U$9055 ( \9370 , \9369 , \8770 );
and \U$9056 ( \9371 , \9367 , \9370 );
and \U$9057 ( \9372 , \9365 , \9370 );
or \U$9058 ( \9373 , \9368 , \9371 , \9372 );
and \U$9059 ( \9374 , \9075 , \9373 );
xor \U$9060 ( \9375 , \9075 , \9373 );
xor \U$9061 ( \9376 , \9365 , \9367 );
xor \U$9062 ( \9377 , \9376 , \9370 );
and \U$9063 ( \9378 , \5248 , \1160 );
and \U$9064 ( \9379 , \4779 , \1158 );
nor \U$9065 ( \9380 , \9378 , \9379 );
xnor \U$9066 ( \9381 , \9380 , \1082 );
and \U$9067 ( \9382 , \5517 , \996 );
and \U$9068 ( \9383 , \5253 , \994 );
nor \U$9069 ( \9384 , \9382 , \9383 );
xnor \U$9070 ( \9385 , \9384 , \902 );
and \U$9071 ( \9386 , \9381 , \9385 );
and \U$9072 ( \9387 , \6148 , \826 );
and \U$9073 ( \9388 , \5776 , \824 );
nor \U$9074 ( \9389 , \9387 , \9388 );
xnor \U$9075 ( \9390 , \9389 , \754 );
and \U$9076 ( \9391 , \9385 , \9390 );
and \U$9077 ( \9392 , \9381 , \9390 );
or \U$9078 ( \9393 , \9386 , \9391 , \9392 );
and \U$9079 ( \9394 , \4011 , \1826 );
and \U$9080 ( \9395 , \3889 , \1824 );
nor \U$9081 ( \9396 , \9394 , \9395 );
xnor \U$9082 ( \9397 , \9396 , \1670 );
and \U$9083 ( \9398 , \4272 , \1554 );
and \U$9084 ( \9399 , \4016 , \1552 );
nor \U$9085 ( \9400 , \9398 , \9399 );
xnor \U$9086 ( \9401 , \9400 , \1441 );
and \U$9087 ( \9402 , \9397 , \9401 );
and \U$9088 ( \9403 , \4771 , \1360 );
and \U$9089 ( \9404 , \4469 , \1358 );
nor \U$9090 ( \9405 , \9403 , \9404 );
xnor \U$9091 ( \9406 , \9405 , \1224 );
and \U$9092 ( \9407 , \9401 , \9406 );
and \U$9093 ( \9408 , \9397 , \9406 );
or \U$9094 ( \9409 , \9402 , \9407 , \9408 );
and \U$9095 ( \9410 , \9393 , \9409 );
and \U$9096 ( \9411 , \6500 , \692 );
and \U$9097 ( \9412 , \6157 , \690 );
nor \U$9098 ( \9413 , \9411 , \9412 );
xnor \U$9099 ( \9414 , \9413 , \649 );
and \U$9100 ( \9415 , \7005 , \579 );
and \U$9101 ( \9416 , \6702 , \577 );
nor \U$9102 ( \9417 , \9415 , \9416 );
xnor \U$9103 ( \9418 , \9417 , \530 );
and \U$9104 ( \9419 , \9414 , \9418 );
and \U$9105 ( \9420 , \7703 , \478 );
and \U$9106 ( \9421 , \7177 , \476 );
nor \U$9107 ( \9422 , \9420 , \9421 );
xnor \U$9108 ( \9423 , \9422 , \437 );
and \U$9109 ( \9424 , \9418 , \9423 );
and \U$9110 ( \9425 , \9414 , \9423 );
or \U$9111 ( \9426 , \9419 , \9424 , \9425 );
and \U$9112 ( \9427 , \9409 , \9426 );
and \U$9113 ( \9428 , \9393 , \9426 );
or \U$9114 ( \9429 , \9410 , \9427 , \9428 );
xor \U$9115 ( \9430 , \8522 , \9119 );
xor \U$9116 ( \9431 , \9119 , \9120 );
not \U$9117 ( \9432 , \9431 );
and \U$9118 ( \9433 , \9430 , \9432 );
and \U$9119 ( \9434 , \316 , \9433 );
not \U$9120 ( \9435 , \9434 );
xnor \U$9121 ( \9436 , \9435 , \9123 );
and \U$9122 ( \9437 , \348 , \8896 );
and \U$9123 ( \9438 , \330 , \8894 );
nor \U$9124 ( \9439 , \9437 , \9438 );
xnor \U$9125 ( \9440 , \9439 , \8525 );
and \U$9126 ( \9441 , \9436 , \9440 );
and \U$9127 ( \9442 , \417 , \8334 );
and \U$9128 ( \9443 , \369 , \8332 );
nor \U$9129 ( \9444 , \9442 , \9443 );
xnor \U$9130 ( \9445 , \9444 , \8016 );
and \U$9131 ( \9446 , \9440 , \9445 );
and \U$9132 ( \9447 , \9436 , \9445 );
or \U$9133 ( \9448 , \9441 , \9446 , \9447 );
and \U$9134 ( \9449 , \789 , \6235 );
and \U$9135 ( \9450 , \709 , \6233 );
nor \U$9136 ( \9451 , \9449 , \9450 );
xnor \U$9137 ( \9452 , \9451 , \5895 );
and \U$9138 ( \9453 , \925 , \5646 );
and \U$9139 ( \9454 , \863 , \5644 );
nor \U$9140 ( \9455 , \9453 , \9454 );
xnor \U$9141 ( \9456 , \9455 , \5405 );
and \U$9142 ( \9457 , \9452 , \9456 );
and \U$9143 ( \9458 , \1186 , \5180 );
and \U$9144 ( \9459 , \988 , \5178 );
nor \U$9145 ( \9460 , \9458 , \9459 );
xnor \U$9146 ( \9461 , \9460 , \4992 );
and \U$9147 ( \9462 , \9456 , \9461 );
and \U$9148 ( \9463 , \9452 , \9461 );
or \U$9149 ( \9464 , \9457 , \9462 , \9463 );
and \U$9150 ( \9465 , \9448 , \9464 );
and \U$9151 ( \9466 , \494 , \7767 );
and \U$9152 ( \9467 , \425 , \7765 );
nor \U$9153 ( \9468 , \9466 , \9467 );
xnor \U$9154 ( \9469 , \9468 , \7518 );
and \U$9155 ( \9470 , \553 , \7238 );
and \U$9156 ( \9471 , \499 , \7236 );
nor \U$9157 ( \9472 , \9470 , \9471 );
xnor \U$9158 ( \9473 , \9472 , \6978 );
and \U$9159 ( \9474 , \9469 , \9473 );
and \U$9160 ( \9475 , \681 , \6744 );
and \U$9161 ( \9476 , \604 , \6742 );
nor \U$9162 ( \9477 , \9475 , \9476 );
xnor \U$9163 ( \9478 , \9477 , \6429 );
and \U$9164 ( \9479 , \9473 , \9478 );
and \U$9165 ( \9480 , \9469 , \9478 );
or \U$9166 ( \9481 , \9474 , \9479 , \9480 );
and \U$9167 ( \9482 , \9464 , \9481 );
and \U$9168 ( \9483 , \9448 , \9481 );
or \U$9169 ( \9484 , \9465 , \9482 , \9483 );
and \U$9170 ( \9485 , \9429 , \9484 );
and \U$9171 ( \9486 , \1379 , \4806 );
and \U$9172 ( \9487 , \1274 , \4804 );
nor \U$9173 ( \9488 , \9486 , \9487 );
xnor \U$9174 ( \9489 , \9488 , \4574 );
and \U$9175 ( \9490 , \1500 , \4355 );
and \U$9176 ( \9491 , \1384 , \4353 );
nor \U$9177 ( \9492 , \9490 , \9491 );
xnor \U$9178 ( \9493 , \9492 , \4212 );
and \U$9179 ( \9494 , \9489 , \9493 );
and \U$9180 ( \9495 , \1791 , \4032 );
and \U$9181 ( \9496 , \1615 , \4030 );
nor \U$9182 ( \9497 , \9495 , \9496 );
xnor \U$9183 ( \9498 , \9497 , \3786 );
and \U$9184 ( \9499 , \9493 , \9498 );
and \U$9185 ( \9500 , \9489 , \9498 );
or \U$9186 ( \9501 , \9494 , \9499 , \9500 );
and \U$9187 ( \9502 , \2840 , \2596 );
and \U$9188 ( \9503 , \2666 , \2594 );
nor \U$9189 ( \9504 , \9502 , \9503 );
xnor \U$9190 ( \9505 , \9504 , \2454 );
and \U$9191 ( \9506 , \3145 , \2300 );
and \U$9192 ( \9507 , \3007 , \2298 );
nor \U$9193 ( \9508 , \9506 , \9507 );
xnor \U$9194 ( \9509 , \9508 , \2163 );
and \U$9195 ( \9510 , \9505 , \9509 );
and \U$9196 ( \9511 , \3681 , \2094 );
and \U$9197 ( \9512 , \3264 , \2092 );
nor \U$9198 ( \9513 , \9511 , \9512 );
xnor \U$9199 ( \9514 , \9513 , \1942 );
and \U$9200 ( \9515 , \9509 , \9514 );
and \U$9201 ( \9516 , \9505 , \9514 );
or \U$9202 ( \9517 , \9510 , \9515 , \9516 );
and \U$9203 ( \9518 , \9501 , \9517 );
and \U$9204 ( \9519 , \2042 , \3637 );
and \U$9205 ( \9520 , \1799 , \3635 );
nor \U$9206 ( \9521 , \9519 , \9520 );
xnor \U$9207 ( \9522 , \9521 , \3450 );
and \U$9208 ( \9523 , \2233 , \3324 );
and \U$9209 ( \9524 , \2047 , \3322 );
nor \U$9210 ( \9525 , \9523 , \9524 );
xnor \U$9211 ( \9526 , \9525 , \3119 );
and \U$9212 ( \9527 , \9522 , \9526 );
and \U$9213 ( \9528 , \2641 , \2918 );
and \U$9214 ( \9529 , \2377 , \2916 );
nor \U$9215 ( \9530 , \9528 , \9529 );
xnor \U$9216 ( \9531 , \9530 , \2769 );
and \U$9217 ( \9532 , \9526 , \9531 );
and \U$9218 ( \9533 , \9522 , \9531 );
or \U$9219 ( \9534 , \9527 , \9532 , \9533 );
and \U$9220 ( \9535 , \9517 , \9534 );
and \U$9221 ( \9536 , \9501 , \9534 );
or \U$9222 ( \9537 , \9518 , \9535 , \9536 );
and \U$9223 ( \9538 , \9484 , \9537 );
and \U$9224 ( \9539 , \9429 , \9537 );
or \U$9225 ( \9540 , \9485 , \9538 , \9539 );
and \U$9226 ( \9541 , \8373 , \408 );
and \U$9227 ( \9542 , \8127 , \406 );
nor \U$9228 ( \9543 , \9541 , \9542 );
xnor \U$9229 ( \9544 , \9543 , \378 );
and \U$9230 ( \9545 , \8697 , \360 );
and \U$9231 ( \9546 , \8378 , \358 );
nor \U$9232 ( \9547 , \9545 , \9546 );
xnor \U$9233 ( \9548 , \9547 , \341 );
and \U$9234 ( \9549 , \9544 , \9548 );
buf \U$9235 ( \9550 , RIc0c5e20_124);
and \U$9236 ( \9551 , \9550 , \323 );
and \U$9237 ( \9552 , \8981 , \321 );
nor \U$9238 ( \9553 , \9551 , \9552 );
xnor \U$9239 ( \9554 , \9553 , \328 );
and \U$9240 ( \9555 , \9548 , \9554 );
and \U$9241 ( \9556 , \9544 , \9554 );
or \U$9242 ( \9557 , \9549 , \9555 , \9556 );
buf \U$9243 ( \9558 , RIc0c5da8_125);
and \U$9244 ( \9559 , \9558 , \317 );
buf \U$9245 ( \9560 , \9559 );
and \U$9246 ( \9561 , \9557 , \9560 );
and \U$9247 ( \9562 , \9550 , \317 );
and \U$9248 ( \9563 , \9560 , \9562 );
and \U$9249 ( \9564 , \9557 , \9562 );
or \U$9250 ( \9565 , \9561 , \9563 , \9564 );
xor \U$9251 ( \9566 , \9100 , \9104 );
xor \U$9252 ( \9567 , \9566 , \9109 );
xor \U$9253 ( \9568 , \9229 , \9233 );
xor \U$9254 ( \9569 , \9568 , \9238 );
and \U$9255 ( \9570 , \9567 , \9569 );
xor \U$9256 ( \9571 , \9245 , \9249 );
xor \U$9257 ( \9572 , \9571 , \9254 );
and \U$9258 ( \9573 , \9569 , \9572 );
and \U$9259 ( \9574 , \9567 , \9572 );
or \U$9260 ( \9575 , \9570 , \9573 , \9574 );
and \U$9261 ( \9576 , \9565 , \9575 );
xor \U$9262 ( \9577 , \9262 , \9266 );
xor \U$9263 ( \9578 , \9577 , \9271 );
xor \U$9264 ( \9579 , \9176 , \9180 );
xor \U$9265 ( \9580 , \9579 , \9185 );
and \U$9266 ( \9581 , \9578 , \9580 );
xor \U$9267 ( \9582 , \9192 , \9196 );
xor \U$9268 ( \9583 , \9582 , \9201 );
and \U$9269 ( \9584 , \9580 , \9583 );
and \U$9270 ( \9585 , \9578 , \9583 );
or \U$9271 ( \9586 , \9581 , \9584 , \9585 );
and \U$9272 ( \9587 , \9575 , \9586 );
and \U$9273 ( \9588 , \9565 , \9586 );
or \U$9274 ( \9589 , \9576 , \9587 , \9588 );
and \U$9275 ( \9590 , \9540 , \9589 );
xor \U$9276 ( \9591 , \9140 , \9144 );
xor \U$9277 ( \9592 , \9591 , \9149 );
xor \U$9278 ( \9593 , \9157 , \9161 );
xor \U$9279 ( \9594 , \9593 , \9166 );
and \U$9280 ( \9595 , \9592 , \9594 );
xor \U$9281 ( \9596 , \9209 , \9213 );
xor \U$9282 ( \9597 , \9596 , \9218 );
and \U$9283 ( \9598 , \9594 , \9597 );
and \U$9284 ( \9599 , \9592 , \9597 );
or \U$9285 ( \9600 , \9595 , \9598 , \9599 );
xor \U$9286 ( \9601 , \9283 , \9285 );
xor \U$9287 ( \9602 , \9601 , \9288 );
and \U$9288 ( \9603 , \9600 , \9602 );
xor \U$9289 ( \9604 , \9087 , \9089 );
xor \U$9290 ( \9605 , \9604 , \9092 );
and \U$9291 ( \9606 , \9602 , \9605 );
and \U$9292 ( \9607 , \9600 , \9605 );
or \U$9293 ( \9608 , \9603 , \9606 , \9607 );
and \U$9294 ( \9609 , \9589 , \9608 );
and \U$9295 ( \9610 , \9540 , \9608 );
or \U$9296 ( \9611 , \9590 , \9609 , \9610 );
xor \U$9297 ( \9612 , \9085 , \9095 );
xor \U$9298 ( \9613 , \9612 , \9115 );
xor \U$9299 ( \9614 , \9172 , \9224 );
xor \U$9300 ( \9615 , \9614 , \9277 );
and \U$9301 ( \9616 , \9613 , \9615 );
xor \U$9302 ( \9617 , \9291 , \9293 );
xor \U$9303 ( \9618 , \9617 , \9296 );
and \U$9304 ( \9619 , \9615 , \9618 );
and \U$9305 ( \9620 , \9613 , \9618 );
or \U$9306 ( \9621 , \9616 , \9619 , \9620 );
and \U$9307 ( \9622 , \9611 , \9621 );
xor \U$9308 ( \9623 , \9241 , \9257 );
xor \U$9309 ( \9624 , \9623 , \9274 );
xor \U$9310 ( \9625 , \9077 , \9079 );
xor \U$9311 ( \9626 , \9625 , \9082 );
and \U$9312 ( \9627 , \9624 , \9626 );
xnor \U$9313 ( \9628 , \9112 , \9114 );
and \U$9314 ( \9629 , \9626 , \9628 );
and \U$9315 ( \9630 , \9624 , \9628 );
or \U$9316 ( \9631 , \9627 , \9629 , \9630 );
xor \U$9317 ( \9632 , \9304 , \9306 );
xor \U$9318 ( \9633 , \9632 , \9309 );
and \U$9319 ( \9634 , \9631 , \9633 );
xor \U$9320 ( \9635 , \9314 , \9316 );
xor \U$9321 ( \9636 , \9635 , \9319 );
and \U$9322 ( \9637 , \9633 , \9636 );
and \U$9323 ( \9638 , \9631 , \9636 );
or \U$9324 ( \9639 , \9634 , \9637 , \9638 );
and \U$9325 ( \9640 , \9621 , \9639 );
and \U$9326 ( \9641 , \9611 , \9639 );
or \U$9327 ( \9642 , \9622 , \9640 , \9641 );
xor \U$9328 ( \9643 , \8839 , \8891 );
xor \U$9329 ( \9644 , \9643 , \8947 );
xor \U$9330 ( \9645 , \8960 , \8970 );
xor \U$9331 ( \9646 , \9645 , \8993 );
and \U$9332 ( \9647 , \9644 , \9646 );
xor \U$9333 ( \9648 , \9331 , \9333 );
xor \U$9334 ( \9649 , \9648 , \9336 );
and \U$9335 ( \9650 , \9646 , \9649 );
and \U$9336 ( \9651 , \9644 , \9649 );
or \U$9337 ( \9652 , \9647 , \9650 , \9651 );
and \U$9338 ( \9653 , \9642 , \9652 );
xor \U$9339 ( \9654 , \9344 , \9346 );
xor \U$9340 ( \9655 , \9654 , \9349 );
and \U$9341 ( \9656 , \9652 , \9655 );
and \U$9342 ( \9657 , \9642 , \9655 );
or \U$9343 ( \9658 , \9653 , \9656 , \9657 );
xor \U$9344 ( \9659 , \9010 , \9028 );
xor \U$9345 ( \9660 , \9659 , \9039 );
and \U$9346 ( \9661 , \9658 , \9660 );
xor \U$9347 ( \9662 , \9342 , \9352 );
xor \U$9348 ( \9663 , \9662 , \9355 );
and \U$9349 ( \9664 , \9660 , \9663 );
and \U$9350 ( \9665 , \9658 , \9663 );
or \U$9351 ( \9666 , \9661 , \9664 , \9665 );
xor \U$9352 ( \9667 , \9358 , \9360 );
xor \U$9353 ( \9668 , \9667 , \9362 );
and \U$9354 ( \9669 , \9666 , \9668 );
and \U$9355 ( \9670 , \9377 , \9669 );
xor \U$9356 ( \9671 , \9377 , \9669 );
xor \U$9357 ( \9672 , \9666 , \9668 );
and \U$9358 ( \9673 , \2666 , \2918 );
and \U$9359 ( \9674 , \2641 , \2916 );
nor \U$9360 ( \9675 , \9673 , \9674 );
xnor \U$9361 ( \9676 , \9675 , \2769 );
and \U$9362 ( \9677 , \3007 , \2596 );
and \U$9363 ( \9678 , \2840 , \2594 );
nor \U$9364 ( \9679 , \9677 , \9678 );
xnor \U$9365 ( \9680 , \9679 , \2454 );
and \U$9366 ( \9681 , \9676 , \9680 );
and \U$9367 ( \9682 , \3264 , \2300 );
and \U$9368 ( \9683 , \3145 , \2298 );
nor \U$9369 ( \9684 , \9682 , \9683 );
xnor \U$9370 ( \9685 , \9684 , \2163 );
and \U$9371 ( \9686 , \9680 , \9685 );
and \U$9372 ( \9687 , \9676 , \9685 );
or \U$9373 ( \9688 , \9681 , \9686 , \9687 );
and \U$9374 ( \9689 , \1799 , \4032 );
and \U$9375 ( \9690 , \1791 , \4030 );
nor \U$9376 ( \9691 , \9689 , \9690 );
xnor \U$9377 ( \9692 , \9691 , \3786 );
and \U$9378 ( \9693 , \2047 , \3637 );
and \U$9379 ( \9694 , \2042 , \3635 );
nor \U$9380 ( \9695 , \9693 , \9694 );
xnor \U$9381 ( \9696 , \9695 , \3450 );
and \U$9382 ( \9697 , \9692 , \9696 );
and \U$9383 ( \9698 , \2377 , \3324 );
and \U$9384 ( \9699 , \2233 , \3322 );
nor \U$9385 ( \9700 , \9698 , \9699 );
xnor \U$9386 ( \9701 , \9700 , \3119 );
and \U$9387 ( \9702 , \9696 , \9701 );
and \U$9388 ( \9703 , \9692 , \9701 );
or \U$9389 ( \9704 , \9697 , \9702 , \9703 );
and \U$9390 ( \9705 , \9688 , \9704 );
and \U$9391 ( \9706 , \1274 , \5180 );
and \U$9392 ( \9707 , \1186 , \5178 );
nor \U$9393 ( \9708 , \9706 , \9707 );
xnor \U$9394 ( \9709 , \9708 , \4992 );
and \U$9395 ( \9710 , \1384 , \4806 );
and \U$9396 ( \9711 , \1379 , \4804 );
nor \U$9397 ( \9712 , \9710 , \9711 );
xnor \U$9398 ( \9713 , \9712 , \4574 );
and \U$9399 ( \9714 , \9709 , \9713 );
and \U$9400 ( \9715 , \1615 , \4355 );
and \U$9401 ( \9716 , \1500 , \4353 );
nor \U$9402 ( \9717 , \9715 , \9716 );
xnor \U$9403 ( \9718 , \9717 , \4212 );
and \U$9404 ( \9719 , \9713 , \9718 );
and \U$9405 ( \9720 , \9709 , \9718 );
or \U$9406 ( \9721 , \9714 , \9719 , \9720 );
and \U$9407 ( \9722 , \9704 , \9721 );
and \U$9408 ( \9723 , \9688 , \9721 );
or \U$9409 ( \9724 , \9705 , \9722 , \9723 );
and \U$9410 ( \9725 , \709 , \6744 );
and \U$9411 ( \9726 , \681 , \6742 );
nor \U$9412 ( \9727 , \9725 , \9726 );
xnor \U$9413 ( \9728 , \9727 , \6429 );
and \U$9414 ( \9729 , \863 , \6235 );
and \U$9415 ( \9730 , \789 , \6233 );
nor \U$9416 ( \9731 , \9729 , \9730 );
xnor \U$9417 ( \9732 , \9731 , \5895 );
and \U$9418 ( \9733 , \9728 , \9732 );
and \U$9419 ( \9734 , \988 , \5646 );
and \U$9420 ( \9735 , \925 , \5644 );
nor \U$9421 ( \9736 , \9734 , \9735 );
xnor \U$9422 ( \9737 , \9736 , \5405 );
and \U$9423 ( \9738 , \9732 , \9737 );
and \U$9424 ( \9739 , \9728 , \9737 );
or \U$9425 ( \9740 , \9733 , \9738 , \9739 );
and \U$9426 ( \9741 , \425 , \8334 );
and \U$9427 ( \9742 , \417 , \8332 );
nor \U$9428 ( \9743 , \9741 , \9742 );
xnor \U$9429 ( \9744 , \9743 , \8016 );
and \U$9430 ( \9745 , \499 , \7767 );
and \U$9431 ( \9746 , \494 , \7765 );
nor \U$9432 ( \9747 , \9745 , \9746 );
xnor \U$9433 ( \9748 , \9747 , \7518 );
and \U$9434 ( \9749 , \9744 , \9748 );
and \U$9435 ( \9750 , \604 , \7238 );
and \U$9436 ( \9751 , \553 , \7236 );
nor \U$9437 ( \9752 , \9750 , \9751 );
xnor \U$9438 ( \9753 , \9752 , \6978 );
and \U$9439 ( \9754 , \9748 , \9753 );
and \U$9440 ( \9755 , \9744 , \9753 );
or \U$9441 ( \9756 , \9749 , \9754 , \9755 );
and \U$9442 ( \9757 , \9740 , \9756 );
buf \U$9443 ( \9758 , RIc0c7ab8_63);
buf \U$9444 ( \9759 , RIc0c7a40_64);
and \U$9445 ( \9760 , \9758 , \9759 );
not \U$9446 ( \9761 , \9760 );
and \U$9447 ( \9762 , \9120 , \9761 );
not \U$9448 ( \9763 , \9762 );
and \U$9449 ( \9764 , \330 , \9433 );
and \U$9450 ( \9765 , \316 , \9431 );
nor \U$9451 ( \9766 , \9764 , \9765 );
xnor \U$9452 ( \9767 , \9766 , \9123 );
and \U$9453 ( \9768 , \9763 , \9767 );
and \U$9454 ( \9769 , \369 , \8896 );
and \U$9455 ( \9770 , \348 , \8894 );
nor \U$9456 ( \9771 , \9769 , \9770 );
xnor \U$9457 ( \9772 , \9771 , \8525 );
and \U$9458 ( \9773 , \9767 , \9772 );
and \U$9459 ( \9774 , \9763 , \9772 );
or \U$9460 ( \9775 , \9768 , \9773 , \9774 );
and \U$9461 ( \9776 , \9756 , \9775 );
and \U$9462 ( \9777 , \9740 , \9775 );
or \U$9463 ( \9778 , \9757 , \9776 , \9777 );
and \U$9464 ( \9779 , \9724 , \9778 );
and \U$9465 ( \9780 , \6157 , \826 );
and \U$9466 ( \9781 , \6148 , \824 );
nor \U$9467 ( \9782 , \9780 , \9781 );
xnor \U$9468 ( \9783 , \9782 , \754 );
and \U$9469 ( \9784 , \6702 , \692 );
and \U$9470 ( \9785 , \6500 , \690 );
nor \U$9471 ( \9786 , \9784 , \9785 );
xnor \U$9472 ( \9787 , \9786 , \649 );
and \U$9473 ( \9788 , \9783 , \9787 );
and \U$9474 ( \9789 , \7177 , \579 );
and \U$9475 ( \9790 , \7005 , \577 );
nor \U$9476 ( \9791 , \9789 , \9790 );
xnor \U$9477 ( \9792 , \9791 , \530 );
and \U$9478 ( \9793 , \9787 , \9792 );
and \U$9479 ( \9794 , \9783 , \9792 );
or \U$9480 ( \9795 , \9788 , \9793 , \9794 );
and \U$9481 ( \9796 , \4779 , \1360 );
and \U$9482 ( \9797 , \4771 , \1358 );
nor \U$9483 ( \9798 , \9796 , \9797 );
xnor \U$9484 ( \9799 , \9798 , \1224 );
and \U$9485 ( \9800 , \5253 , \1160 );
and \U$9486 ( \9801 , \5248 , \1158 );
nor \U$9487 ( \9802 , \9800 , \9801 );
xnor \U$9488 ( \9803 , \9802 , \1082 );
and \U$9489 ( \9804 , \9799 , \9803 );
and \U$9490 ( \9805 , \5776 , \996 );
and \U$9491 ( \9806 , \5517 , \994 );
nor \U$9492 ( \9807 , \9805 , \9806 );
xnor \U$9493 ( \9808 , \9807 , \902 );
and \U$9494 ( \9809 , \9803 , \9808 );
and \U$9495 ( \9810 , \9799 , \9808 );
or \U$9496 ( \9811 , \9804 , \9809 , \9810 );
and \U$9497 ( \9812 , \9795 , \9811 );
and \U$9498 ( \9813 , \3889 , \2094 );
and \U$9499 ( \9814 , \3681 , \2092 );
nor \U$9500 ( \9815 , \9813 , \9814 );
xnor \U$9501 ( \9816 , \9815 , \1942 );
and \U$9502 ( \9817 , \4016 , \1826 );
and \U$9503 ( \9818 , \4011 , \1824 );
nor \U$9504 ( \9819 , \9817 , \9818 );
xnor \U$9505 ( \9820 , \9819 , \1670 );
and \U$9506 ( \9821 , \9816 , \9820 );
and \U$9507 ( \9822 , \4469 , \1554 );
and \U$9508 ( \9823 , \4272 , \1552 );
nor \U$9509 ( \9824 , \9822 , \9823 );
xnor \U$9510 ( \9825 , \9824 , \1441 );
and \U$9511 ( \9826 , \9820 , \9825 );
and \U$9512 ( \9827 , \9816 , \9825 );
or \U$9513 ( \9828 , \9821 , \9826 , \9827 );
and \U$9514 ( \9829 , \9811 , \9828 );
and \U$9515 ( \9830 , \9795 , \9828 );
or \U$9516 ( \9831 , \9812 , \9829 , \9830 );
and \U$9517 ( \9832 , \9778 , \9831 );
and \U$9518 ( \9833 , \9724 , \9831 );
or \U$9519 ( \9834 , \9779 , \9832 , \9833 );
xor \U$9520 ( \9835 , \9489 , \9493 );
xor \U$9521 ( \9836 , \9835 , \9498 );
xor \U$9522 ( \9837 , \9505 , \9509 );
xor \U$9523 ( \9838 , \9837 , \9514 );
and \U$9524 ( \9839 , \9836 , \9838 );
xor \U$9525 ( \9840 , \9522 , \9526 );
xor \U$9526 ( \9841 , \9840 , \9531 );
and \U$9527 ( \9842 , \9838 , \9841 );
and \U$9528 ( \9843 , \9836 , \9841 );
or \U$9529 ( \9844 , \9839 , \9842 , \9843 );
xor \U$9530 ( \9845 , \9381 , \9385 );
xor \U$9531 ( \9846 , \9845 , \9390 );
xor \U$9532 ( \9847 , \9397 , \9401 );
xor \U$9533 ( \9848 , \9847 , \9406 );
and \U$9534 ( \9849 , \9846 , \9848 );
xor \U$9535 ( \9850 , \9414 , \9418 );
xor \U$9536 ( \9851 , \9850 , \9423 );
and \U$9537 ( \9852 , \9848 , \9851 );
and \U$9538 ( \9853 , \9846 , \9851 );
or \U$9539 ( \9854 , \9849 , \9852 , \9853 );
and \U$9540 ( \9855 , \9844 , \9854 );
and \U$9541 ( \9856 , \8127 , \478 );
and \U$9542 ( \9857 , \7703 , \476 );
nor \U$9543 ( \9858 , \9856 , \9857 );
xnor \U$9544 ( \9859 , \9858 , \437 );
and \U$9545 ( \9860 , \8378 , \408 );
and \U$9546 ( \9861 , \8373 , \406 );
nor \U$9547 ( \9862 , \9860 , \9861 );
xnor \U$9548 ( \9863 , \9862 , \378 );
and \U$9549 ( \9864 , \9859 , \9863 );
and \U$9550 ( \9865 , \8981 , \360 );
and \U$9551 ( \9866 , \8697 , \358 );
nor \U$9552 ( \9867 , \9865 , \9866 );
xnor \U$9553 ( \9868 , \9867 , \341 );
and \U$9554 ( \9869 , \9863 , \9868 );
and \U$9555 ( \9870 , \9859 , \9868 );
or \U$9556 ( \9871 , \9864 , \9869 , \9870 );
xor \U$9557 ( \9872 , \9544 , \9548 );
xor \U$9558 ( \9873 , \9872 , \9554 );
and \U$9559 ( \9874 , \9871 , \9873 );
not \U$9560 ( \9875 , \9559 );
and \U$9561 ( \9876 , \9873 , \9875 );
and \U$9562 ( \9877 , \9871 , \9875 );
or \U$9563 ( \9878 , \9874 , \9876 , \9877 );
and \U$9564 ( \9879 , \9854 , \9878 );
and \U$9565 ( \9880 , \9844 , \9878 );
or \U$9566 ( \9881 , \9855 , \9879 , \9880 );
and \U$9567 ( \9882 , \9834 , \9881 );
xor \U$9568 ( \9883 , \9436 , \9440 );
xor \U$9569 ( \9884 , \9883 , \9445 );
xor \U$9570 ( \9885 , \9452 , \9456 );
xor \U$9571 ( \9886 , \9885 , \9461 );
and \U$9572 ( \9887 , \9884 , \9886 );
xor \U$9573 ( \9888 , \9469 , \9473 );
xor \U$9574 ( \9889 , \9888 , \9478 );
and \U$9575 ( \9890 , \9886 , \9889 );
and \U$9576 ( \9891 , \9884 , \9889 );
or \U$9577 ( \9892 , \9887 , \9890 , \9891 );
xor \U$9578 ( \9893 , \9124 , \9128 );
xor \U$9579 ( \9894 , \9893 , \9133 );
and \U$9580 ( \9895 , \9892 , \9894 );
xor \U$9581 ( \9896 , \9592 , \9594 );
xor \U$9582 ( \9897 , \9896 , \9597 );
and \U$9583 ( \9898 , \9894 , \9897 );
and \U$9584 ( \9899 , \9892 , \9897 );
or \U$9585 ( \9900 , \9895 , \9898 , \9899 );
and \U$9586 ( \9901 , \9881 , \9900 );
and \U$9587 ( \9902 , \9834 , \9900 );
or \U$9588 ( \9903 , \9882 , \9901 , \9902 );
xor \U$9589 ( \9904 , \9393 , \9409 );
xor \U$9590 ( \9905 , \9904 , \9426 );
xor \U$9591 ( \9906 , \9448 , \9464 );
xor \U$9592 ( \9907 , \9906 , \9481 );
and \U$9593 ( \9908 , \9905 , \9907 );
xor \U$9594 ( \9909 , \9501 , \9517 );
xor \U$9595 ( \9910 , \9909 , \9534 );
and \U$9596 ( \9911 , \9907 , \9910 );
and \U$9597 ( \9912 , \9905 , \9910 );
or \U$9598 ( \9913 , \9908 , \9911 , \9912 );
xor \U$9599 ( \9914 , \9557 , \9560 );
xor \U$9600 ( \9915 , \9914 , \9562 );
xor \U$9601 ( \9916 , \9567 , \9569 );
xor \U$9602 ( \9917 , \9916 , \9572 );
and \U$9603 ( \9918 , \9915 , \9917 );
xor \U$9604 ( \9919 , \9578 , \9580 );
xor \U$9605 ( \9920 , \9919 , \9583 );
and \U$9606 ( \9921 , \9917 , \9920 );
and \U$9607 ( \9922 , \9915 , \9920 );
or \U$9608 ( \9923 , \9918 , \9921 , \9922 );
and \U$9609 ( \9924 , \9913 , \9923 );
xor \U$9610 ( \9925 , \9188 , \9204 );
xor \U$9611 ( \9926 , \9925 , \9221 );
and \U$9612 ( \9927 , \9923 , \9926 );
and \U$9613 ( \9928 , \9913 , \9926 );
or \U$9614 ( \9929 , \9924 , \9927 , \9928 );
and \U$9615 ( \9930 , \9903 , \9929 );
xor \U$9616 ( \9931 , \9136 , \9152 );
xor \U$9617 ( \9932 , \9931 , \9169 );
xor \U$9618 ( \9933 , \9600 , \9602 );
xor \U$9619 ( \9934 , \9933 , \9605 );
and \U$9620 ( \9935 , \9932 , \9934 );
xor \U$9621 ( \9936 , \9624 , \9626 );
xor \U$9622 ( \9937 , \9936 , \9628 );
and \U$9623 ( \9938 , \9934 , \9937 );
and \U$9624 ( \9939 , \9932 , \9937 );
or \U$9625 ( \9940 , \9935 , \9938 , \9939 );
and \U$9626 ( \9941 , \9929 , \9940 );
and \U$9627 ( \9942 , \9903 , \9940 );
or \U$9628 ( \9943 , \9930 , \9941 , \9942 );
xor \U$9629 ( \9944 , \9540 , \9589 );
xor \U$9630 ( \9945 , \9944 , \9608 );
xor \U$9631 ( \9946 , \9613 , \9615 );
xor \U$9632 ( \9947 , \9946 , \9618 );
and \U$9633 ( \9948 , \9945 , \9947 );
xor \U$9634 ( \9949 , \9631 , \9633 );
xor \U$9635 ( \9950 , \9949 , \9636 );
and \U$9636 ( \9951 , \9947 , \9950 );
and \U$9637 ( \9952 , \9945 , \9950 );
or \U$9638 ( \9953 , \9948 , \9951 , \9952 );
and \U$9639 ( \9954 , \9943 , \9953 );
xor \U$9640 ( \9955 , \9312 , \9322 );
xor \U$9641 ( \9956 , \9955 , \9325 );
and \U$9642 ( \9957 , \9953 , \9956 );
and \U$9643 ( \9958 , \9943 , \9956 );
or \U$9644 ( \9959 , \9954 , \9957 , \9958 );
xor \U$9645 ( \9960 , \9118 , \9280 );
xor \U$9646 ( \9961 , \9960 , \9299 );
xor \U$9647 ( \9962 , \9611 , \9621 );
xor \U$9648 ( \9963 , \9962 , \9639 );
and \U$9649 ( \9964 , \9961 , \9963 );
xor \U$9650 ( \9965 , \9644 , \9646 );
xor \U$9651 ( \9966 , \9965 , \9649 );
and \U$9652 ( \9967 , \9963 , \9966 );
and \U$9653 ( \9968 , \9961 , \9966 );
or \U$9654 ( \9969 , \9964 , \9967 , \9968 );
and \U$9655 ( \9970 , \9959 , \9969 );
xor \U$9656 ( \9971 , \9302 , \9328 );
xor \U$9657 ( \9972 , \9971 , \9339 );
and \U$9658 ( \9973 , \9969 , \9972 );
and \U$9659 ( \9974 , \9959 , \9972 );
or \U$9660 ( \9975 , \9970 , \9973 , \9974 );
xor \U$9661 ( \9976 , \9658 , \9660 );
xor \U$9662 ( \9977 , \9976 , \9663 );
and \U$9663 ( \9978 , \9975 , \9977 );
and \U$9664 ( \9979 , \9672 , \9978 );
xor \U$9665 ( \9980 , \9672 , \9978 );
xor \U$9666 ( \9981 , \9975 , \9977 );
and \U$9667 ( \9982 , \789 , \6744 );
and \U$9668 ( \9983 , \709 , \6742 );
nor \U$9669 ( \9984 , \9982 , \9983 );
xnor \U$9670 ( \9985 , \9984 , \6429 );
and \U$9671 ( \9986 , \925 , \6235 );
and \U$9672 ( \9987 , \863 , \6233 );
nor \U$9673 ( \9988 , \9986 , \9987 );
xnor \U$9674 ( \9989 , \9988 , \5895 );
and \U$9675 ( \9990 , \9985 , \9989 );
and \U$9676 ( \9991 , \1186 , \5646 );
and \U$9677 ( \9992 , \988 , \5644 );
nor \U$9678 ( \9993 , \9991 , \9992 );
xnor \U$9679 ( \9994 , \9993 , \5405 );
and \U$9680 ( \9995 , \9989 , \9994 );
and \U$9681 ( \9996 , \9985 , \9994 );
or \U$9682 ( \9997 , \9990 , \9995 , \9996 );
xor \U$9683 ( \9998 , \9120 , \9758 );
xor \U$9684 ( \9999 , \9758 , \9759 );
not \U$9685 ( \10000 , \9999 );
and \U$9686 ( \10001 , \9998 , \10000 );
and \U$9687 ( \10002 , \316 , \10001 );
not \U$9688 ( \10003 , \10002 );
xnor \U$9689 ( \10004 , \10003 , \9762 );
and \U$9690 ( \10005 , \348 , \9433 );
and \U$9691 ( \10006 , \330 , \9431 );
nor \U$9692 ( \10007 , \10005 , \10006 );
xnor \U$9693 ( \10008 , \10007 , \9123 );
and \U$9694 ( \10009 , \10004 , \10008 );
and \U$9695 ( \10010 , \417 , \8896 );
and \U$9696 ( \10011 , \369 , \8894 );
nor \U$9697 ( \10012 , \10010 , \10011 );
xnor \U$9698 ( \10013 , \10012 , \8525 );
and \U$9699 ( \10014 , \10008 , \10013 );
and \U$9700 ( \10015 , \10004 , \10013 );
or \U$9701 ( \10016 , \10009 , \10014 , \10015 );
and \U$9702 ( \10017 , \9997 , \10016 );
and \U$9703 ( \10018 , \494 , \8334 );
and \U$9704 ( \10019 , \425 , \8332 );
nor \U$9705 ( \10020 , \10018 , \10019 );
xnor \U$9706 ( \10021 , \10020 , \8016 );
and \U$9707 ( \10022 , \553 , \7767 );
and \U$9708 ( \10023 , \499 , \7765 );
nor \U$9709 ( \10024 , \10022 , \10023 );
xnor \U$9710 ( \10025 , \10024 , \7518 );
and \U$9711 ( \10026 , \10021 , \10025 );
and \U$9712 ( \10027 , \681 , \7238 );
and \U$9713 ( \10028 , \604 , \7236 );
nor \U$9714 ( \10029 , \10027 , \10028 );
xnor \U$9715 ( \10030 , \10029 , \6978 );
and \U$9716 ( \10031 , \10025 , \10030 );
and \U$9717 ( \10032 , \10021 , \10030 );
or \U$9718 ( \10033 , \10026 , \10031 , \10032 );
and \U$9719 ( \10034 , \10016 , \10033 );
and \U$9720 ( \10035 , \9997 , \10033 );
or \U$9721 ( \10036 , \10017 , \10034 , \10035 );
and \U$9722 ( \10037 , \6500 , \826 );
and \U$9723 ( \10038 , \6157 , \824 );
nor \U$9724 ( \10039 , \10037 , \10038 );
xnor \U$9725 ( \10040 , \10039 , \754 );
and \U$9726 ( \10041 , \7005 , \692 );
and \U$9727 ( \10042 , \6702 , \690 );
nor \U$9728 ( \10043 , \10041 , \10042 );
xnor \U$9729 ( \10044 , \10043 , \649 );
and \U$9730 ( \10045 , \10040 , \10044 );
and \U$9731 ( \10046 , \7703 , \579 );
and \U$9732 ( \10047 , \7177 , \577 );
nor \U$9733 ( \10048 , \10046 , \10047 );
xnor \U$9734 ( \10049 , \10048 , \530 );
and \U$9735 ( \10050 , \10044 , \10049 );
and \U$9736 ( \10051 , \10040 , \10049 );
or \U$9737 ( \10052 , \10045 , \10050 , \10051 );
and \U$9738 ( \10053 , \4011 , \2094 );
and \U$9739 ( \10054 , \3889 , \2092 );
nor \U$9740 ( \10055 , \10053 , \10054 );
xnor \U$9741 ( \10056 , \10055 , \1942 );
and \U$9742 ( \10057 , \4272 , \1826 );
and \U$9743 ( \10058 , \4016 , \1824 );
nor \U$9744 ( \10059 , \10057 , \10058 );
xnor \U$9745 ( \10060 , \10059 , \1670 );
and \U$9746 ( \10061 , \10056 , \10060 );
and \U$9747 ( \10062 , \4771 , \1554 );
and \U$9748 ( \10063 , \4469 , \1552 );
nor \U$9749 ( \10064 , \10062 , \10063 );
xnor \U$9750 ( \10065 , \10064 , \1441 );
and \U$9751 ( \10066 , \10060 , \10065 );
and \U$9752 ( \10067 , \10056 , \10065 );
or \U$9753 ( \10068 , \10061 , \10066 , \10067 );
and \U$9754 ( \10069 , \10052 , \10068 );
and \U$9755 ( \10070 , \5248 , \1360 );
and \U$9756 ( \10071 , \4779 , \1358 );
nor \U$9757 ( \10072 , \10070 , \10071 );
xnor \U$9758 ( \10073 , \10072 , \1224 );
and \U$9759 ( \10074 , \5517 , \1160 );
and \U$9760 ( \10075 , \5253 , \1158 );
nor \U$9761 ( \10076 , \10074 , \10075 );
xnor \U$9762 ( \10077 , \10076 , \1082 );
and \U$9763 ( \10078 , \10073 , \10077 );
and \U$9764 ( \10079 , \6148 , \996 );
and \U$9765 ( \10080 , \5776 , \994 );
nor \U$9766 ( \10081 , \10079 , \10080 );
xnor \U$9767 ( \10082 , \10081 , \902 );
and \U$9768 ( \10083 , \10077 , \10082 );
and \U$9769 ( \10084 , \10073 , \10082 );
or \U$9770 ( \10085 , \10078 , \10083 , \10084 );
and \U$9771 ( \10086 , \10068 , \10085 );
and \U$9772 ( \10087 , \10052 , \10085 );
or \U$9773 ( \10088 , \10069 , \10086 , \10087 );
and \U$9774 ( \10089 , \10036 , \10088 );
and \U$9775 ( \10090 , \1379 , \5180 );
and \U$9776 ( \10091 , \1274 , \5178 );
nor \U$9777 ( \10092 , \10090 , \10091 );
xnor \U$9778 ( \10093 , \10092 , \4992 );
and \U$9779 ( \10094 , \1500 , \4806 );
and \U$9780 ( \10095 , \1384 , \4804 );
nor \U$9781 ( \10096 , \10094 , \10095 );
xnor \U$9782 ( \10097 , \10096 , \4574 );
and \U$9783 ( \10098 , \10093 , \10097 );
and \U$9784 ( \10099 , \1791 , \4355 );
and \U$9785 ( \10100 , \1615 , \4353 );
nor \U$9786 ( \10101 , \10099 , \10100 );
xnor \U$9787 ( \10102 , \10101 , \4212 );
and \U$9788 ( \10103 , \10097 , \10102 );
and \U$9789 ( \10104 , \10093 , \10102 );
or \U$9790 ( \10105 , \10098 , \10103 , \10104 );
and \U$9791 ( \10106 , \2840 , \2918 );
and \U$9792 ( \10107 , \2666 , \2916 );
nor \U$9793 ( \10108 , \10106 , \10107 );
xnor \U$9794 ( \10109 , \10108 , \2769 );
and \U$9795 ( \10110 , \3145 , \2596 );
and \U$9796 ( \10111 , \3007 , \2594 );
nor \U$9797 ( \10112 , \10110 , \10111 );
xnor \U$9798 ( \10113 , \10112 , \2454 );
and \U$9799 ( \10114 , \10109 , \10113 );
and \U$9800 ( \10115 , \3681 , \2300 );
and \U$9801 ( \10116 , \3264 , \2298 );
nor \U$9802 ( \10117 , \10115 , \10116 );
xnor \U$9803 ( \10118 , \10117 , \2163 );
and \U$9804 ( \10119 , \10113 , \10118 );
and \U$9805 ( \10120 , \10109 , \10118 );
or \U$9806 ( \10121 , \10114 , \10119 , \10120 );
and \U$9807 ( \10122 , \10105 , \10121 );
and \U$9808 ( \10123 , \2042 , \4032 );
and \U$9809 ( \10124 , \1799 , \4030 );
nor \U$9810 ( \10125 , \10123 , \10124 );
xnor \U$9811 ( \10126 , \10125 , \3786 );
and \U$9812 ( \10127 , \2233 , \3637 );
and \U$9813 ( \10128 , \2047 , \3635 );
nor \U$9814 ( \10129 , \10127 , \10128 );
xnor \U$9815 ( \10130 , \10129 , \3450 );
and \U$9816 ( \10131 , \10126 , \10130 );
and \U$9817 ( \10132 , \2641 , \3324 );
and \U$9818 ( \10133 , \2377 , \3322 );
nor \U$9819 ( \10134 , \10132 , \10133 );
xnor \U$9820 ( \10135 , \10134 , \3119 );
and \U$9821 ( \10136 , \10130 , \10135 );
and \U$9822 ( \10137 , \10126 , \10135 );
or \U$9823 ( \10138 , \10131 , \10136 , \10137 );
and \U$9824 ( \10139 , \10121 , \10138 );
and \U$9825 ( \10140 , \10105 , \10138 );
or \U$9826 ( \10141 , \10122 , \10139 , \10140 );
and \U$9827 ( \10142 , \10088 , \10141 );
and \U$9828 ( \10143 , \10036 , \10141 );
or \U$9829 ( \10144 , \10089 , \10142 , \10143 );
and \U$9830 ( \10145 , \8373 , \478 );
and \U$9831 ( \10146 , \8127 , \476 );
nor \U$9832 ( \10147 , \10145 , \10146 );
xnor \U$9833 ( \10148 , \10147 , \437 );
and \U$9834 ( \10149 , \8697 , \408 );
and \U$9835 ( \10150 , \8378 , \406 );
nor \U$9836 ( \10151 , \10149 , \10150 );
xnor \U$9837 ( \10152 , \10151 , \378 );
and \U$9838 ( \10153 , \10148 , \10152 );
and \U$9839 ( \10154 , \9550 , \360 );
and \U$9840 ( \10155 , \8981 , \358 );
nor \U$9841 ( \10156 , \10154 , \10155 );
xnor \U$9842 ( \10157 , \10156 , \341 );
and \U$9843 ( \10158 , \10152 , \10157 );
and \U$9844 ( \10159 , \10148 , \10157 );
or \U$9845 ( \10160 , \10153 , \10158 , \10159 );
buf \U$9846 ( \10161 , RIc0c5d30_126);
and \U$9847 ( \10162 , \10161 , \323 );
and \U$9848 ( \10163 , \9558 , \321 );
nor \U$9849 ( \10164 , \10162 , \10163 );
xnor \U$9850 ( \10165 , \10164 , \328 );
buf \U$9851 ( \10166 , RIc340530_127);
and \U$9852 ( \10167 , \10166 , \317 );
or \U$9853 ( \10168 , \10165 , \10167 );
and \U$9854 ( \10169 , \10160 , \10168 );
and \U$9855 ( \10170 , \9558 , \323 );
and \U$9856 ( \10171 , \9550 , \321 );
nor \U$9857 ( \10172 , \10170 , \10171 );
xnor \U$9858 ( \10173 , \10172 , \328 );
and \U$9859 ( \10174 , \10168 , \10173 );
and \U$9860 ( \10175 , \10160 , \10173 );
or \U$9861 ( \10176 , \10169 , \10174 , \10175 );
and \U$9862 ( \10177 , \10161 , \317 );
xor \U$9863 ( \10178 , \9783 , \9787 );
xor \U$9864 ( \10179 , \10178 , \9792 );
and \U$9865 ( \10180 , \10177 , \10179 );
xor \U$9866 ( \10181 , \9859 , \9863 );
xor \U$9867 ( \10182 , \10181 , \9868 );
and \U$9868 ( \10183 , \10179 , \10182 );
and \U$9869 ( \10184 , \10177 , \10182 );
or \U$9870 ( \10185 , \10180 , \10183 , \10184 );
and \U$9871 ( \10186 , \10176 , \10185 );
xor \U$9872 ( \10187 , \9676 , \9680 );
xor \U$9873 ( \10188 , \10187 , \9685 );
xor \U$9874 ( \10189 , \9799 , \9803 );
xor \U$9875 ( \10190 , \10189 , \9808 );
and \U$9876 ( \10191 , \10188 , \10190 );
xor \U$9877 ( \10192 , \9816 , \9820 );
xor \U$9878 ( \10193 , \10192 , \9825 );
and \U$9879 ( \10194 , \10190 , \10193 );
and \U$9880 ( \10195 , \10188 , \10193 );
or \U$9881 ( \10196 , \10191 , \10194 , \10195 );
and \U$9882 ( \10197 , \10185 , \10196 );
and \U$9883 ( \10198 , \10176 , \10196 );
or \U$9884 ( \10199 , \10186 , \10197 , \10198 );
and \U$9885 ( \10200 , \10144 , \10199 );
xor \U$9886 ( \10201 , \9728 , \9732 );
xor \U$9887 ( \10202 , \10201 , \9737 );
xor \U$9888 ( \10203 , \9692 , \9696 );
xor \U$9889 ( \10204 , \10203 , \9701 );
and \U$9890 ( \10205 , \10202 , \10204 );
xor \U$9891 ( \10206 , \9709 , \9713 );
xor \U$9892 ( \10207 , \10206 , \9718 );
and \U$9893 ( \10208 , \10204 , \10207 );
and \U$9894 ( \10209 , \10202 , \10207 );
or \U$9895 ( \10210 , \10205 , \10208 , \10209 );
xor \U$9896 ( \10211 , \9744 , \9748 );
xor \U$9897 ( \10212 , \10211 , \9753 );
xor \U$9898 ( \10213 , \9763 , \9767 );
xor \U$9899 ( \10214 , \10213 , \9772 );
and \U$9900 ( \10215 , \10212 , \10214 );
and \U$9901 ( \10216 , \10210 , \10215 );
xor \U$9902 ( \10217 , \9884 , \9886 );
xor \U$9903 ( \10218 , \10217 , \9889 );
and \U$9904 ( \10219 , \10215 , \10218 );
and \U$9905 ( \10220 , \10210 , \10218 );
or \U$9906 ( \10221 , \10216 , \10219 , \10220 );
and \U$9907 ( \10222 , \10199 , \10221 );
and \U$9908 ( \10223 , \10144 , \10221 );
or \U$9909 ( \10224 , \10200 , \10222 , \10223 );
xor \U$9910 ( \10225 , \9688 , \9704 );
xor \U$9911 ( \10226 , \10225 , \9721 );
xor \U$9912 ( \10227 , \9740 , \9756 );
xor \U$9913 ( \10228 , \10227 , \9775 );
and \U$9914 ( \10229 , \10226 , \10228 );
xor \U$9915 ( \10230 , \9795 , \9811 );
xor \U$9916 ( \10231 , \10230 , \9828 );
and \U$9917 ( \10232 , \10228 , \10231 );
and \U$9918 ( \10233 , \10226 , \10231 );
or \U$9919 ( \10234 , \10229 , \10232 , \10233 );
xor \U$9920 ( \10235 , \9836 , \9838 );
xor \U$9921 ( \10236 , \10235 , \9841 );
xor \U$9922 ( \10237 , \9846 , \9848 );
xor \U$9923 ( \10238 , \10237 , \9851 );
and \U$9924 ( \10239 , \10236 , \10238 );
xor \U$9925 ( \10240 , \9871 , \9873 );
xor \U$9926 ( \10241 , \10240 , \9875 );
and \U$9927 ( \10242 , \10238 , \10241 );
and \U$9928 ( \10243 , \10236 , \10241 );
or \U$9929 ( \10244 , \10239 , \10242 , \10243 );
and \U$9930 ( \10245 , \10234 , \10244 );
xor \U$9931 ( \10246 , \9905 , \9907 );
xor \U$9932 ( \10247 , \10246 , \9910 );
and \U$9933 ( \10248 , \10244 , \10247 );
and \U$9934 ( \10249 , \10234 , \10247 );
or \U$9935 ( \10250 , \10245 , \10248 , \10249 );
and \U$9936 ( \10251 , \10224 , \10250 );
xor \U$9937 ( \10252 , \9844 , \9854 );
xor \U$9938 ( \10253 , \10252 , \9878 );
xor \U$9939 ( \10254 , \9915 , \9917 );
xor \U$9940 ( \10255 , \10254 , \9920 );
and \U$9941 ( \10256 , \10253 , \10255 );
xor \U$9942 ( \10257 , \9892 , \9894 );
xor \U$9943 ( \10258 , \10257 , \9897 );
and \U$9944 ( \10259 , \10255 , \10258 );
and \U$9945 ( \10260 , \10253 , \10258 );
or \U$9946 ( \10261 , \10256 , \10259 , \10260 );
and \U$9947 ( \10262 , \10250 , \10261 );
and \U$9948 ( \10263 , \10224 , \10261 );
or \U$9949 ( \10264 , \10251 , \10262 , \10263 );
xor \U$9950 ( \10265 , \9429 , \9484 );
xor \U$9951 ( \10266 , \10265 , \9537 );
xor \U$9952 ( \10267 , \9565 , \9575 );
xor \U$9953 ( \10268 , \10267 , \9586 );
and \U$9954 ( \10269 , \10266 , \10268 );
xor \U$9955 ( \10270 , \9932 , \9934 );
xor \U$9956 ( \10271 , \10270 , \9937 );
and \U$9957 ( \10272 , \10268 , \10271 );
and \U$9958 ( \10273 , \10266 , \10271 );
or \U$9959 ( \10274 , \10269 , \10272 , \10273 );
and \U$9960 ( \10275 , \10264 , \10274 );
xor \U$9961 ( \10276 , \9945 , \9947 );
xor \U$9962 ( \10277 , \10276 , \9950 );
and \U$9963 ( \10278 , \10274 , \10277 );
and \U$9964 ( \10279 , \10264 , \10277 );
or \U$9965 ( \10280 , \10275 , \10278 , \10279 );
xor \U$9966 ( \10281 , \9943 , \9953 );
xor \U$9967 ( \10282 , \10281 , \9956 );
and \U$9968 ( \10283 , \10280 , \10282 );
xor \U$9969 ( \10284 , \9961 , \9963 );
xor \U$9970 ( \10285 , \10284 , \9966 );
and \U$9971 ( \10286 , \10282 , \10285 );
and \U$9972 ( \10287 , \10280 , \10285 );
or \U$9973 ( \10288 , \10283 , \10286 , \10287 );
xor \U$9974 ( \10289 , \9959 , \9969 );
xor \U$9975 ( \10290 , \10289 , \9972 );
and \U$9976 ( \10291 , \10288 , \10290 );
xor \U$9977 ( \10292 , \9642 , \9652 );
xor \U$9978 ( \10293 , \10292 , \9655 );
and \U$9979 ( \10294 , \10290 , \10293 );
and \U$9980 ( \10295 , \10288 , \10293 );
or \U$9981 ( \10296 , \10291 , \10294 , \10295 );
and \U$9982 ( \10297 , \9981 , \10296 );
xor \U$9983 ( \10298 , \9981 , \10296 );
xor \U$9984 ( \10299 , \10288 , \10290 );
xor \U$9985 ( \10300 , \10299 , \10293 );
xor \U$9986 ( \10301 , \10109 , \10113 );
xor \U$9987 ( \10302 , \10301 , \10118 );
xor \U$9988 ( \10303 , \10126 , \10130 );
xor \U$9989 ( \10304 , \10303 , \10135 );
and \U$9990 ( \10305 , \10302 , \10304 );
xor \U$9991 ( \10306 , \10056 , \10060 );
xor \U$9992 ( \10307 , \10306 , \10065 );
and \U$9993 ( \10308 , \10304 , \10307 );
and \U$9994 ( \10309 , \10302 , \10307 );
or \U$9995 ( \10310 , \10305 , \10308 , \10309 );
xor \U$9996 ( \10311 , \10040 , \10044 );
xor \U$9997 ( \10312 , \10311 , \10049 );
xor \U$9998 ( \10313 , \10148 , \10152 );
xor \U$9999 ( \10314 , \10313 , \10157 );
and \U$10000 ( \10315 , \10312 , \10314 );
xor \U$10001 ( \10316 , \10073 , \10077 );
xor \U$10002 ( \10317 , \10316 , \10082 );
and \U$10003 ( \10318 , \10314 , \10317 );
and \U$10004 ( \10319 , \10312 , \10317 );
or \U$10005 ( \10320 , \10315 , \10318 , \10319 );
and \U$10006 ( \10321 , \10310 , \10320 );
and \U$10007 ( \10322 , \8127 , \579 );
and \U$10008 ( \10323 , \7703 , \577 );
nor \U$10009 ( \10324 , \10322 , \10323 );
xnor \U$10010 ( \10325 , \10324 , \530 );
and \U$10011 ( \10326 , \8378 , \478 );
and \U$10012 ( \10327 , \8373 , \476 );
nor \U$10013 ( \10328 , \10326 , \10327 );
xnor \U$10014 ( \10329 , \10328 , \437 );
and \U$10015 ( \10330 , \10325 , \10329 );
and \U$10016 ( \10331 , \8981 , \408 );
and \U$10017 ( \10332 , \8697 , \406 );
nor \U$10018 ( \10333 , \10331 , \10332 );
xnor \U$10019 ( \10334 , \10333 , \378 );
and \U$10020 ( \10335 , \10329 , \10334 );
and \U$10021 ( \10336 , \10325 , \10334 );
or \U$10022 ( \10337 , \10330 , \10335 , \10336 );
and \U$10023 ( \10338 , \9558 , \360 );
and \U$10024 ( \10339 , \9550 , \358 );
nor \U$10025 ( \10340 , \10338 , \10339 );
xnor \U$10026 ( \10341 , \10340 , \341 );
and \U$10027 ( \10342 , \10166 , \323 );
and \U$10028 ( \10343 , \10161 , \321 );
nor \U$10029 ( \10344 , \10342 , \10343 );
xnor \U$10030 ( \10345 , \10344 , \328 );
and \U$10031 ( \10346 , \10341 , \10345 );
buf \U$10032 ( \10347 , RIc3405a8_128);
and \U$10033 ( \10348 , \10347 , \317 );
and \U$10034 ( \10349 , \10345 , \10348 );
and \U$10035 ( \10350 , \10341 , \10348 );
or \U$10036 ( \10351 , \10346 , \10349 , \10350 );
and \U$10037 ( \10352 , \10337 , \10351 );
xnor \U$10038 ( \10353 , \10165 , \10167 );
and \U$10039 ( \10354 , \10351 , \10353 );
and \U$10040 ( \10355 , \10337 , \10353 );
or \U$10041 ( \10356 , \10352 , \10354 , \10355 );
and \U$10042 ( \10357 , \10320 , \10356 );
and \U$10043 ( \10358 , \10310 , \10356 );
or \U$10044 ( \10359 , \10321 , \10357 , \10358 );
not \U$10045 ( \10360 , \9759 );
and \U$10046 ( \10361 , \330 , \10001 );
and \U$10047 ( \10362 , \316 , \9999 );
nor \U$10048 ( \10363 , \10361 , \10362 );
xnor \U$10049 ( \10364 , \10363 , \9762 );
and \U$10050 ( \10365 , \10360 , \10364 );
and \U$10051 ( \10366 , \369 , \9433 );
and \U$10052 ( \10367 , \348 , \9431 );
nor \U$10053 ( \10368 , \10366 , \10367 );
xnor \U$10054 ( \10369 , \10368 , \9123 );
and \U$10055 ( \10370 , \10364 , \10369 );
and \U$10056 ( \10371 , \10360 , \10369 );
or \U$10057 ( \10372 , \10365 , \10370 , \10371 );
and \U$10058 ( \10373 , \425 , \8896 );
and \U$10059 ( \10374 , \417 , \8894 );
nor \U$10060 ( \10375 , \10373 , \10374 );
xnor \U$10061 ( \10376 , \10375 , \8525 );
and \U$10062 ( \10377 , \499 , \8334 );
and \U$10063 ( \10378 , \494 , \8332 );
nor \U$10064 ( \10379 , \10377 , \10378 );
xnor \U$10065 ( \10380 , \10379 , \8016 );
and \U$10066 ( \10381 , \10376 , \10380 );
and \U$10067 ( \10382 , \604 , \7767 );
and \U$10068 ( \10383 , \553 , \7765 );
nor \U$10069 ( \10384 , \10382 , \10383 );
xnor \U$10070 ( \10385 , \10384 , \7518 );
and \U$10071 ( \10386 , \10380 , \10385 );
and \U$10072 ( \10387 , \10376 , \10385 );
or \U$10073 ( \10388 , \10381 , \10386 , \10387 );
and \U$10074 ( \10389 , \10372 , \10388 );
and \U$10075 ( \10390 , \709 , \7238 );
and \U$10076 ( \10391 , \681 , \7236 );
nor \U$10077 ( \10392 , \10390 , \10391 );
xnor \U$10078 ( \10393 , \10392 , \6978 );
and \U$10079 ( \10394 , \863 , \6744 );
and \U$10080 ( \10395 , \789 , \6742 );
nor \U$10081 ( \10396 , \10394 , \10395 );
xnor \U$10082 ( \10397 , \10396 , \6429 );
and \U$10083 ( \10398 , \10393 , \10397 );
and \U$10084 ( \10399 , \988 , \6235 );
and \U$10085 ( \10400 , \925 , \6233 );
nor \U$10086 ( \10401 , \10399 , \10400 );
xnor \U$10087 ( \10402 , \10401 , \5895 );
and \U$10088 ( \10403 , \10397 , \10402 );
and \U$10089 ( \10404 , \10393 , \10402 );
or \U$10090 ( \10405 , \10398 , \10403 , \10404 );
and \U$10091 ( \10406 , \10388 , \10405 );
and \U$10092 ( \10407 , \10372 , \10405 );
or \U$10093 ( \10408 , \10389 , \10406 , \10407 );
and \U$10094 ( \10409 , \4779 , \1554 );
and \U$10095 ( \10410 , \4771 , \1552 );
nor \U$10096 ( \10411 , \10409 , \10410 );
xnor \U$10097 ( \10412 , \10411 , \1441 );
and \U$10098 ( \10413 , \5253 , \1360 );
and \U$10099 ( \10414 , \5248 , \1358 );
nor \U$10100 ( \10415 , \10413 , \10414 );
xnor \U$10101 ( \10416 , \10415 , \1224 );
and \U$10102 ( \10417 , \10412 , \10416 );
and \U$10103 ( \10418 , \5776 , \1160 );
and \U$10104 ( \10419 , \5517 , \1158 );
nor \U$10105 ( \10420 , \10418 , \10419 );
xnor \U$10106 ( \10421 , \10420 , \1082 );
and \U$10107 ( \10422 , \10416 , \10421 );
and \U$10108 ( \10423 , \10412 , \10421 );
or \U$10109 ( \10424 , \10417 , \10422 , \10423 );
and \U$10110 ( \10425 , \3889 , \2300 );
and \U$10111 ( \10426 , \3681 , \2298 );
nor \U$10112 ( \10427 , \10425 , \10426 );
xnor \U$10113 ( \10428 , \10427 , \2163 );
and \U$10114 ( \10429 , \4016 , \2094 );
and \U$10115 ( \10430 , \4011 , \2092 );
nor \U$10116 ( \10431 , \10429 , \10430 );
xnor \U$10117 ( \10432 , \10431 , \1942 );
and \U$10118 ( \10433 , \10428 , \10432 );
and \U$10119 ( \10434 , \4469 , \1826 );
and \U$10120 ( \10435 , \4272 , \1824 );
nor \U$10121 ( \10436 , \10434 , \10435 );
xnor \U$10122 ( \10437 , \10436 , \1670 );
and \U$10123 ( \10438 , \10432 , \10437 );
and \U$10124 ( \10439 , \10428 , \10437 );
or \U$10125 ( \10440 , \10433 , \10438 , \10439 );
and \U$10126 ( \10441 , \10424 , \10440 );
and \U$10127 ( \10442 , \6157 , \996 );
and \U$10128 ( \10443 , \6148 , \994 );
nor \U$10129 ( \10444 , \10442 , \10443 );
xnor \U$10130 ( \10445 , \10444 , \902 );
and \U$10131 ( \10446 , \6702 , \826 );
and \U$10132 ( \10447 , \6500 , \824 );
nor \U$10133 ( \10448 , \10446 , \10447 );
xnor \U$10134 ( \10449 , \10448 , \754 );
and \U$10135 ( \10450 , \10445 , \10449 );
and \U$10136 ( \10451 , \7177 , \692 );
and \U$10137 ( \10452 , \7005 , \690 );
nor \U$10138 ( \10453 , \10451 , \10452 );
xnor \U$10139 ( \10454 , \10453 , \649 );
and \U$10140 ( \10455 , \10449 , \10454 );
and \U$10141 ( \10456 , \10445 , \10454 );
or \U$10142 ( \10457 , \10450 , \10455 , \10456 );
and \U$10143 ( \10458 , \10440 , \10457 );
and \U$10144 ( \10459 , \10424 , \10457 );
or \U$10145 ( \10460 , \10441 , \10458 , \10459 );
and \U$10146 ( \10461 , \10408 , \10460 );
and \U$10147 ( \10462 , \1799 , \4355 );
and \U$10148 ( \10463 , \1791 , \4353 );
nor \U$10149 ( \10464 , \10462 , \10463 );
xnor \U$10150 ( \10465 , \10464 , \4212 );
and \U$10151 ( \10466 , \2047 , \4032 );
and \U$10152 ( \10467 , \2042 , \4030 );
nor \U$10153 ( \10468 , \10466 , \10467 );
xnor \U$10154 ( \10469 , \10468 , \3786 );
and \U$10155 ( \10470 , \10465 , \10469 );
and \U$10156 ( \10471 , \2377 , \3637 );
and \U$10157 ( \10472 , \2233 , \3635 );
nor \U$10158 ( \10473 , \10471 , \10472 );
xnor \U$10159 ( \10474 , \10473 , \3450 );
and \U$10160 ( \10475 , \10469 , \10474 );
and \U$10161 ( \10476 , \10465 , \10474 );
or \U$10162 ( \10477 , \10470 , \10475 , \10476 );
and \U$10163 ( \10478 , \2666 , \3324 );
and \U$10164 ( \10479 , \2641 , \3322 );
nor \U$10165 ( \10480 , \10478 , \10479 );
xnor \U$10166 ( \10481 , \10480 , \3119 );
and \U$10167 ( \10482 , \3007 , \2918 );
and \U$10168 ( \10483 , \2840 , \2916 );
nor \U$10169 ( \10484 , \10482 , \10483 );
xnor \U$10170 ( \10485 , \10484 , \2769 );
and \U$10171 ( \10486 , \10481 , \10485 );
and \U$10172 ( \10487 , \3264 , \2596 );
and \U$10173 ( \10488 , \3145 , \2594 );
nor \U$10174 ( \10489 , \10487 , \10488 );
xnor \U$10175 ( \10490 , \10489 , \2454 );
and \U$10176 ( \10491 , \10485 , \10490 );
and \U$10177 ( \10492 , \10481 , \10490 );
or \U$10178 ( \10493 , \10486 , \10491 , \10492 );
and \U$10179 ( \10494 , \10477 , \10493 );
and \U$10180 ( \10495 , \1274 , \5646 );
and \U$10181 ( \10496 , \1186 , \5644 );
nor \U$10182 ( \10497 , \10495 , \10496 );
xnor \U$10183 ( \10498 , \10497 , \5405 );
and \U$10184 ( \10499 , \1384 , \5180 );
and \U$10185 ( \10500 , \1379 , \5178 );
nor \U$10186 ( \10501 , \10499 , \10500 );
xnor \U$10187 ( \10502 , \10501 , \4992 );
and \U$10188 ( \10503 , \10498 , \10502 );
and \U$10189 ( \10504 , \1615 , \4806 );
and \U$10190 ( \10505 , \1500 , \4804 );
nor \U$10191 ( \10506 , \10504 , \10505 );
xnor \U$10192 ( \10507 , \10506 , \4574 );
and \U$10193 ( \10508 , \10502 , \10507 );
and \U$10194 ( \10509 , \10498 , \10507 );
or \U$10195 ( \10510 , \10503 , \10508 , \10509 );
and \U$10196 ( \10511 , \10493 , \10510 );
and \U$10197 ( \10512 , \10477 , \10510 );
or \U$10198 ( \10513 , \10494 , \10511 , \10512 );
and \U$10199 ( \10514 , \10460 , \10513 );
and \U$10200 ( \10515 , \10408 , \10513 );
or \U$10201 ( \10516 , \10461 , \10514 , \10515 );
and \U$10202 ( \10517 , \10359 , \10516 );
xor \U$10203 ( \10518 , \10093 , \10097 );
xor \U$10204 ( \10519 , \10518 , \10102 );
xor \U$10205 ( \10520 , \9985 , \9989 );
xor \U$10206 ( \10521 , \10520 , \9994 );
and \U$10207 ( \10522 , \10519 , \10521 );
xor \U$10208 ( \10523 , \10021 , \10025 );
xor \U$10209 ( \10524 , \10523 , \10030 );
and \U$10210 ( \10525 , \10521 , \10524 );
and \U$10211 ( \10526 , \10519 , \10524 );
or \U$10212 ( \10527 , \10522 , \10525 , \10526 );
xor \U$10213 ( \10528 , \10202 , \10204 );
xor \U$10214 ( \10529 , \10528 , \10207 );
and \U$10215 ( \10530 , \10527 , \10529 );
xor \U$10216 ( \10531 , \10212 , \10214 );
and \U$10217 ( \10532 , \10529 , \10531 );
and \U$10218 ( \10533 , \10527 , \10531 );
or \U$10219 ( \10534 , \10530 , \10532 , \10533 );
and \U$10220 ( \10535 , \10516 , \10534 );
and \U$10221 ( \10536 , \10359 , \10534 );
or \U$10222 ( \10537 , \10517 , \10535 , \10536 );
xor \U$10223 ( \10538 , \9997 , \10016 );
xor \U$10224 ( \10539 , \10538 , \10033 );
xor \U$10225 ( \10540 , \10052 , \10068 );
xor \U$10226 ( \10541 , \10540 , \10085 );
and \U$10227 ( \10542 , \10539 , \10541 );
xor \U$10228 ( \10543 , \10105 , \10121 );
xor \U$10229 ( \10544 , \10543 , \10138 );
and \U$10230 ( \10545 , \10541 , \10544 );
and \U$10231 ( \10546 , \10539 , \10544 );
or \U$10232 ( \10547 , \10542 , \10545 , \10546 );
xor \U$10233 ( \10548 , \10160 , \10168 );
xor \U$10234 ( \10549 , \10548 , \10173 );
xor \U$10235 ( \10550 , \10177 , \10179 );
xor \U$10236 ( \10551 , \10550 , \10182 );
and \U$10237 ( \10552 , \10549 , \10551 );
xor \U$10238 ( \10553 , \10188 , \10190 );
xor \U$10239 ( \10554 , \10553 , \10193 );
and \U$10240 ( \10555 , \10551 , \10554 );
and \U$10241 ( \10556 , \10549 , \10554 );
or \U$10242 ( \10557 , \10552 , \10555 , \10556 );
and \U$10243 ( \10558 , \10547 , \10557 );
xor \U$10244 ( \10559 , \10226 , \10228 );
xor \U$10245 ( \10560 , \10559 , \10231 );
and \U$10246 ( \10561 , \10557 , \10560 );
and \U$10247 ( \10562 , \10547 , \10560 );
or \U$10248 ( \10563 , \10558 , \10561 , \10562 );
and \U$10249 ( \10564 , \10537 , \10563 );
xor \U$10250 ( \10565 , \10176 , \10185 );
xor \U$10251 ( \10566 , \10565 , \10196 );
xor \U$10252 ( \10567 , \10210 , \10215 );
xor \U$10253 ( \10568 , \10567 , \10218 );
and \U$10254 ( \10569 , \10566 , \10568 );
xor \U$10255 ( \10570 , \10236 , \10238 );
xor \U$10256 ( \10571 , \10570 , \10241 );
and \U$10257 ( \10572 , \10568 , \10571 );
and \U$10258 ( \10573 , \10566 , \10571 );
or \U$10259 ( \10574 , \10569 , \10572 , \10573 );
and \U$10260 ( \10575 , \10563 , \10574 );
and \U$10261 ( \10576 , \10537 , \10574 );
or \U$10262 ( \10577 , \10564 , \10575 , \10576 );
xor \U$10263 ( \10578 , \9724 , \9778 );
xor \U$10264 ( \10579 , \10578 , \9831 );
xor \U$10265 ( \10580 , \10234 , \10244 );
xor \U$10266 ( \10581 , \10580 , \10247 );
and \U$10267 ( \10582 , \10579 , \10581 );
xor \U$10268 ( \10583 , \10253 , \10255 );
xor \U$10269 ( \10584 , \10583 , \10258 );
and \U$10270 ( \10585 , \10581 , \10584 );
and \U$10271 ( \10586 , \10579 , \10584 );
or \U$10272 ( \10587 , \10582 , \10585 , \10586 );
and \U$10273 ( \10588 , \10577 , \10587 );
xor \U$10274 ( \10589 , \9913 , \9923 );
xor \U$10275 ( \10590 , \10589 , \9926 );
and \U$10276 ( \10591 , \10587 , \10590 );
and \U$10277 ( \10592 , \10577 , \10590 );
or \U$10278 ( \10593 , \10588 , \10591 , \10592 );
xor \U$10279 ( \10594 , \9834 , \9881 );
xor \U$10280 ( \10595 , \10594 , \9900 );
xor \U$10281 ( \10596 , \10224 , \10250 );
xor \U$10282 ( \10597 , \10596 , \10261 );
and \U$10283 ( \10598 , \10595 , \10597 );
xor \U$10284 ( \10599 , \10266 , \10268 );
xor \U$10285 ( \10600 , \10599 , \10271 );
and \U$10286 ( \10601 , \10597 , \10600 );
and \U$10287 ( \10602 , \10595 , \10600 );
or \U$10288 ( \10603 , \10598 , \10601 , \10602 );
and \U$10289 ( \10604 , \10593 , \10603 );
xor \U$10290 ( \10605 , \9903 , \9929 );
xor \U$10291 ( \10606 , \10605 , \9940 );
and \U$10292 ( \10607 , \10603 , \10606 );
and \U$10293 ( \10608 , \10593 , \10606 );
or \U$10294 ( \10609 , \10604 , \10607 , \10608 );
xor \U$10295 ( \10610 , \10280 , \10282 );
xor \U$10296 ( \10611 , \10610 , \10285 );
and \U$10297 ( \10612 , \10609 , \10611 );
and \U$10298 ( \10613 , \10300 , \10612 );
xor \U$10299 ( \10614 , \10300 , \10612 );
xor \U$10300 ( \10615 , \10609 , \10611 );
xor \U$10301 ( \10616 , \10412 , \10416 );
xor \U$10302 ( \10617 , \10616 , \10421 );
xor \U$10303 ( \10618 , \10428 , \10432 );
xor \U$10304 ( \10619 , \10618 , \10437 );
and \U$10305 ( \10620 , \10617 , \10619 );
xor \U$10306 ( \10621 , \10481 , \10485 );
xor \U$10307 ( \10622 , \10621 , \10490 );
and \U$10308 ( \10623 , \10619 , \10622 );
and \U$10309 ( \10624 , \10617 , \10622 );
or \U$10310 ( \10625 , \10620 , \10623 , \10624 );
xor \U$10311 ( \10626 , \10325 , \10329 );
xor \U$10312 ( \10627 , \10626 , \10334 );
xor \U$10313 ( \10628 , \10341 , \10345 );
xor \U$10314 ( \10629 , \10628 , \10348 );
and \U$10315 ( \10630 , \10627 , \10629 );
xor \U$10316 ( \10631 , \10445 , \10449 );
xor \U$10317 ( \10632 , \10631 , \10454 );
and \U$10318 ( \10633 , \10629 , \10632 );
and \U$10319 ( \10634 , \10627 , \10632 );
or \U$10320 ( \10635 , \10630 , \10633 , \10634 );
and \U$10321 ( \10636 , \10625 , \10635 );
and \U$10322 ( \10637 , \7703 , \692 );
and \U$10323 ( \10638 , \7177 , \690 );
nor \U$10324 ( \10639 , \10637 , \10638 );
xnor \U$10325 ( \10640 , \10639 , \649 );
and \U$10326 ( \10641 , \8373 , \579 );
and \U$10327 ( \10642 , \8127 , \577 );
nor \U$10328 ( \10643 , \10641 , \10642 );
xnor \U$10329 ( \10644 , \10643 , \530 );
and \U$10330 ( \10645 , \10640 , \10644 );
and \U$10331 ( \10646 , \8697 , \478 );
and \U$10332 ( \10647 , \8378 , \476 );
nor \U$10333 ( \10648 , \10646 , \10647 );
xnor \U$10334 ( \10649 , \10648 , \437 );
and \U$10335 ( \10650 , \10644 , \10649 );
and \U$10336 ( \10651 , \10640 , \10649 );
or \U$10337 ( \10652 , \10645 , \10650 , \10651 );
and \U$10338 ( \10653 , \9550 , \408 );
and \U$10339 ( \10654 , \8981 , \406 );
nor \U$10340 ( \10655 , \10653 , \10654 );
xnor \U$10341 ( \10656 , \10655 , \378 );
and \U$10342 ( \10657 , \10161 , \360 );
and \U$10343 ( \10658 , \9558 , \358 );
nor \U$10344 ( \10659 , \10657 , \10658 );
xnor \U$10345 ( \10660 , \10659 , \341 );
and \U$10346 ( \10661 , \10656 , \10660 );
and \U$10347 ( \10662 , \10347 , \323 );
and \U$10348 ( \10663 , \10166 , \321 );
nor \U$10349 ( \10664 , \10662 , \10663 );
xnor \U$10350 ( \10665 , \10664 , \328 );
and \U$10351 ( \10666 , \10660 , \10665 );
and \U$10352 ( \10667 , \10656 , \10665 );
or \U$10353 ( \10668 , \10661 , \10666 , \10667 );
or \U$10354 ( \10669 , \10652 , \10668 );
and \U$10355 ( \10670 , \10635 , \10669 );
and \U$10356 ( \10671 , \10625 , \10669 );
or \U$10357 ( \10672 , \10636 , \10670 , \10671 );
and \U$10358 ( \10673 , \4771 , \1826 );
and \U$10359 ( \10674 , \4469 , \1824 );
nor \U$10360 ( \10675 , \10673 , \10674 );
xnor \U$10361 ( \10676 , \10675 , \1670 );
and \U$10362 ( \10677 , \5248 , \1554 );
and \U$10363 ( \10678 , \4779 , \1552 );
nor \U$10364 ( \10679 , \10677 , \10678 );
xnor \U$10365 ( \10680 , \10679 , \1441 );
and \U$10366 ( \10681 , \10676 , \10680 );
and \U$10367 ( \10682 , \5517 , \1360 );
and \U$10368 ( \10683 , \5253 , \1358 );
nor \U$10369 ( \10684 , \10682 , \10683 );
xnor \U$10370 ( \10685 , \10684 , \1224 );
and \U$10371 ( \10686 , \10680 , \10685 );
and \U$10372 ( \10687 , \10676 , \10685 );
or \U$10373 ( \10688 , \10681 , \10686 , \10687 );
and \U$10374 ( \10689 , \6148 , \1160 );
and \U$10375 ( \10690 , \5776 , \1158 );
nor \U$10376 ( \10691 , \10689 , \10690 );
xnor \U$10377 ( \10692 , \10691 , \1082 );
and \U$10378 ( \10693 , \6500 , \996 );
and \U$10379 ( \10694 , \6157 , \994 );
nor \U$10380 ( \10695 , \10693 , \10694 );
xnor \U$10381 ( \10696 , \10695 , \902 );
and \U$10382 ( \10697 , \10692 , \10696 );
and \U$10383 ( \10698 , \7005 , \826 );
and \U$10384 ( \10699 , \6702 , \824 );
nor \U$10385 ( \10700 , \10698 , \10699 );
xnor \U$10386 ( \10701 , \10700 , \754 );
and \U$10387 ( \10702 , \10696 , \10701 );
and \U$10388 ( \10703 , \10692 , \10701 );
or \U$10389 ( \10704 , \10697 , \10702 , \10703 );
and \U$10390 ( \10705 , \10688 , \10704 );
and \U$10391 ( \10706 , \3681 , \2596 );
and \U$10392 ( \10707 , \3264 , \2594 );
nor \U$10393 ( \10708 , \10706 , \10707 );
xnor \U$10394 ( \10709 , \10708 , \2454 );
and \U$10395 ( \10710 , \4011 , \2300 );
and \U$10396 ( \10711 , \3889 , \2298 );
nor \U$10397 ( \10712 , \10710 , \10711 );
xnor \U$10398 ( \10713 , \10712 , \2163 );
and \U$10399 ( \10714 , \10709 , \10713 );
and \U$10400 ( \10715 , \4272 , \2094 );
and \U$10401 ( \10716 , \4016 , \2092 );
nor \U$10402 ( \10717 , \10715 , \10716 );
xnor \U$10403 ( \10718 , \10717 , \1942 );
and \U$10404 ( \10719 , \10713 , \10718 );
and \U$10405 ( \10720 , \10709 , \10718 );
or \U$10406 ( \10721 , \10714 , \10719 , \10720 );
and \U$10407 ( \10722 , \10704 , \10721 );
and \U$10408 ( \10723 , \10688 , \10721 );
or \U$10409 ( \10724 , \10705 , \10722 , \10723 );
and \U$10410 ( \10725 , \1791 , \4806 );
and \U$10411 ( \10726 , \1615 , \4804 );
nor \U$10412 ( \10727 , \10725 , \10726 );
xnor \U$10413 ( \10728 , \10727 , \4574 );
and \U$10414 ( \10729 , \2042 , \4355 );
and \U$10415 ( \10730 , \1799 , \4353 );
nor \U$10416 ( \10731 , \10729 , \10730 );
xnor \U$10417 ( \10732 , \10731 , \4212 );
and \U$10418 ( \10733 , \10728 , \10732 );
and \U$10419 ( \10734 , \2233 , \4032 );
and \U$10420 ( \10735 , \2047 , \4030 );
nor \U$10421 ( \10736 , \10734 , \10735 );
xnor \U$10422 ( \10737 , \10736 , \3786 );
and \U$10423 ( \10738 , \10732 , \10737 );
and \U$10424 ( \10739 , \10728 , \10737 );
or \U$10425 ( \10740 , \10733 , \10738 , \10739 );
and \U$10426 ( \10741 , \2641 , \3637 );
and \U$10427 ( \10742 , \2377 , \3635 );
nor \U$10428 ( \10743 , \10741 , \10742 );
xnor \U$10429 ( \10744 , \10743 , \3450 );
and \U$10430 ( \10745 , \2840 , \3324 );
and \U$10431 ( \10746 , \2666 , \3322 );
nor \U$10432 ( \10747 , \10745 , \10746 );
xnor \U$10433 ( \10748 , \10747 , \3119 );
and \U$10434 ( \10749 , \10744 , \10748 );
and \U$10435 ( \10750 , \3145 , \2918 );
and \U$10436 ( \10751 , \3007 , \2916 );
nor \U$10437 ( \10752 , \10750 , \10751 );
xnor \U$10438 ( \10753 , \10752 , \2769 );
and \U$10439 ( \10754 , \10748 , \10753 );
and \U$10440 ( \10755 , \10744 , \10753 );
or \U$10441 ( \10756 , \10749 , \10754 , \10755 );
and \U$10442 ( \10757 , \10740 , \10756 );
and \U$10443 ( \10758 , \1186 , \6235 );
and \U$10444 ( \10759 , \988 , \6233 );
nor \U$10445 ( \10760 , \10758 , \10759 );
xnor \U$10446 ( \10761 , \10760 , \5895 );
and \U$10447 ( \10762 , \1379 , \5646 );
and \U$10448 ( \10763 , \1274 , \5644 );
nor \U$10449 ( \10764 , \10762 , \10763 );
xnor \U$10450 ( \10765 , \10764 , \5405 );
and \U$10451 ( \10766 , \10761 , \10765 );
and \U$10452 ( \10767 , \1500 , \5180 );
and \U$10453 ( \10768 , \1384 , \5178 );
nor \U$10454 ( \10769 , \10767 , \10768 );
xnor \U$10455 ( \10770 , \10769 , \4992 );
and \U$10456 ( \10771 , \10765 , \10770 );
and \U$10457 ( \10772 , \10761 , \10770 );
or \U$10458 ( \10773 , \10766 , \10771 , \10772 );
and \U$10459 ( \10774 , \10756 , \10773 );
and \U$10460 ( \10775 , \10740 , \10773 );
or \U$10461 ( \10776 , \10757 , \10774 , \10775 );
and \U$10462 ( \10777 , \10724 , \10776 );
and \U$10463 ( \10778 , \417 , \9433 );
and \U$10464 ( \10779 , \369 , \9431 );
nor \U$10465 ( \10780 , \10778 , \10779 );
xnor \U$10466 ( \10781 , \10780 , \9123 );
and \U$10467 ( \10782 , \494 , \8896 );
and \U$10468 ( \10783 , \425 , \8894 );
nor \U$10469 ( \10784 , \10782 , \10783 );
xnor \U$10470 ( \10785 , \10784 , \8525 );
and \U$10471 ( \10786 , \10781 , \10785 );
and \U$10472 ( \10787 , \553 , \8334 );
and \U$10473 ( \10788 , \499 , \8332 );
nor \U$10474 ( \10789 , \10787 , \10788 );
xnor \U$10475 ( \10790 , \10789 , \8016 );
and \U$10476 ( \10791 , \10785 , \10790 );
and \U$10477 ( \10792 , \10781 , \10790 );
or \U$10478 ( \10793 , \10786 , \10791 , \10792 );
and \U$10479 ( \10794 , \681 , \7767 );
and \U$10480 ( \10795 , \604 , \7765 );
nor \U$10481 ( \10796 , \10794 , \10795 );
xnor \U$10482 ( \10797 , \10796 , \7518 );
and \U$10483 ( \10798 , \789 , \7238 );
and \U$10484 ( \10799 , \709 , \7236 );
nor \U$10485 ( \10800 , \10798 , \10799 );
xnor \U$10486 ( \10801 , \10800 , \6978 );
and \U$10487 ( \10802 , \10797 , \10801 );
and \U$10488 ( \10803 , \925 , \6744 );
and \U$10489 ( \10804 , \863 , \6742 );
nor \U$10490 ( \10805 , \10803 , \10804 );
xnor \U$10491 ( \10806 , \10805 , \6429 );
and \U$10492 ( \10807 , \10801 , \10806 );
and \U$10493 ( \10808 , \10797 , \10806 );
or \U$10494 ( \10809 , \10802 , \10807 , \10808 );
and \U$10495 ( \10810 , \10793 , \10809 );
buf \U$10496 ( \10811 , RIc0c79c8_65);
xor \U$10497 ( \10812 , \9759 , \10811 );
not \U$10498 ( \10813 , \10811 );
and \U$10499 ( \10814 , \10812 , \10813 );
and \U$10500 ( \10815 , \316 , \10814 );
not \U$10501 ( \10816 , \10815 );
xnor \U$10502 ( \10817 , \10816 , \9759 );
and \U$10503 ( \10818 , \348 , \10001 );
and \U$10504 ( \10819 , \330 , \9999 );
nor \U$10505 ( \10820 , \10818 , \10819 );
xnor \U$10506 ( \10821 , \10820 , \9762 );
and \U$10507 ( \10822 , \10817 , \10821 );
and \U$10508 ( \10823 , \10809 , \10822 );
and \U$10509 ( \10824 , \10793 , \10822 );
or \U$10510 ( \10825 , \10810 , \10823 , \10824 );
and \U$10511 ( \10826 , \10776 , \10825 );
and \U$10512 ( \10827 , \10724 , \10825 );
or \U$10513 ( \10828 , \10777 , \10826 , \10827 );
and \U$10514 ( \10829 , \10672 , \10828 );
xor \U$10515 ( \10830 , \10465 , \10469 );
xor \U$10516 ( \10831 , \10830 , \10474 );
xor \U$10517 ( \10832 , \10393 , \10397 );
xor \U$10518 ( \10833 , \10832 , \10402 );
and \U$10519 ( \10834 , \10831 , \10833 );
xor \U$10520 ( \10835 , \10498 , \10502 );
xor \U$10521 ( \10836 , \10835 , \10507 );
and \U$10522 ( \10837 , \10833 , \10836 );
and \U$10523 ( \10838 , \10831 , \10836 );
or \U$10524 ( \10839 , \10834 , \10837 , \10838 );
xor \U$10525 ( \10840 , \10360 , \10364 );
xor \U$10526 ( \10841 , \10840 , \10369 );
xor \U$10527 ( \10842 , \10376 , \10380 );
xor \U$10528 ( \10843 , \10842 , \10385 );
and \U$10529 ( \10844 , \10841 , \10843 );
and \U$10530 ( \10845 , \10839 , \10844 );
xor \U$10531 ( \10846 , \10004 , \10008 );
xor \U$10532 ( \10847 , \10846 , \10013 );
and \U$10533 ( \10848 , \10844 , \10847 );
and \U$10534 ( \10849 , \10839 , \10847 );
or \U$10535 ( \10850 , \10845 , \10848 , \10849 );
and \U$10536 ( \10851 , \10828 , \10850 );
and \U$10537 ( \10852 , \10672 , \10850 );
or \U$10538 ( \10853 , \10829 , \10851 , \10852 );
xor \U$10539 ( \10854 , \10519 , \10521 );
xor \U$10540 ( \10855 , \10854 , \10524 );
xor \U$10541 ( \10856 , \10302 , \10304 );
xor \U$10542 ( \10857 , \10856 , \10307 );
and \U$10543 ( \10858 , \10855 , \10857 );
xor \U$10544 ( \10859 , \10312 , \10314 );
xor \U$10545 ( \10860 , \10859 , \10317 );
and \U$10546 ( \10861 , \10857 , \10860 );
and \U$10547 ( \10862 , \10855 , \10860 );
or \U$10548 ( \10863 , \10858 , \10861 , \10862 );
xor \U$10549 ( \10864 , \10424 , \10440 );
xor \U$10550 ( \10865 , \10864 , \10457 );
xor \U$10551 ( \10866 , \10477 , \10493 );
xor \U$10552 ( \10867 , \10866 , \10510 );
and \U$10553 ( \10868 , \10865 , \10867 );
xor \U$10554 ( \10869 , \10337 , \10351 );
xor \U$10555 ( \10870 , \10869 , \10353 );
and \U$10556 ( \10871 , \10867 , \10870 );
and \U$10557 ( \10872 , \10865 , \10870 );
or \U$10558 ( \10873 , \10868 , \10871 , \10872 );
and \U$10559 ( \10874 , \10863 , \10873 );
xor \U$10560 ( \10875 , \10539 , \10541 );
xor \U$10561 ( \10876 , \10875 , \10544 );
and \U$10562 ( \10877 , \10873 , \10876 );
and \U$10563 ( \10878 , \10863 , \10876 );
or \U$10564 ( \10879 , \10874 , \10877 , \10878 );
and \U$10565 ( \10880 , \10853 , \10879 );
xor \U$10566 ( \10881 , \10310 , \10320 );
xor \U$10567 ( \10882 , \10881 , \10356 );
xor \U$10568 ( \10883 , \10549 , \10551 );
xor \U$10569 ( \10884 , \10883 , \10554 );
and \U$10570 ( \10885 , \10882 , \10884 );
xor \U$10571 ( \10886 , \10527 , \10529 );
xor \U$10572 ( \10887 , \10886 , \10531 );
and \U$10573 ( \10888 , \10884 , \10887 );
and \U$10574 ( \10889 , \10882 , \10887 );
or \U$10575 ( \10890 , \10885 , \10888 , \10889 );
and \U$10576 ( \10891 , \10879 , \10890 );
and \U$10577 ( \10892 , \10853 , \10890 );
or \U$10578 ( \10893 , \10880 , \10891 , \10892 );
xor \U$10579 ( \10894 , \10036 , \10088 );
xor \U$10580 ( \10895 , \10894 , \10141 );
xor \U$10581 ( \10896 , \10547 , \10557 );
xor \U$10582 ( \10897 , \10896 , \10560 );
and \U$10583 ( \10898 , \10895 , \10897 );
xor \U$10584 ( \10899 , \10566 , \10568 );
xor \U$10585 ( \10900 , \10899 , \10571 );
and \U$10586 ( \10901 , \10897 , \10900 );
and \U$10587 ( \10902 , \10895 , \10900 );
or \U$10588 ( \10903 , \10898 , \10901 , \10902 );
and \U$10589 ( \10904 , \10893 , \10903 );
xor \U$10590 ( \10905 , \10144 , \10199 );
xor \U$10591 ( \10906 , \10905 , \10221 );
and \U$10592 ( \10907 , \10903 , \10906 );
and \U$10593 ( \10908 , \10893 , \10906 );
or \U$10594 ( \10909 , \10904 , \10907 , \10908 );
xor \U$10595 ( \10910 , \10577 , \10587 );
xor \U$10596 ( \10911 , \10910 , \10590 );
and \U$10597 ( \10912 , \10909 , \10911 );
xor \U$10598 ( \10913 , \10595 , \10597 );
xor \U$10599 ( \10914 , \10913 , \10600 );
and \U$10600 ( \10915 , \10911 , \10914 );
and \U$10601 ( \10916 , \10909 , \10914 );
or \U$10602 ( \10917 , \10912 , \10915 , \10916 );
xor \U$10603 ( \10918 , \10593 , \10603 );
xor \U$10604 ( \10919 , \10918 , \10606 );
and \U$10605 ( \10920 , \10917 , \10919 );
xor \U$10606 ( \10921 , \10264 , \10274 );
xor \U$10607 ( \10922 , \10921 , \10277 );
and \U$10608 ( \10923 , \10919 , \10922 );
and \U$10609 ( \10924 , \10917 , \10922 );
or \U$10610 ( \10925 , \10920 , \10923 , \10924 );
and \U$10611 ( \10926 , \10615 , \10925 );
xor \U$10612 ( \10927 , \10615 , \10925 );
xor \U$10613 ( \10928 , \10917 , \10919 );
xor \U$10614 ( \10929 , \10928 , \10922 );
xor \U$10615 ( \10930 , \10676 , \10680 );
xor \U$10616 ( \10931 , \10930 , \10685 );
xor \U$10617 ( \10932 , \10640 , \10644 );
xor \U$10618 ( \10933 , \10932 , \10649 );
and \U$10619 ( \10934 , \10931 , \10933 );
xor \U$10620 ( \10935 , \10692 , \10696 );
xor \U$10621 ( \10936 , \10935 , \10701 );
and \U$10622 ( \10937 , \10933 , \10936 );
and \U$10623 ( \10938 , \10931 , \10936 );
or \U$10624 ( \10939 , \10934 , \10937 , \10938 );
xor \U$10625 ( \10940 , \10728 , \10732 );
xor \U$10626 ( \10941 , \10940 , \10737 );
xor \U$10627 ( \10942 , \10744 , \10748 );
xor \U$10628 ( \10943 , \10942 , \10753 );
and \U$10629 ( \10944 , \10941 , \10943 );
xor \U$10630 ( \10945 , \10709 , \10713 );
xor \U$10631 ( \10946 , \10945 , \10718 );
and \U$10632 ( \10947 , \10943 , \10946 );
and \U$10633 ( \10948 , \10941 , \10946 );
or \U$10634 ( \10949 , \10944 , \10947 , \10948 );
and \U$10635 ( \10950 , \10939 , \10949 );
and \U$10636 ( \10951 , \8378 , \579 );
and \U$10637 ( \10952 , \8373 , \577 );
nor \U$10638 ( \10953 , \10951 , \10952 );
xnor \U$10639 ( \10954 , \10953 , \530 );
and \U$10640 ( \10955 , \8981 , \478 );
and \U$10641 ( \10956 , \8697 , \476 );
nor \U$10642 ( \10957 , \10955 , \10956 );
xnor \U$10643 ( \10958 , \10957 , \437 );
and \U$10644 ( \10959 , \10954 , \10958 );
and \U$10645 ( \10960 , \9558 , \408 );
and \U$10646 ( \10961 , \9550 , \406 );
nor \U$10647 ( \10962 , \10960 , \10961 );
xnor \U$10648 ( \10963 , \10962 , \378 );
and \U$10649 ( \10964 , \10958 , \10963 );
and \U$10650 ( \10965 , \10954 , \10963 );
or \U$10651 ( \10966 , \10959 , \10964 , \10965 );
buf \U$10652 ( \10967 , RIc340620_129);
nand \U$10653 ( \10968 , \10967 , \317 );
not \U$10654 ( \10969 , \10968 );
and \U$10655 ( \10970 , \10966 , \10969 );
xor \U$10656 ( \10971 , \10656 , \10660 );
xor \U$10657 ( \10972 , \10971 , \10665 );
and \U$10658 ( \10973 , \10969 , \10972 );
and \U$10659 ( \10974 , \10966 , \10972 );
or \U$10660 ( \10975 , \10970 , \10973 , \10974 );
and \U$10661 ( \10976 , \10949 , \10975 );
and \U$10662 ( \10977 , \10939 , \10975 );
or \U$10663 ( \10978 , \10950 , \10976 , \10977 );
and \U$10664 ( \10979 , \2047 , \4355 );
and \U$10665 ( \10980 , \2042 , \4353 );
nor \U$10666 ( \10981 , \10979 , \10980 );
xnor \U$10667 ( \10982 , \10981 , \4212 );
and \U$10668 ( \10983 , \2377 , \4032 );
and \U$10669 ( \10984 , \2233 , \4030 );
nor \U$10670 ( \10985 , \10983 , \10984 );
xnor \U$10671 ( \10986 , \10985 , \3786 );
and \U$10672 ( \10987 , \10982 , \10986 );
and \U$10673 ( \10988 , \2666 , \3637 );
and \U$10674 ( \10989 , \2641 , \3635 );
nor \U$10675 ( \10990 , \10988 , \10989 );
xnor \U$10676 ( \10991 , \10990 , \3450 );
and \U$10677 ( \10992 , \10986 , \10991 );
and \U$10678 ( \10993 , \10982 , \10991 );
or \U$10679 ( \10994 , \10987 , \10992 , \10993 );
and \U$10680 ( \10995 , \1384 , \5646 );
and \U$10681 ( \10996 , \1379 , \5644 );
nor \U$10682 ( \10997 , \10995 , \10996 );
xnor \U$10683 ( \10998 , \10997 , \5405 );
and \U$10684 ( \10999 , \1615 , \5180 );
and \U$10685 ( \11000 , \1500 , \5178 );
nor \U$10686 ( \11001 , \10999 , \11000 );
xnor \U$10687 ( \11002 , \11001 , \4992 );
and \U$10688 ( \11003 , \10998 , \11002 );
and \U$10689 ( \11004 , \1799 , \4806 );
and \U$10690 ( \11005 , \1791 , \4804 );
nor \U$10691 ( \11006 , \11004 , \11005 );
xnor \U$10692 ( \11007 , \11006 , \4574 );
and \U$10693 ( \11008 , \11002 , \11007 );
and \U$10694 ( \11009 , \10998 , \11007 );
or \U$10695 ( \11010 , \11003 , \11008 , \11009 );
and \U$10696 ( \11011 , \10994 , \11010 );
and \U$10697 ( \11012 , \3007 , \3324 );
and \U$10698 ( \11013 , \2840 , \3322 );
nor \U$10699 ( \11014 , \11012 , \11013 );
xnor \U$10700 ( \11015 , \11014 , \3119 );
and \U$10701 ( \11016 , \3264 , \2918 );
and \U$10702 ( \11017 , \3145 , \2916 );
nor \U$10703 ( \11018 , \11016 , \11017 );
xnor \U$10704 ( \11019 , \11018 , \2769 );
and \U$10705 ( \11020 , \11015 , \11019 );
and \U$10706 ( \11021 , \3889 , \2596 );
and \U$10707 ( \11022 , \3681 , \2594 );
nor \U$10708 ( \11023 , \11021 , \11022 );
xnor \U$10709 ( \11024 , \11023 , \2454 );
and \U$10710 ( \11025 , \11019 , \11024 );
and \U$10711 ( \11026 , \11015 , \11024 );
or \U$10712 ( \11027 , \11020 , \11025 , \11026 );
and \U$10713 ( \11028 , \11010 , \11027 );
and \U$10714 ( \11029 , \10994 , \11027 );
or \U$10715 ( \11030 , \11011 , \11028 , \11029 );
and \U$10716 ( \11031 , \863 , \7238 );
and \U$10717 ( \11032 , \789 , \7236 );
nor \U$10718 ( \11033 , \11031 , \11032 );
xnor \U$10719 ( \11034 , \11033 , \6978 );
and \U$10720 ( \11035 , \988 , \6744 );
and \U$10721 ( \11036 , \925 , \6742 );
nor \U$10722 ( \11037 , \11035 , \11036 );
xnor \U$10723 ( \11038 , \11037 , \6429 );
and \U$10724 ( \11039 , \11034 , \11038 );
and \U$10725 ( \11040 , \1274 , \6235 );
and \U$10726 ( \11041 , \1186 , \6233 );
nor \U$10727 ( \11042 , \11040 , \11041 );
xnor \U$10728 ( \11043 , \11042 , \5895 );
and \U$10729 ( \11044 , \11038 , \11043 );
and \U$10730 ( \11045 , \11034 , \11043 );
or \U$10731 ( \11046 , \11039 , \11044 , \11045 );
and \U$10732 ( \11047 , \499 , \8896 );
and \U$10733 ( \11048 , \494 , \8894 );
nor \U$10734 ( \11049 , \11047 , \11048 );
xnor \U$10735 ( \11050 , \11049 , \8525 );
and \U$10736 ( \11051 , \604 , \8334 );
and \U$10737 ( \11052 , \553 , \8332 );
nor \U$10738 ( \11053 , \11051 , \11052 );
xnor \U$10739 ( \11054 , \11053 , \8016 );
and \U$10740 ( \11055 , \11050 , \11054 );
and \U$10741 ( \11056 , \709 , \7767 );
and \U$10742 ( \11057 , \681 , \7765 );
nor \U$10743 ( \11058 , \11056 , \11057 );
xnor \U$10744 ( \11059 , \11058 , \7518 );
and \U$10745 ( \11060 , \11054 , \11059 );
and \U$10746 ( \11061 , \11050 , \11059 );
or \U$10747 ( \11062 , \11055 , \11060 , \11061 );
and \U$10748 ( \11063 , \11046 , \11062 );
and \U$10749 ( \11064 , \330 , \10814 );
and \U$10750 ( \11065 , \316 , \10811 );
nor \U$10751 ( \11066 , \11064 , \11065 );
xnor \U$10752 ( \11067 , \11066 , \9759 );
and \U$10753 ( \11068 , \369 , \10001 );
and \U$10754 ( \11069 , \348 , \9999 );
nor \U$10755 ( \11070 , \11068 , \11069 );
xnor \U$10756 ( \11071 , \11070 , \9762 );
and \U$10757 ( \11072 , \11067 , \11071 );
and \U$10758 ( \11073 , \425 , \9433 );
and \U$10759 ( \11074 , \417 , \9431 );
nor \U$10760 ( \11075 , \11073 , \11074 );
xnor \U$10761 ( \11076 , \11075 , \9123 );
and \U$10762 ( \11077 , \11071 , \11076 );
and \U$10763 ( \11078 , \11067 , \11076 );
or \U$10764 ( \11079 , \11072 , \11077 , \11078 );
and \U$10765 ( \11080 , \11062 , \11079 );
and \U$10766 ( \11081 , \11046 , \11079 );
or \U$10767 ( \11082 , \11063 , \11080 , \11081 );
and \U$10768 ( \11083 , \11030 , \11082 );
and \U$10769 ( \11084 , \5253 , \1554 );
and \U$10770 ( \11085 , \5248 , \1552 );
nor \U$10771 ( \11086 , \11084 , \11085 );
xnor \U$10772 ( \11087 , \11086 , \1441 );
and \U$10773 ( \11088 , \5776 , \1360 );
and \U$10774 ( \11089 , \5517 , \1358 );
nor \U$10775 ( \11090 , \11088 , \11089 );
xnor \U$10776 ( \11091 , \11090 , \1224 );
and \U$10777 ( \11092 , \11087 , \11091 );
and \U$10778 ( \11093 , \6157 , \1160 );
and \U$10779 ( \11094 , \6148 , \1158 );
nor \U$10780 ( \11095 , \11093 , \11094 );
xnor \U$10781 ( \11096 , \11095 , \1082 );
and \U$10782 ( \11097 , \11091 , \11096 );
and \U$10783 ( \11098 , \11087 , \11096 );
or \U$10784 ( \11099 , \11092 , \11097 , \11098 );
and \U$10785 ( \11100 , \4016 , \2300 );
and \U$10786 ( \11101 , \4011 , \2298 );
nor \U$10787 ( \11102 , \11100 , \11101 );
xnor \U$10788 ( \11103 , \11102 , \2163 );
and \U$10789 ( \11104 , \4469 , \2094 );
and \U$10790 ( \11105 , \4272 , \2092 );
nor \U$10791 ( \11106 , \11104 , \11105 );
xnor \U$10792 ( \11107 , \11106 , \1942 );
and \U$10793 ( \11108 , \11103 , \11107 );
and \U$10794 ( \11109 , \4779 , \1826 );
and \U$10795 ( \11110 , \4771 , \1824 );
nor \U$10796 ( \11111 , \11109 , \11110 );
xnor \U$10797 ( \11112 , \11111 , \1670 );
and \U$10798 ( \11113 , \11107 , \11112 );
and \U$10799 ( \11114 , \11103 , \11112 );
or \U$10800 ( \11115 , \11108 , \11113 , \11114 );
and \U$10801 ( \11116 , \11099 , \11115 );
and \U$10802 ( \11117 , \6702 , \996 );
and \U$10803 ( \11118 , \6500 , \994 );
nor \U$10804 ( \11119 , \11117 , \11118 );
xnor \U$10805 ( \11120 , \11119 , \902 );
and \U$10806 ( \11121 , \7177 , \826 );
and \U$10807 ( \11122 , \7005 , \824 );
nor \U$10808 ( \11123 , \11121 , \11122 );
xnor \U$10809 ( \11124 , \11123 , \754 );
and \U$10810 ( \11125 , \11120 , \11124 );
and \U$10811 ( \11126 , \8127 , \692 );
and \U$10812 ( \11127 , \7703 , \690 );
nor \U$10813 ( \11128 , \11126 , \11127 );
xnor \U$10814 ( \11129 , \11128 , \649 );
and \U$10815 ( \11130 , \11124 , \11129 );
and \U$10816 ( \11131 , \11120 , \11129 );
or \U$10817 ( \11132 , \11125 , \11130 , \11131 );
and \U$10818 ( \11133 , \11115 , \11132 );
and \U$10819 ( \11134 , \11099 , \11132 );
or \U$10820 ( \11135 , \11116 , \11133 , \11134 );
and \U$10821 ( \11136 , \11082 , \11135 );
and \U$10822 ( \11137 , \11030 , \11135 );
or \U$10823 ( \11138 , \11083 , \11136 , \11137 );
and \U$10824 ( \11139 , \10978 , \11138 );
xor \U$10825 ( \11140 , \10781 , \10785 );
xor \U$10826 ( \11141 , \11140 , \10790 );
xor \U$10827 ( \11142 , \10797 , \10801 );
xor \U$10828 ( \11143 , \11142 , \10806 );
and \U$10829 ( \11144 , \11141 , \11143 );
xor \U$10830 ( \11145 , \10761 , \10765 );
xor \U$10831 ( \11146 , \11145 , \10770 );
and \U$10832 ( \11147 , \11143 , \11146 );
and \U$10833 ( \11148 , \11141 , \11146 );
or \U$10834 ( \11149 , \11144 , \11147 , \11148 );
xor \U$10835 ( \11150 , \10831 , \10833 );
xor \U$10836 ( \11151 , \11150 , \10836 );
and \U$10837 ( \11152 , \11149 , \11151 );
xor \U$10838 ( \11153 , \10841 , \10843 );
and \U$10839 ( \11154 , \11151 , \11153 );
and \U$10840 ( \11155 , \11149 , \11153 );
or \U$10841 ( \11156 , \11152 , \11154 , \11155 );
and \U$10842 ( \11157 , \11138 , \11156 );
and \U$10843 ( \11158 , \10978 , \11156 );
or \U$10844 ( \11159 , \11139 , \11157 , \11158 );
xor \U$10845 ( \11160 , \10688 , \10704 );
xor \U$10846 ( \11161 , \11160 , \10721 );
xor \U$10847 ( \11162 , \10740 , \10756 );
xor \U$10848 ( \11163 , \11162 , \10773 );
and \U$10849 ( \11164 , \11161 , \11163 );
xor \U$10850 ( \11165 , \10793 , \10809 );
xor \U$10851 ( \11166 , \11165 , \10822 );
and \U$10852 ( \11167 , \11163 , \11166 );
and \U$10853 ( \11168 , \11161 , \11166 );
or \U$10854 ( \11169 , \11164 , \11167 , \11168 );
xor \U$10855 ( \11170 , \10617 , \10619 );
xor \U$10856 ( \11171 , \11170 , \10622 );
xor \U$10857 ( \11172 , \10627 , \10629 );
xor \U$10858 ( \11173 , \11172 , \10632 );
and \U$10859 ( \11174 , \11171 , \11173 );
xnor \U$10860 ( \11175 , \10652 , \10668 );
and \U$10861 ( \11176 , \11173 , \11175 );
and \U$10862 ( \11177 , \11171 , \11175 );
or \U$10863 ( \11178 , \11174 , \11176 , \11177 );
and \U$10864 ( \11179 , \11169 , \11178 );
xor \U$10865 ( \11180 , \10372 , \10388 );
xor \U$10866 ( \11181 , \11180 , \10405 );
and \U$10867 ( \11182 , \11178 , \11181 );
and \U$10868 ( \11183 , \11169 , \11181 );
or \U$10869 ( \11184 , \11179 , \11182 , \11183 );
and \U$10870 ( \11185 , \11159 , \11184 );
xor \U$10871 ( \11186 , \10839 , \10844 );
xor \U$10872 ( \11187 , \11186 , \10847 );
xor \U$10873 ( \11188 , \10855 , \10857 );
xor \U$10874 ( \11189 , \11188 , \10860 );
and \U$10875 ( \11190 , \11187 , \11189 );
xor \U$10876 ( \11191 , \10865 , \10867 );
xor \U$10877 ( \11192 , \11191 , \10870 );
and \U$10878 ( \11193 , \11189 , \11192 );
and \U$10879 ( \11194 , \11187 , \11192 );
or \U$10880 ( \11195 , \11190 , \11193 , \11194 );
and \U$10881 ( \11196 , \11184 , \11195 );
and \U$10882 ( \11197 , \11159 , \11195 );
or \U$10883 ( \11198 , \11185 , \11196 , \11197 );
xor \U$10884 ( \11199 , \10408 , \10460 );
xor \U$10885 ( \11200 , \11199 , \10513 );
xor \U$10886 ( \11201 , \10863 , \10873 );
xor \U$10887 ( \11202 , \11201 , \10876 );
and \U$10888 ( \11203 , \11200 , \11202 );
xor \U$10889 ( \11204 , \10882 , \10884 );
xor \U$10890 ( \11205 , \11204 , \10887 );
and \U$10891 ( \11206 , \11202 , \11205 );
and \U$10892 ( \11207 , \11200 , \11205 );
or \U$10893 ( \11208 , \11203 , \11206 , \11207 );
and \U$10894 ( \11209 , \11198 , \11208 );
xor \U$10895 ( \11210 , \10359 , \10516 );
xor \U$10896 ( \11211 , \11210 , \10534 );
and \U$10897 ( \11212 , \11208 , \11211 );
and \U$10898 ( \11213 , \11198 , \11211 );
or \U$10899 ( \11214 , \11209 , \11212 , \11213 );
xor \U$10900 ( \11215 , \10853 , \10879 );
xor \U$10901 ( \11216 , \11215 , \10890 );
xor \U$10902 ( \11217 , \10895 , \10897 );
xor \U$10903 ( \11218 , \11217 , \10900 );
and \U$10904 ( \11219 , \11216 , \11218 );
and \U$10905 ( \11220 , \11214 , \11219 );
xor \U$10906 ( \11221 , \10579 , \10581 );
xor \U$10907 ( \11222 , \11221 , \10584 );
and \U$10908 ( \11223 , \11219 , \11222 );
and \U$10909 ( \11224 , \11214 , \11222 );
or \U$10910 ( \11225 , \11220 , \11223 , \11224 );
xor \U$10911 ( \11226 , \10537 , \10563 );
xor \U$10912 ( \11227 , \11226 , \10574 );
xor \U$10913 ( \11228 , \10893 , \10903 );
xor \U$10914 ( \11229 , \11228 , \10906 );
and \U$10915 ( \11230 , \11227 , \11229 );
and \U$10916 ( \11231 , \11225 , \11230 );
xor \U$10917 ( \11232 , \10909 , \10911 );
xor \U$10918 ( \11233 , \11232 , \10914 );
and \U$10919 ( \11234 , \11230 , \11233 );
and \U$10920 ( \11235 , \11225 , \11233 );
or \U$10921 ( \11236 , \11231 , \11234 , \11235 );
and \U$10922 ( \11237 , \10929 , \11236 );
xor \U$10923 ( \11238 , \10929 , \11236 );
xor \U$10924 ( \11239 , \11225 , \11230 );
xor \U$10925 ( \11240 , \11239 , \11233 );
and \U$10926 ( \11241 , \10161 , \408 );
and \U$10927 ( \11242 , \9558 , \406 );
nor \U$10928 ( \11243 , \11241 , \11242 );
xnor \U$10929 ( \11244 , \11243 , \378 );
and \U$10930 ( \11245 , \10347 , \360 );
and \U$10931 ( \11246 , \10166 , \358 );
nor \U$10932 ( \11247 , \11245 , \11246 );
xnor \U$10933 ( \11248 , \11247 , \341 );
and \U$10934 ( \11249 , \11244 , \11248 );
nand \U$10935 ( \11250 , \10967 , \321 );
xnor \U$10936 ( \11251 , \11250 , \328 );
and \U$10937 ( \11252 , \11248 , \11251 );
and \U$10938 ( \11253 , \11244 , \11251 );
or \U$10939 ( \11254 , \11249 , \11252 , \11253 );
and \U$10940 ( \11255 , \8373 , \692 );
and \U$10941 ( \11256 , \8127 , \690 );
nor \U$10942 ( \11257 , \11255 , \11256 );
xnor \U$10943 ( \11258 , \11257 , \649 );
and \U$10944 ( \11259 , \8697 , \579 );
and \U$10945 ( \11260 , \8378 , \577 );
nor \U$10946 ( \11261 , \11259 , \11260 );
xnor \U$10947 ( \11262 , \11261 , \530 );
and \U$10948 ( \11263 , \11258 , \11262 );
and \U$10949 ( \11264 , \9550 , \478 );
and \U$10950 ( \11265 , \8981 , \476 );
nor \U$10951 ( \11266 , \11264 , \11265 );
xnor \U$10952 ( \11267 , \11266 , \437 );
and \U$10953 ( \11268 , \11262 , \11267 );
and \U$10954 ( \11269 , \11258 , \11267 );
or \U$10955 ( \11270 , \11263 , \11268 , \11269 );
and \U$10956 ( \11271 , \11254 , \11270 );
and \U$10957 ( \11272 , \10166 , \360 );
and \U$10958 ( \11273 , \10161 , \358 );
nor \U$10959 ( \11274 , \11272 , \11273 );
xnor \U$10960 ( \11275 , \11274 , \341 );
and \U$10961 ( \11276 , \11270 , \11275 );
and \U$10962 ( \11277 , \11254 , \11275 );
or \U$10963 ( \11278 , \11271 , \11276 , \11277 );
and \U$10964 ( \11279 , \10967 , \323 );
and \U$10965 ( \11280 , \10347 , \321 );
nor \U$10966 ( \11281 , \11279 , \11280 );
xnor \U$10967 ( \11282 , \11281 , \328 );
xor \U$10968 ( \11283 , \11120 , \11124 );
xor \U$10969 ( \11284 , \11283 , \11129 );
and \U$10970 ( \11285 , \11282 , \11284 );
xor \U$10971 ( \11286 , \10954 , \10958 );
xor \U$10972 ( \11287 , \11286 , \10963 );
and \U$10973 ( \11288 , \11284 , \11287 );
and \U$10974 ( \11289 , \11282 , \11287 );
or \U$10975 ( \11290 , \11285 , \11288 , \11289 );
and \U$10976 ( \11291 , \11278 , \11290 );
xor \U$10977 ( \11292 , \11087 , \11091 );
xor \U$10978 ( \11293 , \11292 , \11096 );
xor \U$10979 ( \11294 , \11103 , \11107 );
xor \U$10980 ( \11295 , \11294 , \11112 );
and \U$10981 ( \11296 , \11293 , \11295 );
xor \U$10982 ( \11297 , \11015 , \11019 );
xor \U$10983 ( \11298 , \11297 , \11024 );
and \U$10984 ( \11299 , \11295 , \11298 );
and \U$10985 ( \11300 , \11293 , \11298 );
or \U$10986 ( \11301 , \11296 , \11299 , \11300 );
and \U$10987 ( \11302 , \11290 , \11301 );
and \U$10988 ( \11303 , \11278 , \11301 );
or \U$10989 ( \11304 , \11291 , \11302 , \11303 );
and \U$10990 ( \11305 , \5248 , \1826 );
and \U$10991 ( \11306 , \4779 , \1824 );
nor \U$10992 ( \11307 , \11305 , \11306 );
xnor \U$10993 ( \11308 , \11307 , \1670 );
and \U$10994 ( \11309 , \5517 , \1554 );
and \U$10995 ( \11310 , \5253 , \1552 );
nor \U$10996 ( \11311 , \11309 , \11310 );
xnor \U$10997 ( \11312 , \11311 , \1441 );
and \U$10998 ( \11313 , \11308 , \11312 );
and \U$10999 ( \11314 , \6148 , \1360 );
and \U$11000 ( \11315 , \5776 , \1358 );
nor \U$11001 ( \11316 , \11314 , \11315 );
xnor \U$11002 ( \11317 , \11316 , \1224 );
and \U$11003 ( \11318 , \11312 , \11317 );
and \U$11004 ( \11319 , \11308 , \11317 );
or \U$11005 ( \11320 , \11313 , \11318 , \11319 );
and \U$11006 ( \11321 , \4011 , \2596 );
and \U$11007 ( \11322 , \3889 , \2594 );
nor \U$11008 ( \11323 , \11321 , \11322 );
xnor \U$11009 ( \11324 , \11323 , \2454 );
and \U$11010 ( \11325 , \4272 , \2300 );
and \U$11011 ( \11326 , \4016 , \2298 );
nor \U$11012 ( \11327 , \11325 , \11326 );
xnor \U$11013 ( \11328 , \11327 , \2163 );
and \U$11014 ( \11329 , \11324 , \11328 );
and \U$11015 ( \11330 , \4771 , \2094 );
and \U$11016 ( \11331 , \4469 , \2092 );
nor \U$11017 ( \11332 , \11330 , \11331 );
xnor \U$11018 ( \11333 , \11332 , \1942 );
and \U$11019 ( \11334 , \11328 , \11333 );
and \U$11020 ( \11335 , \11324 , \11333 );
or \U$11021 ( \11336 , \11329 , \11334 , \11335 );
and \U$11022 ( \11337 , \11320 , \11336 );
and \U$11023 ( \11338 , \6500 , \1160 );
and \U$11024 ( \11339 , \6157 , \1158 );
nor \U$11025 ( \11340 , \11338 , \11339 );
xnor \U$11026 ( \11341 , \11340 , \1082 );
and \U$11027 ( \11342 , \7005 , \996 );
and \U$11028 ( \11343 , \6702 , \994 );
nor \U$11029 ( \11344 , \11342 , \11343 );
xnor \U$11030 ( \11345 , \11344 , \902 );
and \U$11031 ( \11346 , \11341 , \11345 );
and \U$11032 ( \11347 , \7703 , \826 );
and \U$11033 ( \11348 , \7177 , \824 );
nor \U$11034 ( \11349 , \11347 , \11348 );
xnor \U$11035 ( \11350 , \11349 , \754 );
and \U$11036 ( \11351 , \11345 , \11350 );
and \U$11037 ( \11352 , \11341 , \11350 );
or \U$11038 ( \11353 , \11346 , \11351 , \11352 );
and \U$11039 ( \11354 , \11336 , \11353 );
and \U$11040 ( \11355 , \11320 , \11353 );
or \U$11041 ( \11356 , \11337 , \11354 , \11355 );
and \U$11042 ( \11357 , \789 , \7767 );
and \U$11043 ( \11358 , \709 , \7765 );
nor \U$11044 ( \11359 , \11357 , \11358 );
xnor \U$11045 ( \11360 , \11359 , \7518 );
and \U$11046 ( \11361 , \925 , \7238 );
and \U$11047 ( \11362 , \863 , \7236 );
nor \U$11048 ( \11363 , \11361 , \11362 );
xnor \U$11049 ( \11364 , \11363 , \6978 );
and \U$11050 ( \11365 , \11360 , \11364 );
and \U$11051 ( \11366 , \1186 , \6744 );
and \U$11052 ( \11367 , \988 , \6742 );
nor \U$11053 ( \11368 , \11366 , \11367 );
xnor \U$11054 ( \11369 , \11368 , \6429 );
and \U$11055 ( \11370 , \11364 , \11369 );
and \U$11056 ( \11371 , \11360 , \11369 );
or \U$11057 ( \11372 , \11365 , \11370 , \11371 );
and \U$11058 ( \11373 , \348 , \10814 );
and \U$11059 ( \11374 , \330 , \10811 );
nor \U$11060 ( \11375 , \11373 , \11374 );
xnor \U$11061 ( \11376 , \11375 , \9759 );
and \U$11062 ( \11377 , \417 , \10001 );
and \U$11063 ( \11378 , \369 , \9999 );
nor \U$11064 ( \11379 , \11377 , \11378 );
xnor \U$11065 ( \11380 , \11379 , \9762 );
and \U$11066 ( \11381 , \11376 , \11380 );
and \U$11067 ( \11382 , \11380 , \328 );
and \U$11068 ( \11383 , \11376 , \328 );
or \U$11069 ( \11384 , \11381 , \11382 , \11383 );
and \U$11070 ( \11385 , \11372 , \11384 );
and \U$11071 ( \11386 , \494 , \9433 );
and \U$11072 ( \11387 , \425 , \9431 );
nor \U$11073 ( \11388 , \11386 , \11387 );
xnor \U$11074 ( \11389 , \11388 , \9123 );
and \U$11075 ( \11390 , \553 , \8896 );
and \U$11076 ( \11391 , \499 , \8894 );
nor \U$11077 ( \11392 , \11390 , \11391 );
xnor \U$11078 ( \11393 , \11392 , \8525 );
and \U$11079 ( \11394 , \11389 , \11393 );
and \U$11080 ( \11395 , \681 , \8334 );
and \U$11081 ( \11396 , \604 , \8332 );
nor \U$11082 ( \11397 , \11395 , \11396 );
xnor \U$11083 ( \11398 , \11397 , \8016 );
and \U$11084 ( \11399 , \11393 , \11398 );
and \U$11085 ( \11400 , \11389 , \11398 );
or \U$11086 ( \11401 , \11394 , \11399 , \11400 );
and \U$11087 ( \11402 , \11384 , \11401 );
and \U$11088 ( \11403 , \11372 , \11401 );
or \U$11089 ( \11404 , \11385 , \11402 , \11403 );
and \U$11090 ( \11405 , \11356 , \11404 );
and \U$11091 ( \11406 , \2042 , \4806 );
and \U$11092 ( \11407 , \1799 , \4804 );
nor \U$11093 ( \11408 , \11406 , \11407 );
xnor \U$11094 ( \11409 , \11408 , \4574 );
and \U$11095 ( \11410 , \2233 , \4355 );
and \U$11096 ( \11411 , \2047 , \4353 );
nor \U$11097 ( \11412 , \11410 , \11411 );
xnor \U$11098 ( \11413 , \11412 , \4212 );
and \U$11099 ( \11414 , \11409 , \11413 );
and \U$11100 ( \11415 , \2641 , \4032 );
and \U$11101 ( \11416 , \2377 , \4030 );
nor \U$11102 ( \11417 , \11415 , \11416 );
xnor \U$11103 ( \11418 , \11417 , \3786 );
and \U$11104 ( \11419 , \11413 , \11418 );
and \U$11105 ( \11420 , \11409 , \11418 );
or \U$11106 ( \11421 , \11414 , \11419 , \11420 );
and \U$11107 ( \11422 , \1379 , \6235 );
and \U$11108 ( \11423 , \1274 , \6233 );
nor \U$11109 ( \11424 , \11422 , \11423 );
xnor \U$11110 ( \11425 , \11424 , \5895 );
and \U$11111 ( \11426 , \1500 , \5646 );
and \U$11112 ( \11427 , \1384 , \5644 );
nor \U$11113 ( \11428 , \11426 , \11427 );
xnor \U$11114 ( \11429 , \11428 , \5405 );
and \U$11115 ( \11430 , \11425 , \11429 );
and \U$11116 ( \11431 , \1791 , \5180 );
and \U$11117 ( \11432 , \1615 , \5178 );
nor \U$11118 ( \11433 , \11431 , \11432 );
xnor \U$11119 ( \11434 , \11433 , \4992 );
and \U$11120 ( \11435 , \11429 , \11434 );
and \U$11121 ( \11436 , \11425 , \11434 );
or \U$11122 ( \11437 , \11430 , \11435 , \11436 );
and \U$11123 ( \11438 , \11421 , \11437 );
and \U$11124 ( \11439 , \2840 , \3637 );
and \U$11125 ( \11440 , \2666 , \3635 );
nor \U$11126 ( \11441 , \11439 , \11440 );
xnor \U$11127 ( \11442 , \11441 , \3450 );
and \U$11128 ( \11443 , \3145 , \3324 );
and \U$11129 ( \11444 , \3007 , \3322 );
nor \U$11130 ( \11445 , \11443 , \11444 );
xnor \U$11131 ( \11446 , \11445 , \3119 );
and \U$11132 ( \11447 , \11442 , \11446 );
and \U$11133 ( \11448 , \3681 , \2918 );
and \U$11134 ( \11449 , \3264 , \2916 );
nor \U$11135 ( \11450 , \11448 , \11449 );
xnor \U$11136 ( \11451 , \11450 , \2769 );
and \U$11137 ( \11452 , \11446 , \11451 );
and \U$11138 ( \11453 , \11442 , \11451 );
or \U$11139 ( \11454 , \11447 , \11452 , \11453 );
and \U$11140 ( \11455 , \11437 , \11454 );
and \U$11141 ( \11456 , \11421 , \11454 );
or \U$11142 ( \11457 , \11438 , \11455 , \11456 );
and \U$11143 ( \11458 , \11404 , \11457 );
and \U$11144 ( \11459 , \11356 , \11457 );
or \U$11145 ( \11460 , \11405 , \11458 , \11459 );
and \U$11146 ( \11461 , \11304 , \11460 );
xor \U$11147 ( \11462 , \10982 , \10986 );
xor \U$11148 ( \11463 , \11462 , \10991 );
xor \U$11149 ( \11464 , \10998 , \11002 );
xor \U$11150 ( \11465 , \11464 , \11007 );
and \U$11151 ( \11466 , \11463 , \11465 );
xor \U$11152 ( \11467 , \11034 , \11038 );
xor \U$11153 ( \11468 , \11467 , \11043 );
and \U$11154 ( \11469 , \11465 , \11468 );
and \U$11155 ( \11470 , \11463 , \11468 );
or \U$11156 ( \11471 , \11466 , \11469 , \11470 );
xor \U$11157 ( \11472 , \11050 , \11054 );
xor \U$11158 ( \11473 , \11472 , \11059 );
xor \U$11159 ( \11474 , \11067 , \11071 );
xor \U$11160 ( \11475 , \11474 , \11076 );
and \U$11161 ( \11476 , \11473 , \11475 );
and \U$11162 ( \11477 , \11471 , \11476 );
xor \U$11163 ( \11478 , \10817 , \10821 );
and \U$11164 ( \11479 , \11476 , \11478 );
and \U$11165 ( \11480 , \11471 , \11478 );
or \U$11166 ( \11481 , \11477 , \11479 , \11480 );
and \U$11167 ( \11482 , \11460 , \11481 );
and \U$11168 ( \11483 , \11304 , \11481 );
or \U$11169 ( \11484 , \11461 , \11482 , \11483 );
xor \U$11170 ( \11485 , \10994 , \11010 );
xor \U$11171 ( \11486 , \11485 , \11027 );
xor \U$11172 ( \11487 , \11099 , \11115 );
xor \U$11173 ( \11488 , \11487 , \11132 );
and \U$11174 ( \11489 , \11486 , \11488 );
xor \U$11175 ( \11490 , \10966 , \10969 );
xor \U$11176 ( \11491 , \11490 , \10972 );
and \U$11177 ( \11492 , \11488 , \11491 );
and \U$11178 ( \11493 , \11486 , \11491 );
or \U$11179 ( \11494 , \11489 , \11492 , \11493 );
xor \U$11180 ( \11495 , \11141 , \11143 );
xor \U$11181 ( \11496 , \11495 , \11146 );
xor \U$11182 ( \11497 , \10931 , \10933 );
xor \U$11183 ( \11498 , \11497 , \10936 );
and \U$11184 ( \11499 , \11496 , \11498 );
xor \U$11185 ( \11500 , \10941 , \10943 );
xor \U$11186 ( \11501 , \11500 , \10946 );
and \U$11187 ( \11502 , \11498 , \11501 );
and \U$11188 ( \11503 , \11496 , \11501 );
or \U$11189 ( \11504 , \11499 , \11502 , \11503 );
and \U$11190 ( \11505 , \11494 , \11504 );
xor \U$11191 ( \11506 , \11161 , \11163 );
xor \U$11192 ( \11507 , \11506 , \11166 );
and \U$11193 ( \11508 , \11504 , \11507 );
and \U$11194 ( \11509 , \11494 , \11507 );
or \U$11195 ( \11510 , \11505 , \11508 , \11509 );
and \U$11196 ( \11511 , \11484 , \11510 );
xor \U$11197 ( \11512 , \10939 , \10949 );
xor \U$11198 ( \11513 , \11512 , \10975 );
xor \U$11199 ( \11514 , \11171 , \11173 );
xor \U$11200 ( \11515 , \11514 , \11175 );
and \U$11201 ( \11516 , \11513 , \11515 );
xor \U$11202 ( \11517 , \11149 , \11151 );
xor \U$11203 ( \11518 , \11517 , \11153 );
and \U$11204 ( \11519 , \11515 , \11518 );
and \U$11205 ( \11520 , \11513 , \11518 );
or \U$11206 ( \11521 , \11516 , \11519 , \11520 );
and \U$11207 ( \11522 , \11510 , \11521 );
and \U$11208 ( \11523 , \11484 , \11521 );
or \U$11209 ( \11524 , \11511 , \11522 , \11523 );
xor \U$11210 ( \11525 , \10625 , \10635 );
xor \U$11211 ( \11526 , \11525 , \10669 );
xor \U$11212 ( \11527 , \10724 , \10776 );
xor \U$11213 ( \11528 , \11527 , \10825 );
and \U$11214 ( \11529 , \11526 , \11528 );
xor \U$11215 ( \11530 , \11187 , \11189 );
xor \U$11216 ( \11531 , \11530 , \11192 );
and \U$11217 ( \11532 , \11528 , \11531 );
and \U$11218 ( \11533 , \11526 , \11531 );
or \U$11219 ( \11534 , \11529 , \11532 , \11533 );
and \U$11220 ( \11535 , \11524 , \11534 );
xor \U$11221 ( \11536 , \10672 , \10828 );
xor \U$11222 ( \11537 , \11536 , \10850 );
and \U$11223 ( \11538 , \11534 , \11537 );
and \U$11224 ( \11539 , \11524 , \11537 );
or \U$11225 ( \11540 , \11535 , \11538 , \11539 );
xor \U$11226 ( \11541 , \11198 , \11208 );
xor \U$11227 ( \11542 , \11541 , \11211 );
and \U$11228 ( \11543 , \11540 , \11542 );
xor \U$11229 ( \11544 , \11216 , \11218 );
and \U$11230 ( \11545 , \11542 , \11544 );
and \U$11231 ( \11546 , \11540 , \11544 );
or \U$11232 ( \11547 , \11543 , \11545 , \11546 );
xor \U$11233 ( \11548 , \11214 , \11219 );
xor \U$11234 ( \11549 , \11548 , \11222 );
and \U$11235 ( \11550 , \11547 , \11549 );
xor \U$11236 ( \11551 , \11227 , \11229 );
and \U$11237 ( \11552 , \11549 , \11551 );
and \U$11238 ( \11553 , \11547 , \11551 );
or \U$11239 ( \11554 , \11550 , \11552 , \11553 );
and \U$11240 ( \11555 , \11240 , \11554 );
xor \U$11241 ( \11556 , \11240 , \11554 );
xor \U$11242 ( \11557 , \11547 , \11549 );
xor \U$11243 ( \11558 , \11557 , \11551 );
and \U$11244 ( \11559 , \604 , \8896 );
and \U$11245 ( \11560 , \553 , \8894 );
nor \U$11246 ( \11561 , \11559 , \11560 );
xnor \U$11247 ( \11562 , \11561 , \8525 );
and \U$11248 ( \11563 , \709 , \8334 );
and \U$11249 ( \11564 , \681 , \8332 );
nor \U$11250 ( \11565 , \11563 , \11564 );
xnor \U$11251 ( \11566 , \11565 , \8016 );
and \U$11252 ( \11567 , \11562 , \11566 );
and \U$11253 ( \11568 , \863 , \7767 );
and \U$11254 ( \11569 , \789 , \7765 );
nor \U$11255 ( \11570 , \11568 , \11569 );
xnor \U$11256 ( \11571 , \11570 , \7518 );
and \U$11257 ( \11572 , \11566 , \11571 );
and \U$11258 ( \11573 , \11562 , \11571 );
or \U$11259 ( \11574 , \11567 , \11572 , \11573 );
and \U$11260 ( \11575 , \369 , \10814 );
and \U$11261 ( \11576 , \348 , \10811 );
nor \U$11262 ( \11577 , \11575 , \11576 );
xnor \U$11263 ( \11578 , \11577 , \9759 );
and \U$11264 ( \11579 , \425 , \10001 );
and \U$11265 ( \11580 , \417 , \9999 );
nor \U$11266 ( \11581 , \11579 , \11580 );
xnor \U$11267 ( \11582 , \11581 , \9762 );
and \U$11268 ( \11583 , \11578 , \11582 );
and \U$11269 ( \11584 , \499 , \9433 );
and \U$11270 ( \11585 , \494 , \9431 );
nor \U$11271 ( \11586 , \11584 , \11585 );
xnor \U$11272 ( \11587 , \11586 , \9123 );
and \U$11273 ( \11588 , \11582 , \11587 );
and \U$11274 ( \11589 , \11578 , \11587 );
or \U$11275 ( \11590 , \11583 , \11588 , \11589 );
and \U$11276 ( \11591 , \11574 , \11590 );
and \U$11277 ( \11592 , \988 , \7238 );
and \U$11278 ( \11593 , \925 , \7236 );
nor \U$11279 ( \11594 , \11592 , \11593 );
xnor \U$11280 ( \11595 , \11594 , \6978 );
and \U$11281 ( \11596 , \1274 , \6744 );
and \U$11282 ( \11597 , \1186 , \6742 );
nor \U$11283 ( \11598 , \11596 , \11597 );
xnor \U$11284 ( \11599 , \11598 , \6429 );
and \U$11285 ( \11600 , \11595 , \11599 );
and \U$11286 ( \11601 , \1384 , \6235 );
and \U$11287 ( \11602 , \1379 , \6233 );
nor \U$11288 ( \11603 , \11601 , \11602 );
xnor \U$11289 ( \11604 , \11603 , \5895 );
and \U$11290 ( \11605 , \11599 , \11604 );
and \U$11291 ( \11606 , \11595 , \11604 );
or \U$11292 ( \11607 , \11600 , \11605 , \11606 );
and \U$11293 ( \11608 , \11590 , \11607 );
and \U$11294 ( \11609 , \11574 , \11607 );
or \U$11295 ( \11610 , \11591 , \11608 , \11609 );
and \U$11296 ( \11611 , \5776 , \1554 );
and \U$11297 ( \11612 , \5517 , \1552 );
nor \U$11298 ( \11613 , \11611 , \11612 );
xnor \U$11299 ( \11614 , \11613 , \1441 );
and \U$11300 ( \11615 , \6157 , \1360 );
and \U$11301 ( \11616 , \6148 , \1358 );
nor \U$11302 ( \11617 , \11615 , \11616 );
xnor \U$11303 ( \11618 , \11617 , \1224 );
and \U$11304 ( \11619 , \11614 , \11618 );
and \U$11305 ( \11620 , \6702 , \1160 );
and \U$11306 ( \11621 , \6500 , \1158 );
nor \U$11307 ( \11622 , \11620 , \11621 );
xnor \U$11308 ( \11623 , \11622 , \1082 );
and \U$11309 ( \11624 , \11618 , \11623 );
and \U$11310 ( \11625 , \11614 , \11623 );
or \U$11311 ( \11626 , \11619 , \11624 , \11625 );
and \U$11312 ( \11627 , \7177 , \996 );
and \U$11313 ( \11628 , \7005 , \994 );
nor \U$11314 ( \11629 , \11627 , \11628 );
xnor \U$11315 ( \11630 , \11629 , \902 );
and \U$11316 ( \11631 , \8127 , \826 );
and \U$11317 ( \11632 , \7703 , \824 );
nor \U$11318 ( \11633 , \11631 , \11632 );
xnor \U$11319 ( \11634 , \11633 , \754 );
and \U$11320 ( \11635 , \11630 , \11634 );
and \U$11321 ( \11636 , \8378 , \692 );
and \U$11322 ( \11637 , \8373 , \690 );
nor \U$11323 ( \11638 , \11636 , \11637 );
xnor \U$11324 ( \11639 , \11638 , \649 );
and \U$11325 ( \11640 , \11634 , \11639 );
and \U$11326 ( \11641 , \11630 , \11639 );
or \U$11327 ( \11642 , \11635 , \11640 , \11641 );
and \U$11328 ( \11643 , \11626 , \11642 );
and \U$11329 ( \11644 , \4469 , \2300 );
and \U$11330 ( \11645 , \4272 , \2298 );
nor \U$11331 ( \11646 , \11644 , \11645 );
xnor \U$11332 ( \11647 , \11646 , \2163 );
and \U$11333 ( \11648 , \4779 , \2094 );
and \U$11334 ( \11649 , \4771 , \2092 );
nor \U$11335 ( \11650 , \11648 , \11649 );
xnor \U$11336 ( \11651 , \11650 , \1942 );
and \U$11337 ( \11652 , \11647 , \11651 );
and \U$11338 ( \11653 , \5253 , \1826 );
and \U$11339 ( \11654 , \5248 , \1824 );
nor \U$11340 ( \11655 , \11653 , \11654 );
xnor \U$11341 ( \11656 , \11655 , \1670 );
and \U$11342 ( \11657 , \11651 , \11656 );
and \U$11343 ( \11658 , \11647 , \11656 );
or \U$11344 ( \11659 , \11652 , \11657 , \11658 );
and \U$11345 ( \11660 , \11642 , \11659 );
and \U$11346 ( \11661 , \11626 , \11659 );
or \U$11347 ( \11662 , \11643 , \11660 , \11661 );
and \U$11348 ( \11663 , \11610 , \11662 );
and \U$11349 ( \11664 , \1615 , \5646 );
and \U$11350 ( \11665 , \1500 , \5644 );
nor \U$11351 ( \11666 , \11664 , \11665 );
xnor \U$11352 ( \11667 , \11666 , \5405 );
and \U$11353 ( \11668 , \1799 , \5180 );
and \U$11354 ( \11669 , \1791 , \5178 );
nor \U$11355 ( \11670 , \11668 , \11669 );
xnor \U$11356 ( \11671 , \11670 , \4992 );
and \U$11357 ( \11672 , \11667 , \11671 );
and \U$11358 ( \11673 , \2047 , \4806 );
and \U$11359 ( \11674 , \2042 , \4804 );
nor \U$11360 ( \11675 , \11673 , \11674 );
xnor \U$11361 ( \11676 , \11675 , \4574 );
and \U$11362 ( \11677 , \11671 , \11676 );
and \U$11363 ( \11678 , \11667 , \11676 );
or \U$11364 ( \11679 , \11672 , \11677 , \11678 );
and \U$11365 ( \11680 , \3264 , \3324 );
and \U$11366 ( \11681 , \3145 , \3322 );
nor \U$11367 ( \11682 , \11680 , \11681 );
xnor \U$11368 ( \11683 , \11682 , \3119 );
and \U$11369 ( \11684 , \3889 , \2918 );
and \U$11370 ( \11685 , \3681 , \2916 );
nor \U$11371 ( \11686 , \11684 , \11685 );
xnor \U$11372 ( \11687 , \11686 , \2769 );
and \U$11373 ( \11688 , \11683 , \11687 );
and \U$11374 ( \11689 , \4016 , \2596 );
and \U$11375 ( \11690 , \4011 , \2594 );
nor \U$11376 ( \11691 , \11689 , \11690 );
xnor \U$11377 ( \11692 , \11691 , \2454 );
and \U$11378 ( \11693 , \11687 , \11692 );
and \U$11379 ( \11694 , \11683 , \11692 );
or \U$11380 ( \11695 , \11688 , \11693 , \11694 );
and \U$11381 ( \11696 , \11679 , \11695 );
and \U$11382 ( \11697 , \2377 , \4355 );
and \U$11383 ( \11698 , \2233 , \4353 );
nor \U$11384 ( \11699 , \11697 , \11698 );
xnor \U$11385 ( \11700 , \11699 , \4212 );
and \U$11386 ( \11701 , \2666 , \4032 );
and \U$11387 ( \11702 , \2641 , \4030 );
nor \U$11388 ( \11703 , \11701 , \11702 );
xnor \U$11389 ( \11704 , \11703 , \3786 );
and \U$11390 ( \11705 , \11700 , \11704 );
and \U$11391 ( \11706 , \3007 , \3637 );
and \U$11392 ( \11707 , \2840 , \3635 );
nor \U$11393 ( \11708 , \11706 , \11707 );
xnor \U$11394 ( \11709 , \11708 , \3450 );
and \U$11395 ( \11710 , \11704 , \11709 );
and \U$11396 ( \11711 , \11700 , \11709 );
or \U$11397 ( \11712 , \11705 , \11710 , \11711 );
and \U$11398 ( \11713 , \11695 , \11712 );
and \U$11399 ( \11714 , \11679 , \11712 );
or \U$11400 ( \11715 , \11696 , \11713 , \11714 );
and \U$11401 ( \11716 , \11662 , \11715 );
and \U$11402 ( \11717 , \11610 , \11715 );
or \U$11403 ( \11718 , \11663 , \11716 , \11717 );
xor \U$11404 ( \11719 , \11409 , \11413 );
xor \U$11405 ( \11720 , \11719 , \11418 );
xor \U$11406 ( \11721 , \11425 , \11429 );
xor \U$11407 ( \11722 , \11721 , \11434 );
and \U$11408 ( \11723 , \11720 , \11722 );
xor \U$11409 ( \11724 , \11442 , \11446 );
xor \U$11410 ( \11725 , \11724 , \11451 );
and \U$11411 ( \11726 , \11722 , \11725 );
and \U$11412 ( \11727 , \11720 , \11725 );
or \U$11413 ( \11728 , \11723 , \11726 , \11727 );
and \U$11414 ( \11729 , \8981 , \579 );
and \U$11415 ( \11730 , \8697 , \577 );
nor \U$11416 ( \11731 , \11729 , \11730 );
xnor \U$11417 ( \11732 , \11731 , \530 );
and \U$11418 ( \11733 , \9558 , \478 );
and \U$11419 ( \11734 , \9550 , \476 );
nor \U$11420 ( \11735 , \11733 , \11734 );
xnor \U$11421 ( \11736 , \11735 , \437 );
and \U$11422 ( \11737 , \11732 , \11736 );
and \U$11423 ( \11738 , \10166 , \408 );
and \U$11424 ( \11739 , \10161 , \406 );
nor \U$11425 ( \11740 , \11738 , \11739 );
xnor \U$11426 ( \11741 , \11740 , \378 );
and \U$11427 ( \11742 , \11736 , \11741 );
and \U$11428 ( \11743 , \11732 , \11741 );
or \U$11429 ( \11744 , \11737 , \11742 , \11743 );
xor \U$11430 ( \11745 , \11244 , \11248 );
xor \U$11431 ( \11746 , \11745 , \11251 );
and \U$11432 ( \11747 , \11744 , \11746 );
xor \U$11433 ( \11748 , \11258 , \11262 );
xor \U$11434 ( \11749 , \11748 , \11267 );
and \U$11435 ( \11750 , \11746 , \11749 );
and \U$11436 ( \11751 , \11744 , \11749 );
or \U$11437 ( \11752 , \11747 , \11750 , \11751 );
and \U$11438 ( \11753 , \11728 , \11752 );
xor \U$11439 ( \11754 , \11308 , \11312 );
xor \U$11440 ( \11755 , \11754 , \11317 );
xor \U$11441 ( \11756 , \11324 , \11328 );
xor \U$11442 ( \11757 , \11756 , \11333 );
and \U$11443 ( \11758 , \11755 , \11757 );
xor \U$11444 ( \11759 , \11341 , \11345 );
xor \U$11445 ( \11760 , \11759 , \11350 );
and \U$11446 ( \11761 , \11757 , \11760 );
and \U$11447 ( \11762 , \11755 , \11760 );
or \U$11448 ( \11763 , \11758 , \11761 , \11762 );
and \U$11449 ( \11764 , \11752 , \11763 );
and \U$11450 ( \11765 , \11728 , \11763 );
or \U$11451 ( \11766 , \11753 , \11764 , \11765 );
and \U$11452 ( \11767 , \11718 , \11766 );
xor \U$11453 ( \11768 , \11360 , \11364 );
xor \U$11454 ( \11769 , \11768 , \11369 );
xor \U$11455 ( \11770 , \11376 , \11380 );
xor \U$11456 ( \11771 , \11770 , \328 );
and \U$11457 ( \11772 , \11769 , \11771 );
xor \U$11458 ( \11773 , \11389 , \11393 );
xor \U$11459 ( \11774 , \11773 , \11398 );
and \U$11460 ( \11775 , \11771 , \11774 );
and \U$11461 ( \11776 , \11769 , \11774 );
or \U$11462 ( \11777 , \11772 , \11775 , \11776 );
xor \U$11463 ( \11778 , \11463 , \11465 );
xor \U$11464 ( \11779 , \11778 , \11468 );
and \U$11465 ( \11780 , \11777 , \11779 );
xor \U$11466 ( \11781 , \11473 , \11475 );
and \U$11467 ( \11782 , \11779 , \11781 );
and \U$11468 ( \11783 , \11777 , \11781 );
or \U$11469 ( \11784 , \11780 , \11782 , \11783 );
and \U$11470 ( \11785 , \11766 , \11784 );
and \U$11471 ( \11786 , \11718 , \11784 );
or \U$11472 ( \11787 , \11767 , \11785 , \11786 );
xor \U$11473 ( \11788 , \11320 , \11336 );
xor \U$11474 ( \11789 , \11788 , \11353 );
xor \U$11475 ( \11790 , \11372 , \11384 );
xor \U$11476 ( \11791 , \11790 , \11401 );
and \U$11477 ( \11792 , \11789 , \11791 );
xor \U$11478 ( \11793 , \11421 , \11437 );
xor \U$11479 ( \11794 , \11793 , \11454 );
and \U$11480 ( \11795 , \11791 , \11794 );
and \U$11481 ( \11796 , \11789 , \11794 );
or \U$11482 ( \11797 , \11792 , \11795 , \11796 );
xor \U$11483 ( \11798 , \11254 , \11270 );
xor \U$11484 ( \11799 , \11798 , \11275 );
xor \U$11485 ( \11800 , \11282 , \11284 );
xor \U$11486 ( \11801 , \11800 , \11287 );
and \U$11487 ( \11802 , \11799 , \11801 );
xor \U$11488 ( \11803 , \11293 , \11295 );
xor \U$11489 ( \11804 , \11803 , \11298 );
and \U$11490 ( \11805 , \11801 , \11804 );
and \U$11491 ( \11806 , \11799 , \11804 );
or \U$11492 ( \11807 , \11802 , \11805 , \11806 );
and \U$11493 ( \11808 , \11797 , \11807 );
xor \U$11494 ( \11809 , \11046 , \11062 );
xor \U$11495 ( \11810 , \11809 , \11079 );
and \U$11496 ( \11811 , \11807 , \11810 );
and \U$11497 ( \11812 , \11797 , \11810 );
or \U$11498 ( \11813 , \11808 , \11811 , \11812 );
and \U$11499 ( \11814 , \11787 , \11813 );
xor \U$11500 ( \11815 , \11486 , \11488 );
xor \U$11501 ( \11816 , \11815 , \11491 );
xor \U$11502 ( \11817 , \11496 , \11498 );
xor \U$11503 ( \11818 , \11817 , \11501 );
and \U$11504 ( \11819 , \11816 , \11818 );
xor \U$11505 ( \11820 , \11471 , \11476 );
xor \U$11506 ( \11821 , \11820 , \11478 );
and \U$11507 ( \11822 , \11818 , \11821 );
and \U$11508 ( \11823 , \11816 , \11821 );
or \U$11509 ( \11824 , \11819 , \11822 , \11823 );
and \U$11510 ( \11825 , \11813 , \11824 );
and \U$11511 ( \11826 , \11787 , \11824 );
or \U$11512 ( \11827 , \11814 , \11825 , \11826 );
xor \U$11513 ( \11828 , \11030 , \11082 );
xor \U$11514 ( \11829 , \11828 , \11135 );
xor \U$11515 ( \11830 , \11494 , \11504 );
xor \U$11516 ( \11831 , \11830 , \11507 );
and \U$11517 ( \11832 , \11829 , \11831 );
xor \U$11518 ( \11833 , \11513 , \11515 );
xor \U$11519 ( \11834 , \11833 , \11518 );
and \U$11520 ( \11835 , \11831 , \11834 );
and \U$11521 ( \11836 , \11829 , \11834 );
or \U$11522 ( \11837 , \11832 , \11835 , \11836 );
and \U$11523 ( \11838 , \11827 , \11837 );
xor \U$11524 ( \11839 , \11169 , \11178 );
xor \U$11525 ( \11840 , \11839 , \11181 );
and \U$11526 ( \11841 , \11837 , \11840 );
and \U$11527 ( \11842 , \11827 , \11840 );
or \U$11528 ( \11843 , \11838 , \11841 , \11842 );
xor \U$11529 ( \11844 , \10978 , \11138 );
xor \U$11530 ( \11845 , \11844 , \11156 );
xor \U$11531 ( \11846 , \11484 , \11510 );
xor \U$11532 ( \11847 , \11846 , \11521 );
and \U$11533 ( \11848 , \11845 , \11847 );
xor \U$11534 ( \11849 , \11526 , \11528 );
xor \U$11535 ( \11850 , \11849 , \11531 );
and \U$11536 ( \11851 , \11847 , \11850 );
and \U$11537 ( \11852 , \11845 , \11850 );
or \U$11538 ( \11853 , \11848 , \11851 , \11852 );
and \U$11539 ( \11854 , \11843 , \11853 );
xor \U$11540 ( \11855 , \11200 , \11202 );
xor \U$11541 ( \11856 , \11855 , \11205 );
and \U$11542 ( \11857 , \11853 , \11856 );
and \U$11543 ( \11858 , \11843 , \11856 );
or \U$11544 ( \11859 , \11854 , \11857 , \11858 );
xor \U$11545 ( \11860 , \11159 , \11184 );
xor \U$11546 ( \11861 , \11860 , \11195 );
xor \U$11547 ( \11862 , \11524 , \11534 );
xor \U$11548 ( \11863 , \11862 , \11537 );
and \U$11549 ( \11864 , \11861 , \11863 );
and \U$11550 ( \11865 , \11859 , \11864 );
xor \U$11551 ( \11866 , \11540 , \11542 );
xor \U$11552 ( \11867 , \11866 , \11544 );
and \U$11553 ( \11868 , \11864 , \11867 );
and \U$11554 ( \11869 , \11859 , \11867 );
or \U$11555 ( \11870 , \11865 , \11868 , \11869 );
and \U$11556 ( \11871 , \11558 , \11870 );
xor \U$11557 ( \11872 , \11558 , \11870 );
xor \U$11558 ( \11873 , \11859 , \11864 );
xor \U$11559 ( \11874 , \11873 , \11867 );
and \U$11560 ( \11875 , \7005 , \1160 );
and \U$11561 ( \11876 , \6702 , \1158 );
nor \U$11562 ( \11877 , \11875 , \11876 );
xnor \U$11563 ( \11878 , \11877 , \1082 );
and \U$11564 ( \11879 , \7703 , \996 );
and \U$11565 ( \11880 , \7177 , \994 );
nor \U$11566 ( \11881 , \11879 , \11880 );
xnor \U$11567 ( \11882 , \11881 , \902 );
and \U$11568 ( \11883 , \11878 , \11882 );
and \U$11569 ( \11884 , \8373 , \826 );
and \U$11570 ( \11885 , \8127 , \824 );
nor \U$11571 ( \11886 , \11884 , \11885 );
xnor \U$11572 ( \11887 , \11886 , \754 );
and \U$11573 ( \11888 , \11882 , \11887 );
and \U$11574 ( \11889 , \11878 , \11887 );
or \U$11575 ( \11890 , \11883 , \11888 , \11889 );
and \U$11576 ( \11891 , \4272 , \2596 );
and \U$11577 ( \11892 , \4016 , \2594 );
nor \U$11578 ( \11893 , \11891 , \11892 );
xnor \U$11579 ( \11894 , \11893 , \2454 );
and \U$11580 ( \11895 , \4771 , \2300 );
and \U$11581 ( \11896 , \4469 , \2298 );
nor \U$11582 ( \11897 , \11895 , \11896 );
xnor \U$11583 ( \11898 , \11897 , \2163 );
and \U$11584 ( \11899 , \11894 , \11898 );
and \U$11585 ( \11900 , \5248 , \2094 );
and \U$11586 ( \11901 , \4779 , \2092 );
nor \U$11587 ( \11902 , \11900 , \11901 );
xnor \U$11588 ( \11903 , \11902 , \1942 );
and \U$11589 ( \11904 , \11898 , \11903 );
and \U$11590 ( \11905 , \11894 , \11903 );
or \U$11591 ( \11906 , \11899 , \11904 , \11905 );
and \U$11592 ( \11907 , \11890 , \11906 );
and \U$11593 ( \11908 , \5517 , \1826 );
and \U$11594 ( \11909 , \5253 , \1824 );
nor \U$11595 ( \11910 , \11908 , \11909 );
xnor \U$11596 ( \11911 , \11910 , \1670 );
and \U$11597 ( \11912 , \6148 , \1554 );
and \U$11598 ( \11913 , \5776 , \1552 );
nor \U$11599 ( \11914 , \11912 , \11913 );
xnor \U$11600 ( \11915 , \11914 , \1441 );
and \U$11601 ( \11916 , \11911 , \11915 );
and \U$11602 ( \11917 , \6500 , \1360 );
and \U$11603 ( \11918 , \6157 , \1358 );
nor \U$11604 ( \11919 , \11917 , \11918 );
xnor \U$11605 ( \11920 , \11919 , \1224 );
and \U$11606 ( \11921 , \11915 , \11920 );
and \U$11607 ( \11922 , \11911 , \11920 );
or \U$11608 ( \11923 , \11916 , \11921 , \11922 );
and \U$11609 ( \11924 , \11906 , \11923 );
and \U$11610 ( \11925 , \11890 , \11923 );
or \U$11611 ( \11926 , \11907 , \11924 , \11925 );
and \U$11612 ( \11927 , \925 , \7767 );
and \U$11613 ( \11928 , \863 , \7765 );
nor \U$11614 ( \11929 , \11927 , \11928 );
xnor \U$11615 ( \11930 , \11929 , \7518 );
and \U$11616 ( \11931 , \1186 , \7238 );
and \U$11617 ( \11932 , \988 , \7236 );
nor \U$11618 ( \11933 , \11931 , \11932 );
xnor \U$11619 ( \11934 , \11933 , \6978 );
and \U$11620 ( \11935 , \11930 , \11934 );
and \U$11621 ( \11936 , \1379 , \6744 );
and \U$11622 ( \11937 , \1274 , \6742 );
nor \U$11623 ( \11938 , \11936 , \11937 );
xnor \U$11624 ( \11939 , \11938 , \6429 );
and \U$11625 ( \11940 , \11934 , \11939 );
and \U$11626 ( \11941 , \11930 , \11939 );
or \U$11627 ( \11942 , \11935 , \11940 , \11941 );
and \U$11628 ( \11943 , \553 , \9433 );
and \U$11629 ( \11944 , \499 , \9431 );
nor \U$11630 ( \11945 , \11943 , \11944 );
xnor \U$11631 ( \11946 , \11945 , \9123 );
and \U$11632 ( \11947 , \681 , \8896 );
and \U$11633 ( \11948 , \604 , \8894 );
nor \U$11634 ( \11949 , \11947 , \11948 );
xnor \U$11635 ( \11950 , \11949 , \8525 );
and \U$11636 ( \11951 , \11946 , \11950 );
and \U$11637 ( \11952 , \789 , \8334 );
and \U$11638 ( \11953 , \709 , \8332 );
nor \U$11639 ( \11954 , \11952 , \11953 );
xnor \U$11640 ( \11955 , \11954 , \8016 );
and \U$11641 ( \11956 , \11950 , \11955 );
and \U$11642 ( \11957 , \11946 , \11955 );
or \U$11643 ( \11958 , \11951 , \11956 , \11957 );
and \U$11644 ( \11959 , \11942 , \11958 );
and \U$11645 ( \11960 , \417 , \10814 );
and \U$11646 ( \11961 , \369 , \10811 );
nor \U$11647 ( \11962 , \11960 , \11961 );
xnor \U$11648 ( \11963 , \11962 , \9759 );
and \U$11649 ( \11964 , \494 , \10001 );
and \U$11650 ( \11965 , \425 , \9999 );
nor \U$11651 ( \11966 , \11964 , \11965 );
xnor \U$11652 ( \11967 , \11966 , \9762 );
and \U$11653 ( \11968 , \11963 , \11967 );
and \U$11654 ( \11969 , \11967 , \341 );
and \U$11655 ( \11970 , \11963 , \341 );
or \U$11656 ( \11971 , \11968 , \11969 , \11970 );
and \U$11657 ( \11972 , \11958 , \11971 );
and \U$11658 ( \11973 , \11942 , \11971 );
or \U$11659 ( \11974 , \11959 , \11972 , \11973 );
and \U$11660 ( \11975 , \11926 , \11974 );
and \U$11661 ( \11976 , \1500 , \6235 );
and \U$11662 ( \11977 , \1384 , \6233 );
nor \U$11663 ( \11978 , \11976 , \11977 );
xnor \U$11664 ( \11979 , \11978 , \5895 );
and \U$11665 ( \11980 , \1791 , \5646 );
and \U$11666 ( \11981 , \1615 , \5644 );
nor \U$11667 ( \11982 , \11980 , \11981 );
xnor \U$11668 ( \11983 , \11982 , \5405 );
and \U$11669 ( \11984 , \11979 , \11983 );
and \U$11670 ( \11985 , \2042 , \5180 );
and \U$11671 ( \11986 , \1799 , \5178 );
nor \U$11672 ( \11987 , \11985 , \11986 );
xnor \U$11673 ( \11988 , \11987 , \4992 );
and \U$11674 ( \11989 , \11983 , \11988 );
and \U$11675 ( \11990 , \11979 , \11988 );
or \U$11676 ( \11991 , \11984 , \11989 , \11990 );
and \U$11677 ( \11992 , \2233 , \4806 );
and \U$11678 ( \11993 , \2047 , \4804 );
nor \U$11679 ( \11994 , \11992 , \11993 );
xnor \U$11680 ( \11995 , \11994 , \4574 );
and \U$11681 ( \11996 , \2641 , \4355 );
and \U$11682 ( \11997 , \2377 , \4353 );
nor \U$11683 ( \11998 , \11996 , \11997 );
xnor \U$11684 ( \11999 , \11998 , \4212 );
and \U$11685 ( \12000 , \11995 , \11999 );
and \U$11686 ( \12001 , \2840 , \4032 );
and \U$11687 ( \12002 , \2666 , \4030 );
nor \U$11688 ( \12003 , \12001 , \12002 );
xnor \U$11689 ( \12004 , \12003 , \3786 );
and \U$11690 ( \12005 , \11999 , \12004 );
and \U$11691 ( \12006 , \11995 , \12004 );
or \U$11692 ( \12007 , \12000 , \12005 , \12006 );
and \U$11693 ( \12008 , \11991 , \12007 );
and \U$11694 ( \12009 , \3145 , \3637 );
and \U$11695 ( \12010 , \3007 , \3635 );
nor \U$11696 ( \12011 , \12009 , \12010 );
xnor \U$11697 ( \12012 , \12011 , \3450 );
and \U$11698 ( \12013 , \3681 , \3324 );
and \U$11699 ( \12014 , \3264 , \3322 );
nor \U$11700 ( \12015 , \12013 , \12014 );
xnor \U$11701 ( \12016 , \12015 , \3119 );
and \U$11702 ( \12017 , \12012 , \12016 );
and \U$11703 ( \12018 , \4011 , \2918 );
and \U$11704 ( \12019 , \3889 , \2916 );
nor \U$11705 ( \12020 , \12018 , \12019 );
xnor \U$11706 ( \12021 , \12020 , \2769 );
and \U$11707 ( \12022 , \12016 , \12021 );
and \U$11708 ( \12023 , \12012 , \12021 );
or \U$11709 ( \12024 , \12017 , \12022 , \12023 );
and \U$11710 ( \12025 , \12007 , \12024 );
and \U$11711 ( \12026 , \11991 , \12024 );
or \U$11712 ( \12027 , \12008 , \12025 , \12026 );
and \U$11713 ( \12028 , \11974 , \12027 );
and \U$11714 ( \12029 , \11926 , \12027 );
or \U$11715 ( \12030 , \11975 , \12028 , \12029 );
and \U$11716 ( \12031 , \8697 , \692 );
and \U$11717 ( \12032 , \8378 , \690 );
nor \U$11718 ( \12033 , \12031 , \12032 );
xnor \U$11719 ( \12034 , \12033 , \649 );
and \U$11720 ( \12035 , \9550 , \579 );
and \U$11721 ( \12036 , \8981 , \577 );
nor \U$11722 ( \12037 , \12035 , \12036 );
xnor \U$11723 ( \12038 , \12037 , \530 );
and \U$11724 ( \12039 , \12034 , \12038 );
and \U$11725 ( \12040 , \10161 , \478 );
and \U$11726 ( \12041 , \9558 , \476 );
nor \U$11727 ( \12042 , \12040 , \12041 );
xnor \U$11728 ( \12043 , \12042 , \437 );
and \U$11729 ( \12044 , \12038 , \12043 );
and \U$11730 ( \12045 , \12034 , \12043 );
or \U$11731 ( \12046 , \12039 , \12044 , \12045 );
and \U$11732 ( \12047 , \10347 , \408 );
and \U$11733 ( \12048 , \10166 , \406 );
nor \U$11734 ( \12049 , \12047 , \12048 );
xnor \U$11735 ( \12050 , \12049 , \378 );
nand \U$11736 ( \12051 , \10967 , \358 );
xnor \U$11737 ( \12052 , \12051 , \341 );
and \U$11738 ( \12053 , \12050 , \12052 );
and \U$11739 ( \12054 , \12046 , \12053 );
and \U$11740 ( \12055 , \10967 , \360 );
and \U$11741 ( \12056 , \10347 , \358 );
nor \U$11742 ( \12057 , \12055 , \12056 );
xnor \U$11743 ( \12058 , \12057 , \341 );
and \U$11744 ( \12059 , \12053 , \12058 );
and \U$11745 ( \12060 , \12046 , \12058 );
or \U$11746 ( \12061 , \12054 , \12059 , \12060 );
xor \U$11747 ( \12062 , \11647 , \11651 );
xor \U$11748 ( \12063 , \12062 , \11656 );
xor \U$11749 ( \12064 , \11683 , \11687 );
xor \U$11750 ( \12065 , \12064 , \11692 );
and \U$11751 ( \12066 , \12063 , \12065 );
xor \U$11752 ( \12067 , \11700 , \11704 );
xor \U$11753 ( \12068 , \12067 , \11709 );
and \U$11754 ( \12069 , \12065 , \12068 );
and \U$11755 ( \12070 , \12063 , \12068 );
or \U$11756 ( \12071 , \12066 , \12069 , \12070 );
and \U$11757 ( \12072 , \12061 , \12071 );
xor \U$11758 ( \12073 , \11614 , \11618 );
xor \U$11759 ( \12074 , \12073 , \11623 );
xor \U$11760 ( \12075 , \11630 , \11634 );
xor \U$11761 ( \12076 , \12075 , \11639 );
and \U$11762 ( \12077 , \12074 , \12076 );
xor \U$11763 ( \12078 , \11732 , \11736 );
xor \U$11764 ( \12079 , \12078 , \11741 );
and \U$11765 ( \12080 , \12076 , \12079 );
and \U$11766 ( \12081 , \12074 , \12079 );
or \U$11767 ( \12082 , \12077 , \12080 , \12081 );
and \U$11768 ( \12083 , \12071 , \12082 );
and \U$11769 ( \12084 , \12061 , \12082 );
or \U$11770 ( \12085 , \12072 , \12083 , \12084 );
and \U$11771 ( \12086 , \12030 , \12085 );
xor \U$11772 ( \12087 , \11562 , \11566 );
xor \U$11773 ( \12088 , \12087 , \11571 );
xor \U$11774 ( \12089 , \11667 , \11671 );
xor \U$11775 ( \12090 , \12089 , \11676 );
and \U$11776 ( \12091 , \12088 , \12090 );
xor \U$11777 ( \12092 , \11595 , \11599 );
xor \U$11778 ( \12093 , \12092 , \11604 );
and \U$11779 ( \12094 , \12090 , \12093 );
and \U$11780 ( \12095 , \12088 , \12093 );
or \U$11781 ( \12096 , \12091 , \12094 , \12095 );
xor \U$11782 ( \12097 , \11769 , \11771 );
xor \U$11783 ( \12098 , \12097 , \11774 );
and \U$11784 ( \12099 , \12096 , \12098 );
xor \U$11785 ( \12100 , \11720 , \11722 );
xor \U$11786 ( \12101 , \12100 , \11725 );
and \U$11787 ( \12102 , \12098 , \12101 );
and \U$11788 ( \12103 , \12096 , \12101 );
or \U$11789 ( \12104 , \12099 , \12102 , \12103 );
and \U$11790 ( \12105 , \12085 , \12104 );
and \U$11791 ( \12106 , \12030 , \12104 );
or \U$11792 ( \12107 , \12086 , \12105 , \12106 );
xor \U$11793 ( \12108 , \11626 , \11642 );
xor \U$11794 ( \12109 , \12108 , \11659 );
xor \U$11795 ( \12110 , \11744 , \11746 );
xor \U$11796 ( \12111 , \12110 , \11749 );
and \U$11797 ( \12112 , \12109 , \12111 );
xor \U$11798 ( \12113 , \11755 , \11757 );
xor \U$11799 ( \12114 , \12113 , \11760 );
and \U$11800 ( \12115 , \12111 , \12114 );
and \U$11801 ( \12116 , \12109 , \12114 );
or \U$11802 ( \12117 , \12112 , \12115 , \12116 );
xor \U$11803 ( \12118 , \11789 , \11791 );
xor \U$11804 ( \12119 , \12118 , \11794 );
and \U$11805 ( \12120 , \12117 , \12119 );
xor \U$11806 ( \12121 , \11799 , \11801 );
xor \U$11807 ( \12122 , \12121 , \11804 );
and \U$11808 ( \12123 , \12119 , \12122 );
and \U$11809 ( \12124 , \12117 , \12122 );
or \U$11810 ( \12125 , \12120 , \12123 , \12124 );
and \U$11811 ( \12126 , \12107 , \12125 );
xor \U$11812 ( \12127 , \11610 , \11662 );
xor \U$11813 ( \12128 , \12127 , \11715 );
xor \U$11814 ( \12129 , \11728 , \11752 );
xor \U$11815 ( \12130 , \12129 , \11763 );
and \U$11816 ( \12131 , \12128 , \12130 );
xor \U$11817 ( \12132 , \11777 , \11779 );
xor \U$11818 ( \12133 , \12132 , \11781 );
and \U$11819 ( \12134 , \12130 , \12133 );
and \U$11820 ( \12135 , \12128 , \12133 );
or \U$11821 ( \12136 , \12131 , \12134 , \12135 );
and \U$11822 ( \12137 , \12125 , \12136 );
and \U$11823 ( \12138 , \12107 , \12136 );
or \U$11824 ( \12139 , \12126 , \12137 , \12138 );
xor \U$11825 ( \12140 , \11278 , \11290 );
xor \U$11826 ( \12141 , \12140 , \11301 );
xor \U$11827 ( \12142 , \11356 , \11404 );
xor \U$11828 ( \12143 , \12142 , \11457 );
and \U$11829 ( \12144 , \12141 , \12143 );
xor \U$11830 ( \12145 , \11816 , \11818 );
xor \U$11831 ( \12146 , \12145 , \11821 );
and \U$11832 ( \12147 , \12143 , \12146 );
and \U$11833 ( \12148 , \12141 , \12146 );
or \U$11834 ( \12149 , \12144 , \12147 , \12148 );
and \U$11835 ( \12150 , \12139 , \12149 );
xor \U$11836 ( \12151 , \11304 , \11460 );
xor \U$11837 ( \12152 , \12151 , \11481 );
and \U$11838 ( \12153 , \12149 , \12152 );
and \U$11839 ( \12154 , \12139 , \12152 );
or \U$11840 ( \12155 , \12150 , \12153 , \12154 );
xor \U$11841 ( \12156 , \11827 , \11837 );
xor \U$11842 ( \12157 , \12156 , \11840 );
and \U$11843 ( \12158 , \12155 , \12157 );
xor \U$11844 ( \12159 , \11845 , \11847 );
xor \U$11845 ( \12160 , \12159 , \11850 );
and \U$11846 ( \12161 , \12157 , \12160 );
and \U$11847 ( \12162 , \12155 , \12160 );
or \U$11848 ( \12163 , \12158 , \12161 , \12162 );
xor \U$11849 ( \12164 , \11843 , \11853 );
xor \U$11850 ( \12165 , \12164 , \11856 );
and \U$11851 ( \12166 , \12163 , \12165 );
xor \U$11852 ( \12167 , \11861 , \11863 );
and \U$11853 ( \12168 , \12165 , \12167 );
and \U$11854 ( \12169 , \12163 , \12167 );
or \U$11855 ( \12170 , \12166 , \12168 , \12169 );
and \U$11856 ( \12171 , \11874 , \12170 );
xor \U$11857 ( \12172 , \11874 , \12170 );
xor \U$11858 ( \12173 , \12163 , \12165 );
xor \U$11859 ( \12174 , \12173 , \12167 );
xor \U$11860 ( \12175 , \11878 , \11882 );
xor \U$11861 ( \12176 , \12175 , \11887 );
xor \U$11862 ( \12177 , \11894 , \11898 );
xor \U$11863 ( \12178 , \12177 , \11903 );
and \U$11864 ( \12179 , \12176 , \12178 );
xor \U$11865 ( \12180 , \11911 , \11915 );
xor \U$11866 ( \12181 , \12180 , \11920 );
and \U$11867 ( \12182 , \12178 , \12181 );
and \U$11868 ( \12183 , \12176 , \12181 );
or \U$11869 ( \12184 , \12179 , \12182 , \12183 );
xor \U$11870 ( \12185 , \11979 , \11983 );
xor \U$11871 ( \12186 , \12185 , \11988 );
xor \U$11872 ( \12187 , \11995 , \11999 );
xor \U$11873 ( \12188 , \12187 , \12004 );
and \U$11874 ( \12189 , \12186 , \12188 );
xor \U$11875 ( \12190 , \12012 , \12016 );
xor \U$11876 ( \12191 , \12190 , \12021 );
and \U$11877 ( \12192 , \12188 , \12191 );
and \U$11878 ( \12193 , \12186 , \12191 );
or \U$11879 ( \12194 , \12189 , \12192 , \12193 );
and \U$11880 ( \12195 , \12184 , \12194 );
and \U$11881 ( \12196 , \9558 , \579 );
and \U$11882 ( \12197 , \9550 , \577 );
nor \U$11883 ( \12198 , \12196 , \12197 );
xnor \U$11884 ( \12199 , \12198 , \530 );
and \U$11885 ( \12200 , \10166 , \478 );
and \U$11886 ( \12201 , \10161 , \476 );
nor \U$11887 ( \12202 , \12200 , \12201 );
xnor \U$11888 ( \12203 , \12202 , \437 );
and \U$11889 ( \12204 , \12199 , \12203 );
and \U$11890 ( \12205 , \10967 , \408 );
and \U$11891 ( \12206 , \10347 , \406 );
nor \U$11892 ( \12207 , \12205 , \12206 );
xnor \U$11893 ( \12208 , \12207 , \378 );
and \U$11894 ( \12209 , \12203 , \12208 );
and \U$11895 ( \12210 , \12199 , \12208 );
or \U$11896 ( \12211 , \12204 , \12209 , \12210 );
xor \U$11897 ( \12212 , \12034 , \12038 );
xor \U$11898 ( \12213 , \12212 , \12043 );
and \U$11899 ( \12214 , \12211 , \12213 );
xor \U$11900 ( \12215 , \12050 , \12052 );
and \U$11901 ( \12216 , \12213 , \12215 );
and \U$11902 ( \12217 , \12211 , \12215 );
or \U$11903 ( \12218 , \12214 , \12216 , \12217 );
and \U$11904 ( \12219 , \12194 , \12218 );
and \U$11905 ( \12220 , \12184 , \12218 );
or \U$11906 ( \12221 , \12195 , \12219 , \12220 );
and \U$11907 ( \12222 , \3889 , \3324 );
and \U$11908 ( \12223 , \3681 , \3322 );
nor \U$11909 ( \12224 , \12222 , \12223 );
xnor \U$11910 ( \12225 , \12224 , \3119 );
and \U$11911 ( \12226 , \4016 , \2918 );
and \U$11912 ( \12227 , \4011 , \2916 );
nor \U$11913 ( \12228 , \12226 , \12227 );
xnor \U$11914 ( \12229 , \12228 , \2769 );
and \U$11915 ( \12230 , \12225 , \12229 );
and \U$11916 ( \12231 , \4469 , \2596 );
and \U$11917 ( \12232 , \4272 , \2594 );
nor \U$11918 ( \12233 , \12231 , \12232 );
xnor \U$11919 ( \12234 , \12233 , \2454 );
and \U$11920 ( \12235 , \12229 , \12234 );
and \U$11921 ( \12236 , \12225 , \12234 );
or \U$11922 ( \12237 , \12230 , \12235 , \12236 );
and \U$11923 ( \12238 , \1799 , \5646 );
and \U$11924 ( \12239 , \1791 , \5644 );
nor \U$11925 ( \12240 , \12238 , \12239 );
xnor \U$11926 ( \12241 , \12240 , \5405 );
and \U$11927 ( \12242 , \2047 , \5180 );
and \U$11928 ( \12243 , \2042 , \5178 );
nor \U$11929 ( \12244 , \12242 , \12243 );
xnor \U$11930 ( \12245 , \12244 , \4992 );
and \U$11931 ( \12246 , \12241 , \12245 );
and \U$11932 ( \12247 , \2377 , \4806 );
and \U$11933 ( \12248 , \2233 , \4804 );
nor \U$11934 ( \12249 , \12247 , \12248 );
xnor \U$11935 ( \12250 , \12249 , \4574 );
and \U$11936 ( \12251 , \12245 , \12250 );
and \U$11937 ( \12252 , \12241 , \12250 );
or \U$11938 ( \12253 , \12246 , \12251 , \12252 );
and \U$11939 ( \12254 , \12237 , \12253 );
and \U$11940 ( \12255 , \2666 , \4355 );
and \U$11941 ( \12256 , \2641 , \4353 );
nor \U$11942 ( \12257 , \12255 , \12256 );
xnor \U$11943 ( \12258 , \12257 , \4212 );
and \U$11944 ( \12259 , \3007 , \4032 );
and \U$11945 ( \12260 , \2840 , \4030 );
nor \U$11946 ( \12261 , \12259 , \12260 );
xnor \U$11947 ( \12262 , \12261 , \3786 );
and \U$11948 ( \12263 , \12258 , \12262 );
and \U$11949 ( \12264 , \3264 , \3637 );
and \U$11950 ( \12265 , \3145 , \3635 );
nor \U$11951 ( \12266 , \12264 , \12265 );
xnor \U$11952 ( \12267 , \12266 , \3450 );
and \U$11953 ( \12268 , \12262 , \12267 );
and \U$11954 ( \12269 , \12258 , \12267 );
or \U$11955 ( \12270 , \12263 , \12268 , \12269 );
and \U$11956 ( \12271 , \12253 , \12270 );
and \U$11957 ( \12272 , \12237 , \12270 );
or \U$11958 ( \12273 , \12254 , \12271 , \12272 );
and \U$11959 ( \12274 , \1274 , \7238 );
and \U$11960 ( \12275 , \1186 , \7236 );
nor \U$11961 ( \12276 , \12274 , \12275 );
xnor \U$11962 ( \12277 , \12276 , \6978 );
and \U$11963 ( \12278 , \1384 , \6744 );
and \U$11964 ( \12279 , \1379 , \6742 );
nor \U$11965 ( \12280 , \12278 , \12279 );
xnor \U$11966 ( \12281 , \12280 , \6429 );
and \U$11967 ( \12282 , \12277 , \12281 );
and \U$11968 ( \12283 , \1615 , \6235 );
and \U$11969 ( \12284 , \1500 , \6233 );
nor \U$11970 ( \12285 , \12283 , \12284 );
xnor \U$11971 ( \12286 , \12285 , \5895 );
and \U$11972 ( \12287 , \12281 , \12286 );
and \U$11973 ( \12288 , \12277 , \12286 );
or \U$11974 ( \12289 , \12282 , \12287 , \12288 );
and \U$11975 ( \12290 , \425 , \10814 );
and \U$11976 ( \12291 , \417 , \10811 );
nor \U$11977 ( \12292 , \12290 , \12291 );
xnor \U$11978 ( \12293 , \12292 , \9759 );
and \U$11979 ( \12294 , \499 , \10001 );
and \U$11980 ( \12295 , \494 , \9999 );
nor \U$11981 ( \12296 , \12294 , \12295 );
xnor \U$11982 ( \12297 , \12296 , \9762 );
and \U$11983 ( \12298 , \12293 , \12297 );
and \U$11984 ( \12299 , \604 , \9433 );
and \U$11985 ( \12300 , \553 , \9431 );
nor \U$11986 ( \12301 , \12299 , \12300 );
xnor \U$11987 ( \12302 , \12301 , \9123 );
and \U$11988 ( \12303 , \12297 , \12302 );
and \U$11989 ( \12304 , \12293 , \12302 );
or \U$11990 ( \12305 , \12298 , \12303 , \12304 );
and \U$11991 ( \12306 , \12289 , \12305 );
and \U$11992 ( \12307 , \709 , \8896 );
and \U$11993 ( \12308 , \681 , \8894 );
nor \U$11994 ( \12309 , \12307 , \12308 );
xnor \U$11995 ( \12310 , \12309 , \8525 );
and \U$11996 ( \12311 , \863 , \8334 );
and \U$11997 ( \12312 , \789 , \8332 );
nor \U$11998 ( \12313 , \12311 , \12312 );
xnor \U$11999 ( \12314 , \12313 , \8016 );
and \U$12000 ( \12315 , \12310 , \12314 );
and \U$12001 ( \12316 , \988 , \7767 );
and \U$12002 ( \12317 , \925 , \7765 );
nor \U$12003 ( \12318 , \12316 , \12317 );
xnor \U$12004 ( \12319 , \12318 , \7518 );
and \U$12005 ( \12320 , \12314 , \12319 );
and \U$12006 ( \12321 , \12310 , \12319 );
or \U$12007 ( \12322 , \12315 , \12320 , \12321 );
and \U$12008 ( \12323 , \12305 , \12322 );
and \U$12009 ( \12324 , \12289 , \12322 );
or \U$12010 ( \12325 , \12306 , \12323 , \12324 );
and \U$12011 ( \12326 , \12273 , \12325 );
and \U$12012 ( \12327 , \4779 , \2300 );
and \U$12013 ( \12328 , \4771 , \2298 );
nor \U$12014 ( \12329 , \12327 , \12328 );
xnor \U$12015 ( \12330 , \12329 , \2163 );
and \U$12016 ( \12331 , \5253 , \2094 );
and \U$12017 ( \12332 , \5248 , \2092 );
nor \U$12018 ( \12333 , \12331 , \12332 );
xnor \U$12019 ( \12334 , \12333 , \1942 );
and \U$12020 ( \12335 , \12330 , \12334 );
and \U$12021 ( \12336 , \5776 , \1826 );
and \U$12022 ( \12337 , \5517 , \1824 );
nor \U$12023 ( \12338 , \12336 , \12337 );
xnor \U$12024 ( \12339 , \12338 , \1670 );
and \U$12025 ( \12340 , \12334 , \12339 );
and \U$12026 ( \12341 , \12330 , \12339 );
or \U$12027 ( \12342 , \12335 , \12340 , \12341 );
and \U$12028 ( \12343 , \8127 , \996 );
and \U$12029 ( \12344 , \7703 , \994 );
nor \U$12030 ( \12345 , \12343 , \12344 );
xnor \U$12031 ( \12346 , \12345 , \902 );
and \U$12032 ( \12347 , \8378 , \826 );
and \U$12033 ( \12348 , \8373 , \824 );
nor \U$12034 ( \12349 , \12347 , \12348 );
xnor \U$12035 ( \12350 , \12349 , \754 );
and \U$12036 ( \12351 , \12346 , \12350 );
and \U$12037 ( \12352 , \8981 , \692 );
and \U$12038 ( \12353 , \8697 , \690 );
nor \U$12039 ( \12354 , \12352 , \12353 );
xnor \U$12040 ( \12355 , \12354 , \649 );
and \U$12041 ( \12356 , \12350 , \12355 );
and \U$12042 ( \12357 , \12346 , \12355 );
or \U$12043 ( \12358 , \12351 , \12356 , \12357 );
and \U$12044 ( \12359 , \12342 , \12358 );
and \U$12045 ( \12360 , \6157 , \1554 );
and \U$12046 ( \12361 , \6148 , \1552 );
nor \U$12047 ( \12362 , \12360 , \12361 );
xnor \U$12048 ( \12363 , \12362 , \1441 );
and \U$12049 ( \12364 , \6702 , \1360 );
and \U$12050 ( \12365 , \6500 , \1358 );
nor \U$12051 ( \12366 , \12364 , \12365 );
xnor \U$12052 ( \12367 , \12366 , \1224 );
and \U$12053 ( \12368 , \12363 , \12367 );
and \U$12054 ( \12369 , \7177 , \1160 );
and \U$12055 ( \12370 , \7005 , \1158 );
nor \U$12056 ( \12371 , \12369 , \12370 );
xnor \U$12057 ( \12372 , \12371 , \1082 );
and \U$12058 ( \12373 , \12367 , \12372 );
and \U$12059 ( \12374 , \12363 , \12372 );
or \U$12060 ( \12375 , \12368 , \12373 , \12374 );
and \U$12061 ( \12376 , \12358 , \12375 );
and \U$12062 ( \12377 , \12342 , \12375 );
or \U$12063 ( \12378 , \12359 , \12376 , \12377 );
and \U$12064 ( \12379 , \12325 , \12378 );
and \U$12065 ( \12380 , \12273 , \12378 );
or \U$12066 ( \12381 , \12326 , \12379 , \12380 );
and \U$12067 ( \12382 , \12221 , \12381 );
xor \U$12068 ( \12383 , \11930 , \11934 );
xor \U$12069 ( \12384 , \12383 , \11939 );
xor \U$12070 ( \12385 , \11946 , \11950 );
xor \U$12071 ( \12386 , \12385 , \11955 );
and \U$12072 ( \12387 , \12384 , \12386 );
xor \U$12073 ( \12388 , \11963 , \11967 );
xor \U$12074 ( \12389 , \12388 , \341 );
and \U$12075 ( \12390 , \12386 , \12389 );
and \U$12076 ( \12391 , \12384 , \12389 );
or \U$12077 ( \12392 , \12387 , \12390 , \12391 );
xor \U$12078 ( \12393 , \11578 , \11582 );
xor \U$12079 ( \12394 , \12393 , \11587 );
and \U$12080 ( \12395 , \12392 , \12394 );
xor \U$12081 ( \12396 , \12088 , \12090 );
xor \U$12082 ( \12397 , \12396 , \12093 );
and \U$12083 ( \12398 , \12394 , \12397 );
and \U$12084 ( \12399 , \12392 , \12397 );
or \U$12085 ( \12400 , \12395 , \12398 , \12399 );
and \U$12086 ( \12401 , \12381 , \12400 );
and \U$12087 ( \12402 , \12221 , \12400 );
or \U$12088 ( \12403 , \12382 , \12401 , \12402 );
xor \U$12089 ( \12404 , \11890 , \11906 );
xor \U$12090 ( \12405 , \12404 , \11923 );
xor \U$12091 ( \12406 , \11942 , \11958 );
xor \U$12092 ( \12407 , \12406 , \11971 );
and \U$12093 ( \12408 , \12405 , \12407 );
xor \U$12094 ( \12409 , \11991 , \12007 );
xor \U$12095 ( \12410 , \12409 , \12024 );
and \U$12096 ( \12411 , \12407 , \12410 );
and \U$12097 ( \12412 , \12405 , \12410 );
or \U$12098 ( \12413 , \12408 , \12411 , \12412 );
xor \U$12099 ( \12414 , \12046 , \12053 );
xor \U$12100 ( \12415 , \12414 , \12058 );
xor \U$12101 ( \12416 , \12063 , \12065 );
xor \U$12102 ( \12417 , \12416 , \12068 );
and \U$12103 ( \12418 , \12415 , \12417 );
xor \U$12104 ( \12419 , \12074 , \12076 );
xor \U$12105 ( \12420 , \12419 , \12079 );
and \U$12106 ( \12421 , \12417 , \12420 );
and \U$12107 ( \12422 , \12415 , \12420 );
or \U$12108 ( \12423 , \12418 , \12421 , \12422 );
and \U$12109 ( \12424 , \12413 , \12423 );
xor \U$12110 ( \12425 , \11679 , \11695 );
xor \U$12111 ( \12426 , \12425 , \11712 );
and \U$12112 ( \12427 , \12423 , \12426 );
and \U$12113 ( \12428 , \12413 , \12426 );
or \U$12114 ( \12429 , \12424 , \12427 , \12428 );
and \U$12115 ( \12430 , \12403 , \12429 );
xor \U$12116 ( \12431 , \11574 , \11590 );
xor \U$12117 ( \12432 , \12431 , \11607 );
xor \U$12118 ( \12433 , \12109 , \12111 );
xor \U$12119 ( \12434 , \12433 , \12114 );
and \U$12120 ( \12435 , \12432 , \12434 );
xor \U$12121 ( \12436 , \12096 , \12098 );
xor \U$12122 ( \12437 , \12436 , \12101 );
and \U$12123 ( \12438 , \12434 , \12437 );
and \U$12124 ( \12439 , \12432 , \12437 );
or \U$12125 ( \12440 , \12435 , \12438 , \12439 );
and \U$12126 ( \12441 , \12429 , \12440 );
and \U$12127 ( \12442 , \12403 , \12440 );
or \U$12128 ( \12443 , \12430 , \12441 , \12442 );
xor \U$12129 ( \12444 , \12030 , \12085 );
xor \U$12130 ( \12445 , \12444 , \12104 );
xor \U$12131 ( \12446 , \12117 , \12119 );
xor \U$12132 ( \12447 , \12446 , \12122 );
and \U$12133 ( \12448 , \12445 , \12447 );
xor \U$12134 ( \12449 , \12128 , \12130 );
xor \U$12135 ( \12450 , \12449 , \12133 );
and \U$12136 ( \12451 , \12447 , \12450 );
and \U$12137 ( \12452 , \12445 , \12450 );
or \U$12138 ( \12453 , \12448 , \12451 , \12452 );
and \U$12139 ( \12454 , \12443 , \12453 );
xor \U$12140 ( \12455 , \11797 , \11807 );
xor \U$12141 ( \12456 , \12455 , \11810 );
and \U$12142 ( \12457 , \12453 , \12456 );
and \U$12143 ( \12458 , \12443 , \12456 );
or \U$12144 ( \12459 , \12454 , \12457 , \12458 );
xor \U$12145 ( \12460 , \11718 , \11766 );
xor \U$12146 ( \12461 , \12460 , \11784 );
xor \U$12147 ( \12462 , \12107 , \12125 );
xor \U$12148 ( \12463 , \12462 , \12136 );
and \U$12149 ( \12464 , \12461 , \12463 );
xor \U$12150 ( \12465 , \12141 , \12143 );
xor \U$12151 ( \12466 , \12465 , \12146 );
and \U$12152 ( \12467 , \12463 , \12466 );
and \U$12153 ( \12468 , \12461 , \12466 );
or \U$12154 ( \12469 , \12464 , \12467 , \12468 );
and \U$12155 ( \12470 , \12459 , \12469 );
xor \U$12156 ( \12471 , \11829 , \11831 );
xor \U$12157 ( \12472 , \12471 , \11834 );
and \U$12158 ( \12473 , \12469 , \12472 );
and \U$12159 ( \12474 , \12459 , \12472 );
or \U$12160 ( \12475 , \12470 , \12473 , \12474 );
xor \U$12161 ( \12476 , \11787 , \11813 );
xor \U$12162 ( \12477 , \12476 , \11824 );
xor \U$12163 ( \12478 , \12139 , \12149 );
xor \U$12164 ( \12479 , \12478 , \12152 );
and \U$12165 ( \12480 , \12477 , \12479 );
and \U$12166 ( \12481 , \12475 , \12480 );
xor \U$12167 ( \12482 , \12155 , \12157 );
xor \U$12168 ( \12483 , \12482 , \12160 );
and \U$12169 ( \12484 , \12480 , \12483 );
and \U$12170 ( \12485 , \12475 , \12483 );
or \U$12171 ( \12486 , \12481 , \12484 , \12485 );
and \U$12172 ( \12487 , \12174 , \12486 );
xor \U$12173 ( \12488 , \12174 , \12486 );
xor \U$12174 ( \12489 , \12475 , \12480 );
xor \U$12175 ( \12490 , \12489 , \12483 );
xor \U$12176 ( \12491 , \12225 , \12229 );
xor \U$12177 ( \12492 , \12491 , \12234 );
xor \U$12178 ( \12493 , \12330 , \12334 );
xor \U$12179 ( \12494 , \12493 , \12339 );
and \U$12180 ( \12495 , \12492 , \12494 );
xor \U$12181 ( \12496 , \12363 , \12367 );
xor \U$12182 ( \12497 , \12496 , \12372 );
and \U$12183 ( \12498 , \12494 , \12497 );
and \U$12184 ( \12499 , \12492 , \12497 );
or \U$12185 ( \12500 , \12495 , \12498 , \12499 );
and \U$12186 ( \12501 , \9550 , \692 );
and \U$12187 ( \12502 , \8981 , \690 );
nor \U$12188 ( \12503 , \12501 , \12502 );
xnor \U$12189 ( \12504 , \12503 , \649 );
and \U$12190 ( \12505 , \10161 , \579 );
and \U$12191 ( \12506 , \9558 , \577 );
nor \U$12192 ( \12507 , \12505 , \12506 );
xnor \U$12193 ( \12508 , \12507 , \530 );
and \U$12194 ( \12509 , \12504 , \12508 );
and \U$12195 ( \12510 , \10347 , \478 );
and \U$12196 ( \12511 , \10166 , \476 );
nor \U$12197 ( \12512 , \12510 , \12511 );
xnor \U$12198 ( \12513 , \12512 , \437 );
and \U$12199 ( \12514 , \12508 , \12513 );
and \U$12200 ( \12515 , \12504 , \12513 );
or \U$12201 ( \12516 , \12509 , \12514 , \12515 );
xor \U$12202 ( \12517 , \12346 , \12350 );
xor \U$12203 ( \12518 , \12517 , \12355 );
and \U$12204 ( \12519 , \12516 , \12518 );
xor \U$12205 ( \12520 , \12199 , \12203 );
xor \U$12206 ( \12521 , \12520 , \12208 );
and \U$12207 ( \12522 , \12518 , \12521 );
and \U$12208 ( \12523 , \12516 , \12521 );
or \U$12209 ( \12524 , \12519 , \12522 , \12523 );
and \U$12210 ( \12525 , \12500 , \12524 );
xor \U$12211 ( \12526 , \12277 , \12281 );
xor \U$12212 ( \12527 , \12526 , \12286 );
xor \U$12213 ( \12528 , \12241 , \12245 );
xor \U$12214 ( \12529 , \12528 , \12250 );
and \U$12215 ( \12530 , \12527 , \12529 );
xor \U$12216 ( \12531 , \12258 , \12262 );
xor \U$12217 ( \12532 , \12531 , \12267 );
and \U$12218 ( \12533 , \12529 , \12532 );
and \U$12219 ( \12534 , \12527 , \12532 );
or \U$12220 ( \12535 , \12530 , \12533 , \12534 );
and \U$12221 ( \12536 , \12524 , \12535 );
and \U$12222 ( \12537 , \12500 , \12535 );
or \U$12223 ( \12538 , \12525 , \12536 , \12537 );
and \U$12224 ( \12539 , \1186 , \7767 );
and \U$12225 ( \12540 , \988 , \7765 );
nor \U$12226 ( \12541 , \12539 , \12540 );
xnor \U$12227 ( \12542 , \12541 , \7518 );
and \U$12228 ( \12543 , \1379 , \7238 );
and \U$12229 ( \12544 , \1274 , \7236 );
nor \U$12230 ( \12545 , \12543 , \12544 );
xnor \U$12231 ( \12546 , \12545 , \6978 );
and \U$12232 ( \12547 , \12542 , \12546 );
and \U$12233 ( \12548 , \1500 , \6744 );
and \U$12234 ( \12549 , \1384 , \6742 );
nor \U$12235 ( \12550 , \12548 , \12549 );
xnor \U$12236 ( \12551 , \12550 , \6429 );
and \U$12237 ( \12552 , \12546 , \12551 );
and \U$12238 ( \12553 , \12542 , \12551 );
or \U$12239 ( \12554 , \12547 , \12552 , \12553 );
and \U$12240 ( \12555 , \494 , \10814 );
and \U$12241 ( \12556 , \425 , \10811 );
nor \U$12242 ( \12557 , \12555 , \12556 );
xnor \U$12243 ( \12558 , \12557 , \9759 );
and \U$12244 ( \12559 , \553 , \10001 );
and \U$12245 ( \12560 , \499 , \9999 );
nor \U$12246 ( \12561 , \12559 , \12560 );
xnor \U$12247 ( \12562 , \12561 , \9762 );
and \U$12248 ( \12563 , \12558 , \12562 );
and \U$12249 ( \12564 , \12562 , \378 );
and \U$12250 ( \12565 , \12558 , \378 );
or \U$12251 ( \12566 , \12563 , \12564 , \12565 );
and \U$12252 ( \12567 , \12554 , \12566 );
and \U$12253 ( \12568 , \681 , \9433 );
and \U$12254 ( \12569 , \604 , \9431 );
nor \U$12255 ( \12570 , \12568 , \12569 );
xnor \U$12256 ( \12571 , \12570 , \9123 );
and \U$12257 ( \12572 , \789 , \8896 );
and \U$12258 ( \12573 , \709 , \8894 );
nor \U$12259 ( \12574 , \12572 , \12573 );
xnor \U$12260 ( \12575 , \12574 , \8525 );
and \U$12261 ( \12576 , \12571 , \12575 );
and \U$12262 ( \12577 , \925 , \8334 );
and \U$12263 ( \12578 , \863 , \8332 );
nor \U$12264 ( \12579 , \12577 , \12578 );
xnor \U$12265 ( \12580 , \12579 , \8016 );
and \U$12266 ( \12581 , \12575 , \12580 );
and \U$12267 ( \12582 , \12571 , \12580 );
or \U$12268 ( \12583 , \12576 , \12581 , \12582 );
and \U$12269 ( \12584 , \12566 , \12583 );
and \U$12270 ( \12585 , \12554 , \12583 );
or \U$12271 ( \12586 , \12567 , \12584 , \12585 );
and \U$12272 ( \12587 , \3681 , \3637 );
and \U$12273 ( \12588 , \3264 , \3635 );
nor \U$12274 ( \12589 , \12587 , \12588 );
xnor \U$12275 ( \12590 , \12589 , \3450 );
and \U$12276 ( \12591 , \4011 , \3324 );
and \U$12277 ( \12592 , \3889 , \3322 );
nor \U$12278 ( \12593 , \12591 , \12592 );
xnor \U$12279 ( \12594 , \12593 , \3119 );
and \U$12280 ( \12595 , \12590 , \12594 );
and \U$12281 ( \12596 , \4272 , \2918 );
and \U$12282 ( \12597 , \4016 , \2916 );
nor \U$12283 ( \12598 , \12596 , \12597 );
xnor \U$12284 ( \12599 , \12598 , \2769 );
and \U$12285 ( \12600 , \12594 , \12599 );
and \U$12286 ( \12601 , \12590 , \12599 );
or \U$12287 ( \12602 , \12595 , \12600 , \12601 );
and \U$12288 ( \12603 , \2641 , \4806 );
and \U$12289 ( \12604 , \2377 , \4804 );
nor \U$12290 ( \12605 , \12603 , \12604 );
xnor \U$12291 ( \12606 , \12605 , \4574 );
and \U$12292 ( \12607 , \2840 , \4355 );
and \U$12293 ( \12608 , \2666 , \4353 );
nor \U$12294 ( \12609 , \12607 , \12608 );
xnor \U$12295 ( \12610 , \12609 , \4212 );
and \U$12296 ( \12611 , \12606 , \12610 );
and \U$12297 ( \12612 , \3145 , \4032 );
and \U$12298 ( \12613 , \3007 , \4030 );
nor \U$12299 ( \12614 , \12612 , \12613 );
xnor \U$12300 ( \12615 , \12614 , \3786 );
and \U$12301 ( \12616 , \12610 , \12615 );
and \U$12302 ( \12617 , \12606 , \12615 );
or \U$12303 ( \12618 , \12611 , \12616 , \12617 );
and \U$12304 ( \12619 , \12602 , \12618 );
and \U$12305 ( \12620 , \1791 , \6235 );
and \U$12306 ( \12621 , \1615 , \6233 );
nor \U$12307 ( \12622 , \12620 , \12621 );
xnor \U$12308 ( \12623 , \12622 , \5895 );
and \U$12309 ( \12624 , \2042 , \5646 );
and \U$12310 ( \12625 , \1799 , \5644 );
nor \U$12311 ( \12626 , \12624 , \12625 );
xnor \U$12312 ( \12627 , \12626 , \5405 );
and \U$12313 ( \12628 , \12623 , \12627 );
and \U$12314 ( \12629 , \2233 , \5180 );
and \U$12315 ( \12630 , \2047 , \5178 );
nor \U$12316 ( \12631 , \12629 , \12630 );
xnor \U$12317 ( \12632 , \12631 , \4992 );
and \U$12318 ( \12633 , \12627 , \12632 );
and \U$12319 ( \12634 , \12623 , \12632 );
or \U$12320 ( \12635 , \12628 , \12633 , \12634 );
and \U$12321 ( \12636 , \12618 , \12635 );
and \U$12322 ( \12637 , \12602 , \12635 );
or \U$12323 ( \12638 , \12619 , \12636 , \12637 );
and \U$12324 ( \12639 , \12586 , \12638 );
and \U$12325 ( \12640 , \4771 , \2596 );
and \U$12326 ( \12641 , \4469 , \2594 );
nor \U$12327 ( \12642 , \12640 , \12641 );
xnor \U$12328 ( \12643 , \12642 , \2454 );
and \U$12329 ( \12644 , \5248 , \2300 );
and \U$12330 ( \12645 , \4779 , \2298 );
nor \U$12331 ( \12646 , \12644 , \12645 );
xnor \U$12332 ( \12647 , \12646 , \2163 );
and \U$12333 ( \12648 , \12643 , \12647 );
and \U$12334 ( \12649 , \5517 , \2094 );
and \U$12335 ( \12650 , \5253 , \2092 );
nor \U$12336 ( \12651 , \12649 , \12650 );
xnor \U$12337 ( \12652 , \12651 , \1942 );
and \U$12338 ( \12653 , \12647 , \12652 );
and \U$12339 ( \12654 , \12643 , \12652 );
or \U$12340 ( \12655 , \12648 , \12653 , \12654 );
and \U$12341 ( \12656 , \6148 , \1826 );
and \U$12342 ( \12657 , \5776 , \1824 );
nor \U$12343 ( \12658 , \12656 , \12657 );
xnor \U$12344 ( \12659 , \12658 , \1670 );
and \U$12345 ( \12660 , \6500 , \1554 );
and \U$12346 ( \12661 , \6157 , \1552 );
nor \U$12347 ( \12662 , \12660 , \12661 );
xnor \U$12348 ( \12663 , \12662 , \1441 );
and \U$12349 ( \12664 , \12659 , \12663 );
and \U$12350 ( \12665 , \7005 , \1360 );
and \U$12351 ( \12666 , \6702 , \1358 );
nor \U$12352 ( \12667 , \12665 , \12666 );
xnor \U$12353 ( \12668 , \12667 , \1224 );
and \U$12354 ( \12669 , \12663 , \12668 );
and \U$12355 ( \12670 , \12659 , \12668 );
or \U$12356 ( \12671 , \12664 , \12669 , \12670 );
and \U$12357 ( \12672 , \12655 , \12671 );
and \U$12358 ( \12673 , \7703 , \1160 );
and \U$12359 ( \12674 , \7177 , \1158 );
nor \U$12360 ( \12675 , \12673 , \12674 );
xnor \U$12361 ( \12676 , \12675 , \1082 );
and \U$12362 ( \12677 , \8373 , \996 );
and \U$12363 ( \12678 , \8127 , \994 );
nor \U$12364 ( \12679 , \12677 , \12678 );
xnor \U$12365 ( \12680 , \12679 , \902 );
and \U$12366 ( \12681 , \12676 , \12680 );
and \U$12367 ( \12682 , \8697 , \826 );
and \U$12368 ( \12683 , \8378 , \824 );
nor \U$12369 ( \12684 , \12682 , \12683 );
xnor \U$12370 ( \12685 , \12684 , \754 );
and \U$12371 ( \12686 , \12680 , \12685 );
and \U$12372 ( \12687 , \12676 , \12685 );
or \U$12373 ( \12688 , \12681 , \12686 , \12687 );
and \U$12374 ( \12689 , \12671 , \12688 );
and \U$12375 ( \12690 , \12655 , \12688 );
or \U$12376 ( \12691 , \12672 , \12689 , \12690 );
and \U$12377 ( \12692 , \12638 , \12691 );
and \U$12378 ( \12693 , \12586 , \12691 );
or \U$12379 ( \12694 , \12639 , \12692 , \12693 );
and \U$12380 ( \12695 , \12538 , \12694 );
xor \U$12381 ( \12696 , \12384 , \12386 );
xor \U$12382 ( \12697 , \12696 , \12389 );
xor \U$12383 ( \12698 , \12176 , \12178 );
xor \U$12384 ( \12699 , \12698 , \12181 );
and \U$12385 ( \12700 , \12697 , \12699 );
xor \U$12386 ( \12701 , \12186 , \12188 );
xor \U$12387 ( \12702 , \12701 , \12191 );
and \U$12388 ( \12703 , \12699 , \12702 );
and \U$12389 ( \12704 , \12697 , \12702 );
or \U$12390 ( \12705 , \12700 , \12703 , \12704 );
and \U$12391 ( \12706 , \12694 , \12705 );
and \U$12392 ( \12707 , \12538 , \12705 );
or \U$12393 ( \12708 , \12695 , \12706 , \12707 );
xor \U$12394 ( \12709 , \12237 , \12253 );
xor \U$12395 ( \12710 , \12709 , \12270 );
xor \U$12396 ( \12711 , \12342 , \12358 );
xor \U$12397 ( \12712 , \12711 , \12375 );
and \U$12398 ( \12713 , \12710 , \12712 );
xor \U$12399 ( \12714 , \12211 , \12213 );
xor \U$12400 ( \12715 , \12714 , \12215 );
and \U$12401 ( \12716 , \12712 , \12715 );
and \U$12402 ( \12717 , \12710 , \12715 );
or \U$12403 ( \12718 , \12713 , \12716 , \12717 );
xor \U$12404 ( \12719 , \12405 , \12407 );
xor \U$12405 ( \12720 , \12719 , \12410 );
and \U$12406 ( \12721 , \12718 , \12720 );
xor \U$12407 ( \12722 , \12415 , \12417 );
xor \U$12408 ( \12723 , \12722 , \12420 );
and \U$12409 ( \12724 , \12720 , \12723 );
and \U$12410 ( \12725 , \12718 , \12723 );
or \U$12411 ( \12726 , \12721 , \12724 , \12725 );
and \U$12412 ( \12727 , \12708 , \12726 );
xor \U$12413 ( \12728 , \12184 , \12194 );
xor \U$12414 ( \12729 , \12728 , \12218 );
xor \U$12415 ( \12730 , \12273 , \12325 );
xor \U$12416 ( \12731 , \12730 , \12378 );
and \U$12417 ( \12732 , \12729 , \12731 );
xor \U$12418 ( \12733 , \12392 , \12394 );
xor \U$12419 ( \12734 , \12733 , \12397 );
and \U$12420 ( \12735 , \12731 , \12734 );
and \U$12421 ( \12736 , \12729 , \12734 );
or \U$12422 ( \12737 , \12732 , \12735 , \12736 );
and \U$12423 ( \12738 , \12726 , \12737 );
and \U$12424 ( \12739 , \12708 , \12737 );
or \U$12425 ( \12740 , \12727 , \12738 , \12739 );
xor \U$12426 ( \12741 , \11926 , \11974 );
xor \U$12427 ( \12742 , \12741 , \12027 );
xor \U$12428 ( \12743 , \12061 , \12071 );
xor \U$12429 ( \12744 , \12743 , \12082 );
and \U$12430 ( \12745 , \12742 , \12744 );
xor \U$12431 ( \12746 , \12432 , \12434 );
xor \U$12432 ( \12747 , \12746 , \12437 );
and \U$12433 ( \12748 , \12744 , \12747 );
and \U$12434 ( \12749 , \12742 , \12747 );
or \U$12435 ( \12750 , \12745 , \12748 , \12749 );
and \U$12436 ( \12751 , \12740 , \12750 );
xor \U$12437 ( \12752 , \12445 , \12447 );
xor \U$12438 ( \12753 , \12752 , \12450 );
and \U$12439 ( \12754 , \12750 , \12753 );
and \U$12440 ( \12755 , \12740 , \12753 );
or \U$12441 ( \12756 , \12751 , \12754 , \12755 );
xor \U$12442 ( \12757 , \12443 , \12453 );
xor \U$12443 ( \12758 , \12757 , \12456 );
and \U$12444 ( \12759 , \12756 , \12758 );
xor \U$12445 ( \12760 , \12461 , \12463 );
xor \U$12446 ( \12761 , \12760 , \12466 );
and \U$12447 ( \12762 , \12758 , \12761 );
and \U$12448 ( \12763 , \12756 , \12761 );
or \U$12449 ( \12764 , \12759 , \12762 , \12763 );
xor \U$12450 ( \12765 , \12459 , \12469 );
xor \U$12451 ( \12766 , \12765 , \12472 );
and \U$12452 ( \12767 , \12764 , \12766 );
xor \U$12453 ( \12768 , \12477 , \12479 );
and \U$12454 ( \12769 , \12766 , \12768 );
and \U$12455 ( \12770 , \12764 , \12768 );
or \U$12456 ( \12771 , \12767 , \12769 , \12770 );
and \U$12457 ( \12772 , \12490 , \12771 );
xor \U$12458 ( \12773 , \12490 , \12771 );
xor \U$12459 ( \12774 , \12764 , \12766 );
xor \U$12460 ( \12775 , \12774 , \12768 );
and \U$12461 ( \12776 , \3007 , \4355 );
and \U$12462 ( \12777 , \2840 , \4353 );
nor \U$12463 ( \12778 , \12776 , \12777 );
xnor \U$12464 ( \12779 , \12778 , \4212 );
and \U$12465 ( \12780 , \3264 , \4032 );
and \U$12466 ( \12781 , \3145 , \4030 );
nor \U$12467 ( \12782 , \12780 , \12781 );
xnor \U$12468 ( \12783 , \12782 , \3786 );
and \U$12469 ( \12784 , \12779 , \12783 );
and \U$12470 ( \12785 , \3889 , \3637 );
and \U$12471 ( \12786 , \3681 , \3635 );
nor \U$12472 ( \12787 , \12785 , \12786 );
xnor \U$12473 ( \12788 , \12787 , \3450 );
and \U$12474 ( \12789 , \12783 , \12788 );
and \U$12475 ( \12790 , \12779 , \12788 );
or \U$12476 ( \12791 , \12784 , \12789 , \12790 );
and \U$12477 ( \12792 , \4016 , \3324 );
and \U$12478 ( \12793 , \4011 , \3322 );
nor \U$12479 ( \12794 , \12792 , \12793 );
xnor \U$12480 ( \12795 , \12794 , \3119 );
and \U$12481 ( \12796 , \4469 , \2918 );
and \U$12482 ( \12797 , \4272 , \2916 );
nor \U$12483 ( \12798 , \12796 , \12797 );
xnor \U$12484 ( \12799 , \12798 , \2769 );
and \U$12485 ( \12800 , \12795 , \12799 );
and \U$12486 ( \12801 , \4779 , \2596 );
and \U$12487 ( \12802 , \4771 , \2594 );
nor \U$12488 ( \12803 , \12801 , \12802 );
xnor \U$12489 ( \12804 , \12803 , \2454 );
and \U$12490 ( \12805 , \12799 , \12804 );
and \U$12491 ( \12806 , \12795 , \12804 );
or \U$12492 ( \12807 , \12800 , \12805 , \12806 );
and \U$12493 ( \12808 , \12791 , \12807 );
and \U$12494 ( \12809 , \2047 , \5646 );
and \U$12495 ( \12810 , \2042 , \5644 );
nor \U$12496 ( \12811 , \12809 , \12810 );
xnor \U$12497 ( \12812 , \12811 , \5405 );
and \U$12498 ( \12813 , \2377 , \5180 );
and \U$12499 ( \12814 , \2233 , \5178 );
nor \U$12500 ( \12815 , \12813 , \12814 );
xnor \U$12501 ( \12816 , \12815 , \4992 );
and \U$12502 ( \12817 , \12812 , \12816 );
and \U$12503 ( \12818 , \2666 , \4806 );
and \U$12504 ( \12819 , \2641 , \4804 );
nor \U$12505 ( \12820 , \12818 , \12819 );
xnor \U$12506 ( \12821 , \12820 , \4574 );
and \U$12507 ( \12822 , \12816 , \12821 );
and \U$12508 ( \12823 , \12812 , \12821 );
or \U$12509 ( \12824 , \12817 , \12822 , \12823 );
and \U$12510 ( \12825 , \12807 , \12824 );
and \U$12511 ( \12826 , \12791 , \12824 );
or \U$12512 ( \12827 , \12808 , \12825 , \12826 );
and \U$12513 ( \12828 , \6702 , \1554 );
and \U$12514 ( \12829 , \6500 , \1552 );
nor \U$12515 ( \12830 , \12828 , \12829 );
xnor \U$12516 ( \12831 , \12830 , \1441 );
and \U$12517 ( \12832 , \7177 , \1360 );
and \U$12518 ( \12833 , \7005 , \1358 );
nor \U$12519 ( \12834 , \12832 , \12833 );
xnor \U$12520 ( \12835 , \12834 , \1224 );
and \U$12521 ( \12836 , \12831 , \12835 );
and \U$12522 ( \12837 , \8127 , \1160 );
and \U$12523 ( \12838 , \7703 , \1158 );
nor \U$12524 ( \12839 , \12837 , \12838 );
xnor \U$12525 ( \12840 , \12839 , \1082 );
and \U$12526 ( \12841 , \12835 , \12840 );
and \U$12527 ( \12842 , \12831 , \12840 );
or \U$12528 ( \12843 , \12836 , \12841 , \12842 );
and \U$12529 ( \12844 , \8378 , \996 );
and \U$12530 ( \12845 , \8373 , \994 );
nor \U$12531 ( \12846 , \12844 , \12845 );
xnor \U$12532 ( \12847 , \12846 , \902 );
and \U$12533 ( \12848 , \8981 , \826 );
and \U$12534 ( \12849 , \8697 , \824 );
nor \U$12535 ( \12850 , \12848 , \12849 );
xnor \U$12536 ( \12851 , \12850 , \754 );
and \U$12537 ( \12852 , \12847 , \12851 );
and \U$12538 ( \12853 , \9558 , \692 );
and \U$12539 ( \12854 , \9550 , \690 );
nor \U$12540 ( \12855 , \12853 , \12854 );
xnor \U$12541 ( \12856 , \12855 , \649 );
and \U$12542 ( \12857 , \12851 , \12856 );
and \U$12543 ( \12858 , \12847 , \12856 );
or \U$12544 ( \12859 , \12852 , \12857 , \12858 );
and \U$12545 ( \12860 , \12843 , \12859 );
and \U$12546 ( \12861 , \5253 , \2300 );
and \U$12547 ( \12862 , \5248 , \2298 );
nor \U$12548 ( \12863 , \12861 , \12862 );
xnor \U$12549 ( \12864 , \12863 , \2163 );
and \U$12550 ( \12865 , \5776 , \2094 );
and \U$12551 ( \12866 , \5517 , \2092 );
nor \U$12552 ( \12867 , \12865 , \12866 );
xnor \U$12553 ( \12868 , \12867 , \1942 );
and \U$12554 ( \12869 , \12864 , \12868 );
and \U$12555 ( \12870 , \6157 , \1826 );
and \U$12556 ( \12871 , \6148 , \1824 );
nor \U$12557 ( \12872 , \12870 , \12871 );
xnor \U$12558 ( \12873 , \12872 , \1670 );
and \U$12559 ( \12874 , \12868 , \12873 );
and \U$12560 ( \12875 , \12864 , \12873 );
or \U$12561 ( \12876 , \12869 , \12874 , \12875 );
and \U$12562 ( \12877 , \12859 , \12876 );
and \U$12563 ( \12878 , \12843 , \12876 );
or \U$12564 ( \12879 , \12860 , \12877 , \12878 );
and \U$12565 ( \12880 , \12827 , \12879 );
and \U$12566 ( \12881 , \499 , \10814 );
and \U$12567 ( \12882 , \494 , \10811 );
nor \U$12568 ( \12883 , \12881 , \12882 );
xnor \U$12569 ( \12884 , \12883 , \9759 );
and \U$12570 ( \12885 , \604 , \10001 );
and \U$12571 ( \12886 , \553 , \9999 );
nor \U$12572 ( \12887 , \12885 , \12886 );
xnor \U$12573 ( \12888 , \12887 , \9762 );
and \U$12574 ( \12889 , \12884 , \12888 );
and \U$12575 ( \12890 , \709 , \9433 );
and \U$12576 ( \12891 , \681 , \9431 );
nor \U$12577 ( \12892 , \12890 , \12891 );
xnor \U$12578 ( \12893 , \12892 , \9123 );
and \U$12579 ( \12894 , \12888 , \12893 );
and \U$12580 ( \12895 , \12884 , \12893 );
or \U$12581 ( \12896 , \12889 , \12894 , \12895 );
and \U$12582 ( \12897 , \863 , \8896 );
and \U$12583 ( \12898 , \789 , \8894 );
nor \U$12584 ( \12899 , \12897 , \12898 );
xnor \U$12585 ( \12900 , \12899 , \8525 );
and \U$12586 ( \12901 , \988 , \8334 );
and \U$12587 ( \12902 , \925 , \8332 );
nor \U$12588 ( \12903 , \12901 , \12902 );
xnor \U$12589 ( \12904 , \12903 , \8016 );
and \U$12590 ( \12905 , \12900 , \12904 );
and \U$12591 ( \12906 , \1274 , \7767 );
and \U$12592 ( \12907 , \1186 , \7765 );
nor \U$12593 ( \12908 , \12906 , \12907 );
xnor \U$12594 ( \12909 , \12908 , \7518 );
and \U$12595 ( \12910 , \12904 , \12909 );
and \U$12596 ( \12911 , \12900 , \12909 );
or \U$12597 ( \12912 , \12905 , \12910 , \12911 );
and \U$12598 ( \12913 , \12896 , \12912 );
and \U$12599 ( \12914 , \1384 , \7238 );
and \U$12600 ( \12915 , \1379 , \7236 );
nor \U$12601 ( \12916 , \12914 , \12915 );
xnor \U$12602 ( \12917 , \12916 , \6978 );
and \U$12603 ( \12918 , \1615 , \6744 );
and \U$12604 ( \12919 , \1500 , \6742 );
nor \U$12605 ( \12920 , \12918 , \12919 );
xnor \U$12606 ( \12921 , \12920 , \6429 );
and \U$12607 ( \12922 , \12917 , \12921 );
and \U$12608 ( \12923 , \1799 , \6235 );
and \U$12609 ( \12924 , \1791 , \6233 );
nor \U$12610 ( \12925 , \12923 , \12924 );
xnor \U$12611 ( \12926 , \12925 , \5895 );
and \U$12612 ( \12927 , \12921 , \12926 );
and \U$12613 ( \12928 , \12917 , \12926 );
or \U$12614 ( \12929 , \12922 , \12927 , \12928 );
and \U$12615 ( \12930 , \12912 , \12929 );
and \U$12616 ( \12931 , \12896 , \12929 );
or \U$12617 ( \12932 , \12913 , \12930 , \12931 );
and \U$12618 ( \12933 , \12879 , \12932 );
and \U$12619 ( \12934 , \12827 , \12932 );
or \U$12620 ( \12935 , \12880 , \12933 , \12934 );
xor \U$12621 ( \12936 , \12542 , \12546 );
xor \U$12622 ( \12937 , \12936 , \12551 );
xor \U$12623 ( \12938 , \12606 , \12610 );
xor \U$12624 ( \12939 , \12938 , \12615 );
and \U$12625 ( \12940 , \12937 , \12939 );
xor \U$12626 ( \12941 , \12623 , \12627 );
xor \U$12627 ( \12942 , \12941 , \12632 );
and \U$12628 ( \12943 , \12939 , \12942 );
and \U$12629 ( \12944 , \12937 , \12942 );
or \U$12630 ( \12945 , \12940 , \12943 , \12944 );
xor \U$12631 ( \12946 , \12590 , \12594 );
xor \U$12632 ( \12947 , \12946 , \12599 );
xor \U$12633 ( \12948 , \12643 , \12647 );
xor \U$12634 ( \12949 , \12948 , \12652 );
and \U$12635 ( \12950 , \12947 , \12949 );
xor \U$12636 ( \12951 , \12659 , \12663 );
xor \U$12637 ( \12952 , \12951 , \12668 );
and \U$12638 ( \12953 , \12949 , \12952 );
and \U$12639 ( \12954 , \12947 , \12952 );
or \U$12640 ( \12955 , \12950 , \12953 , \12954 );
and \U$12641 ( \12956 , \12945 , \12955 );
nand \U$12642 ( \12957 , \10967 , \406 );
xnor \U$12643 ( \12958 , \12957 , \378 );
xor \U$12644 ( \12959 , \12676 , \12680 );
xor \U$12645 ( \12960 , \12959 , \12685 );
and \U$12646 ( \12961 , \12958 , \12960 );
xor \U$12647 ( \12962 , \12504 , \12508 );
xor \U$12648 ( \12963 , \12962 , \12513 );
and \U$12649 ( \12964 , \12960 , \12963 );
and \U$12650 ( \12965 , \12958 , \12963 );
or \U$12651 ( \12966 , \12961 , \12964 , \12965 );
and \U$12652 ( \12967 , \12955 , \12966 );
and \U$12653 ( \12968 , \12945 , \12966 );
or \U$12654 ( \12969 , \12956 , \12967 , \12968 );
and \U$12655 ( \12970 , \12935 , \12969 );
xor \U$12656 ( \12971 , \12293 , \12297 );
xor \U$12657 ( \12972 , \12971 , \12302 );
xor \U$12658 ( \12973 , \12310 , \12314 );
xor \U$12659 ( \12974 , \12973 , \12319 );
and \U$12660 ( \12975 , \12972 , \12974 );
xor \U$12661 ( \12976 , \12527 , \12529 );
xor \U$12662 ( \12977 , \12976 , \12532 );
and \U$12663 ( \12978 , \12974 , \12977 );
and \U$12664 ( \12979 , \12972 , \12977 );
or \U$12665 ( \12980 , \12975 , \12978 , \12979 );
and \U$12666 ( \12981 , \12969 , \12980 );
and \U$12667 ( \12982 , \12935 , \12980 );
or \U$12668 ( \12983 , \12970 , \12981 , \12982 );
xor \U$12669 ( \12984 , \12500 , \12524 );
xor \U$12670 ( \12985 , \12984 , \12535 );
xor \U$12671 ( \12986 , \12586 , \12638 );
xor \U$12672 ( \12987 , \12986 , \12691 );
and \U$12673 ( \12988 , \12985 , \12987 );
xor \U$12674 ( \12989 , \12697 , \12699 );
xor \U$12675 ( \12990 , \12989 , \12702 );
and \U$12676 ( \12991 , \12987 , \12990 );
and \U$12677 ( \12992 , \12985 , \12990 );
or \U$12678 ( \12993 , \12988 , \12991 , \12992 );
and \U$12679 ( \12994 , \12983 , \12993 );
xor \U$12680 ( \12995 , \12655 , \12671 );
xor \U$12681 ( \12996 , \12995 , \12688 );
xor \U$12682 ( \12997 , \12492 , \12494 );
xor \U$12683 ( \12998 , \12997 , \12497 );
and \U$12684 ( \12999 , \12996 , \12998 );
xor \U$12685 ( \13000 , \12516 , \12518 );
xor \U$12686 ( \13001 , \13000 , \12521 );
and \U$12687 ( \13002 , \12998 , \13001 );
and \U$12688 ( \13003 , \12996 , \13001 );
or \U$12689 ( \13004 , \12999 , \13002 , \13003 );
xor \U$12690 ( \13005 , \12289 , \12305 );
xor \U$12691 ( \13006 , \13005 , \12322 );
and \U$12692 ( \13007 , \13004 , \13006 );
xor \U$12693 ( \13008 , \12710 , \12712 );
xor \U$12694 ( \13009 , \13008 , \12715 );
and \U$12695 ( \13010 , \13006 , \13009 );
and \U$12696 ( \13011 , \13004 , \13009 );
or \U$12697 ( \13012 , \13007 , \13010 , \13011 );
and \U$12698 ( \13013 , \12993 , \13012 );
and \U$12699 ( \13014 , \12983 , \13012 );
or \U$12700 ( \13015 , \12994 , \13013 , \13014 );
xor \U$12701 ( \13016 , \12538 , \12694 );
xor \U$12702 ( \13017 , \13016 , \12705 );
xor \U$12703 ( \13018 , \12718 , \12720 );
xor \U$12704 ( \13019 , \13018 , \12723 );
and \U$12705 ( \13020 , \13017 , \13019 );
xor \U$12706 ( \13021 , \12729 , \12731 );
xor \U$12707 ( \13022 , \13021 , \12734 );
and \U$12708 ( \13023 , \13019 , \13022 );
and \U$12709 ( \13024 , \13017 , \13022 );
or \U$12710 ( \13025 , \13020 , \13023 , \13024 );
and \U$12711 ( \13026 , \13015 , \13025 );
xor \U$12712 ( \13027 , \12413 , \12423 );
xor \U$12713 ( \13028 , \13027 , \12426 );
and \U$12714 ( \13029 , \13025 , \13028 );
and \U$12715 ( \13030 , \13015 , \13028 );
or \U$12716 ( \13031 , \13026 , \13029 , \13030 );
xor \U$12717 ( \13032 , \12221 , \12381 );
xor \U$12718 ( \13033 , \13032 , \12400 );
xor \U$12719 ( \13034 , \12708 , \12726 );
xor \U$12720 ( \13035 , \13034 , \12737 );
and \U$12721 ( \13036 , \13033 , \13035 );
xor \U$12722 ( \13037 , \12742 , \12744 );
xor \U$12723 ( \13038 , \13037 , \12747 );
and \U$12724 ( \13039 , \13035 , \13038 );
and \U$12725 ( \13040 , \13033 , \13038 );
or \U$12726 ( \13041 , \13036 , \13039 , \13040 );
and \U$12727 ( \13042 , \13031 , \13041 );
xor \U$12728 ( \13043 , \12403 , \12429 );
xor \U$12729 ( \13044 , \13043 , \12440 );
and \U$12730 ( \13045 , \13041 , \13044 );
and \U$12731 ( \13046 , \13031 , \13044 );
or \U$12732 ( \13047 , \13042 , \13045 , \13046 );
xor \U$12733 ( \13048 , \12756 , \12758 );
xor \U$12734 ( \13049 , \13048 , \12761 );
and \U$12735 ( \13050 , \13047 , \13049 );
and \U$12736 ( \13051 , \12775 , \13050 );
xor \U$12737 ( \13052 , \12775 , \13050 );
xor \U$12738 ( \13053 , \13047 , \13049 );
and \U$12739 ( \13054 , \10161 , \692 );
and \U$12740 ( \13055 , \9558 , \690 );
nor \U$12741 ( \13056 , \13054 , \13055 );
xnor \U$12742 ( \13057 , \13056 , \649 );
and \U$12743 ( \13058 , \10347 , \579 );
and \U$12744 ( \13059 , \10166 , \577 );
nor \U$12745 ( \13060 , \13058 , \13059 );
xnor \U$12746 ( \13061 , \13060 , \530 );
and \U$12747 ( \13062 , \13057 , \13061 );
nand \U$12748 ( \13063 , \10967 , \476 );
xnor \U$12749 ( \13064 , \13063 , \437 );
and \U$12750 ( \13065 , \13061 , \13064 );
and \U$12751 ( \13066 , \13057 , \13064 );
or \U$12752 ( \13067 , \13062 , \13065 , \13066 );
and \U$12753 ( \13068 , \10166 , \579 );
and \U$12754 ( \13069 , \10161 , \577 );
nor \U$12755 ( \13070 , \13068 , \13069 );
xnor \U$12756 ( \13071 , \13070 , \530 );
and \U$12757 ( \13072 , \13067 , \13071 );
and \U$12758 ( \13073 , \10967 , \478 );
and \U$12759 ( \13074 , \10347 , \476 );
nor \U$12760 ( \13075 , \13073 , \13074 );
xnor \U$12761 ( \13076 , \13075 , \437 );
and \U$12762 ( \13077 , \13071 , \13076 );
and \U$12763 ( \13078 , \13067 , \13076 );
or \U$12764 ( \13079 , \13072 , \13077 , \13078 );
xor \U$12765 ( \13080 , \12831 , \12835 );
xor \U$12766 ( \13081 , \13080 , \12840 );
xor \U$12767 ( \13082 , \12847 , \12851 );
xor \U$12768 ( \13083 , \13082 , \12856 );
and \U$12769 ( \13084 , \13081 , \13083 );
xor \U$12770 ( \13085 , \12864 , \12868 );
xor \U$12771 ( \13086 , \13085 , \12873 );
and \U$12772 ( \13087 , \13083 , \13086 );
and \U$12773 ( \13088 , \13081 , \13086 );
or \U$12774 ( \13089 , \13084 , \13087 , \13088 );
and \U$12775 ( \13090 , \13079 , \13089 );
xor \U$12776 ( \13091 , \12779 , \12783 );
xor \U$12777 ( \13092 , \13091 , \12788 );
xor \U$12778 ( \13093 , \12795 , \12799 );
xor \U$12779 ( \13094 , \13093 , \12804 );
and \U$12780 ( \13095 , \13092 , \13094 );
xor \U$12781 ( \13096 , \12812 , \12816 );
xor \U$12782 ( \13097 , \13096 , \12821 );
and \U$12783 ( \13098 , \13094 , \13097 );
and \U$12784 ( \13099 , \13092 , \13097 );
or \U$12785 ( \13100 , \13095 , \13098 , \13099 );
and \U$12786 ( \13101 , \13089 , \13100 );
and \U$12787 ( \13102 , \13079 , \13100 );
or \U$12788 ( \13103 , \13090 , \13101 , \13102 );
and \U$12789 ( \13104 , \789 , \9433 );
and \U$12790 ( \13105 , \709 , \9431 );
nor \U$12791 ( \13106 , \13104 , \13105 );
xnor \U$12792 ( \13107 , \13106 , \9123 );
and \U$12793 ( \13108 , \925 , \8896 );
and \U$12794 ( \13109 , \863 , \8894 );
nor \U$12795 ( \13110 , \13108 , \13109 );
xnor \U$12796 ( \13111 , \13110 , \8525 );
and \U$12797 ( \13112 , \13107 , \13111 );
and \U$12798 ( \13113 , \1186 , \8334 );
and \U$12799 ( \13114 , \988 , \8332 );
nor \U$12800 ( \13115 , \13113 , \13114 );
xnor \U$12801 ( \13116 , \13115 , \8016 );
and \U$12802 ( \13117 , \13111 , \13116 );
and \U$12803 ( \13118 , \13107 , \13116 );
or \U$12804 ( \13119 , \13112 , \13117 , \13118 );
and \U$12805 ( \13120 , \1379 , \7767 );
and \U$12806 ( \13121 , \1274 , \7765 );
nor \U$12807 ( \13122 , \13120 , \13121 );
xnor \U$12808 ( \13123 , \13122 , \7518 );
and \U$12809 ( \13124 , \1500 , \7238 );
and \U$12810 ( \13125 , \1384 , \7236 );
nor \U$12811 ( \13126 , \13124 , \13125 );
xnor \U$12812 ( \13127 , \13126 , \6978 );
and \U$12813 ( \13128 , \13123 , \13127 );
and \U$12814 ( \13129 , \1791 , \6744 );
and \U$12815 ( \13130 , \1615 , \6742 );
nor \U$12816 ( \13131 , \13129 , \13130 );
xnor \U$12817 ( \13132 , \13131 , \6429 );
and \U$12818 ( \13133 , \13127 , \13132 );
and \U$12819 ( \13134 , \13123 , \13132 );
or \U$12820 ( \13135 , \13128 , \13133 , \13134 );
and \U$12821 ( \13136 , \13119 , \13135 );
and \U$12822 ( \13137 , \553 , \10814 );
and \U$12823 ( \13138 , \499 , \10811 );
nor \U$12824 ( \13139 , \13137 , \13138 );
xnor \U$12825 ( \13140 , \13139 , \9759 );
and \U$12826 ( \13141 , \681 , \10001 );
and \U$12827 ( \13142 , \604 , \9999 );
nor \U$12828 ( \13143 , \13141 , \13142 );
xnor \U$12829 ( \13144 , \13143 , \9762 );
and \U$12830 ( \13145 , \13140 , \13144 );
and \U$12831 ( \13146 , \13144 , \437 );
and \U$12832 ( \13147 , \13140 , \437 );
or \U$12833 ( \13148 , \13145 , \13146 , \13147 );
and \U$12834 ( \13149 , \13135 , \13148 );
and \U$12835 ( \13150 , \13119 , \13148 );
or \U$12836 ( \13151 , \13136 , \13149 , \13150 );
and \U$12837 ( \13152 , \4011 , \3637 );
and \U$12838 ( \13153 , \3889 , \3635 );
nor \U$12839 ( \13154 , \13152 , \13153 );
xnor \U$12840 ( \13155 , \13154 , \3450 );
and \U$12841 ( \13156 , \4272 , \3324 );
and \U$12842 ( \13157 , \4016 , \3322 );
nor \U$12843 ( \13158 , \13156 , \13157 );
xnor \U$12844 ( \13159 , \13158 , \3119 );
and \U$12845 ( \13160 , \13155 , \13159 );
and \U$12846 ( \13161 , \4771 , \2918 );
and \U$12847 ( \13162 , \4469 , \2916 );
nor \U$12848 ( \13163 , \13161 , \13162 );
xnor \U$12849 ( \13164 , \13163 , \2769 );
and \U$12850 ( \13165 , \13159 , \13164 );
and \U$12851 ( \13166 , \13155 , \13164 );
or \U$12852 ( \13167 , \13160 , \13165 , \13166 );
and \U$12853 ( \13168 , \2042 , \6235 );
and \U$12854 ( \13169 , \1799 , \6233 );
nor \U$12855 ( \13170 , \13168 , \13169 );
xnor \U$12856 ( \13171 , \13170 , \5895 );
and \U$12857 ( \13172 , \2233 , \5646 );
and \U$12858 ( \13173 , \2047 , \5644 );
nor \U$12859 ( \13174 , \13172 , \13173 );
xnor \U$12860 ( \13175 , \13174 , \5405 );
and \U$12861 ( \13176 , \13171 , \13175 );
and \U$12862 ( \13177 , \2641 , \5180 );
and \U$12863 ( \13178 , \2377 , \5178 );
nor \U$12864 ( \13179 , \13177 , \13178 );
xnor \U$12865 ( \13180 , \13179 , \4992 );
and \U$12866 ( \13181 , \13175 , \13180 );
and \U$12867 ( \13182 , \13171 , \13180 );
or \U$12868 ( \13183 , \13176 , \13181 , \13182 );
and \U$12869 ( \13184 , \13167 , \13183 );
and \U$12870 ( \13185 , \2840 , \4806 );
and \U$12871 ( \13186 , \2666 , \4804 );
nor \U$12872 ( \13187 , \13185 , \13186 );
xnor \U$12873 ( \13188 , \13187 , \4574 );
and \U$12874 ( \13189 , \3145 , \4355 );
and \U$12875 ( \13190 , \3007 , \4353 );
nor \U$12876 ( \13191 , \13189 , \13190 );
xnor \U$12877 ( \13192 , \13191 , \4212 );
and \U$12878 ( \13193 , \13188 , \13192 );
and \U$12879 ( \13194 , \3681 , \4032 );
and \U$12880 ( \13195 , \3264 , \4030 );
nor \U$12881 ( \13196 , \13194 , \13195 );
xnor \U$12882 ( \13197 , \13196 , \3786 );
and \U$12883 ( \13198 , \13192 , \13197 );
and \U$12884 ( \13199 , \13188 , \13197 );
or \U$12885 ( \13200 , \13193 , \13198 , \13199 );
and \U$12886 ( \13201 , \13183 , \13200 );
and \U$12887 ( \13202 , \13167 , \13200 );
or \U$12888 ( \13203 , \13184 , \13201 , \13202 );
and \U$12889 ( \13204 , \13151 , \13203 );
and \U$12890 ( \13205 , \6500 , \1826 );
and \U$12891 ( \13206 , \6157 , \1824 );
nor \U$12892 ( \13207 , \13205 , \13206 );
xnor \U$12893 ( \13208 , \13207 , \1670 );
and \U$12894 ( \13209 , \7005 , \1554 );
and \U$12895 ( \13210 , \6702 , \1552 );
nor \U$12896 ( \13211 , \13209 , \13210 );
xnor \U$12897 ( \13212 , \13211 , \1441 );
and \U$12898 ( \13213 , \13208 , \13212 );
and \U$12899 ( \13214 , \7703 , \1360 );
and \U$12900 ( \13215 , \7177 , \1358 );
nor \U$12901 ( \13216 , \13214 , \13215 );
xnor \U$12902 ( \13217 , \13216 , \1224 );
and \U$12903 ( \13218 , \13212 , \13217 );
and \U$12904 ( \13219 , \13208 , \13217 );
or \U$12905 ( \13220 , \13213 , \13218 , \13219 );
and \U$12906 ( \13221 , \8373 , \1160 );
and \U$12907 ( \13222 , \8127 , \1158 );
nor \U$12908 ( \13223 , \13221 , \13222 );
xnor \U$12909 ( \13224 , \13223 , \1082 );
and \U$12910 ( \13225 , \8697 , \996 );
and \U$12911 ( \13226 , \8378 , \994 );
nor \U$12912 ( \13227 , \13225 , \13226 );
xnor \U$12913 ( \13228 , \13227 , \902 );
and \U$12914 ( \13229 , \13224 , \13228 );
and \U$12915 ( \13230 , \9550 , \826 );
and \U$12916 ( \13231 , \8981 , \824 );
nor \U$12917 ( \13232 , \13230 , \13231 );
xnor \U$12918 ( \13233 , \13232 , \754 );
and \U$12919 ( \13234 , \13228 , \13233 );
and \U$12920 ( \13235 , \13224 , \13233 );
or \U$12921 ( \13236 , \13229 , \13234 , \13235 );
and \U$12922 ( \13237 , \13220 , \13236 );
and \U$12923 ( \13238 , \5248 , \2596 );
and \U$12924 ( \13239 , \4779 , \2594 );
nor \U$12925 ( \13240 , \13238 , \13239 );
xnor \U$12926 ( \13241 , \13240 , \2454 );
and \U$12927 ( \13242 , \5517 , \2300 );
and \U$12928 ( \13243 , \5253 , \2298 );
nor \U$12929 ( \13244 , \13242 , \13243 );
xnor \U$12930 ( \13245 , \13244 , \2163 );
and \U$12931 ( \13246 , \13241 , \13245 );
and \U$12932 ( \13247 , \6148 , \2094 );
and \U$12933 ( \13248 , \5776 , \2092 );
nor \U$12934 ( \13249 , \13247 , \13248 );
xnor \U$12935 ( \13250 , \13249 , \1942 );
and \U$12936 ( \13251 , \13245 , \13250 );
and \U$12937 ( \13252 , \13241 , \13250 );
or \U$12938 ( \13253 , \13246 , \13251 , \13252 );
and \U$12939 ( \13254 , \13236 , \13253 );
and \U$12940 ( \13255 , \13220 , \13253 );
or \U$12941 ( \13256 , \13237 , \13254 , \13255 );
and \U$12942 ( \13257 , \13203 , \13256 );
and \U$12943 ( \13258 , \13151 , \13256 );
or \U$12944 ( \13259 , \13204 , \13257 , \13258 );
and \U$12945 ( \13260 , \13103 , \13259 );
xor \U$12946 ( \13261 , \12884 , \12888 );
xor \U$12947 ( \13262 , \13261 , \12893 );
xor \U$12948 ( \13263 , \12900 , \12904 );
xor \U$12949 ( \13264 , \13263 , \12909 );
and \U$12950 ( \13265 , \13262 , \13264 );
xor \U$12951 ( \13266 , \12917 , \12921 );
xor \U$12952 ( \13267 , \13266 , \12926 );
and \U$12953 ( \13268 , \13264 , \13267 );
and \U$12954 ( \13269 , \13262 , \13267 );
or \U$12955 ( \13270 , \13265 , \13268 , \13269 );
xor \U$12956 ( \13271 , \12558 , \12562 );
xor \U$12957 ( \13272 , \13271 , \378 );
and \U$12958 ( \13273 , \13270 , \13272 );
xor \U$12959 ( \13274 , \12571 , \12575 );
xor \U$12960 ( \13275 , \13274 , \12580 );
and \U$12961 ( \13276 , \13272 , \13275 );
and \U$12962 ( \13277 , \13270 , \13275 );
or \U$12963 ( \13278 , \13273 , \13276 , \13277 );
and \U$12964 ( \13279 , \13259 , \13278 );
and \U$12965 ( \13280 , \13103 , \13278 );
or \U$12966 ( \13281 , \13260 , \13279 , \13280 );
xor \U$12967 ( \13282 , \12791 , \12807 );
xor \U$12968 ( \13283 , \13282 , \12824 );
xor \U$12969 ( \13284 , \12843 , \12859 );
xor \U$12970 ( \13285 , \13284 , \12876 );
and \U$12971 ( \13286 , \13283 , \13285 );
xor \U$12972 ( \13287 , \12896 , \12912 );
xor \U$12973 ( \13288 , \13287 , \12929 );
and \U$12974 ( \13289 , \13285 , \13288 );
and \U$12975 ( \13290 , \13283 , \13288 );
or \U$12976 ( \13291 , \13286 , \13289 , \13290 );
xor \U$12977 ( \13292 , \12937 , \12939 );
xor \U$12978 ( \13293 , \13292 , \12942 );
xor \U$12979 ( \13294 , \12947 , \12949 );
xor \U$12980 ( \13295 , \13294 , \12952 );
and \U$12981 ( \13296 , \13293 , \13295 );
xor \U$12982 ( \13297 , \12958 , \12960 );
xor \U$12983 ( \13298 , \13297 , \12963 );
and \U$12984 ( \13299 , \13295 , \13298 );
and \U$12985 ( \13300 , \13293 , \13298 );
or \U$12986 ( \13301 , \13296 , \13299 , \13300 );
and \U$12987 ( \13302 , \13291 , \13301 );
xor \U$12988 ( \13303 , \12602 , \12618 );
xor \U$12989 ( \13304 , \13303 , \12635 );
and \U$12990 ( \13305 , \13301 , \13304 );
and \U$12991 ( \13306 , \13291 , \13304 );
or \U$12992 ( \13307 , \13302 , \13305 , \13306 );
and \U$12993 ( \13308 , \13281 , \13307 );
xor \U$12994 ( \13309 , \12554 , \12566 );
xor \U$12995 ( \13310 , \13309 , \12583 );
xor \U$12996 ( \13311 , \12972 , \12974 );
xor \U$12997 ( \13312 , \13311 , \12977 );
and \U$12998 ( \13313 , \13310 , \13312 );
xor \U$12999 ( \13314 , \12996 , \12998 );
xor \U$13000 ( \13315 , \13314 , \13001 );
and \U$13001 ( \13316 , \13312 , \13315 );
and \U$13002 ( \13317 , \13310 , \13315 );
or \U$13003 ( \13318 , \13313 , \13316 , \13317 );
and \U$13004 ( \13319 , \13307 , \13318 );
and \U$13005 ( \13320 , \13281 , \13318 );
or \U$13006 ( \13321 , \13308 , \13319 , \13320 );
xor \U$13007 ( \13322 , \12935 , \12969 );
xor \U$13008 ( \13323 , \13322 , \12980 );
xor \U$13009 ( \13324 , \12985 , \12987 );
xor \U$13010 ( \13325 , \13324 , \12990 );
and \U$13011 ( \13326 , \13323 , \13325 );
xor \U$13012 ( \13327 , \13004 , \13006 );
xor \U$13013 ( \13328 , \13327 , \13009 );
and \U$13014 ( \13329 , \13325 , \13328 );
and \U$13015 ( \13330 , \13323 , \13328 );
or \U$13016 ( \13331 , \13326 , \13329 , \13330 );
and \U$13017 ( \13332 , \13321 , \13331 );
xor \U$13018 ( \13333 , \13017 , \13019 );
xor \U$13019 ( \13334 , \13333 , \13022 );
and \U$13020 ( \13335 , \13331 , \13334 );
and \U$13021 ( \13336 , \13321 , \13334 );
or \U$13022 ( \13337 , \13332 , \13335 , \13336 );
xor \U$13023 ( \13338 , \13015 , \13025 );
xor \U$13024 ( \13339 , \13338 , \13028 );
and \U$13025 ( \13340 , \13337 , \13339 );
xor \U$13026 ( \13341 , \13033 , \13035 );
xor \U$13027 ( \13342 , \13341 , \13038 );
and \U$13028 ( \13343 , \13339 , \13342 );
and \U$13029 ( \13344 , \13337 , \13342 );
or \U$13030 ( \13345 , \13340 , \13343 , \13344 );
xor \U$13031 ( \13346 , \13031 , \13041 );
xor \U$13032 ( \13347 , \13346 , \13044 );
and \U$13033 ( \13348 , \13345 , \13347 );
xor \U$13034 ( \13349 , \12740 , \12750 );
xor \U$13035 ( \13350 , \13349 , \12753 );
and \U$13036 ( \13351 , \13347 , \13350 );
and \U$13037 ( \13352 , \13345 , \13350 );
or \U$13038 ( \13353 , \13348 , \13351 , \13352 );
and \U$13039 ( \13354 , \13053 , \13353 );
xor \U$13040 ( \13355 , \13053 , \13353 );
xor \U$13041 ( \13356 , \13345 , \13347 );
xor \U$13042 ( \13357 , \13356 , \13350 );
xor \U$13043 ( \13358 , \13107 , \13111 );
xor \U$13044 ( \13359 , \13358 , \13116 );
xor \U$13045 ( \13360 , \13123 , \13127 );
xor \U$13046 ( \13361 , \13360 , \13132 );
and \U$13047 ( \13362 , \13359 , \13361 );
xor \U$13048 ( \13363 , \13171 , \13175 );
xor \U$13049 ( \13364 , \13363 , \13180 );
and \U$13050 ( \13365 , \13361 , \13364 );
and \U$13051 ( \13366 , \13359 , \13364 );
or \U$13052 ( \13367 , \13362 , \13365 , \13366 );
xor \U$13053 ( \13368 , \13155 , \13159 );
xor \U$13054 ( \13369 , \13368 , \13164 );
xor \U$13055 ( \13370 , \13188 , \13192 );
xor \U$13056 ( \13371 , \13370 , \13197 );
and \U$13057 ( \13372 , \13369 , \13371 );
xor \U$13058 ( \13373 , \13241 , \13245 );
xor \U$13059 ( \13374 , \13373 , \13250 );
and \U$13060 ( \13375 , \13371 , \13374 );
and \U$13061 ( \13376 , \13369 , \13374 );
or \U$13062 ( \13377 , \13372 , \13375 , \13376 );
and \U$13063 ( \13378 , \13367 , \13377 );
xor \U$13064 ( \13379 , \13208 , \13212 );
xor \U$13065 ( \13380 , \13379 , \13217 );
xor \U$13066 ( \13381 , \13057 , \13061 );
xor \U$13067 ( \13382 , \13381 , \13064 );
and \U$13068 ( \13383 , \13380 , \13382 );
xor \U$13069 ( \13384 , \13224 , \13228 );
xor \U$13070 ( \13385 , \13384 , \13233 );
and \U$13071 ( \13386 , \13382 , \13385 );
and \U$13072 ( \13387 , \13380 , \13385 );
or \U$13073 ( \13388 , \13383 , \13386 , \13387 );
and \U$13074 ( \13389 , \13377 , \13388 );
and \U$13075 ( \13390 , \13367 , \13388 );
or \U$13076 ( \13391 , \13378 , \13389 , \13390 );
and \U$13077 ( \13392 , \2377 , \5646 );
and \U$13078 ( \13393 , \2233 , \5644 );
nor \U$13079 ( \13394 , \13392 , \13393 );
xnor \U$13080 ( \13395 , \13394 , \5405 );
and \U$13081 ( \13396 , \2666 , \5180 );
and \U$13082 ( \13397 , \2641 , \5178 );
nor \U$13083 ( \13398 , \13396 , \13397 );
xnor \U$13084 ( \13399 , \13398 , \4992 );
and \U$13085 ( \13400 , \13395 , \13399 );
and \U$13086 ( \13401 , \3007 , \4806 );
and \U$13087 ( \13402 , \2840 , \4804 );
nor \U$13088 ( \13403 , \13401 , \13402 );
xnor \U$13089 ( \13404 , \13403 , \4574 );
and \U$13090 ( \13405 , \13399 , \13404 );
and \U$13091 ( \13406 , \13395 , \13404 );
or \U$13092 ( \13407 , \13400 , \13405 , \13406 );
and \U$13093 ( \13408 , \4469 , \3324 );
and \U$13094 ( \13409 , \4272 , \3322 );
nor \U$13095 ( \13410 , \13408 , \13409 );
xnor \U$13096 ( \13411 , \13410 , \3119 );
and \U$13097 ( \13412 , \4779 , \2918 );
and \U$13098 ( \13413 , \4771 , \2916 );
nor \U$13099 ( \13414 , \13412 , \13413 );
xnor \U$13100 ( \13415 , \13414 , \2769 );
and \U$13101 ( \13416 , \13411 , \13415 );
and \U$13102 ( \13417 , \5253 , \2596 );
and \U$13103 ( \13418 , \5248 , \2594 );
nor \U$13104 ( \13419 , \13417 , \13418 );
xnor \U$13105 ( \13420 , \13419 , \2454 );
and \U$13106 ( \13421 , \13415 , \13420 );
and \U$13107 ( \13422 , \13411 , \13420 );
or \U$13108 ( \13423 , \13416 , \13421 , \13422 );
and \U$13109 ( \13424 , \13407 , \13423 );
and \U$13110 ( \13425 , \3264 , \4355 );
and \U$13111 ( \13426 , \3145 , \4353 );
nor \U$13112 ( \13427 , \13425 , \13426 );
xnor \U$13113 ( \13428 , \13427 , \4212 );
and \U$13114 ( \13429 , \3889 , \4032 );
and \U$13115 ( \13430 , \3681 , \4030 );
nor \U$13116 ( \13431 , \13429 , \13430 );
xnor \U$13117 ( \13432 , \13431 , \3786 );
and \U$13118 ( \13433 , \13428 , \13432 );
and \U$13119 ( \13434 , \4016 , \3637 );
and \U$13120 ( \13435 , \4011 , \3635 );
nor \U$13121 ( \13436 , \13434 , \13435 );
xnor \U$13122 ( \13437 , \13436 , \3450 );
and \U$13123 ( \13438 , \13432 , \13437 );
and \U$13124 ( \13439 , \13428 , \13437 );
or \U$13125 ( \13440 , \13433 , \13438 , \13439 );
and \U$13126 ( \13441 , \13423 , \13440 );
and \U$13127 ( \13442 , \13407 , \13440 );
or \U$13128 ( \13443 , \13424 , \13441 , \13442 );
and \U$13129 ( \13444 , \8981 , \996 );
and \U$13130 ( \13445 , \8697 , \994 );
nor \U$13131 ( \13446 , \13444 , \13445 );
xnor \U$13132 ( \13447 , \13446 , \902 );
and \U$13133 ( \13448 , \9558 , \826 );
and \U$13134 ( \13449 , \9550 , \824 );
nor \U$13135 ( \13450 , \13448 , \13449 );
xnor \U$13136 ( \13451 , \13450 , \754 );
and \U$13137 ( \13452 , \13447 , \13451 );
and \U$13138 ( \13453 , \10166 , \692 );
and \U$13139 ( \13454 , \10161 , \690 );
nor \U$13140 ( \13455 , \13453 , \13454 );
xnor \U$13141 ( \13456 , \13455 , \649 );
and \U$13142 ( \13457 , \13451 , \13456 );
and \U$13143 ( \13458 , \13447 , \13456 );
or \U$13144 ( \13459 , \13452 , \13457 , \13458 );
and \U$13145 ( \13460 , \7177 , \1554 );
and \U$13146 ( \13461 , \7005 , \1552 );
nor \U$13147 ( \13462 , \13460 , \13461 );
xnor \U$13148 ( \13463 , \13462 , \1441 );
and \U$13149 ( \13464 , \8127 , \1360 );
and \U$13150 ( \13465 , \7703 , \1358 );
nor \U$13151 ( \13466 , \13464 , \13465 );
xnor \U$13152 ( \13467 , \13466 , \1224 );
and \U$13153 ( \13468 , \13463 , \13467 );
and \U$13154 ( \13469 , \8378 , \1160 );
and \U$13155 ( \13470 , \8373 , \1158 );
nor \U$13156 ( \13471 , \13469 , \13470 );
xnor \U$13157 ( \13472 , \13471 , \1082 );
and \U$13158 ( \13473 , \13467 , \13472 );
and \U$13159 ( \13474 , \13463 , \13472 );
or \U$13160 ( \13475 , \13468 , \13473 , \13474 );
and \U$13161 ( \13476 , \13459 , \13475 );
and \U$13162 ( \13477 , \5776 , \2300 );
and \U$13163 ( \13478 , \5517 , \2298 );
nor \U$13164 ( \13479 , \13477 , \13478 );
xnor \U$13165 ( \13480 , \13479 , \2163 );
and \U$13166 ( \13481 , \6157 , \2094 );
and \U$13167 ( \13482 , \6148 , \2092 );
nor \U$13168 ( \13483 , \13481 , \13482 );
xnor \U$13169 ( \13484 , \13483 , \1942 );
and \U$13170 ( \13485 , \13480 , \13484 );
and \U$13171 ( \13486 , \6702 , \1826 );
and \U$13172 ( \13487 , \6500 , \1824 );
nor \U$13173 ( \13488 , \13486 , \13487 );
xnor \U$13174 ( \13489 , \13488 , \1670 );
and \U$13175 ( \13490 , \13484 , \13489 );
and \U$13176 ( \13491 , \13480 , \13489 );
or \U$13177 ( \13492 , \13485 , \13490 , \13491 );
and \U$13178 ( \13493 , \13475 , \13492 );
and \U$13179 ( \13494 , \13459 , \13492 );
or \U$13180 ( \13495 , \13476 , \13493 , \13494 );
and \U$13181 ( \13496 , \13443 , \13495 );
and \U$13182 ( \13497 , \1615 , \7238 );
and \U$13183 ( \13498 , \1500 , \7236 );
nor \U$13184 ( \13499 , \13497 , \13498 );
xnor \U$13185 ( \13500 , \13499 , \6978 );
and \U$13186 ( \13501 , \1799 , \6744 );
and \U$13187 ( \13502 , \1791 , \6742 );
nor \U$13188 ( \13503 , \13501 , \13502 );
xnor \U$13189 ( \13504 , \13503 , \6429 );
and \U$13190 ( \13505 , \13500 , \13504 );
and \U$13191 ( \13506 , \2047 , \6235 );
and \U$13192 ( \13507 , \2042 , \6233 );
nor \U$13193 ( \13508 , \13506 , \13507 );
xnor \U$13194 ( \13509 , \13508 , \5895 );
and \U$13195 ( \13510 , \13504 , \13509 );
and \U$13196 ( \13511 , \13500 , \13509 );
or \U$13197 ( \13512 , \13505 , \13510 , \13511 );
and \U$13198 ( \13513 , \604 , \10814 );
and \U$13199 ( \13514 , \553 , \10811 );
nor \U$13200 ( \13515 , \13513 , \13514 );
xnor \U$13201 ( \13516 , \13515 , \9759 );
and \U$13202 ( \13517 , \709 , \10001 );
and \U$13203 ( \13518 , \681 , \9999 );
nor \U$13204 ( \13519 , \13517 , \13518 );
xnor \U$13205 ( \13520 , \13519 , \9762 );
and \U$13206 ( \13521 , \13516 , \13520 );
and \U$13207 ( \13522 , \863 , \9433 );
and \U$13208 ( \13523 , \789 , \9431 );
nor \U$13209 ( \13524 , \13522 , \13523 );
xnor \U$13210 ( \13525 , \13524 , \9123 );
and \U$13211 ( \13526 , \13520 , \13525 );
and \U$13212 ( \13527 , \13516 , \13525 );
or \U$13213 ( \13528 , \13521 , \13526 , \13527 );
and \U$13214 ( \13529 , \13512 , \13528 );
and \U$13215 ( \13530 , \988 , \8896 );
and \U$13216 ( \13531 , \925 , \8894 );
nor \U$13217 ( \13532 , \13530 , \13531 );
xnor \U$13218 ( \13533 , \13532 , \8525 );
and \U$13219 ( \13534 , \1274 , \8334 );
and \U$13220 ( \13535 , \1186 , \8332 );
nor \U$13221 ( \13536 , \13534 , \13535 );
xnor \U$13222 ( \13537 , \13536 , \8016 );
and \U$13223 ( \13538 , \13533 , \13537 );
and \U$13224 ( \13539 , \1384 , \7767 );
and \U$13225 ( \13540 , \1379 , \7765 );
nor \U$13226 ( \13541 , \13539 , \13540 );
xnor \U$13227 ( \13542 , \13541 , \7518 );
and \U$13228 ( \13543 , \13537 , \13542 );
and \U$13229 ( \13544 , \13533 , \13542 );
or \U$13230 ( \13545 , \13538 , \13543 , \13544 );
and \U$13231 ( \13546 , \13528 , \13545 );
and \U$13232 ( \13547 , \13512 , \13545 );
or \U$13233 ( \13548 , \13529 , \13546 , \13547 );
and \U$13234 ( \13549 , \13495 , \13548 );
and \U$13235 ( \13550 , \13443 , \13548 );
or \U$13236 ( \13551 , \13496 , \13549 , \13550 );
and \U$13237 ( \13552 , \13391 , \13551 );
xor \U$13238 ( \13553 , \13081 , \13083 );
xor \U$13239 ( \13554 , \13553 , \13086 );
xor \U$13240 ( \13555 , \13262 , \13264 );
xor \U$13241 ( \13556 , \13555 , \13267 );
and \U$13242 ( \13557 , \13554 , \13556 );
xor \U$13243 ( \13558 , \13092 , \13094 );
xor \U$13244 ( \13559 , \13558 , \13097 );
and \U$13245 ( \13560 , \13556 , \13559 );
and \U$13246 ( \13561 , \13554 , \13559 );
or \U$13247 ( \13562 , \13557 , \13560 , \13561 );
and \U$13248 ( \13563 , \13551 , \13562 );
and \U$13249 ( \13564 , \13391 , \13562 );
or \U$13250 ( \13565 , \13552 , \13563 , \13564 );
xor \U$13251 ( \13566 , \13079 , \13089 );
xor \U$13252 ( \13567 , \13566 , \13100 );
xor \U$13253 ( \13568 , \13151 , \13203 );
xor \U$13254 ( \13569 , \13568 , \13256 );
and \U$13255 ( \13570 , \13567 , \13569 );
xor \U$13256 ( \13571 , \13270 , \13272 );
xor \U$13257 ( \13572 , \13571 , \13275 );
and \U$13258 ( \13573 , \13569 , \13572 );
and \U$13259 ( \13574 , \13567 , \13572 );
or \U$13260 ( \13575 , \13570 , \13573 , \13574 );
and \U$13261 ( \13576 , \13565 , \13575 );
xor \U$13262 ( \13577 , \13067 , \13071 );
xor \U$13263 ( \13578 , \13577 , \13076 );
xor \U$13264 ( \13579 , \13167 , \13183 );
xor \U$13265 ( \13580 , \13579 , \13200 );
and \U$13266 ( \13581 , \13578 , \13580 );
xor \U$13267 ( \13582 , \13220 , \13236 );
xor \U$13268 ( \13583 , \13582 , \13253 );
and \U$13269 ( \13584 , \13580 , \13583 );
and \U$13270 ( \13585 , \13578 , \13583 );
or \U$13271 ( \13586 , \13581 , \13584 , \13585 );
xor \U$13272 ( \13587 , \13283 , \13285 );
xor \U$13273 ( \13588 , \13587 , \13288 );
and \U$13274 ( \13589 , \13586 , \13588 );
xor \U$13275 ( \13590 , \13293 , \13295 );
xor \U$13276 ( \13591 , \13590 , \13298 );
and \U$13277 ( \13592 , \13588 , \13591 );
and \U$13278 ( \13593 , \13586 , \13591 );
or \U$13279 ( \13594 , \13589 , \13592 , \13593 );
and \U$13280 ( \13595 , \13575 , \13594 );
and \U$13281 ( \13596 , \13565 , \13594 );
or \U$13282 ( \13597 , \13576 , \13595 , \13596 );
xor \U$13283 ( \13598 , \12827 , \12879 );
xor \U$13284 ( \13599 , \13598 , \12932 );
xor \U$13285 ( \13600 , \12945 , \12955 );
xor \U$13286 ( \13601 , \13600 , \12966 );
and \U$13287 ( \13602 , \13599 , \13601 );
xor \U$13288 ( \13603 , \13310 , \13312 );
xor \U$13289 ( \13604 , \13603 , \13315 );
and \U$13290 ( \13605 , \13601 , \13604 );
and \U$13291 ( \13606 , \13599 , \13604 );
or \U$13292 ( \13607 , \13602 , \13605 , \13606 );
and \U$13293 ( \13608 , \13597 , \13607 );
xor \U$13294 ( \13609 , \13323 , \13325 );
xor \U$13295 ( \13610 , \13609 , \13328 );
and \U$13296 ( \13611 , \13607 , \13610 );
and \U$13297 ( \13612 , \13597 , \13610 );
or \U$13298 ( \13613 , \13608 , \13611 , \13612 );
xor \U$13299 ( \13614 , \12983 , \12993 );
xor \U$13300 ( \13615 , \13614 , \13012 );
and \U$13301 ( \13616 , \13613 , \13615 );
xor \U$13302 ( \13617 , \13321 , \13331 );
xor \U$13303 ( \13618 , \13617 , \13334 );
and \U$13304 ( \13619 , \13615 , \13618 );
and \U$13305 ( \13620 , \13613 , \13618 );
or \U$13306 ( \13621 , \13616 , \13619 , \13620 );
xor \U$13307 ( \13622 , \13337 , \13339 );
xor \U$13308 ( \13623 , \13622 , \13342 );
and \U$13309 ( \13624 , \13621 , \13623 );
and \U$13310 ( \13625 , \13357 , \13624 );
xor \U$13311 ( \13626 , \13357 , \13624 );
xor \U$13312 ( \13627 , \13621 , \13623 );
xor \U$13313 ( \13628 , \13411 , \13415 );
xor \U$13314 ( \13629 , \13628 , \13420 );
xor \U$13315 ( \13630 , \13428 , \13432 );
xor \U$13316 ( \13631 , \13630 , \13437 );
and \U$13317 ( \13632 , \13629 , \13631 );
xor \U$13318 ( \13633 , \13480 , \13484 );
xor \U$13319 ( \13634 , \13633 , \13489 );
and \U$13320 ( \13635 , \13631 , \13634 );
and \U$13321 ( \13636 , \13629 , \13634 );
or \U$13322 ( \13637 , \13632 , \13635 , \13636 );
xor \U$13323 ( \13638 , \13395 , \13399 );
xor \U$13324 ( \13639 , \13638 , \13404 );
xor \U$13325 ( \13640 , \13500 , \13504 );
xor \U$13326 ( \13641 , \13640 , \13509 );
and \U$13327 ( \13642 , \13639 , \13641 );
xor \U$13328 ( \13643 , \13533 , \13537 );
xor \U$13329 ( \13644 , \13643 , \13542 );
and \U$13330 ( \13645 , \13641 , \13644 );
and \U$13331 ( \13646 , \13639 , \13644 );
or \U$13332 ( \13647 , \13642 , \13645 , \13646 );
and \U$13333 ( \13648 , \13637 , \13647 );
and \U$13334 ( \13649 , \10967 , \579 );
and \U$13335 ( \13650 , \10347 , \577 );
nor \U$13336 ( \13651 , \13649 , \13650 );
xnor \U$13337 ( \13652 , \13651 , \530 );
xor \U$13338 ( \13653 , \13447 , \13451 );
xor \U$13339 ( \13654 , \13653 , \13456 );
and \U$13340 ( \13655 , \13652 , \13654 );
xor \U$13341 ( \13656 , \13463 , \13467 );
xor \U$13342 ( \13657 , \13656 , \13472 );
and \U$13343 ( \13658 , \13654 , \13657 );
and \U$13344 ( \13659 , \13652 , \13657 );
or \U$13345 ( \13660 , \13655 , \13658 , \13659 );
and \U$13346 ( \13661 , \13647 , \13660 );
and \U$13347 ( \13662 , \13637 , \13660 );
or \U$13348 ( \13663 , \13648 , \13661 , \13662 );
and \U$13349 ( \13664 , \1500 , \7767 );
and \U$13350 ( \13665 , \1384 , \7765 );
nor \U$13351 ( \13666 , \13664 , \13665 );
xnor \U$13352 ( \13667 , \13666 , \7518 );
and \U$13353 ( \13668 , \1791 , \7238 );
and \U$13354 ( \13669 , \1615 , \7236 );
nor \U$13355 ( \13670 , \13668 , \13669 );
xnor \U$13356 ( \13671 , \13670 , \6978 );
and \U$13357 ( \13672 , \13667 , \13671 );
and \U$13358 ( \13673 , \2042 , \6744 );
and \U$13359 ( \13674 , \1799 , \6742 );
nor \U$13360 ( \13675 , \13673 , \13674 );
xnor \U$13361 ( \13676 , \13675 , \6429 );
and \U$13362 ( \13677 , \13671 , \13676 );
and \U$13363 ( \13678 , \13667 , \13676 );
or \U$13364 ( \13679 , \13672 , \13677 , \13678 );
and \U$13365 ( \13680 , \925 , \9433 );
and \U$13366 ( \13681 , \863 , \9431 );
nor \U$13367 ( \13682 , \13680 , \13681 );
xnor \U$13368 ( \13683 , \13682 , \9123 );
and \U$13369 ( \13684 , \1186 , \8896 );
and \U$13370 ( \13685 , \988 , \8894 );
nor \U$13371 ( \13686 , \13684 , \13685 );
xnor \U$13372 ( \13687 , \13686 , \8525 );
and \U$13373 ( \13688 , \13683 , \13687 );
and \U$13374 ( \13689 , \1379 , \8334 );
and \U$13375 ( \13690 , \1274 , \8332 );
nor \U$13376 ( \13691 , \13689 , \13690 );
xnor \U$13377 ( \13692 , \13691 , \8016 );
and \U$13378 ( \13693 , \13687 , \13692 );
and \U$13379 ( \13694 , \13683 , \13692 );
or \U$13380 ( \13695 , \13688 , \13693 , \13694 );
and \U$13381 ( \13696 , \13679 , \13695 );
and \U$13382 ( \13697 , \681 , \10814 );
and \U$13383 ( \13698 , \604 , \10811 );
nor \U$13384 ( \13699 , \13697 , \13698 );
xnor \U$13385 ( \13700 , \13699 , \9759 );
and \U$13386 ( \13701 , \789 , \10001 );
and \U$13387 ( \13702 , \709 , \9999 );
nor \U$13388 ( \13703 , \13701 , \13702 );
xnor \U$13389 ( \13704 , \13703 , \9762 );
and \U$13390 ( \13705 , \13700 , \13704 );
and \U$13391 ( \13706 , \13704 , \530 );
and \U$13392 ( \13707 , \13700 , \530 );
or \U$13393 ( \13708 , \13705 , \13706 , \13707 );
and \U$13394 ( \13709 , \13695 , \13708 );
and \U$13395 ( \13710 , \13679 , \13708 );
or \U$13396 ( \13711 , \13696 , \13709 , \13710 );
and \U$13397 ( \13712 , \8697 , \1160 );
and \U$13398 ( \13713 , \8378 , \1158 );
nor \U$13399 ( \13714 , \13712 , \13713 );
xnor \U$13400 ( \13715 , \13714 , \1082 );
and \U$13401 ( \13716 , \9550 , \996 );
and \U$13402 ( \13717 , \8981 , \994 );
nor \U$13403 ( \13718 , \13716 , \13717 );
xnor \U$13404 ( \13719 , \13718 , \902 );
and \U$13405 ( \13720 , \13715 , \13719 );
and \U$13406 ( \13721 , \10161 , \826 );
and \U$13407 ( \13722 , \9558 , \824 );
nor \U$13408 ( \13723 , \13721 , \13722 );
xnor \U$13409 ( \13724 , \13723 , \754 );
and \U$13410 ( \13725 , \13719 , \13724 );
and \U$13411 ( \13726 , \13715 , \13724 );
or \U$13412 ( \13727 , \13720 , \13725 , \13726 );
and \U$13413 ( \13728 , \5517 , \2596 );
and \U$13414 ( \13729 , \5253 , \2594 );
nor \U$13415 ( \13730 , \13728 , \13729 );
xnor \U$13416 ( \13731 , \13730 , \2454 );
and \U$13417 ( \13732 , \6148 , \2300 );
and \U$13418 ( \13733 , \5776 , \2298 );
nor \U$13419 ( \13734 , \13732 , \13733 );
xnor \U$13420 ( \13735 , \13734 , \2163 );
and \U$13421 ( \13736 , \13731 , \13735 );
and \U$13422 ( \13737 , \6500 , \2094 );
and \U$13423 ( \13738 , \6157 , \2092 );
nor \U$13424 ( \13739 , \13737 , \13738 );
xnor \U$13425 ( \13740 , \13739 , \1942 );
and \U$13426 ( \13741 , \13735 , \13740 );
and \U$13427 ( \13742 , \13731 , \13740 );
or \U$13428 ( \13743 , \13736 , \13741 , \13742 );
and \U$13429 ( \13744 , \13727 , \13743 );
and \U$13430 ( \13745 , \7005 , \1826 );
and \U$13431 ( \13746 , \6702 , \1824 );
nor \U$13432 ( \13747 , \13745 , \13746 );
xnor \U$13433 ( \13748 , \13747 , \1670 );
and \U$13434 ( \13749 , \7703 , \1554 );
and \U$13435 ( \13750 , \7177 , \1552 );
nor \U$13436 ( \13751 , \13749 , \13750 );
xnor \U$13437 ( \13752 , \13751 , \1441 );
and \U$13438 ( \13753 , \13748 , \13752 );
and \U$13439 ( \13754 , \8373 , \1360 );
and \U$13440 ( \13755 , \8127 , \1358 );
nor \U$13441 ( \13756 , \13754 , \13755 );
xnor \U$13442 ( \13757 , \13756 , \1224 );
and \U$13443 ( \13758 , \13752 , \13757 );
and \U$13444 ( \13759 , \13748 , \13757 );
or \U$13445 ( \13760 , \13753 , \13758 , \13759 );
and \U$13446 ( \13761 , \13743 , \13760 );
and \U$13447 ( \13762 , \13727 , \13760 );
or \U$13448 ( \13763 , \13744 , \13761 , \13762 );
and \U$13449 ( \13764 , \13711 , \13763 );
and \U$13450 ( \13765 , \4272 , \3637 );
and \U$13451 ( \13766 , \4016 , \3635 );
nor \U$13452 ( \13767 , \13765 , \13766 );
xnor \U$13453 ( \13768 , \13767 , \3450 );
and \U$13454 ( \13769 , \4771 , \3324 );
and \U$13455 ( \13770 , \4469 , \3322 );
nor \U$13456 ( \13771 , \13769 , \13770 );
xnor \U$13457 ( \13772 , \13771 , \3119 );
and \U$13458 ( \13773 , \13768 , \13772 );
and \U$13459 ( \13774 , \5248 , \2918 );
and \U$13460 ( \13775 , \4779 , \2916 );
nor \U$13461 ( \13776 , \13774 , \13775 );
xnor \U$13462 ( \13777 , \13776 , \2769 );
and \U$13463 ( \13778 , \13772 , \13777 );
and \U$13464 ( \13779 , \13768 , \13777 );
or \U$13465 ( \13780 , \13773 , \13778 , \13779 );
and \U$13466 ( \13781 , \3145 , \4806 );
and \U$13467 ( \13782 , \3007 , \4804 );
nor \U$13468 ( \13783 , \13781 , \13782 );
xnor \U$13469 ( \13784 , \13783 , \4574 );
and \U$13470 ( \13785 , \3681 , \4355 );
and \U$13471 ( \13786 , \3264 , \4353 );
nor \U$13472 ( \13787 , \13785 , \13786 );
xnor \U$13473 ( \13788 , \13787 , \4212 );
and \U$13474 ( \13789 , \13784 , \13788 );
and \U$13475 ( \13790 , \4011 , \4032 );
and \U$13476 ( \13791 , \3889 , \4030 );
nor \U$13477 ( \13792 , \13790 , \13791 );
xnor \U$13478 ( \13793 , \13792 , \3786 );
and \U$13479 ( \13794 , \13788 , \13793 );
and \U$13480 ( \13795 , \13784 , \13793 );
or \U$13481 ( \13796 , \13789 , \13794 , \13795 );
and \U$13482 ( \13797 , \13780 , \13796 );
and \U$13483 ( \13798 , \2233 , \6235 );
and \U$13484 ( \13799 , \2047 , \6233 );
nor \U$13485 ( \13800 , \13798 , \13799 );
xnor \U$13486 ( \13801 , \13800 , \5895 );
and \U$13487 ( \13802 , \2641 , \5646 );
and \U$13488 ( \13803 , \2377 , \5644 );
nor \U$13489 ( \13804 , \13802 , \13803 );
xnor \U$13490 ( \13805 , \13804 , \5405 );
and \U$13491 ( \13806 , \13801 , \13805 );
and \U$13492 ( \13807 , \2840 , \5180 );
and \U$13493 ( \13808 , \2666 , \5178 );
nor \U$13494 ( \13809 , \13807 , \13808 );
xnor \U$13495 ( \13810 , \13809 , \4992 );
and \U$13496 ( \13811 , \13805 , \13810 );
and \U$13497 ( \13812 , \13801 , \13810 );
or \U$13498 ( \13813 , \13806 , \13811 , \13812 );
and \U$13499 ( \13814 , \13796 , \13813 );
and \U$13500 ( \13815 , \13780 , \13813 );
or \U$13501 ( \13816 , \13797 , \13814 , \13815 );
and \U$13502 ( \13817 , \13763 , \13816 );
and \U$13503 ( \13818 , \13711 , \13816 );
or \U$13504 ( \13819 , \13764 , \13817 , \13818 );
and \U$13505 ( \13820 , \13663 , \13819 );
xor \U$13506 ( \13821 , \13140 , \13144 );
xor \U$13507 ( \13822 , \13821 , \437 );
xor \U$13508 ( \13823 , \13359 , \13361 );
xor \U$13509 ( \13824 , \13823 , \13364 );
and \U$13510 ( \13825 , \13822 , \13824 );
xor \U$13511 ( \13826 , \13369 , \13371 );
xor \U$13512 ( \13827 , \13826 , \13374 );
and \U$13513 ( \13828 , \13824 , \13827 );
and \U$13514 ( \13829 , \13822 , \13827 );
or \U$13515 ( \13830 , \13825 , \13828 , \13829 );
and \U$13516 ( \13831 , \13819 , \13830 );
and \U$13517 ( \13832 , \13663 , \13830 );
or \U$13518 ( \13833 , \13820 , \13831 , \13832 );
xor \U$13519 ( \13834 , \13407 , \13423 );
xor \U$13520 ( \13835 , \13834 , \13440 );
xor \U$13521 ( \13836 , \13459 , \13475 );
xor \U$13522 ( \13837 , \13836 , \13492 );
and \U$13523 ( \13838 , \13835 , \13837 );
xor \U$13524 ( \13839 , \13380 , \13382 );
xor \U$13525 ( \13840 , \13839 , \13385 );
and \U$13526 ( \13841 , \13837 , \13840 );
and \U$13527 ( \13842 , \13835 , \13840 );
or \U$13528 ( \13843 , \13838 , \13841 , \13842 );
xor \U$13529 ( \13844 , \13119 , \13135 );
xor \U$13530 ( \13845 , \13844 , \13148 );
and \U$13531 ( \13846 , \13843 , \13845 );
xor \U$13532 ( \13847 , \13578 , \13580 );
xor \U$13533 ( \13848 , \13847 , \13583 );
and \U$13534 ( \13849 , \13845 , \13848 );
and \U$13535 ( \13850 , \13843 , \13848 );
or \U$13536 ( \13851 , \13846 , \13849 , \13850 );
and \U$13537 ( \13852 , \13833 , \13851 );
xor \U$13538 ( \13853 , \13367 , \13377 );
xor \U$13539 ( \13854 , \13853 , \13388 );
xor \U$13540 ( \13855 , \13443 , \13495 );
xor \U$13541 ( \13856 , \13855 , \13548 );
and \U$13542 ( \13857 , \13854 , \13856 );
xor \U$13543 ( \13858 , \13554 , \13556 );
xor \U$13544 ( \13859 , \13858 , \13559 );
and \U$13545 ( \13860 , \13856 , \13859 );
and \U$13546 ( \13861 , \13854 , \13859 );
or \U$13547 ( \13862 , \13857 , \13860 , \13861 );
and \U$13548 ( \13863 , \13851 , \13862 );
and \U$13549 ( \13864 , \13833 , \13862 );
or \U$13550 ( \13865 , \13852 , \13863 , \13864 );
xor \U$13551 ( \13866 , \13391 , \13551 );
xor \U$13552 ( \13867 , \13866 , \13562 );
xor \U$13553 ( \13868 , \13567 , \13569 );
xor \U$13554 ( \13869 , \13868 , \13572 );
and \U$13555 ( \13870 , \13867 , \13869 );
xor \U$13556 ( \13871 , \13586 , \13588 );
xor \U$13557 ( \13872 , \13871 , \13591 );
and \U$13558 ( \13873 , \13869 , \13872 );
and \U$13559 ( \13874 , \13867 , \13872 );
or \U$13560 ( \13875 , \13870 , \13873 , \13874 );
and \U$13561 ( \13876 , \13865 , \13875 );
xor \U$13562 ( \13877 , \13291 , \13301 );
xor \U$13563 ( \13878 , \13877 , \13304 );
and \U$13564 ( \13879 , \13875 , \13878 );
and \U$13565 ( \13880 , \13865 , \13878 );
or \U$13566 ( \13881 , \13876 , \13879 , \13880 );
xor \U$13567 ( \13882 , \13103 , \13259 );
xor \U$13568 ( \13883 , \13882 , \13278 );
xor \U$13569 ( \13884 , \13565 , \13575 );
xor \U$13570 ( \13885 , \13884 , \13594 );
and \U$13571 ( \13886 , \13883 , \13885 );
xor \U$13572 ( \13887 , \13599 , \13601 );
xor \U$13573 ( \13888 , \13887 , \13604 );
and \U$13574 ( \13889 , \13885 , \13888 );
and \U$13575 ( \13890 , \13883 , \13888 );
or \U$13576 ( \13891 , \13886 , \13889 , \13890 );
and \U$13577 ( \13892 , \13881 , \13891 );
xor \U$13578 ( \13893 , \13281 , \13307 );
xor \U$13579 ( \13894 , \13893 , \13318 );
and \U$13580 ( \13895 , \13891 , \13894 );
and \U$13581 ( \13896 , \13881 , \13894 );
or \U$13582 ( \13897 , \13892 , \13895 , \13896 );
xor \U$13583 ( \13898 , \13613 , \13615 );
xor \U$13584 ( \13899 , \13898 , \13618 );
and \U$13585 ( \13900 , \13897 , \13899 );
and \U$13586 ( \13901 , \13627 , \13900 );
xor \U$13587 ( \13902 , \13627 , \13900 );
xor \U$13588 ( \13903 , \13897 , \13899 );
xor \U$13589 ( \13904 , \13768 , \13772 );
xor \U$13590 ( \13905 , \13904 , \13777 );
xor \U$13591 ( \13906 , \13731 , \13735 );
xor \U$13592 ( \13907 , \13906 , \13740 );
and \U$13593 ( \13908 , \13905 , \13907 );
xor \U$13594 ( \13909 , \13748 , \13752 );
xor \U$13595 ( \13910 , \13909 , \13757 );
and \U$13596 ( \13911 , \13907 , \13910 );
and \U$13597 ( \13912 , \13905 , \13910 );
or \U$13598 ( \13913 , \13908 , \13911 , \13912 );
and \U$13599 ( \13914 , \10347 , \692 );
and \U$13600 ( \13915 , \10166 , \690 );
nor \U$13601 ( \13916 , \13914 , \13915 );
xnor \U$13602 ( \13917 , \13916 , \649 );
nand \U$13603 ( \13918 , \10967 , \577 );
xnor \U$13604 ( \13919 , \13918 , \530 );
and \U$13605 ( \13920 , \13917 , \13919 );
xor \U$13606 ( \13921 , \13715 , \13719 );
xor \U$13607 ( \13922 , \13921 , \13724 );
and \U$13608 ( \13923 , \13919 , \13922 );
and \U$13609 ( \13924 , \13917 , \13922 );
or \U$13610 ( \13925 , \13920 , \13923 , \13924 );
and \U$13611 ( \13926 , \13913 , \13925 );
xor \U$13612 ( \13927 , \13667 , \13671 );
xor \U$13613 ( \13928 , \13927 , \13676 );
xor \U$13614 ( \13929 , \13784 , \13788 );
xor \U$13615 ( \13930 , \13929 , \13793 );
and \U$13616 ( \13931 , \13928 , \13930 );
xor \U$13617 ( \13932 , \13801 , \13805 );
xor \U$13618 ( \13933 , \13932 , \13810 );
and \U$13619 ( \13934 , \13930 , \13933 );
and \U$13620 ( \13935 , \13928 , \13933 );
or \U$13621 ( \13936 , \13931 , \13934 , \13935 );
and \U$13622 ( \13937 , \13925 , \13936 );
and \U$13623 ( \13938 , \13913 , \13936 );
or \U$13624 ( \13939 , \13926 , \13937 , \13938 );
and \U$13625 ( \13940 , \9558 , \996 );
and \U$13626 ( \13941 , \9550 , \994 );
nor \U$13627 ( \13942 , \13940 , \13941 );
xnor \U$13628 ( \13943 , \13942 , \902 );
and \U$13629 ( \13944 , \10166 , \826 );
and \U$13630 ( \13945 , \10161 , \824 );
nor \U$13631 ( \13946 , \13944 , \13945 );
xnor \U$13632 ( \13947 , \13946 , \754 );
and \U$13633 ( \13948 , \13943 , \13947 );
and \U$13634 ( \13949 , \10967 , \692 );
and \U$13635 ( \13950 , \10347 , \690 );
nor \U$13636 ( \13951 , \13949 , \13950 );
xnor \U$13637 ( \13952 , \13951 , \649 );
and \U$13638 ( \13953 , \13947 , \13952 );
and \U$13639 ( \13954 , \13943 , \13952 );
or \U$13640 ( \13955 , \13948 , \13953 , \13954 );
and \U$13641 ( \13956 , \6157 , \2300 );
and \U$13642 ( \13957 , \6148 , \2298 );
nor \U$13643 ( \13958 , \13956 , \13957 );
xnor \U$13644 ( \13959 , \13958 , \2163 );
and \U$13645 ( \13960 , \6702 , \2094 );
and \U$13646 ( \13961 , \6500 , \2092 );
nor \U$13647 ( \13962 , \13960 , \13961 );
xnor \U$13648 ( \13963 , \13962 , \1942 );
and \U$13649 ( \13964 , \13959 , \13963 );
and \U$13650 ( \13965 , \7177 , \1826 );
and \U$13651 ( \13966 , \7005 , \1824 );
nor \U$13652 ( \13967 , \13965 , \13966 );
xnor \U$13653 ( \13968 , \13967 , \1670 );
and \U$13654 ( \13969 , \13963 , \13968 );
and \U$13655 ( \13970 , \13959 , \13968 );
or \U$13656 ( \13971 , \13964 , \13969 , \13970 );
and \U$13657 ( \13972 , \13955 , \13971 );
and \U$13658 ( \13973 , \8127 , \1554 );
and \U$13659 ( \13974 , \7703 , \1552 );
nor \U$13660 ( \13975 , \13973 , \13974 );
xnor \U$13661 ( \13976 , \13975 , \1441 );
and \U$13662 ( \13977 , \8378 , \1360 );
and \U$13663 ( \13978 , \8373 , \1358 );
nor \U$13664 ( \13979 , \13977 , \13978 );
xnor \U$13665 ( \13980 , \13979 , \1224 );
and \U$13666 ( \13981 , \13976 , \13980 );
and \U$13667 ( \13982 , \8981 , \1160 );
and \U$13668 ( \13983 , \8697 , \1158 );
nor \U$13669 ( \13984 , \13982 , \13983 );
xnor \U$13670 ( \13985 , \13984 , \1082 );
and \U$13671 ( \13986 , \13980 , \13985 );
and \U$13672 ( \13987 , \13976 , \13985 );
or \U$13673 ( \13988 , \13981 , \13986 , \13987 );
and \U$13674 ( \13989 , \13971 , \13988 );
and \U$13675 ( \13990 , \13955 , \13988 );
or \U$13676 ( \13991 , \13972 , \13989 , \13990 );
and \U$13677 ( \13992 , \1274 , \8896 );
and \U$13678 ( \13993 , \1186 , \8894 );
nor \U$13679 ( \13994 , \13992 , \13993 );
xnor \U$13680 ( \13995 , \13994 , \8525 );
and \U$13681 ( \13996 , \1384 , \8334 );
and \U$13682 ( \13997 , \1379 , \8332 );
nor \U$13683 ( \13998 , \13996 , \13997 );
xnor \U$13684 ( \13999 , \13998 , \8016 );
and \U$13685 ( \14000 , \13995 , \13999 );
and \U$13686 ( \14001 , \1615 , \7767 );
and \U$13687 ( \14002 , \1500 , \7765 );
nor \U$13688 ( \14003 , \14001 , \14002 );
xnor \U$13689 ( \14004 , \14003 , \7518 );
and \U$13690 ( \14005 , \13999 , \14004 );
and \U$13691 ( \14006 , \13995 , \14004 );
or \U$13692 ( \14007 , \14000 , \14005 , \14006 );
and \U$13693 ( \14008 , \1799 , \7238 );
and \U$13694 ( \14009 , \1791 , \7236 );
nor \U$13695 ( \14010 , \14008 , \14009 );
xnor \U$13696 ( \14011 , \14010 , \6978 );
and \U$13697 ( \14012 , \2047 , \6744 );
and \U$13698 ( \14013 , \2042 , \6742 );
nor \U$13699 ( \14014 , \14012 , \14013 );
xnor \U$13700 ( \14015 , \14014 , \6429 );
and \U$13701 ( \14016 , \14011 , \14015 );
and \U$13702 ( \14017 , \2377 , \6235 );
and \U$13703 ( \14018 , \2233 , \6233 );
nor \U$13704 ( \14019 , \14017 , \14018 );
xnor \U$13705 ( \14020 , \14019 , \5895 );
and \U$13706 ( \14021 , \14015 , \14020 );
and \U$13707 ( \14022 , \14011 , \14020 );
or \U$13708 ( \14023 , \14016 , \14021 , \14022 );
and \U$13709 ( \14024 , \14007 , \14023 );
and \U$13710 ( \14025 , \709 , \10814 );
and \U$13711 ( \14026 , \681 , \10811 );
nor \U$13712 ( \14027 , \14025 , \14026 );
xnor \U$13713 ( \14028 , \14027 , \9759 );
and \U$13714 ( \14029 , \863 , \10001 );
and \U$13715 ( \14030 , \789 , \9999 );
nor \U$13716 ( \14031 , \14029 , \14030 );
xnor \U$13717 ( \14032 , \14031 , \9762 );
and \U$13718 ( \14033 , \14028 , \14032 );
and \U$13719 ( \14034 , \988 , \9433 );
and \U$13720 ( \14035 , \925 , \9431 );
nor \U$13721 ( \14036 , \14034 , \14035 );
xnor \U$13722 ( \14037 , \14036 , \9123 );
and \U$13723 ( \14038 , \14032 , \14037 );
and \U$13724 ( \14039 , \14028 , \14037 );
or \U$13725 ( \14040 , \14033 , \14038 , \14039 );
and \U$13726 ( \14041 , \14023 , \14040 );
and \U$13727 ( \14042 , \14007 , \14040 );
or \U$13728 ( \14043 , \14024 , \14041 , \14042 );
and \U$13729 ( \14044 , \13991 , \14043 );
and \U$13730 ( \14045 , \4779 , \3324 );
and \U$13731 ( \14046 , \4771 , \3322 );
nor \U$13732 ( \14047 , \14045 , \14046 );
xnor \U$13733 ( \14048 , \14047 , \3119 );
and \U$13734 ( \14049 , \5253 , \2918 );
and \U$13735 ( \14050 , \5248 , \2916 );
nor \U$13736 ( \14051 , \14049 , \14050 );
xnor \U$13737 ( \14052 , \14051 , \2769 );
and \U$13738 ( \14053 , \14048 , \14052 );
and \U$13739 ( \14054 , \5776 , \2596 );
and \U$13740 ( \14055 , \5517 , \2594 );
nor \U$13741 ( \14056 , \14054 , \14055 );
xnor \U$13742 ( \14057 , \14056 , \2454 );
and \U$13743 ( \14058 , \14052 , \14057 );
and \U$13744 ( \14059 , \14048 , \14057 );
or \U$13745 ( \14060 , \14053 , \14058 , \14059 );
and \U$13746 ( \14061 , \3889 , \4355 );
and \U$13747 ( \14062 , \3681 , \4353 );
nor \U$13748 ( \14063 , \14061 , \14062 );
xnor \U$13749 ( \14064 , \14063 , \4212 );
and \U$13750 ( \14065 , \4016 , \4032 );
and \U$13751 ( \14066 , \4011 , \4030 );
nor \U$13752 ( \14067 , \14065 , \14066 );
xnor \U$13753 ( \14068 , \14067 , \3786 );
and \U$13754 ( \14069 , \14064 , \14068 );
and \U$13755 ( \14070 , \4469 , \3637 );
and \U$13756 ( \14071 , \4272 , \3635 );
nor \U$13757 ( \14072 , \14070 , \14071 );
xnor \U$13758 ( \14073 , \14072 , \3450 );
and \U$13759 ( \14074 , \14068 , \14073 );
and \U$13760 ( \14075 , \14064 , \14073 );
or \U$13761 ( \14076 , \14069 , \14074 , \14075 );
and \U$13762 ( \14077 , \14060 , \14076 );
and \U$13763 ( \14078 , \2666 , \5646 );
and \U$13764 ( \14079 , \2641 , \5644 );
nor \U$13765 ( \14080 , \14078 , \14079 );
xnor \U$13766 ( \14081 , \14080 , \5405 );
and \U$13767 ( \14082 , \3007 , \5180 );
and \U$13768 ( \14083 , \2840 , \5178 );
nor \U$13769 ( \14084 , \14082 , \14083 );
xnor \U$13770 ( \14085 , \14084 , \4992 );
and \U$13771 ( \14086 , \14081 , \14085 );
and \U$13772 ( \14087 , \3264 , \4806 );
and \U$13773 ( \14088 , \3145 , \4804 );
nor \U$13774 ( \14089 , \14087 , \14088 );
xnor \U$13775 ( \14090 , \14089 , \4574 );
and \U$13776 ( \14091 , \14085 , \14090 );
and \U$13777 ( \14092 , \14081 , \14090 );
or \U$13778 ( \14093 , \14086 , \14091 , \14092 );
and \U$13779 ( \14094 , \14076 , \14093 );
and \U$13780 ( \14095 , \14060 , \14093 );
or \U$13781 ( \14096 , \14077 , \14094 , \14095 );
and \U$13782 ( \14097 , \14043 , \14096 );
and \U$13783 ( \14098 , \13991 , \14096 );
or \U$13784 ( \14099 , \14044 , \14097 , \14098 );
and \U$13785 ( \14100 , \13939 , \14099 );
xor \U$13786 ( \14101 , \13516 , \13520 );
xor \U$13787 ( \14102 , \14101 , \13525 );
xor \U$13788 ( \14103 , \13629 , \13631 );
xor \U$13789 ( \14104 , \14103 , \13634 );
and \U$13790 ( \14105 , \14102 , \14104 );
xor \U$13791 ( \14106 , \13639 , \13641 );
xor \U$13792 ( \14107 , \14106 , \13644 );
and \U$13793 ( \14108 , \14104 , \14107 );
and \U$13794 ( \14109 , \14102 , \14107 );
or \U$13795 ( \14110 , \14105 , \14108 , \14109 );
and \U$13796 ( \14111 , \14099 , \14110 );
and \U$13797 ( \14112 , \13939 , \14110 );
or \U$13798 ( \14113 , \14100 , \14111 , \14112 );
xor \U$13799 ( \14114 , \13727 , \13743 );
xor \U$13800 ( \14115 , \14114 , \13760 );
xor \U$13801 ( \14116 , \13780 , \13796 );
xor \U$13802 ( \14117 , \14116 , \13813 );
and \U$13803 ( \14118 , \14115 , \14117 );
xor \U$13804 ( \14119 , \13652 , \13654 );
xor \U$13805 ( \14120 , \14119 , \13657 );
and \U$13806 ( \14121 , \14117 , \14120 );
and \U$13807 ( \14122 , \14115 , \14120 );
or \U$13808 ( \14123 , \14118 , \14121 , \14122 );
xor \U$13809 ( \14124 , \13512 , \13528 );
xor \U$13810 ( \14125 , \14124 , \13545 );
and \U$13811 ( \14126 , \14123 , \14125 );
xor \U$13812 ( \14127 , \13835 , \13837 );
xor \U$13813 ( \14128 , \14127 , \13840 );
and \U$13814 ( \14129 , \14125 , \14128 );
and \U$13815 ( \14130 , \14123 , \14128 );
or \U$13816 ( \14131 , \14126 , \14129 , \14130 );
and \U$13817 ( \14132 , \14113 , \14131 );
xor \U$13818 ( \14133 , \13637 , \13647 );
xor \U$13819 ( \14134 , \14133 , \13660 );
xor \U$13820 ( \14135 , \13711 , \13763 );
xor \U$13821 ( \14136 , \14135 , \13816 );
and \U$13822 ( \14137 , \14134 , \14136 );
xor \U$13823 ( \14138 , \13822 , \13824 );
xor \U$13824 ( \14139 , \14138 , \13827 );
and \U$13825 ( \14140 , \14136 , \14139 );
and \U$13826 ( \14141 , \14134 , \14139 );
or \U$13827 ( \14142 , \14137 , \14140 , \14141 );
and \U$13828 ( \14143 , \14131 , \14142 );
and \U$13829 ( \14144 , \14113 , \14142 );
or \U$13830 ( \14145 , \14132 , \14143 , \14144 );
xor \U$13831 ( \14146 , \13663 , \13819 );
xor \U$13832 ( \14147 , \14146 , \13830 );
xor \U$13833 ( \14148 , \13843 , \13845 );
xor \U$13834 ( \14149 , \14148 , \13848 );
and \U$13835 ( \14150 , \14147 , \14149 );
xor \U$13836 ( \14151 , \13854 , \13856 );
xor \U$13837 ( \14152 , \14151 , \13859 );
and \U$13838 ( \14153 , \14149 , \14152 );
and \U$13839 ( \14154 , \14147 , \14152 );
or \U$13840 ( \14155 , \14150 , \14153 , \14154 );
and \U$13841 ( \14156 , \14145 , \14155 );
xor \U$13842 ( \14157 , \13867 , \13869 );
xor \U$13843 ( \14158 , \14157 , \13872 );
and \U$13844 ( \14159 , \14155 , \14158 );
and \U$13845 ( \14160 , \14145 , \14158 );
or \U$13846 ( \14161 , \14156 , \14159 , \14160 );
xor \U$13847 ( \14162 , \13865 , \13875 );
xor \U$13848 ( \14163 , \14162 , \13878 );
and \U$13849 ( \14164 , \14161 , \14163 );
xor \U$13850 ( \14165 , \13883 , \13885 );
xor \U$13851 ( \14166 , \14165 , \13888 );
and \U$13852 ( \14167 , \14163 , \14166 );
and \U$13853 ( \14168 , \14161 , \14166 );
or \U$13854 ( \14169 , \14164 , \14167 , \14168 );
xor \U$13855 ( \14170 , \13881 , \13891 );
xor \U$13856 ( \14171 , \14170 , \13894 );
and \U$13857 ( \14172 , \14169 , \14171 );
xor \U$13858 ( \14173 , \13597 , \13607 );
xor \U$13859 ( \14174 , \14173 , \13610 );
and \U$13860 ( \14175 , \14171 , \14174 );
and \U$13861 ( \14176 , \14169 , \14174 );
or \U$13862 ( \14177 , \14172 , \14175 , \14176 );
and \U$13863 ( \14178 , \13903 , \14177 );
xor \U$13864 ( \14179 , \13903 , \14177 );
xor \U$13865 ( \14180 , \14169 , \14171 );
xor \U$13866 ( \14181 , \14180 , \14174 );
xor \U$13867 ( \14182 , \14048 , \14052 );
xor \U$13868 ( \14183 , \14182 , \14057 );
xor \U$13869 ( \14184 , \14064 , \14068 );
xor \U$13870 ( \14185 , \14184 , \14073 );
and \U$13871 ( \14186 , \14183 , \14185 );
xor \U$13872 ( \14187 , \14081 , \14085 );
xor \U$13873 ( \14188 , \14187 , \14090 );
and \U$13874 ( \14189 , \14185 , \14188 );
and \U$13875 ( \14190 , \14183 , \14188 );
or \U$13876 ( \14191 , \14186 , \14189 , \14190 );
xor \U$13877 ( \14192 , \13943 , \13947 );
xor \U$13878 ( \14193 , \14192 , \13952 );
xor \U$13879 ( \14194 , \13959 , \13963 );
xor \U$13880 ( \14195 , \14194 , \13968 );
and \U$13881 ( \14196 , \14193 , \14195 );
xor \U$13882 ( \14197 , \13976 , \13980 );
xor \U$13883 ( \14198 , \14197 , \13985 );
and \U$13884 ( \14199 , \14195 , \14198 );
and \U$13885 ( \14200 , \14193 , \14198 );
or \U$13886 ( \14201 , \14196 , \14199 , \14200 );
and \U$13887 ( \14202 , \14191 , \14201 );
xor \U$13888 ( \14203 , \13995 , \13999 );
xor \U$13889 ( \14204 , \14203 , \14004 );
xor \U$13890 ( \14205 , \14011 , \14015 );
xor \U$13891 ( \14206 , \14205 , \14020 );
and \U$13892 ( \14207 , \14204 , \14206 );
xor \U$13893 ( \14208 , \14028 , \14032 );
xor \U$13894 ( \14209 , \14208 , \14037 );
and \U$13895 ( \14210 , \14206 , \14209 );
and \U$13896 ( \14211 , \14204 , \14209 );
or \U$13897 ( \14212 , \14207 , \14210 , \14211 );
and \U$13898 ( \14213 , \14201 , \14212 );
and \U$13899 ( \14214 , \14191 , \14212 );
or \U$13900 ( \14215 , \14202 , \14213 , \14214 );
and \U$13901 ( \14216 , \4771 , \3637 );
and \U$13902 ( \14217 , \4469 , \3635 );
nor \U$13903 ( \14218 , \14216 , \14217 );
xnor \U$13904 ( \14219 , \14218 , \3450 );
and \U$13905 ( \14220 , \5248 , \3324 );
and \U$13906 ( \14221 , \4779 , \3322 );
nor \U$13907 ( \14222 , \14220 , \14221 );
xnor \U$13908 ( \14223 , \14222 , \3119 );
and \U$13909 ( \14224 , \14219 , \14223 );
and \U$13910 ( \14225 , \5517 , \2918 );
and \U$13911 ( \14226 , \5253 , \2916 );
nor \U$13912 ( \14227 , \14225 , \14226 );
xnor \U$13913 ( \14228 , \14227 , \2769 );
and \U$13914 ( \14229 , \14223 , \14228 );
and \U$13915 ( \14230 , \14219 , \14228 );
or \U$13916 ( \14231 , \14224 , \14229 , \14230 );
and \U$13917 ( \14232 , \2641 , \6235 );
and \U$13918 ( \14233 , \2377 , \6233 );
nor \U$13919 ( \14234 , \14232 , \14233 );
xnor \U$13920 ( \14235 , \14234 , \5895 );
and \U$13921 ( \14236 , \2840 , \5646 );
and \U$13922 ( \14237 , \2666 , \5644 );
nor \U$13923 ( \14238 , \14236 , \14237 );
xnor \U$13924 ( \14239 , \14238 , \5405 );
and \U$13925 ( \14240 , \14235 , \14239 );
and \U$13926 ( \14241 , \3145 , \5180 );
and \U$13927 ( \14242 , \3007 , \5178 );
nor \U$13928 ( \14243 , \14241 , \14242 );
xnor \U$13929 ( \14244 , \14243 , \4992 );
and \U$13930 ( \14245 , \14239 , \14244 );
and \U$13931 ( \14246 , \14235 , \14244 );
or \U$13932 ( \14247 , \14240 , \14245 , \14246 );
and \U$13933 ( \14248 , \14231 , \14247 );
and \U$13934 ( \14249 , \3681 , \4806 );
and \U$13935 ( \14250 , \3264 , \4804 );
nor \U$13936 ( \14251 , \14249 , \14250 );
xnor \U$13937 ( \14252 , \14251 , \4574 );
and \U$13938 ( \14253 , \4011 , \4355 );
and \U$13939 ( \14254 , \3889 , \4353 );
nor \U$13940 ( \14255 , \14253 , \14254 );
xnor \U$13941 ( \14256 , \14255 , \4212 );
and \U$13942 ( \14257 , \14252 , \14256 );
and \U$13943 ( \14258 , \4272 , \4032 );
and \U$13944 ( \14259 , \4016 , \4030 );
nor \U$13945 ( \14260 , \14258 , \14259 );
xnor \U$13946 ( \14261 , \14260 , \3786 );
and \U$13947 ( \14262 , \14256 , \14261 );
and \U$13948 ( \14263 , \14252 , \14261 );
or \U$13949 ( \14264 , \14257 , \14262 , \14263 );
and \U$13950 ( \14265 , \14247 , \14264 );
and \U$13951 ( \14266 , \14231 , \14264 );
or \U$13952 ( \14267 , \14248 , \14265 , \14266 );
and \U$13953 ( \14268 , \1186 , \9433 );
and \U$13954 ( \14269 , \988 , \9431 );
nor \U$13955 ( \14270 , \14268 , \14269 );
xnor \U$13956 ( \14271 , \14270 , \9123 );
and \U$13957 ( \14272 , \1379 , \8896 );
and \U$13958 ( \14273 , \1274 , \8894 );
nor \U$13959 ( \14274 , \14272 , \14273 );
xnor \U$13960 ( \14275 , \14274 , \8525 );
and \U$13961 ( \14276 , \14271 , \14275 );
and \U$13962 ( \14277 , \1500 , \8334 );
and \U$13963 ( \14278 , \1384 , \8332 );
nor \U$13964 ( \14279 , \14277 , \14278 );
xnor \U$13965 ( \14280 , \14279 , \8016 );
and \U$13966 ( \14281 , \14275 , \14280 );
and \U$13967 ( \14282 , \14271 , \14280 );
or \U$13968 ( \14283 , \14276 , \14281 , \14282 );
and \U$13969 ( \14284 , \789 , \10814 );
and \U$13970 ( \14285 , \709 , \10811 );
nor \U$13971 ( \14286 , \14284 , \14285 );
xnor \U$13972 ( \14287 , \14286 , \9759 );
and \U$13973 ( \14288 , \925 , \10001 );
and \U$13974 ( \14289 , \863 , \9999 );
nor \U$13975 ( \14290 , \14288 , \14289 );
xnor \U$13976 ( \14291 , \14290 , \9762 );
and \U$13977 ( \14292 , \14287 , \14291 );
and \U$13978 ( \14293 , \14291 , \649 );
and \U$13979 ( \14294 , \14287 , \649 );
or \U$13980 ( \14295 , \14292 , \14293 , \14294 );
and \U$13981 ( \14296 , \14283 , \14295 );
and \U$13982 ( \14297 , \1791 , \7767 );
and \U$13983 ( \14298 , \1615 , \7765 );
nor \U$13984 ( \14299 , \14297 , \14298 );
xnor \U$13985 ( \14300 , \14299 , \7518 );
and \U$13986 ( \14301 , \2042 , \7238 );
and \U$13987 ( \14302 , \1799 , \7236 );
nor \U$13988 ( \14303 , \14301 , \14302 );
xnor \U$13989 ( \14304 , \14303 , \6978 );
and \U$13990 ( \14305 , \14300 , \14304 );
and \U$13991 ( \14306 , \2233 , \6744 );
and \U$13992 ( \14307 , \2047 , \6742 );
nor \U$13993 ( \14308 , \14306 , \14307 );
xnor \U$13994 ( \14309 , \14308 , \6429 );
and \U$13995 ( \14310 , \14304 , \14309 );
and \U$13996 ( \14311 , \14300 , \14309 );
or \U$13997 ( \14312 , \14305 , \14310 , \14311 );
and \U$13998 ( \14313 , \14295 , \14312 );
and \U$13999 ( \14314 , \14283 , \14312 );
or \U$14000 ( \14315 , \14296 , \14313 , \14314 );
and \U$14001 ( \14316 , \14267 , \14315 );
and \U$14002 ( \14317 , \9550 , \1160 );
and \U$14003 ( \14318 , \8981 , \1158 );
nor \U$14004 ( \14319 , \14317 , \14318 );
xnor \U$14005 ( \14320 , \14319 , \1082 );
and \U$14006 ( \14321 , \10161 , \996 );
and \U$14007 ( \14322 , \9558 , \994 );
nor \U$14008 ( \14323 , \14321 , \14322 );
xnor \U$14009 ( \14324 , \14323 , \902 );
and \U$14010 ( \14325 , \14320 , \14324 );
and \U$14011 ( \14326 , \10347 , \826 );
and \U$14012 ( \14327 , \10166 , \824 );
nor \U$14013 ( \14328 , \14326 , \14327 );
xnor \U$14014 ( \14329 , \14328 , \754 );
and \U$14015 ( \14330 , \14324 , \14329 );
and \U$14016 ( \14331 , \14320 , \14329 );
or \U$14017 ( \14332 , \14325 , \14330 , \14331 );
and \U$14018 ( \14333 , \6148 , \2596 );
and \U$14019 ( \14334 , \5776 , \2594 );
nor \U$14020 ( \14335 , \14333 , \14334 );
xnor \U$14021 ( \14336 , \14335 , \2454 );
and \U$14022 ( \14337 , \6500 , \2300 );
and \U$14023 ( \14338 , \6157 , \2298 );
nor \U$14024 ( \14339 , \14337 , \14338 );
xnor \U$14025 ( \14340 , \14339 , \2163 );
and \U$14026 ( \14341 , \14336 , \14340 );
and \U$14027 ( \14342 , \7005 , \2094 );
and \U$14028 ( \14343 , \6702 , \2092 );
nor \U$14029 ( \14344 , \14342 , \14343 );
xnor \U$14030 ( \14345 , \14344 , \1942 );
and \U$14031 ( \14346 , \14340 , \14345 );
and \U$14032 ( \14347 , \14336 , \14345 );
or \U$14033 ( \14348 , \14341 , \14346 , \14347 );
and \U$14034 ( \14349 , \14332 , \14348 );
and \U$14035 ( \14350 , \7703 , \1826 );
and \U$14036 ( \14351 , \7177 , \1824 );
nor \U$14037 ( \14352 , \14350 , \14351 );
xnor \U$14038 ( \14353 , \14352 , \1670 );
and \U$14039 ( \14354 , \8373 , \1554 );
and \U$14040 ( \14355 , \8127 , \1552 );
nor \U$14041 ( \14356 , \14354 , \14355 );
xnor \U$14042 ( \14357 , \14356 , \1441 );
and \U$14043 ( \14358 , \14353 , \14357 );
and \U$14044 ( \14359 , \8697 , \1360 );
and \U$14045 ( \14360 , \8378 , \1358 );
nor \U$14046 ( \14361 , \14359 , \14360 );
xnor \U$14047 ( \14362 , \14361 , \1224 );
and \U$14048 ( \14363 , \14357 , \14362 );
and \U$14049 ( \14364 , \14353 , \14362 );
or \U$14050 ( \14365 , \14358 , \14363 , \14364 );
and \U$14051 ( \14366 , \14348 , \14365 );
and \U$14052 ( \14367 , \14332 , \14365 );
or \U$14053 ( \14368 , \14349 , \14366 , \14367 );
and \U$14054 ( \14369 , \14315 , \14368 );
and \U$14055 ( \14370 , \14267 , \14368 );
or \U$14056 ( \14371 , \14316 , \14369 , \14370 );
and \U$14057 ( \14372 , \14215 , \14371 );
xor \U$14058 ( \14373 , \13683 , \13687 );
xor \U$14059 ( \14374 , \14373 , \13692 );
xor \U$14060 ( \14375 , \13700 , \13704 );
xor \U$14061 ( \14376 , \14375 , \530 );
and \U$14062 ( \14377 , \14374 , \14376 );
xor \U$14063 ( \14378 , \13928 , \13930 );
xor \U$14064 ( \14379 , \14378 , \13933 );
and \U$14065 ( \14380 , \14376 , \14379 );
and \U$14066 ( \14381 , \14374 , \14379 );
or \U$14067 ( \14382 , \14377 , \14380 , \14381 );
and \U$14068 ( \14383 , \14371 , \14382 );
and \U$14069 ( \14384 , \14215 , \14382 );
or \U$14070 ( \14385 , \14372 , \14383 , \14384 );
xor \U$14071 ( \14386 , \13955 , \13971 );
xor \U$14072 ( \14387 , \14386 , \13988 );
xor \U$14073 ( \14388 , \13905 , \13907 );
xor \U$14074 ( \14389 , \14388 , \13910 );
and \U$14075 ( \14390 , \14387 , \14389 );
xor \U$14076 ( \14391 , \13917 , \13919 );
xor \U$14077 ( \14392 , \14391 , \13922 );
and \U$14078 ( \14393 , \14389 , \14392 );
and \U$14079 ( \14394 , \14387 , \14392 );
or \U$14080 ( \14395 , \14390 , \14393 , \14394 );
xor \U$14081 ( \14396 , \14007 , \14023 );
xor \U$14082 ( \14397 , \14396 , \14040 );
xor \U$14083 ( \14398 , \14060 , \14076 );
xor \U$14084 ( \14399 , \14398 , \14093 );
and \U$14085 ( \14400 , \14397 , \14399 );
and \U$14086 ( \14401 , \14395 , \14400 );
xor \U$14087 ( \14402 , \13679 , \13695 );
xor \U$14088 ( \14403 , \14402 , \13708 );
and \U$14089 ( \14404 , \14400 , \14403 );
and \U$14090 ( \14405 , \14395 , \14403 );
or \U$14091 ( \14406 , \14401 , \14404 , \14405 );
and \U$14092 ( \14407 , \14385 , \14406 );
xor \U$14093 ( \14408 , \13913 , \13925 );
xor \U$14094 ( \14409 , \14408 , \13936 );
xor \U$14095 ( \14410 , \14115 , \14117 );
xor \U$14096 ( \14411 , \14410 , \14120 );
and \U$14097 ( \14412 , \14409 , \14411 );
xor \U$14098 ( \14413 , \14102 , \14104 );
xor \U$14099 ( \14414 , \14413 , \14107 );
and \U$14100 ( \14415 , \14411 , \14414 );
and \U$14101 ( \14416 , \14409 , \14414 );
or \U$14102 ( \14417 , \14412 , \14415 , \14416 );
and \U$14103 ( \14418 , \14406 , \14417 );
and \U$14104 ( \14419 , \14385 , \14417 );
or \U$14105 ( \14420 , \14407 , \14418 , \14419 );
xor \U$14106 ( \14421 , \13939 , \14099 );
xor \U$14107 ( \14422 , \14421 , \14110 );
xor \U$14108 ( \14423 , \14123 , \14125 );
xor \U$14109 ( \14424 , \14423 , \14128 );
and \U$14110 ( \14425 , \14422 , \14424 );
xor \U$14111 ( \14426 , \14134 , \14136 );
xor \U$14112 ( \14427 , \14426 , \14139 );
and \U$14113 ( \14428 , \14424 , \14427 );
and \U$14114 ( \14429 , \14422 , \14427 );
or \U$14115 ( \14430 , \14425 , \14428 , \14429 );
and \U$14116 ( \14431 , \14420 , \14430 );
xor \U$14117 ( \14432 , \14147 , \14149 );
xor \U$14118 ( \14433 , \14432 , \14152 );
and \U$14119 ( \14434 , \14430 , \14433 );
and \U$14120 ( \14435 , \14420 , \14433 );
or \U$14121 ( \14436 , \14431 , \14434 , \14435 );
xor \U$14122 ( \14437 , \13833 , \13851 );
xor \U$14123 ( \14438 , \14437 , \13862 );
and \U$14124 ( \14439 , \14436 , \14438 );
xor \U$14125 ( \14440 , \14145 , \14155 );
xor \U$14126 ( \14441 , \14440 , \14158 );
and \U$14127 ( \14442 , \14438 , \14441 );
and \U$14128 ( \14443 , \14436 , \14441 );
or \U$14129 ( \14444 , \14439 , \14442 , \14443 );
xor \U$14130 ( \14445 , \14161 , \14163 );
xor \U$14131 ( \14446 , \14445 , \14166 );
and \U$14132 ( \14447 , \14444 , \14446 );
and \U$14133 ( \14448 , \14181 , \14447 );
xor \U$14134 ( \14449 , \14181 , \14447 );
xor \U$14135 ( \14450 , \14444 , \14446 );
and \U$14136 ( \14451 , \4016 , \4355 );
and \U$14137 ( \14452 , \4011 , \4353 );
nor \U$14138 ( \14453 , \14451 , \14452 );
xnor \U$14139 ( \14454 , \14453 , \4212 );
and \U$14140 ( \14455 , \4469 , \4032 );
and \U$14141 ( \14456 , \4272 , \4030 );
nor \U$14142 ( \14457 , \14455 , \14456 );
xnor \U$14143 ( \14458 , \14457 , \3786 );
and \U$14144 ( \14459 , \14454 , \14458 );
and \U$14145 ( \14460 , \4779 , \3637 );
and \U$14146 ( \14461 , \4771 , \3635 );
nor \U$14147 ( \14462 , \14460 , \14461 );
xnor \U$14148 ( \14463 , \14462 , \3450 );
and \U$14149 ( \14464 , \14458 , \14463 );
and \U$14150 ( \14465 , \14454 , \14463 );
or \U$14151 ( \14466 , \14459 , \14464 , \14465 );
and \U$14152 ( \14467 , \3007 , \5646 );
and \U$14153 ( \14468 , \2840 , \5644 );
nor \U$14154 ( \14469 , \14467 , \14468 );
xnor \U$14155 ( \14470 , \14469 , \5405 );
and \U$14156 ( \14471 , \3264 , \5180 );
and \U$14157 ( \14472 , \3145 , \5178 );
nor \U$14158 ( \14473 , \14471 , \14472 );
xnor \U$14159 ( \14474 , \14473 , \4992 );
and \U$14160 ( \14475 , \14470 , \14474 );
and \U$14161 ( \14476 , \3889 , \4806 );
and \U$14162 ( \14477 , \3681 , \4804 );
nor \U$14163 ( \14478 , \14476 , \14477 );
xnor \U$14164 ( \14479 , \14478 , \4574 );
and \U$14165 ( \14480 , \14474 , \14479 );
and \U$14166 ( \14481 , \14470 , \14479 );
or \U$14167 ( \14482 , \14475 , \14480 , \14481 );
and \U$14168 ( \14483 , \14466 , \14482 );
and \U$14169 ( \14484 , \5253 , \3324 );
and \U$14170 ( \14485 , \5248 , \3322 );
nor \U$14171 ( \14486 , \14484 , \14485 );
xnor \U$14172 ( \14487 , \14486 , \3119 );
and \U$14173 ( \14488 , \5776 , \2918 );
and \U$14174 ( \14489 , \5517 , \2916 );
nor \U$14175 ( \14490 , \14488 , \14489 );
xnor \U$14176 ( \14491 , \14490 , \2769 );
and \U$14177 ( \14492 , \14487 , \14491 );
and \U$14178 ( \14493 , \6157 , \2596 );
and \U$14179 ( \14494 , \6148 , \2594 );
nor \U$14180 ( \14495 , \14493 , \14494 );
xnor \U$14181 ( \14496 , \14495 , \2454 );
and \U$14182 ( \14497 , \14491 , \14496 );
and \U$14183 ( \14498 , \14487 , \14496 );
or \U$14184 ( \14499 , \14492 , \14497 , \14498 );
and \U$14185 ( \14500 , \14482 , \14499 );
and \U$14186 ( \14501 , \14466 , \14499 );
or \U$14187 ( \14502 , \14483 , \14500 , \14501 );
and \U$14188 ( \14503 , \8378 , \1554 );
and \U$14189 ( \14504 , \8373 , \1552 );
nor \U$14190 ( \14505 , \14503 , \14504 );
xnor \U$14191 ( \14506 , \14505 , \1441 );
and \U$14192 ( \14507 , \8981 , \1360 );
and \U$14193 ( \14508 , \8697 , \1358 );
nor \U$14194 ( \14509 , \14507 , \14508 );
xnor \U$14195 ( \14510 , \14509 , \1224 );
and \U$14196 ( \14511 , \14506 , \14510 );
and \U$14197 ( \14512 , \9558 , \1160 );
and \U$14198 ( \14513 , \9550 , \1158 );
nor \U$14199 ( \14514 , \14512 , \14513 );
xnor \U$14200 ( \14515 , \14514 , \1082 );
and \U$14201 ( \14516 , \14510 , \14515 );
and \U$14202 ( \14517 , \14506 , \14515 );
or \U$14203 ( \14518 , \14511 , \14516 , \14517 );
and \U$14204 ( \14519 , \6702 , \2300 );
and \U$14205 ( \14520 , \6500 , \2298 );
nor \U$14206 ( \14521 , \14519 , \14520 );
xnor \U$14207 ( \14522 , \14521 , \2163 );
and \U$14208 ( \14523 , \7177 , \2094 );
and \U$14209 ( \14524 , \7005 , \2092 );
nor \U$14210 ( \14525 , \14523 , \14524 );
xnor \U$14211 ( \14526 , \14525 , \1942 );
and \U$14212 ( \14527 , \14522 , \14526 );
and \U$14213 ( \14528 , \8127 , \1826 );
and \U$14214 ( \14529 , \7703 , \1824 );
nor \U$14215 ( \14530 , \14528 , \14529 );
xnor \U$14216 ( \14531 , \14530 , \1670 );
and \U$14217 ( \14532 , \14526 , \14531 );
and \U$14218 ( \14533 , \14522 , \14531 );
or \U$14219 ( \14534 , \14527 , \14532 , \14533 );
and \U$14220 ( \14535 , \14518 , \14534 );
and \U$14221 ( \14536 , \10166 , \996 );
and \U$14222 ( \14537 , \10161 , \994 );
nor \U$14223 ( \14538 , \14536 , \14537 );
xnor \U$14224 ( \14539 , \14538 , \902 );
and \U$14225 ( \14540 , \10967 , \826 );
and \U$14226 ( \14541 , \10347 , \824 );
nor \U$14227 ( \14542 , \14540 , \14541 );
xnor \U$14228 ( \14543 , \14542 , \754 );
and \U$14229 ( \14544 , \14539 , \14543 );
and \U$14230 ( \14545 , \14534 , \14544 );
and \U$14231 ( \14546 , \14518 , \14544 );
or \U$14232 ( \14547 , \14535 , \14545 , \14546 );
and \U$14233 ( \14548 , \14502 , \14547 );
and \U$14234 ( \14549 , \2047 , \7238 );
and \U$14235 ( \14550 , \2042 , \7236 );
nor \U$14236 ( \14551 , \14549 , \14550 );
xnor \U$14237 ( \14552 , \14551 , \6978 );
and \U$14238 ( \14553 , \2377 , \6744 );
and \U$14239 ( \14554 , \2233 , \6742 );
nor \U$14240 ( \14555 , \14553 , \14554 );
xnor \U$14241 ( \14556 , \14555 , \6429 );
and \U$14242 ( \14557 , \14552 , \14556 );
and \U$14243 ( \14558 , \2666 , \6235 );
and \U$14244 ( \14559 , \2641 , \6233 );
nor \U$14245 ( \14560 , \14558 , \14559 );
xnor \U$14246 ( \14561 , \14560 , \5895 );
and \U$14247 ( \14562 , \14556 , \14561 );
and \U$14248 ( \14563 , \14552 , \14561 );
or \U$14249 ( \14564 , \14557 , \14562 , \14563 );
and \U$14250 ( \14565 , \863 , \10814 );
and \U$14251 ( \14566 , \789 , \10811 );
nor \U$14252 ( \14567 , \14565 , \14566 );
xnor \U$14253 ( \14568 , \14567 , \9759 );
and \U$14254 ( \14569 , \988 , \10001 );
and \U$14255 ( \14570 , \925 , \9999 );
nor \U$14256 ( \14571 , \14569 , \14570 );
xnor \U$14257 ( \14572 , \14571 , \9762 );
and \U$14258 ( \14573 , \14568 , \14572 );
and \U$14259 ( \14574 , \1274 , \9433 );
and \U$14260 ( \14575 , \1186 , \9431 );
nor \U$14261 ( \14576 , \14574 , \14575 );
xnor \U$14262 ( \14577 , \14576 , \9123 );
and \U$14263 ( \14578 , \14572 , \14577 );
and \U$14264 ( \14579 , \14568 , \14577 );
or \U$14265 ( \14580 , \14573 , \14578 , \14579 );
and \U$14266 ( \14581 , \14564 , \14580 );
and \U$14267 ( \14582 , \1384 , \8896 );
and \U$14268 ( \14583 , \1379 , \8894 );
nor \U$14269 ( \14584 , \14582 , \14583 );
xnor \U$14270 ( \14585 , \14584 , \8525 );
and \U$14271 ( \14586 , \1615 , \8334 );
and \U$14272 ( \14587 , \1500 , \8332 );
nor \U$14273 ( \14588 , \14586 , \14587 );
xnor \U$14274 ( \14589 , \14588 , \8016 );
and \U$14275 ( \14590 , \14585 , \14589 );
and \U$14276 ( \14591 , \1799 , \7767 );
and \U$14277 ( \14592 , \1791 , \7765 );
nor \U$14278 ( \14593 , \14591 , \14592 );
xnor \U$14279 ( \14594 , \14593 , \7518 );
and \U$14280 ( \14595 , \14589 , \14594 );
and \U$14281 ( \14596 , \14585 , \14594 );
or \U$14282 ( \14597 , \14590 , \14595 , \14596 );
and \U$14283 ( \14598 , \14580 , \14597 );
and \U$14284 ( \14599 , \14564 , \14597 );
or \U$14285 ( \14600 , \14581 , \14598 , \14599 );
and \U$14286 ( \14601 , \14547 , \14600 );
and \U$14287 ( \14602 , \14502 , \14600 );
or \U$14288 ( \14603 , \14548 , \14601 , \14602 );
xor \U$14289 ( \14604 , \14271 , \14275 );
xor \U$14290 ( \14605 , \14604 , \14280 );
xor \U$14291 ( \14606 , \14300 , \14304 );
xor \U$14292 ( \14607 , \14606 , \14309 );
and \U$14293 ( \14608 , \14605 , \14607 );
xor \U$14294 ( \14609 , \14235 , \14239 );
xor \U$14295 ( \14610 , \14609 , \14244 );
and \U$14296 ( \14611 , \14607 , \14610 );
and \U$14297 ( \14612 , \14605 , \14610 );
or \U$14298 ( \14613 , \14608 , \14611 , \14612 );
nand \U$14299 ( \14614 , \10967 , \690 );
xnor \U$14300 ( \14615 , \14614 , \649 );
xor \U$14301 ( \14616 , \14320 , \14324 );
xor \U$14302 ( \14617 , \14616 , \14329 );
and \U$14303 ( \14618 , \14615 , \14617 );
xor \U$14304 ( \14619 , \14353 , \14357 );
xor \U$14305 ( \14620 , \14619 , \14362 );
and \U$14306 ( \14621 , \14617 , \14620 );
and \U$14307 ( \14622 , \14615 , \14620 );
or \U$14308 ( \14623 , \14618 , \14621 , \14622 );
and \U$14309 ( \14624 , \14613 , \14623 );
xor \U$14310 ( \14625 , \14336 , \14340 );
xor \U$14311 ( \14626 , \14625 , \14345 );
xor \U$14312 ( \14627 , \14219 , \14223 );
xor \U$14313 ( \14628 , \14627 , \14228 );
and \U$14314 ( \14629 , \14626 , \14628 );
xor \U$14315 ( \14630 , \14252 , \14256 );
xor \U$14316 ( \14631 , \14630 , \14261 );
and \U$14317 ( \14632 , \14628 , \14631 );
and \U$14318 ( \14633 , \14626 , \14631 );
or \U$14319 ( \14634 , \14629 , \14632 , \14633 );
and \U$14320 ( \14635 , \14623 , \14634 );
and \U$14321 ( \14636 , \14613 , \14634 );
or \U$14322 ( \14637 , \14624 , \14635 , \14636 );
and \U$14323 ( \14638 , \14603 , \14637 );
xor \U$14324 ( \14639 , \14183 , \14185 );
xor \U$14325 ( \14640 , \14639 , \14188 );
xor \U$14326 ( \14641 , \14193 , \14195 );
xor \U$14327 ( \14642 , \14641 , \14198 );
and \U$14328 ( \14643 , \14640 , \14642 );
xor \U$14329 ( \14644 , \14204 , \14206 );
xor \U$14330 ( \14645 , \14644 , \14209 );
and \U$14331 ( \14646 , \14642 , \14645 );
and \U$14332 ( \14647 , \14640 , \14645 );
or \U$14333 ( \14648 , \14643 , \14646 , \14647 );
and \U$14334 ( \14649 , \14637 , \14648 );
and \U$14335 ( \14650 , \14603 , \14648 );
or \U$14336 ( \14651 , \14638 , \14649 , \14650 );
xor \U$14337 ( \14652 , \14191 , \14201 );
xor \U$14338 ( \14653 , \14652 , \14212 );
xor \U$14339 ( \14654 , \14267 , \14315 );
xor \U$14340 ( \14655 , \14654 , \14368 );
and \U$14341 ( \14656 , \14653 , \14655 );
xor \U$14342 ( \14657 , \14374 , \14376 );
xor \U$14343 ( \14658 , \14657 , \14379 );
and \U$14344 ( \14659 , \14655 , \14658 );
and \U$14345 ( \14660 , \14653 , \14658 );
or \U$14346 ( \14661 , \14656 , \14659 , \14660 );
and \U$14347 ( \14662 , \14651 , \14661 );
xor \U$14348 ( \14663 , \14231 , \14247 );
xor \U$14349 ( \14664 , \14663 , \14264 );
xor \U$14350 ( \14665 , \14283 , \14295 );
xor \U$14351 ( \14666 , \14665 , \14312 );
and \U$14352 ( \14667 , \14664 , \14666 );
xor \U$14353 ( \14668 , \14332 , \14348 );
xor \U$14354 ( \14669 , \14668 , \14365 );
and \U$14355 ( \14670 , \14666 , \14669 );
and \U$14356 ( \14671 , \14664 , \14669 );
or \U$14357 ( \14672 , \14667 , \14670 , \14671 );
xor \U$14358 ( \14673 , \14387 , \14389 );
xor \U$14359 ( \14674 , \14673 , \14392 );
and \U$14360 ( \14675 , \14672 , \14674 );
xor \U$14361 ( \14676 , \14397 , \14399 );
and \U$14362 ( \14677 , \14674 , \14676 );
and \U$14363 ( \14678 , \14672 , \14676 );
or \U$14364 ( \14679 , \14675 , \14677 , \14678 );
and \U$14365 ( \14680 , \14661 , \14679 );
and \U$14366 ( \14681 , \14651 , \14679 );
or \U$14367 ( \14682 , \14662 , \14680 , \14681 );
xor \U$14368 ( \14683 , \13991 , \14043 );
xor \U$14369 ( \14684 , \14683 , \14096 );
xor \U$14370 ( \14685 , \14395 , \14400 );
xor \U$14371 ( \14686 , \14685 , \14403 );
and \U$14372 ( \14687 , \14684 , \14686 );
xor \U$14373 ( \14688 , \14409 , \14411 );
xor \U$14374 ( \14689 , \14688 , \14414 );
and \U$14375 ( \14690 , \14686 , \14689 );
and \U$14376 ( \14691 , \14684 , \14689 );
or \U$14377 ( \14692 , \14687 , \14690 , \14691 );
and \U$14378 ( \14693 , \14682 , \14692 );
xor \U$14379 ( \14694 , \14422 , \14424 );
xor \U$14380 ( \14695 , \14694 , \14427 );
and \U$14381 ( \14696 , \14692 , \14695 );
and \U$14382 ( \14697 , \14682 , \14695 );
or \U$14383 ( \14698 , \14693 , \14696 , \14697 );
xor \U$14384 ( \14699 , \14113 , \14131 );
xor \U$14385 ( \14700 , \14699 , \14142 );
and \U$14386 ( \14701 , \14698 , \14700 );
xor \U$14387 ( \14702 , \14420 , \14430 );
xor \U$14388 ( \14703 , \14702 , \14433 );
and \U$14389 ( \14704 , \14700 , \14703 );
and \U$14390 ( \14705 , \14698 , \14703 );
or \U$14391 ( \14706 , \14701 , \14704 , \14705 );
xor \U$14392 ( \14707 , \14436 , \14438 );
xor \U$14393 ( \14708 , \14707 , \14441 );
and \U$14394 ( \14709 , \14706 , \14708 );
and \U$14395 ( \14710 , \14450 , \14709 );
xor \U$14396 ( \14711 , \14450 , \14709 );
xor \U$14397 ( \14712 , \14706 , \14708 );
and \U$14398 ( \14713 , \4011 , \4806 );
and \U$14399 ( \14714 , \3889 , \4804 );
nor \U$14400 ( \14715 , \14713 , \14714 );
xnor \U$14401 ( \14716 , \14715 , \4574 );
and \U$14402 ( \14717 , \4272 , \4355 );
and \U$14403 ( \14718 , \4016 , \4353 );
nor \U$14404 ( \14719 , \14717 , \14718 );
xnor \U$14405 ( \14720 , \14719 , \4212 );
and \U$14406 ( \14721 , \14716 , \14720 );
and \U$14407 ( \14722 , \4771 , \4032 );
and \U$14408 ( \14723 , \4469 , \4030 );
nor \U$14409 ( \14724 , \14722 , \14723 );
xnor \U$14410 ( \14725 , \14724 , \3786 );
and \U$14411 ( \14726 , \14720 , \14725 );
and \U$14412 ( \14727 , \14716 , \14725 );
or \U$14413 ( \14728 , \14721 , \14726 , \14727 );
and \U$14414 ( \14729 , \2840 , \6235 );
and \U$14415 ( \14730 , \2666 , \6233 );
nor \U$14416 ( \14731 , \14729 , \14730 );
xnor \U$14417 ( \14732 , \14731 , \5895 );
and \U$14418 ( \14733 , \3145 , \5646 );
and \U$14419 ( \14734 , \3007 , \5644 );
nor \U$14420 ( \14735 , \14733 , \14734 );
xnor \U$14421 ( \14736 , \14735 , \5405 );
and \U$14422 ( \14737 , \14732 , \14736 );
and \U$14423 ( \14738 , \3681 , \5180 );
and \U$14424 ( \14739 , \3264 , \5178 );
nor \U$14425 ( \14740 , \14738 , \14739 );
xnor \U$14426 ( \14741 , \14740 , \4992 );
and \U$14427 ( \14742 , \14736 , \14741 );
and \U$14428 ( \14743 , \14732 , \14741 );
or \U$14429 ( \14744 , \14737 , \14742 , \14743 );
and \U$14430 ( \14745 , \14728 , \14744 );
and \U$14431 ( \14746 , \5248 , \3637 );
and \U$14432 ( \14747 , \4779 , \3635 );
nor \U$14433 ( \14748 , \14746 , \14747 );
xnor \U$14434 ( \14749 , \14748 , \3450 );
and \U$14435 ( \14750 , \5517 , \3324 );
and \U$14436 ( \14751 , \5253 , \3322 );
nor \U$14437 ( \14752 , \14750 , \14751 );
xnor \U$14438 ( \14753 , \14752 , \3119 );
and \U$14439 ( \14754 , \14749 , \14753 );
and \U$14440 ( \14755 , \6148 , \2918 );
and \U$14441 ( \14756 , \5776 , \2916 );
nor \U$14442 ( \14757 , \14755 , \14756 );
xnor \U$14443 ( \14758 , \14757 , \2769 );
and \U$14444 ( \14759 , \14753 , \14758 );
and \U$14445 ( \14760 , \14749 , \14758 );
or \U$14446 ( \14761 , \14754 , \14759 , \14760 );
and \U$14447 ( \14762 , \14744 , \14761 );
and \U$14448 ( \14763 , \14728 , \14761 );
or \U$14449 ( \14764 , \14745 , \14762 , \14763 );
and \U$14450 ( \14765 , \2042 , \7767 );
and \U$14451 ( \14766 , \1799 , \7765 );
nor \U$14452 ( \14767 , \14765 , \14766 );
xnor \U$14453 ( \14768 , \14767 , \7518 );
and \U$14454 ( \14769 , \2233 , \7238 );
and \U$14455 ( \14770 , \2047 , \7236 );
nor \U$14456 ( \14771 , \14769 , \14770 );
xnor \U$14457 ( \14772 , \14771 , \6978 );
and \U$14458 ( \14773 , \14768 , \14772 );
and \U$14459 ( \14774 , \2641 , \6744 );
and \U$14460 ( \14775 , \2377 , \6742 );
nor \U$14461 ( \14776 , \14774 , \14775 );
xnor \U$14462 ( \14777 , \14776 , \6429 );
and \U$14463 ( \14778 , \14772 , \14777 );
and \U$14464 ( \14779 , \14768 , \14777 );
or \U$14465 ( \14780 , \14773 , \14778 , \14779 );
and \U$14466 ( \14781 , \1379 , \9433 );
and \U$14467 ( \14782 , \1274 , \9431 );
nor \U$14468 ( \14783 , \14781 , \14782 );
xnor \U$14469 ( \14784 , \14783 , \9123 );
and \U$14470 ( \14785 , \1500 , \8896 );
and \U$14471 ( \14786 , \1384 , \8894 );
nor \U$14472 ( \14787 , \14785 , \14786 );
xnor \U$14473 ( \14788 , \14787 , \8525 );
and \U$14474 ( \14789 , \14784 , \14788 );
and \U$14475 ( \14790 , \1791 , \8334 );
and \U$14476 ( \14791 , \1615 , \8332 );
nor \U$14477 ( \14792 , \14790 , \14791 );
xnor \U$14478 ( \14793 , \14792 , \8016 );
and \U$14479 ( \14794 , \14788 , \14793 );
and \U$14480 ( \14795 , \14784 , \14793 );
or \U$14481 ( \14796 , \14789 , \14794 , \14795 );
and \U$14482 ( \14797 , \14780 , \14796 );
and \U$14483 ( \14798 , \925 , \10814 );
and \U$14484 ( \14799 , \863 , \10811 );
nor \U$14485 ( \14800 , \14798 , \14799 );
xnor \U$14486 ( \14801 , \14800 , \9759 );
and \U$14487 ( \14802 , \1186 , \10001 );
and \U$14488 ( \14803 , \988 , \9999 );
nor \U$14489 ( \14804 , \14802 , \14803 );
xnor \U$14490 ( \14805 , \14804 , \9762 );
and \U$14491 ( \14806 , \14801 , \14805 );
and \U$14492 ( \14807 , \14805 , \754 );
and \U$14493 ( \14808 , \14801 , \754 );
or \U$14494 ( \14809 , \14806 , \14807 , \14808 );
and \U$14495 ( \14810 , \14796 , \14809 );
and \U$14496 ( \14811 , \14780 , \14809 );
or \U$14497 ( \14812 , \14797 , \14810 , \14811 );
and \U$14498 ( \14813 , \14764 , \14812 );
and \U$14499 ( \14814 , \6500 , \2596 );
and \U$14500 ( \14815 , \6157 , \2594 );
nor \U$14501 ( \14816 , \14814 , \14815 );
xnor \U$14502 ( \14817 , \14816 , \2454 );
and \U$14503 ( \14818 , \7005 , \2300 );
and \U$14504 ( \14819 , \6702 , \2298 );
nor \U$14505 ( \14820 , \14818 , \14819 );
xnor \U$14506 ( \14821 , \14820 , \2163 );
and \U$14507 ( \14822 , \14817 , \14821 );
and \U$14508 ( \14823 , \7703 , \2094 );
and \U$14509 ( \14824 , \7177 , \2092 );
nor \U$14510 ( \14825 , \14823 , \14824 );
xnor \U$14511 ( \14826 , \14825 , \1942 );
and \U$14512 ( \14827 , \14821 , \14826 );
and \U$14513 ( \14828 , \14817 , \14826 );
or \U$14514 ( \14829 , \14822 , \14827 , \14828 );
and \U$14515 ( \14830 , \10161 , \1160 );
and \U$14516 ( \14831 , \9558 , \1158 );
nor \U$14517 ( \14832 , \14830 , \14831 );
xnor \U$14518 ( \14833 , \14832 , \1082 );
and \U$14519 ( \14834 , \10347 , \996 );
and \U$14520 ( \14835 , \10166 , \994 );
nor \U$14521 ( \14836 , \14834 , \14835 );
xnor \U$14522 ( \14837 , \14836 , \902 );
and \U$14523 ( \14838 , \14833 , \14837 );
nand \U$14524 ( \14839 , \10967 , \824 );
xnor \U$14525 ( \14840 , \14839 , \754 );
and \U$14526 ( \14841 , \14837 , \14840 );
and \U$14527 ( \14842 , \14833 , \14840 );
or \U$14528 ( \14843 , \14838 , \14841 , \14842 );
and \U$14529 ( \14844 , \14829 , \14843 );
and \U$14530 ( \14845 , \8373 , \1826 );
and \U$14531 ( \14846 , \8127 , \1824 );
nor \U$14532 ( \14847 , \14845 , \14846 );
xnor \U$14533 ( \14848 , \14847 , \1670 );
and \U$14534 ( \14849 , \8697 , \1554 );
and \U$14535 ( \14850 , \8378 , \1552 );
nor \U$14536 ( \14851 , \14849 , \14850 );
xnor \U$14537 ( \14852 , \14851 , \1441 );
and \U$14538 ( \14853 , \14848 , \14852 );
and \U$14539 ( \14854 , \9550 , \1360 );
and \U$14540 ( \14855 , \8981 , \1358 );
nor \U$14541 ( \14856 , \14854 , \14855 );
xnor \U$14542 ( \14857 , \14856 , \1224 );
and \U$14543 ( \14858 , \14852 , \14857 );
and \U$14544 ( \14859 , \14848 , \14857 );
or \U$14545 ( \14860 , \14853 , \14858 , \14859 );
and \U$14546 ( \14861 , \14843 , \14860 );
and \U$14547 ( \14862 , \14829 , \14860 );
or \U$14548 ( \14863 , \14844 , \14861 , \14862 );
and \U$14549 ( \14864 , \14812 , \14863 );
and \U$14550 ( \14865 , \14764 , \14863 );
or \U$14551 ( \14866 , \14813 , \14864 , \14865 );
xor \U$14552 ( \14867 , \14552 , \14556 );
xor \U$14553 ( \14868 , \14867 , \14561 );
xor \U$14554 ( \14869 , \14568 , \14572 );
xor \U$14555 ( \14870 , \14869 , \14577 );
and \U$14556 ( \14871 , \14868 , \14870 );
xor \U$14557 ( \14872 , \14585 , \14589 );
xor \U$14558 ( \14873 , \14872 , \14594 );
and \U$14559 ( \14874 , \14870 , \14873 );
and \U$14560 ( \14875 , \14868 , \14873 );
or \U$14561 ( \14876 , \14871 , \14874 , \14875 );
xor \U$14562 ( \14877 , \14454 , \14458 );
xor \U$14563 ( \14878 , \14877 , \14463 );
xor \U$14564 ( \14879 , \14470 , \14474 );
xor \U$14565 ( \14880 , \14879 , \14479 );
and \U$14566 ( \14881 , \14878 , \14880 );
xor \U$14567 ( \14882 , \14487 , \14491 );
xor \U$14568 ( \14883 , \14882 , \14496 );
and \U$14569 ( \14884 , \14880 , \14883 );
and \U$14570 ( \14885 , \14878 , \14883 );
or \U$14571 ( \14886 , \14881 , \14884 , \14885 );
and \U$14572 ( \14887 , \14876 , \14886 );
xor \U$14573 ( \14888 , \14506 , \14510 );
xor \U$14574 ( \14889 , \14888 , \14515 );
xor \U$14575 ( \14890 , \14522 , \14526 );
xor \U$14576 ( \14891 , \14890 , \14531 );
and \U$14577 ( \14892 , \14889 , \14891 );
xor \U$14578 ( \14893 , \14539 , \14543 );
and \U$14579 ( \14894 , \14891 , \14893 );
and \U$14580 ( \14895 , \14889 , \14893 );
or \U$14581 ( \14896 , \14892 , \14894 , \14895 );
and \U$14582 ( \14897 , \14886 , \14896 );
and \U$14583 ( \14898 , \14876 , \14896 );
or \U$14584 ( \14899 , \14887 , \14897 , \14898 );
and \U$14585 ( \14900 , \14866 , \14899 );
xor \U$14586 ( \14901 , \14287 , \14291 );
xor \U$14587 ( \14902 , \14901 , \649 );
xor \U$14588 ( \14903 , \14605 , \14607 );
xor \U$14589 ( \14904 , \14903 , \14610 );
and \U$14590 ( \14905 , \14902 , \14904 );
xor \U$14591 ( \14906 , \14626 , \14628 );
xor \U$14592 ( \14907 , \14906 , \14631 );
and \U$14593 ( \14908 , \14904 , \14907 );
and \U$14594 ( \14909 , \14902 , \14907 );
or \U$14595 ( \14910 , \14905 , \14908 , \14909 );
and \U$14596 ( \14911 , \14899 , \14910 );
and \U$14597 ( \14912 , \14866 , \14910 );
or \U$14598 ( \14913 , \14900 , \14911 , \14912 );
xor \U$14599 ( \14914 , \14466 , \14482 );
xor \U$14600 ( \14915 , \14914 , \14499 );
xor \U$14601 ( \14916 , \14518 , \14534 );
xor \U$14602 ( \14917 , \14916 , \14544 );
and \U$14603 ( \14918 , \14915 , \14917 );
xor \U$14604 ( \14919 , \14615 , \14617 );
xor \U$14605 ( \14920 , \14919 , \14620 );
and \U$14606 ( \14921 , \14917 , \14920 );
and \U$14607 ( \14922 , \14915 , \14920 );
or \U$14608 ( \14923 , \14918 , \14921 , \14922 );
xor \U$14609 ( \14924 , \14664 , \14666 );
xor \U$14610 ( \14925 , \14924 , \14669 );
and \U$14611 ( \14926 , \14923 , \14925 );
xor \U$14612 ( \14927 , \14640 , \14642 );
xor \U$14613 ( \14928 , \14927 , \14645 );
and \U$14614 ( \14929 , \14925 , \14928 );
and \U$14615 ( \14930 , \14923 , \14928 );
or \U$14616 ( \14931 , \14926 , \14929 , \14930 );
and \U$14617 ( \14932 , \14913 , \14931 );
xor \U$14618 ( \14933 , \14502 , \14547 );
xor \U$14619 ( \14934 , \14933 , \14600 );
xor \U$14620 ( \14935 , \14613 , \14623 );
xor \U$14621 ( \14936 , \14935 , \14634 );
and \U$14622 ( \14937 , \14934 , \14936 );
and \U$14623 ( \14938 , \14931 , \14937 );
and \U$14624 ( \14939 , \14913 , \14937 );
or \U$14625 ( \14940 , \14932 , \14938 , \14939 );
xor \U$14626 ( \14941 , \14603 , \14637 );
xor \U$14627 ( \14942 , \14941 , \14648 );
xor \U$14628 ( \14943 , \14653 , \14655 );
xor \U$14629 ( \14944 , \14943 , \14658 );
and \U$14630 ( \14945 , \14942 , \14944 );
xor \U$14631 ( \14946 , \14672 , \14674 );
xor \U$14632 ( \14947 , \14946 , \14676 );
and \U$14633 ( \14948 , \14944 , \14947 );
and \U$14634 ( \14949 , \14942 , \14947 );
or \U$14635 ( \14950 , \14945 , \14948 , \14949 );
and \U$14636 ( \14951 , \14940 , \14950 );
xor \U$14637 ( \14952 , \14215 , \14371 );
xor \U$14638 ( \14953 , \14952 , \14382 );
and \U$14639 ( \14954 , \14950 , \14953 );
and \U$14640 ( \14955 , \14940 , \14953 );
or \U$14641 ( \14956 , \14951 , \14954 , \14955 );
xor \U$14642 ( \14957 , \14651 , \14661 );
xor \U$14643 ( \14958 , \14957 , \14679 );
xor \U$14644 ( \14959 , \14684 , \14686 );
xor \U$14645 ( \14960 , \14959 , \14689 );
and \U$14646 ( \14961 , \14958 , \14960 );
and \U$14647 ( \14962 , \14956 , \14961 );
xor \U$14648 ( \14963 , \14385 , \14406 );
xor \U$14649 ( \14964 , \14963 , \14417 );
and \U$14650 ( \14965 , \14961 , \14964 );
and \U$14651 ( \14966 , \14956 , \14964 );
or \U$14652 ( \14967 , \14962 , \14965 , \14966 );
xor \U$14653 ( \14968 , \14698 , \14700 );
xor \U$14654 ( \14969 , \14968 , \14703 );
and \U$14655 ( \14970 , \14967 , \14969 );
and \U$14656 ( \14971 , \14712 , \14970 );
xor \U$14657 ( \14972 , \14712 , \14970 );
xor \U$14658 ( \14973 , \14967 , \14969 );
xor \U$14659 ( \14974 , \14956 , \14961 );
xor \U$14660 ( \14975 , \14974 , \14964 );
xor \U$14661 ( \14976 , \14682 , \14692 );
xor \U$14662 ( \14977 , \14976 , \14695 );
and \U$14663 ( \14978 , \14975 , \14977 );
and \U$14664 ( \14979 , \14973 , \14978 );
xor \U$14665 ( \14980 , \14973 , \14978 );
xor \U$14666 ( \14981 , \14975 , \14977 );
and \U$14667 ( \14982 , \2377 , \7238 );
and \U$14668 ( \14983 , \2233 , \7236 );
nor \U$14669 ( \14984 , \14982 , \14983 );
xnor \U$14670 ( \14985 , \14984 , \6978 );
and \U$14671 ( \14986 , \2666 , \6744 );
and \U$14672 ( \14987 , \2641 , \6742 );
nor \U$14673 ( \14988 , \14986 , \14987 );
xnor \U$14674 ( \14989 , \14988 , \6429 );
and \U$14675 ( \14990 , \14985 , \14989 );
and \U$14676 ( \14991 , \3007 , \6235 );
and \U$14677 ( \14992 , \2840 , \6233 );
nor \U$14678 ( \14993 , \14991 , \14992 );
xnor \U$14679 ( \14994 , \14993 , \5895 );
and \U$14680 ( \14995 , \14989 , \14994 );
and \U$14681 ( \14996 , \14985 , \14994 );
or \U$14682 ( \14997 , \14990 , \14995 , \14996 );
and \U$14683 ( \14998 , \988 , \10814 );
and \U$14684 ( \14999 , \925 , \10811 );
nor \U$14685 ( \15000 , \14998 , \14999 );
xnor \U$14686 ( \15001 , \15000 , \9759 );
and \U$14687 ( \15002 , \1274 , \10001 );
and \U$14688 ( \15003 , \1186 , \9999 );
nor \U$14689 ( \15004 , \15002 , \15003 );
xnor \U$14690 ( \15005 , \15004 , \9762 );
and \U$14691 ( \15006 , \15001 , \15005 );
and \U$14692 ( \15007 , \1384 , \9433 );
and \U$14693 ( \15008 , \1379 , \9431 );
nor \U$14694 ( \15009 , \15007 , \15008 );
xnor \U$14695 ( \15010 , \15009 , \9123 );
and \U$14696 ( \15011 , \15005 , \15010 );
and \U$14697 ( \15012 , \15001 , \15010 );
or \U$14698 ( \15013 , \15006 , \15011 , \15012 );
and \U$14699 ( \15014 , \14997 , \15013 );
and \U$14700 ( \15015 , \1615 , \8896 );
and \U$14701 ( \15016 , \1500 , \8894 );
nor \U$14702 ( \15017 , \15015 , \15016 );
xnor \U$14703 ( \15018 , \15017 , \8525 );
and \U$14704 ( \15019 , \1799 , \8334 );
and \U$14705 ( \15020 , \1791 , \8332 );
nor \U$14706 ( \15021 , \15019 , \15020 );
xnor \U$14707 ( \15022 , \15021 , \8016 );
and \U$14708 ( \15023 , \15018 , \15022 );
and \U$14709 ( \15024 , \2047 , \7767 );
and \U$14710 ( \15025 , \2042 , \7765 );
nor \U$14711 ( \15026 , \15024 , \15025 );
xnor \U$14712 ( \15027 , \15026 , \7518 );
and \U$14713 ( \15028 , \15022 , \15027 );
and \U$14714 ( \15029 , \15018 , \15027 );
or \U$14715 ( \15030 , \15023 , \15028 , \15029 );
and \U$14716 ( \15031 , \15013 , \15030 );
and \U$14717 ( \15032 , \14997 , \15030 );
or \U$14718 ( \15033 , \15014 , \15031 , \15032 );
and \U$14719 ( \15034 , \4469 , \4355 );
and \U$14720 ( \15035 , \4272 , \4353 );
nor \U$14721 ( \15036 , \15034 , \15035 );
xnor \U$14722 ( \15037 , \15036 , \4212 );
and \U$14723 ( \15038 , \4779 , \4032 );
and \U$14724 ( \15039 , \4771 , \4030 );
nor \U$14725 ( \15040 , \15038 , \15039 );
xnor \U$14726 ( \15041 , \15040 , \3786 );
and \U$14727 ( \15042 , \15037 , \15041 );
and \U$14728 ( \15043 , \5253 , \3637 );
and \U$14729 ( \15044 , \5248 , \3635 );
nor \U$14730 ( \15045 , \15043 , \15044 );
xnor \U$14731 ( \15046 , \15045 , \3450 );
and \U$14732 ( \15047 , \15041 , \15046 );
and \U$14733 ( \15048 , \15037 , \15046 );
or \U$14734 ( \15049 , \15042 , \15047 , \15048 );
and \U$14735 ( \15050 , \3264 , \5646 );
and \U$14736 ( \15051 , \3145 , \5644 );
nor \U$14737 ( \15052 , \15050 , \15051 );
xnor \U$14738 ( \15053 , \15052 , \5405 );
and \U$14739 ( \15054 , \3889 , \5180 );
and \U$14740 ( \15055 , \3681 , \5178 );
nor \U$14741 ( \15056 , \15054 , \15055 );
xnor \U$14742 ( \15057 , \15056 , \4992 );
and \U$14743 ( \15058 , \15053 , \15057 );
and \U$14744 ( \15059 , \4016 , \4806 );
and \U$14745 ( \15060 , \4011 , \4804 );
nor \U$14746 ( \15061 , \15059 , \15060 );
xnor \U$14747 ( \15062 , \15061 , \4574 );
and \U$14748 ( \15063 , \15057 , \15062 );
and \U$14749 ( \15064 , \15053 , \15062 );
or \U$14750 ( \15065 , \15058 , \15063 , \15064 );
and \U$14751 ( \15066 , \15049 , \15065 );
and \U$14752 ( \15067 , \5776 , \3324 );
and \U$14753 ( \15068 , \5517 , \3322 );
nor \U$14754 ( \15069 , \15067 , \15068 );
xnor \U$14755 ( \15070 , \15069 , \3119 );
and \U$14756 ( \15071 , \6157 , \2918 );
and \U$14757 ( \15072 , \6148 , \2916 );
nor \U$14758 ( \15073 , \15071 , \15072 );
xnor \U$14759 ( \15074 , \15073 , \2769 );
and \U$14760 ( \15075 , \15070 , \15074 );
and \U$14761 ( \15076 , \6702 , \2596 );
and \U$14762 ( \15077 , \6500 , \2594 );
nor \U$14763 ( \15078 , \15076 , \15077 );
xnor \U$14764 ( \15079 , \15078 , \2454 );
and \U$14765 ( \15080 , \15074 , \15079 );
and \U$14766 ( \15081 , \15070 , \15079 );
or \U$14767 ( \15082 , \15075 , \15080 , \15081 );
and \U$14768 ( \15083 , \15065 , \15082 );
and \U$14769 ( \15084 , \15049 , \15082 );
or \U$14770 ( \15085 , \15066 , \15083 , \15084 );
and \U$14771 ( \15086 , \15033 , \15085 );
and \U$14772 ( \15087 , \8981 , \1554 );
and \U$14773 ( \15088 , \8697 , \1552 );
nor \U$14774 ( \15089 , \15087 , \15088 );
xnor \U$14775 ( \15090 , \15089 , \1441 );
and \U$14776 ( \15091 , \9558 , \1360 );
and \U$14777 ( \15092 , \9550 , \1358 );
nor \U$14778 ( \15093 , \15091 , \15092 );
xnor \U$14779 ( \15094 , \15093 , \1224 );
and \U$14780 ( \15095 , \15090 , \15094 );
and \U$14781 ( \15096 , \10166 , \1160 );
and \U$14782 ( \15097 , \10161 , \1158 );
nor \U$14783 ( \15098 , \15096 , \15097 );
xnor \U$14784 ( \15099 , \15098 , \1082 );
and \U$14785 ( \15100 , \15094 , \15099 );
and \U$14786 ( \15101 , \15090 , \15099 );
or \U$14787 ( \15102 , \15095 , \15100 , \15101 );
and \U$14788 ( \15103 , \7177 , \2300 );
and \U$14789 ( \15104 , \7005 , \2298 );
nor \U$14790 ( \15105 , \15103 , \15104 );
xnor \U$14791 ( \15106 , \15105 , \2163 );
and \U$14792 ( \15107 , \8127 , \2094 );
and \U$14793 ( \15108 , \7703 , \2092 );
nor \U$14794 ( \15109 , \15107 , \15108 );
xnor \U$14795 ( \15110 , \15109 , \1942 );
and \U$14796 ( \15111 , \15106 , \15110 );
and \U$14797 ( \15112 , \8378 , \1826 );
and \U$14798 ( \15113 , \8373 , \1824 );
nor \U$14799 ( \15114 , \15112 , \15113 );
xnor \U$14800 ( \15115 , \15114 , \1670 );
and \U$14801 ( \15116 , \15110 , \15115 );
and \U$14802 ( \15117 , \15106 , \15115 );
or \U$14803 ( \15118 , \15111 , \15116 , \15117 );
and \U$14804 ( \15119 , \15102 , \15118 );
xor \U$14805 ( \15120 , \14833 , \14837 );
xor \U$14806 ( \15121 , \15120 , \14840 );
and \U$14807 ( \15122 , \15118 , \15121 );
and \U$14808 ( \15123 , \15102 , \15121 );
or \U$14809 ( \15124 , \15119 , \15122 , \15123 );
and \U$14810 ( \15125 , \15085 , \15124 );
and \U$14811 ( \15126 , \15033 , \15124 );
or \U$14812 ( \15127 , \15086 , \15125 , \15126 );
xor \U$14813 ( \15128 , \14817 , \14821 );
xor \U$14814 ( \15129 , \15128 , \14826 );
xor \U$14815 ( \15130 , \14749 , \14753 );
xor \U$14816 ( \15131 , \15130 , \14758 );
and \U$14817 ( \15132 , \15129 , \15131 );
xor \U$14818 ( \15133 , \14848 , \14852 );
xor \U$14819 ( \15134 , \15133 , \14857 );
and \U$14820 ( \15135 , \15131 , \15134 );
and \U$14821 ( \15136 , \15129 , \15134 );
or \U$14822 ( \15137 , \15132 , \15135 , \15136 );
xor \U$14823 ( \15138 , \14716 , \14720 );
xor \U$14824 ( \15139 , \15138 , \14725 );
xor \U$14825 ( \15140 , \14732 , \14736 );
xor \U$14826 ( \15141 , \15140 , \14741 );
and \U$14827 ( \15142 , \15139 , \15141 );
xor \U$14828 ( \15143 , \14768 , \14772 );
xor \U$14829 ( \15144 , \15143 , \14777 );
and \U$14830 ( \15145 , \15141 , \15144 );
and \U$14831 ( \15146 , \15139 , \15144 );
or \U$14832 ( \15147 , \15142 , \15145 , \15146 );
and \U$14833 ( \15148 , \15137 , \15147 );
xor \U$14834 ( \15149 , \14784 , \14788 );
xor \U$14835 ( \15150 , \15149 , \14793 );
xor \U$14836 ( \15151 , \14801 , \14805 );
xor \U$14837 ( \15152 , \15151 , \754 );
and \U$14838 ( \15153 , \15150 , \15152 );
and \U$14839 ( \15154 , \15147 , \15153 );
and \U$14840 ( \15155 , \15137 , \15153 );
or \U$14841 ( \15156 , \15148 , \15154 , \15155 );
and \U$14842 ( \15157 , \15127 , \15156 );
xor \U$14843 ( \15158 , \14868 , \14870 );
xor \U$14844 ( \15159 , \15158 , \14873 );
xor \U$14845 ( \15160 , \14878 , \14880 );
xor \U$14846 ( \15161 , \15160 , \14883 );
and \U$14847 ( \15162 , \15159 , \15161 );
xor \U$14848 ( \15163 , \14889 , \14891 );
xor \U$14849 ( \15164 , \15163 , \14893 );
and \U$14850 ( \15165 , \15161 , \15164 );
and \U$14851 ( \15166 , \15159 , \15164 );
or \U$14852 ( \15167 , \15162 , \15165 , \15166 );
and \U$14853 ( \15168 , \15156 , \15167 );
and \U$14854 ( \15169 , \15127 , \15167 );
or \U$14855 ( \15170 , \15157 , \15168 , \15169 );
xor \U$14856 ( \15171 , \14728 , \14744 );
xor \U$14857 ( \15172 , \15171 , \14761 );
xor \U$14858 ( \15173 , \14780 , \14796 );
xor \U$14859 ( \15174 , \15173 , \14809 );
and \U$14860 ( \15175 , \15172 , \15174 );
xor \U$14861 ( \15176 , \14829 , \14843 );
xor \U$14862 ( \15177 , \15176 , \14860 );
and \U$14863 ( \15178 , \15174 , \15177 );
and \U$14864 ( \15179 , \15172 , \15177 );
or \U$14865 ( \15180 , \15175 , \15178 , \15179 );
xor \U$14866 ( \15181 , \14564 , \14580 );
xor \U$14867 ( \15182 , \15181 , \14597 );
and \U$14868 ( \15183 , \15180 , \15182 );
xor \U$14869 ( \15184 , \14915 , \14917 );
xor \U$14870 ( \15185 , \15184 , \14920 );
and \U$14871 ( \15186 , \15182 , \15185 );
and \U$14872 ( \15187 , \15180 , \15185 );
or \U$14873 ( \15188 , \15183 , \15186 , \15187 );
and \U$14874 ( \15189 , \15170 , \15188 );
xor \U$14875 ( \15190 , \14764 , \14812 );
xor \U$14876 ( \15191 , \15190 , \14863 );
xor \U$14877 ( \15192 , \14876 , \14886 );
xor \U$14878 ( \15193 , \15192 , \14896 );
and \U$14879 ( \15194 , \15191 , \15193 );
xor \U$14880 ( \15195 , \14902 , \14904 );
xor \U$14881 ( \15196 , \15195 , \14907 );
and \U$14882 ( \15197 , \15193 , \15196 );
and \U$14883 ( \15198 , \15191 , \15196 );
or \U$14884 ( \15199 , \15194 , \15197 , \15198 );
and \U$14885 ( \15200 , \15188 , \15199 );
and \U$14886 ( \15201 , \15170 , \15199 );
or \U$14887 ( \15202 , \15189 , \15200 , \15201 );
xor \U$14888 ( \15203 , \14866 , \14899 );
xor \U$14889 ( \15204 , \15203 , \14910 );
xor \U$14890 ( \15205 , \14923 , \14925 );
xor \U$14891 ( \15206 , \15205 , \14928 );
and \U$14892 ( \15207 , \15204 , \15206 );
xor \U$14893 ( \15208 , \14934 , \14936 );
and \U$14894 ( \15209 , \15206 , \15208 );
and \U$14895 ( \15210 , \15204 , \15208 );
or \U$14896 ( \15211 , \15207 , \15209 , \15210 );
and \U$14897 ( \15212 , \15202 , \15211 );
xor \U$14898 ( \15213 , \14942 , \14944 );
xor \U$14899 ( \15214 , \15213 , \14947 );
and \U$14900 ( \15215 , \15211 , \15214 );
and \U$14901 ( \15216 , \15202 , \15214 );
or \U$14902 ( \15217 , \15212 , \15215 , \15216 );
xor \U$14903 ( \15218 , \14940 , \14950 );
xor \U$14904 ( \15219 , \15218 , \14953 );
and \U$14905 ( \15220 , \15217 , \15219 );
xor \U$14906 ( \15221 , \14958 , \14960 );
and \U$14907 ( \15222 , \15219 , \15221 );
and \U$14908 ( \15223 , \15217 , \15221 );
or \U$14909 ( \15224 , \15220 , \15222 , \15223 );
and \U$14910 ( \15225 , \14981 , \15224 );
xor \U$14911 ( \15226 , \14981 , \15224 );
xor \U$14912 ( \15227 , \15217 , \15219 );
xor \U$14913 ( \15228 , \15227 , \15221 );
and \U$14914 ( \15229 , \2233 , \7767 );
and \U$14915 ( \15230 , \2047 , \7765 );
nor \U$14916 ( \15231 , \15229 , \15230 );
xnor \U$14917 ( \15232 , \15231 , \7518 );
and \U$14918 ( \15233 , \2641 , \7238 );
and \U$14919 ( \15234 , \2377 , \7236 );
nor \U$14920 ( \15235 , \15233 , \15234 );
xnor \U$14921 ( \15236 , \15235 , \6978 );
and \U$14922 ( \15237 , \15232 , \15236 );
and \U$14923 ( \15238 , \2840 , \6744 );
and \U$14924 ( \15239 , \2666 , \6742 );
nor \U$14925 ( \15240 , \15238 , \15239 );
xnor \U$14926 ( \15241 , \15240 , \6429 );
and \U$14927 ( \15242 , \15236 , \15241 );
and \U$14928 ( \15243 , \15232 , \15241 );
or \U$14929 ( \15244 , \15237 , \15242 , \15243 );
and \U$14930 ( \15245 , \1500 , \9433 );
and \U$14931 ( \15246 , \1384 , \9431 );
nor \U$14932 ( \15247 , \15245 , \15246 );
xnor \U$14933 ( \15248 , \15247 , \9123 );
and \U$14934 ( \15249 , \1791 , \8896 );
and \U$14935 ( \15250 , \1615 , \8894 );
nor \U$14936 ( \15251 , \15249 , \15250 );
xnor \U$14937 ( \15252 , \15251 , \8525 );
and \U$14938 ( \15253 , \15248 , \15252 );
and \U$14939 ( \15254 , \2042 , \8334 );
and \U$14940 ( \15255 , \1799 , \8332 );
nor \U$14941 ( \15256 , \15254 , \15255 );
xnor \U$14942 ( \15257 , \15256 , \8016 );
and \U$14943 ( \15258 , \15252 , \15257 );
and \U$14944 ( \15259 , \15248 , \15257 );
or \U$14945 ( \15260 , \15253 , \15258 , \15259 );
and \U$14946 ( \15261 , \15244 , \15260 );
and \U$14947 ( \15262 , \1186 , \10814 );
and \U$14948 ( \15263 , \988 , \10811 );
nor \U$14949 ( \15264 , \15262 , \15263 );
xnor \U$14950 ( \15265 , \15264 , \9759 );
and \U$14951 ( \15266 , \1379 , \10001 );
and \U$14952 ( \15267 , \1274 , \9999 );
nor \U$14953 ( \15268 , \15266 , \15267 );
xnor \U$14954 ( \15269 , \15268 , \9762 );
and \U$14955 ( \15270 , \15265 , \15269 );
and \U$14956 ( \15271 , \15269 , \902 );
and \U$14957 ( \15272 , \15265 , \902 );
or \U$14958 ( \15273 , \15270 , \15271 , \15272 );
and \U$14959 ( \15274 , \15260 , \15273 );
and \U$14960 ( \15275 , \15244 , \15273 );
or \U$14961 ( \15276 , \15261 , \15274 , \15275 );
and \U$14962 ( \15277 , \7005 , \2596 );
and \U$14963 ( \15278 , \6702 , \2594 );
nor \U$14964 ( \15279 , \15277 , \15278 );
xnor \U$14965 ( \15280 , \15279 , \2454 );
and \U$14966 ( \15281 , \7703 , \2300 );
and \U$14967 ( \15282 , \7177 , \2298 );
nor \U$14968 ( \15283 , \15281 , \15282 );
xnor \U$14969 ( \15284 , \15283 , \2163 );
and \U$14970 ( \15285 , \15280 , \15284 );
and \U$14971 ( \15286 , \8373 , \2094 );
and \U$14972 ( \15287 , \8127 , \2092 );
nor \U$14973 ( \15288 , \15286 , \15287 );
xnor \U$14974 ( \15289 , \15288 , \1942 );
and \U$14975 ( \15290 , \15284 , \15289 );
and \U$14976 ( \15291 , \15280 , \15289 );
or \U$14977 ( \15292 , \15285 , \15290 , \15291 );
and \U$14978 ( \15293 , \8697 , \1826 );
and \U$14979 ( \15294 , \8378 , \1824 );
nor \U$14980 ( \15295 , \15293 , \15294 );
xnor \U$14981 ( \15296 , \15295 , \1670 );
and \U$14982 ( \15297 , \9550 , \1554 );
and \U$14983 ( \15298 , \8981 , \1552 );
nor \U$14984 ( \15299 , \15297 , \15298 );
xnor \U$14985 ( \15300 , \15299 , \1441 );
and \U$14986 ( \15301 , \15296 , \15300 );
and \U$14987 ( \15302 , \10161 , \1360 );
and \U$14988 ( \15303 , \9558 , \1358 );
nor \U$14989 ( \15304 , \15302 , \15303 );
xnor \U$14990 ( \15305 , \15304 , \1224 );
and \U$14991 ( \15306 , \15300 , \15305 );
and \U$14992 ( \15307 , \15296 , \15305 );
or \U$14993 ( \15308 , \15301 , \15306 , \15307 );
and \U$14994 ( \15309 , \15292 , \15308 );
and \U$14995 ( \15310 , \10967 , \996 );
and \U$14996 ( \15311 , \10347 , \994 );
nor \U$14997 ( \15312 , \15310 , \15311 );
xnor \U$14998 ( \15313 , \15312 , \902 );
and \U$14999 ( \15314 , \15308 , \15313 );
and \U$15000 ( \15315 , \15292 , \15313 );
or \U$15001 ( \15316 , \15309 , \15314 , \15315 );
and \U$15002 ( \15317 , \15276 , \15316 );
and \U$15003 ( \15318 , \4272 , \4806 );
and \U$15004 ( \15319 , \4016 , \4804 );
nor \U$15005 ( \15320 , \15318 , \15319 );
xnor \U$15006 ( \15321 , \15320 , \4574 );
and \U$15007 ( \15322 , \4771 , \4355 );
and \U$15008 ( \15323 , \4469 , \4353 );
nor \U$15009 ( \15324 , \15322 , \15323 );
xnor \U$15010 ( \15325 , \15324 , \4212 );
and \U$15011 ( \15326 , \15321 , \15325 );
and \U$15012 ( \15327 , \5248 , \4032 );
and \U$15013 ( \15328 , \4779 , \4030 );
nor \U$15014 ( \15329 , \15327 , \15328 );
xnor \U$15015 ( \15330 , \15329 , \3786 );
and \U$15016 ( \15331 , \15325 , \15330 );
and \U$15017 ( \15332 , \15321 , \15330 );
or \U$15018 ( \15333 , \15326 , \15331 , \15332 );
and \U$15019 ( \15334 , \3145 , \6235 );
and \U$15020 ( \15335 , \3007 , \6233 );
nor \U$15021 ( \15336 , \15334 , \15335 );
xnor \U$15022 ( \15337 , \15336 , \5895 );
and \U$15023 ( \15338 , \3681 , \5646 );
and \U$15024 ( \15339 , \3264 , \5644 );
nor \U$15025 ( \15340 , \15338 , \15339 );
xnor \U$15026 ( \15341 , \15340 , \5405 );
and \U$15027 ( \15342 , \15337 , \15341 );
and \U$15028 ( \15343 , \4011 , \5180 );
and \U$15029 ( \15344 , \3889 , \5178 );
nor \U$15030 ( \15345 , \15343 , \15344 );
xnor \U$15031 ( \15346 , \15345 , \4992 );
and \U$15032 ( \15347 , \15341 , \15346 );
and \U$15033 ( \15348 , \15337 , \15346 );
or \U$15034 ( \15349 , \15342 , \15347 , \15348 );
and \U$15035 ( \15350 , \15333 , \15349 );
and \U$15036 ( \15351 , \5517 , \3637 );
and \U$15037 ( \15352 , \5253 , \3635 );
nor \U$15038 ( \15353 , \15351 , \15352 );
xnor \U$15039 ( \15354 , \15353 , \3450 );
and \U$15040 ( \15355 , \6148 , \3324 );
and \U$15041 ( \15356 , \5776 , \3322 );
nor \U$15042 ( \15357 , \15355 , \15356 );
xnor \U$15043 ( \15358 , \15357 , \3119 );
and \U$15044 ( \15359 , \15354 , \15358 );
and \U$15045 ( \15360 , \6500 , \2918 );
and \U$15046 ( \15361 , \6157 , \2916 );
nor \U$15047 ( \15362 , \15360 , \15361 );
xnor \U$15048 ( \15363 , \15362 , \2769 );
and \U$15049 ( \15364 , \15358 , \15363 );
and \U$15050 ( \15365 , \15354 , \15363 );
or \U$15051 ( \15366 , \15359 , \15364 , \15365 );
and \U$15052 ( \15367 , \15349 , \15366 );
and \U$15053 ( \15368 , \15333 , \15366 );
or \U$15054 ( \15369 , \15350 , \15367 , \15368 );
and \U$15055 ( \15370 , \15316 , \15369 );
and \U$15056 ( \15371 , \15276 , \15369 );
or \U$15057 ( \15372 , \15317 , \15370 , \15371 );
xor \U$15058 ( \15373 , \15090 , \15094 );
xor \U$15059 ( \15374 , \15373 , \15099 );
xor \U$15060 ( \15375 , \15070 , \15074 );
xor \U$15061 ( \15376 , \15375 , \15079 );
and \U$15062 ( \15377 , \15374 , \15376 );
xor \U$15063 ( \15378 , \15106 , \15110 );
xor \U$15064 ( \15379 , \15378 , \15115 );
and \U$15065 ( \15380 , \15376 , \15379 );
and \U$15066 ( \15381 , \15374 , \15379 );
or \U$15067 ( \15382 , \15377 , \15380 , \15381 );
xor \U$15068 ( \15383 , \15037 , \15041 );
xor \U$15069 ( \15384 , \15383 , \15046 );
xor \U$15070 ( \15385 , \15053 , \15057 );
xor \U$15071 ( \15386 , \15385 , \15062 );
and \U$15072 ( \15387 , \15384 , \15386 );
xor \U$15073 ( \15388 , \14985 , \14989 );
xor \U$15074 ( \15389 , \15388 , \14994 );
and \U$15075 ( \15390 , \15386 , \15389 );
and \U$15076 ( \15391 , \15384 , \15389 );
or \U$15077 ( \15392 , \15387 , \15390 , \15391 );
and \U$15078 ( \15393 , \15382 , \15392 );
xor \U$15079 ( \15394 , \15001 , \15005 );
xor \U$15080 ( \15395 , \15394 , \15010 );
xor \U$15081 ( \15396 , \15018 , \15022 );
xor \U$15082 ( \15397 , \15396 , \15027 );
and \U$15083 ( \15398 , \15395 , \15397 );
and \U$15084 ( \15399 , \15392 , \15398 );
and \U$15085 ( \15400 , \15382 , \15398 );
or \U$15086 ( \15401 , \15393 , \15399 , \15400 );
and \U$15087 ( \15402 , \15372 , \15401 );
xor \U$15088 ( \15403 , \15129 , \15131 );
xor \U$15089 ( \15404 , \15403 , \15134 );
xor \U$15090 ( \15405 , \15139 , \15141 );
xor \U$15091 ( \15406 , \15405 , \15144 );
and \U$15092 ( \15407 , \15404 , \15406 );
xor \U$15093 ( \15408 , \15150 , \15152 );
and \U$15094 ( \15409 , \15406 , \15408 );
and \U$15095 ( \15410 , \15404 , \15408 );
or \U$15096 ( \15411 , \15407 , \15409 , \15410 );
and \U$15097 ( \15412 , \15401 , \15411 );
and \U$15098 ( \15413 , \15372 , \15411 );
or \U$15099 ( \15414 , \15402 , \15412 , \15413 );
xor \U$15100 ( \15415 , \14997 , \15013 );
xor \U$15101 ( \15416 , \15415 , \15030 );
xor \U$15102 ( \15417 , \15049 , \15065 );
xor \U$15103 ( \15418 , \15417 , \15082 );
and \U$15104 ( \15419 , \15416 , \15418 );
xor \U$15105 ( \15420 , \15102 , \15118 );
xor \U$15106 ( \15421 , \15420 , \15121 );
and \U$15107 ( \15422 , \15418 , \15421 );
and \U$15108 ( \15423 , \15416 , \15421 );
or \U$15109 ( \15424 , \15419 , \15422 , \15423 );
xor \U$15110 ( \15425 , \15172 , \15174 );
xor \U$15111 ( \15426 , \15425 , \15177 );
and \U$15112 ( \15427 , \15424 , \15426 );
xor \U$15113 ( \15428 , \15159 , \15161 );
xor \U$15114 ( \15429 , \15428 , \15164 );
and \U$15115 ( \15430 , \15426 , \15429 );
and \U$15116 ( \15431 , \15424 , \15429 );
or \U$15117 ( \15432 , \15427 , \15430 , \15431 );
and \U$15118 ( \15433 , \15414 , \15432 );
xor \U$15119 ( \15434 , \15191 , \15193 );
xor \U$15120 ( \15435 , \15434 , \15196 );
and \U$15121 ( \15436 , \15432 , \15435 );
and \U$15122 ( \15437 , \15414 , \15435 );
or \U$15123 ( \15438 , \15433 , \15436 , \15437 );
xor \U$15124 ( \15439 , \15170 , \15188 );
xor \U$15125 ( \15440 , \15439 , \15199 );
and \U$15126 ( \15441 , \15438 , \15440 );
xor \U$15127 ( \15442 , \15204 , \15206 );
xor \U$15128 ( \15443 , \15442 , \15208 );
and \U$15129 ( \15444 , \15440 , \15443 );
and \U$15130 ( \15445 , \15438 , \15443 );
or \U$15131 ( \15446 , \15441 , \15444 , \15445 );
xor \U$15132 ( \15447 , \14913 , \14931 );
xor \U$15133 ( \15448 , \15447 , \14937 );
and \U$15134 ( \15449 , \15446 , \15448 );
xor \U$15135 ( \15450 , \15202 , \15211 );
xor \U$15136 ( \15451 , \15450 , \15214 );
and \U$15137 ( \15452 , \15448 , \15451 );
and \U$15138 ( \15453 , \15446 , \15451 );
or \U$15139 ( \15454 , \15449 , \15452 , \15453 );
and \U$15140 ( \15455 , \15228 , \15454 );
xor \U$15141 ( \15456 , \15228 , \15454 );
xor \U$15142 ( \15457 , \15446 , \15448 );
xor \U$15143 ( \15458 , \15457 , \15451 );
xor \U$15144 ( \15459 , \15232 , \15236 );
xor \U$15145 ( \15460 , \15459 , \15241 );
xor \U$15146 ( \15461 , \15248 , \15252 );
xor \U$15147 ( \15462 , \15461 , \15257 );
and \U$15148 ( \15463 , \15460 , \15462 );
xor \U$15149 ( \15464 , \15265 , \15269 );
xor \U$15150 ( \15465 , \15464 , \902 );
and \U$15151 ( \15466 , \15462 , \15465 );
and \U$15152 ( \15467 , \15460 , \15465 );
or \U$15153 ( \15468 , \15463 , \15466 , \15467 );
nand \U$15154 ( \15469 , \10967 , \994 );
xnor \U$15155 ( \15470 , \15469 , \902 );
xor \U$15156 ( \15471 , \15280 , \15284 );
xor \U$15157 ( \15472 , \15471 , \15289 );
and \U$15158 ( \15473 , \15470 , \15472 );
xor \U$15159 ( \15474 , \15296 , \15300 );
xor \U$15160 ( \15475 , \15474 , \15305 );
and \U$15161 ( \15476 , \15472 , \15475 );
and \U$15162 ( \15477 , \15470 , \15475 );
or \U$15163 ( \15478 , \15473 , \15476 , \15477 );
and \U$15164 ( \15479 , \15468 , \15478 );
xor \U$15165 ( \15480 , \15321 , \15325 );
xor \U$15166 ( \15481 , \15480 , \15330 );
xor \U$15167 ( \15482 , \15337 , \15341 );
xor \U$15168 ( \15483 , \15482 , \15346 );
and \U$15169 ( \15484 , \15481 , \15483 );
xor \U$15170 ( \15485 , \15354 , \15358 );
xor \U$15171 ( \15486 , \15485 , \15363 );
and \U$15172 ( \15487 , \15483 , \15486 );
and \U$15173 ( \15488 , \15481 , \15486 );
or \U$15174 ( \15489 , \15484 , \15487 , \15488 );
and \U$15175 ( \15490 , \15478 , \15489 );
and \U$15176 ( \15491 , \15468 , \15489 );
or \U$15177 ( \15492 , \15479 , \15490 , \15491 );
and \U$15178 ( \15493 , \8127 , \2300 );
and \U$15179 ( \15494 , \7703 , \2298 );
nor \U$15180 ( \15495 , \15493 , \15494 );
xnor \U$15181 ( \15496 , \15495 , \2163 );
and \U$15182 ( \15497 , \8378 , \2094 );
and \U$15183 ( \15498 , \8373 , \2092 );
nor \U$15184 ( \15499 , \15497 , \15498 );
xnor \U$15185 ( \15500 , \15499 , \1942 );
and \U$15186 ( \15501 , \15496 , \15500 );
and \U$15187 ( \15502 , \8981 , \1826 );
and \U$15188 ( \15503 , \8697 , \1824 );
nor \U$15189 ( \15504 , \15502 , \15503 );
xnor \U$15190 ( \15505 , \15504 , \1670 );
and \U$15191 ( \15506 , \15500 , \15505 );
and \U$15192 ( \15507 , \15496 , \15505 );
or \U$15193 ( \15508 , \15501 , \15506 , \15507 );
and \U$15194 ( \15509 , \9558 , \1554 );
and \U$15195 ( \15510 , \9550 , \1552 );
nor \U$15196 ( \15511 , \15509 , \15510 );
xnor \U$15197 ( \15512 , \15511 , \1441 );
and \U$15198 ( \15513 , \10166 , \1360 );
and \U$15199 ( \15514 , \10161 , \1358 );
nor \U$15200 ( \15515 , \15513 , \15514 );
xnor \U$15201 ( \15516 , \15515 , \1224 );
and \U$15202 ( \15517 , \15512 , \15516 );
and \U$15203 ( \15518 , \10967 , \1160 );
and \U$15204 ( \15519 , \10347 , \1158 );
nor \U$15205 ( \15520 , \15518 , \15519 );
xnor \U$15206 ( \15521 , \15520 , \1082 );
and \U$15207 ( \15522 , \15516 , \15521 );
and \U$15208 ( \15523 , \15512 , \15521 );
or \U$15209 ( \15524 , \15517 , \15522 , \15523 );
and \U$15210 ( \15525 , \15508 , \15524 );
and \U$15211 ( \15526 , \10347 , \1160 );
and \U$15212 ( \15527 , \10166 , \1158 );
nor \U$15213 ( \15528 , \15526 , \15527 );
xnor \U$15214 ( \15529 , \15528 , \1082 );
and \U$15215 ( \15530 , \15524 , \15529 );
and \U$15216 ( \15531 , \15508 , \15529 );
or \U$15217 ( \15532 , \15525 , \15530 , \15531 );
and \U$15218 ( \15533 , \1274 , \10814 );
and \U$15219 ( \15534 , \1186 , \10811 );
nor \U$15220 ( \15535 , \15533 , \15534 );
xnor \U$15221 ( \15536 , \15535 , \9759 );
and \U$15222 ( \15537 , \1384 , \10001 );
and \U$15223 ( \15538 , \1379 , \9999 );
nor \U$15224 ( \15539 , \15537 , \15538 );
xnor \U$15225 ( \15540 , \15539 , \9762 );
and \U$15226 ( \15541 , \15536 , \15540 );
and \U$15227 ( \15542 , \1615 , \9433 );
and \U$15228 ( \15543 , \1500 , \9431 );
nor \U$15229 ( \15544 , \15542 , \15543 );
xnor \U$15230 ( \15545 , \15544 , \9123 );
and \U$15231 ( \15546 , \15540 , \15545 );
and \U$15232 ( \15547 , \15536 , \15545 );
or \U$15233 ( \15548 , \15541 , \15546 , \15547 );
and \U$15234 ( \15549 , \1799 , \8896 );
and \U$15235 ( \15550 , \1791 , \8894 );
nor \U$15236 ( \15551 , \15549 , \15550 );
xnor \U$15237 ( \15552 , \15551 , \8525 );
and \U$15238 ( \15553 , \2047 , \8334 );
and \U$15239 ( \15554 , \2042 , \8332 );
nor \U$15240 ( \15555 , \15553 , \15554 );
xnor \U$15241 ( \15556 , \15555 , \8016 );
and \U$15242 ( \15557 , \15552 , \15556 );
and \U$15243 ( \15558 , \2377 , \7767 );
and \U$15244 ( \15559 , \2233 , \7765 );
nor \U$15245 ( \15560 , \15558 , \15559 );
xnor \U$15246 ( \15561 , \15560 , \7518 );
and \U$15247 ( \15562 , \15556 , \15561 );
and \U$15248 ( \15563 , \15552 , \15561 );
or \U$15249 ( \15564 , \15557 , \15562 , \15563 );
and \U$15250 ( \15565 , \15548 , \15564 );
and \U$15251 ( \15566 , \2666 , \7238 );
and \U$15252 ( \15567 , \2641 , \7236 );
nor \U$15253 ( \15568 , \15566 , \15567 );
xnor \U$15254 ( \15569 , \15568 , \6978 );
and \U$15255 ( \15570 , \3007 , \6744 );
and \U$15256 ( \15571 , \2840 , \6742 );
nor \U$15257 ( \15572 , \15570 , \15571 );
xnor \U$15258 ( \15573 , \15572 , \6429 );
and \U$15259 ( \15574 , \15569 , \15573 );
and \U$15260 ( \15575 , \3264 , \6235 );
and \U$15261 ( \15576 , \3145 , \6233 );
nor \U$15262 ( \15577 , \15575 , \15576 );
xnor \U$15263 ( \15578 , \15577 , \5895 );
and \U$15264 ( \15579 , \15573 , \15578 );
and \U$15265 ( \15580 , \15569 , \15578 );
or \U$15266 ( \15581 , \15574 , \15579 , \15580 );
and \U$15267 ( \15582 , \15564 , \15581 );
and \U$15268 ( \15583 , \15548 , \15581 );
or \U$15269 ( \15584 , \15565 , \15582 , \15583 );
and \U$15270 ( \15585 , \15532 , \15584 );
and \U$15271 ( \15586 , \4779 , \4355 );
and \U$15272 ( \15587 , \4771 , \4353 );
nor \U$15273 ( \15588 , \15586 , \15587 );
xnor \U$15274 ( \15589 , \15588 , \4212 );
and \U$15275 ( \15590 , \5253 , \4032 );
and \U$15276 ( \15591 , \5248 , \4030 );
nor \U$15277 ( \15592 , \15590 , \15591 );
xnor \U$15278 ( \15593 , \15592 , \3786 );
and \U$15279 ( \15594 , \15589 , \15593 );
and \U$15280 ( \15595 , \5776 , \3637 );
and \U$15281 ( \15596 , \5517 , \3635 );
nor \U$15282 ( \15597 , \15595 , \15596 );
xnor \U$15283 ( \15598 , \15597 , \3450 );
and \U$15284 ( \15599 , \15593 , \15598 );
and \U$15285 ( \15600 , \15589 , \15598 );
or \U$15286 ( \15601 , \15594 , \15599 , \15600 );
and \U$15287 ( \15602 , \6157 , \3324 );
and \U$15288 ( \15603 , \6148 , \3322 );
nor \U$15289 ( \15604 , \15602 , \15603 );
xnor \U$15290 ( \15605 , \15604 , \3119 );
and \U$15291 ( \15606 , \6702 , \2918 );
and \U$15292 ( \15607 , \6500 , \2916 );
nor \U$15293 ( \15608 , \15606 , \15607 );
xnor \U$15294 ( \15609 , \15608 , \2769 );
and \U$15295 ( \15610 , \15605 , \15609 );
and \U$15296 ( \15611 , \7177 , \2596 );
and \U$15297 ( \15612 , \7005 , \2594 );
nor \U$15298 ( \15613 , \15611 , \15612 );
xnor \U$15299 ( \15614 , \15613 , \2454 );
and \U$15300 ( \15615 , \15609 , \15614 );
and \U$15301 ( \15616 , \15605 , \15614 );
or \U$15302 ( \15617 , \15610 , \15615 , \15616 );
and \U$15303 ( \15618 , \15601 , \15617 );
and \U$15304 ( \15619 , \3889 , \5646 );
and \U$15305 ( \15620 , \3681 , \5644 );
nor \U$15306 ( \15621 , \15619 , \15620 );
xnor \U$15307 ( \15622 , \15621 , \5405 );
and \U$15308 ( \15623 , \4016 , \5180 );
and \U$15309 ( \15624 , \4011 , \5178 );
nor \U$15310 ( \15625 , \15623 , \15624 );
xnor \U$15311 ( \15626 , \15625 , \4992 );
and \U$15312 ( \15627 , \15622 , \15626 );
and \U$15313 ( \15628 , \4469 , \4806 );
and \U$15314 ( \15629 , \4272 , \4804 );
nor \U$15315 ( \15630 , \15628 , \15629 );
xnor \U$15316 ( \15631 , \15630 , \4574 );
and \U$15317 ( \15632 , \15626 , \15631 );
and \U$15318 ( \15633 , \15622 , \15631 );
or \U$15319 ( \15634 , \15627 , \15632 , \15633 );
and \U$15320 ( \15635 , \15617 , \15634 );
and \U$15321 ( \15636 , \15601 , \15634 );
or \U$15322 ( \15637 , \15618 , \15635 , \15636 );
and \U$15323 ( \15638 , \15584 , \15637 );
and \U$15324 ( \15639 , \15532 , \15637 );
or \U$15325 ( \15640 , \15585 , \15638 , \15639 );
and \U$15326 ( \15641 , \15492 , \15640 );
xor \U$15327 ( \15642 , \15374 , \15376 );
xor \U$15328 ( \15643 , \15642 , \15379 );
xor \U$15329 ( \15644 , \15384 , \15386 );
xor \U$15330 ( \15645 , \15644 , \15389 );
and \U$15331 ( \15646 , \15643 , \15645 );
xor \U$15332 ( \15647 , \15395 , \15397 );
and \U$15333 ( \15648 , \15645 , \15647 );
and \U$15334 ( \15649 , \15643 , \15647 );
or \U$15335 ( \15650 , \15646 , \15648 , \15649 );
and \U$15336 ( \15651 , \15640 , \15650 );
and \U$15337 ( \15652 , \15492 , \15650 );
or \U$15338 ( \15653 , \15641 , \15651 , \15652 );
xor \U$15339 ( \15654 , \15244 , \15260 );
xor \U$15340 ( \15655 , \15654 , \15273 );
xor \U$15341 ( \15656 , \15292 , \15308 );
xor \U$15342 ( \15657 , \15656 , \15313 );
and \U$15343 ( \15658 , \15655 , \15657 );
xor \U$15344 ( \15659 , \15333 , \15349 );
xor \U$15345 ( \15660 , \15659 , \15366 );
and \U$15346 ( \15661 , \15657 , \15660 );
and \U$15347 ( \15662 , \15655 , \15660 );
or \U$15348 ( \15663 , \15658 , \15661 , \15662 );
xor \U$15349 ( \15664 , \15416 , \15418 );
xor \U$15350 ( \15665 , \15664 , \15421 );
and \U$15351 ( \15666 , \15663 , \15665 );
xor \U$15352 ( \15667 , \15404 , \15406 );
xor \U$15353 ( \15668 , \15667 , \15408 );
and \U$15354 ( \15669 , \15665 , \15668 );
and \U$15355 ( \15670 , \15663 , \15668 );
or \U$15356 ( \15671 , \15666 , \15669 , \15670 );
and \U$15357 ( \15672 , \15653 , \15671 );
xor \U$15358 ( \15673 , \15137 , \15147 );
xor \U$15359 ( \15674 , \15673 , \15153 );
and \U$15360 ( \15675 , \15671 , \15674 );
and \U$15361 ( \15676 , \15653 , \15674 );
or \U$15362 ( \15677 , \15672 , \15675 , \15676 );
xor \U$15363 ( \15678 , \15033 , \15085 );
xor \U$15364 ( \15679 , \15678 , \15124 );
xor \U$15365 ( \15680 , \15372 , \15401 );
xor \U$15366 ( \15681 , \15680 , \15411 );
and \U$15367 ( \15682 , \15679 , \15681 );
xor \U$15368 ( \15683 , \15424 , \15426 );
xor \U$15369 ( \15684 , \15683 , \15429 );
and \U$15370 ( \15685 , \15681 , \15684 );
and \U$15371 ( \15686 , \15679 , \15684 );
or \U$15372 ( \15687 , \15682 , \15685 , \15686 );
and \U$15373 ( \15688 , \15677 , \15687 );
xor \U$15374 ( \15689 , \15180 , \15182 );
xor \U$15375 ( \15690 , \15689 , \15185 );
and \U$15376 ( \15691 , \15687 , \15690 );
and \U$15377 ( \15692 , \15677 , \15690 );
or \U$15378 ( \15693 , \15688 , \15691 , \15692 );
xor \U$15379 ( \15694 , \15127 , \15156 );
xor \U$15380 ( \15695 , \15694 , \15167 );
xor \U$15381 ( \15696 , \15414 , \15432 );
xor \U$15382 ( \15697 , \15696 , \15435 );
and \U$15383 ( \15698 , \15695 , \15697 );
and \U$15384 ( \15699 , \15693 , \15698 );
xor \U$15385 ( \15700 , \15438 , \15440 );
xor \U$15386 ( \15701 , \15700 , \15443 );
and \U$15387 ( \15702 , \15698 , \15701 );
and \U$15388 ( \15703 , \15693 , \15701 );
or \U$15389 ( \15704 , \15699 , \15702 , \15703 );
and \U$15390 ( \15705 , \15458 , \15704 );
xor \U$15391 ( \15706 , \15458 , \15704 );
xor \U$15392 ( \15707 , \15693 , \15698 );
xor \U$15393 ( \15708 , \15707 , \15701 );
and \U$15394 ( \15709 , \6148 , \3637 );
and \U$15395 ( \15710 , \5776 , \3635 );
nor \U$15396 ( \15711 , \15709 , \15710 );
xnor \U$15397 ( \15712 , \15711 , \3450 );
and \U$15398 ( \15713 , \6500 , \3324 );
and \U$15399 ( \15714 , \6157 , \3322 );
nor \U$15400 ( \15715 , \15713 , \15714 );
xnor \U$15401 ( \15716 , \15715 , \3119 );
and \U$15402 ( \15717 , \15712 , \15716 );
and \U$15403 ( \15718 , \7005 , \2918 );
and \U$15404 ( \15719 , \6702 , \2916 );
nor \U$15405 ( \15720 , \15718 , \15719 );
xnor \U$15406 ( \15721 , \15720 , \2769 );
and \U$15407 ( \15722 , \15716 , \15721 );
and \U$15408 ( \15723 , \15712 , \15721 );
or \U$15409 ( \15724 , \15717 , \15722 , \15723 );
and \U$15410 ( \15725 , \4771 , \4806 );
and \U$15411 ( \15726 , \4469 , \4804 );
nor \U$15412 ( \15727 , \15725 , \15726 );
xnor \U$15413 ( \15728 , \15727 , \4574 );
and \U$15414 ( \15729 , \5248 , \4355 );
and \U$15415 ( \15730 , \4779 , \4353 );
nor \U$15416 ( \15731 , \15729 , \15730 );
xnor \U$15417 ( \15732 , \15731 , \4212 );
and \U$15418 ( \15733 , \15728 , \15732 );
and \U$15419 ( \15734 , \5517 , \4032 );
and \U$15420 ( \15735 , \5253 , \4030 );
nor \U$15421 ( \15736 , \15734 , \15735 );
xnor \U$15422 ( \15737 , \15736 , \3786 );
and \U$15423 ( \15738 , \15732 , \15737 );
and \U$15424 ( \15739 , \15728 , \15737 );
or \U$15425 ( \15740 , \15733 , \15738 , \15739 );
and \U$15426 ( \15741 , \15724 , \15740 );
and \U$15427 ( \15742 , \3681 , \6235 );
and \U$15428 ( \15743 , \3264 , \6233 );
nor \U$15429 ( \15744 , \15742 , \15743 );
xnor \U$15430 ( \15745 , \15744 , \5895 );
and \U$15431 ( \15746 , \4011 , \5646 );
and \U$15432 ( \15747 , \3889 , \5644 );
nor \U$15433 ( \15748 , \15746 , \15747 );
xnor \U$15434 ( \15749 , \15748 , \5405 );
and \U$15435 ( \15750 , \15745 , \15749 );
and \U$15436 ( \15751 , \4272 , \5180 );
and \U$15437 ( \15752 , \4016 , \5178 );
nor \U$15438 ( \15753 , \15751 , \15752 );
xnor \U$15439 ( \15754 , \15753 , \4992 );
and \U$15440 ( \15755 , \15749 , \15754 );
and \U$15441 ( \15756 , \15745 , \15754 );
or \U$15442 ( \15757 , \15750 , \15755 , \15756 );
and \U$15443 ( \15758 , \15740 , \15757 );
and \U$15444 ( \15759 , \15724 , \15757 );
or \U$15445 ( \15760 , \15741 , \15758 , \15759 );
and \U$15446 ( \15761 , \1791 , \9433 );
and \U$15447 ( \15762 , \1615 , \9431 );
nor \U$15448 ( \15763 , \15761 , \15762 );
xnor \U$15449 ( \15764 , \15763 , \9123 );
and \U$15450 ( \15765 , \2042 , \8896 );
and \U$15451 ( \15766 , \1799 , \8894 );
nor \U$15452 ( \15767 , \15765 , \15766 );
xnor \U$15453 ( \15768 , \15767 , \8525 );
and \U$15454 ( \15769 , \15764 , \15768 );
and \U$15455 ( \15770 , \2233 , \8334 );
and \U$15456 ( \15771 , \2047 , \8332 );
nor \U$15457 ( \15772 , \15770 , \15771 );
xnor \U$15458 ( \15773 , \15772 , \8016 );
and \U$15459 ( \15774 , \15768 , \15773 );
and \U$15460 ( \15775 , \15764 , \15773 );
or \U$15461 ( \15776 , \15769 , \15774 , \15775 );
and \U$15462 ( \15777 , \1379 , \10814 );
and \U$15463 ( \15778 , \1274 , \10811 );
nor \U$15464 ( \15779 , \15777 , \15778 );
xnor \U$15465 ( \15780 , \15779 , \9759 );
and \U$15466 ( \15781 , \1500 , \10001 );
and \U$15467 ( \15782 , \1384 , \9999 );
nor \U$15468 ( \15783 , \15781 , \15782 );
xnor \U$15469 ( \15784 , \15783 , \9762 );
and \U$15470 ( \15785 , \15780 , \15784 );
and \U$15471 ( \15786 , \15784 , \1082 );
and \U$15472 ( \15787 , \15780 , \1082 );
or \U$15473 ( \15788 , \15785 , \15786 , \15787 );
and \U$15474 ( \15789 , \15776 , \15788 );
and \U$15475 ( \15790 , \2641 , \7767 );
and \U$15476 ( \15791 , \2377 , \7765 );
nor \U$15477 ( \15792 , \15790 , \15791 );
xnor \U$15478 ( \15793 , \15792 , \7518 );
and \U$15479 ( \15794 , \2840 , \7238 );
and \U$15480 ( \15795 , \2666 , \7236 );
nor \U$15481 ( \15796 , \15794 , \15795 );
xnor \U$15482 ( \15797 , \15796 , \6978 );
and \U$15483 ( \15798 , \15793 , \15797 );
and \U$15484 ( \15799 , \3145 , \6744 );
and \U$15485 ( \15800 , \3007 , \6742 );
nor \U$15486 ( \15801 , \15799 , \15800 );
xnor \U$15487 ( \15802 , \15801 , \6429 );
and \U$15488 ( \15803 , \15797 , \15802 );
and \U$15489 ( \15804 , \15793 , \15802 );
or \U$15490 ( \15805 , \15798 , \15803 , \15804 );
and \U$15491 ( \15806 , \15788 , \15805 );
and \U$15492 ( \15807 , \15776 , \15805 );
or \U$15493 ( \15808 , \15789 , \15806 , \15807 );
and \U$15494 ( \15809 , \15760 , \15808 );
and \U$15495 ( \15810 , \7703 , \2596 );
and \U$15496 ( \15811 , \7177 , \2594 );
nor \U$15497 ( \15812 , \15810 , \15811 );
xnor \U$15498 ( \15813 , \15812 , \2454 );
and \U$15499 ( \15814 , \8373 , \2300 );
and \U$15500 ( \15815 , \8127 , \2298 );
nor \U$15501 ( \15816 , \15814 , \15815 );
xnor \U$15502 ( \15817 , \15816 , \2163 );
and \U$15503 ( \15818 , \15813 , \15817 );
and \U$15504 ( \15819 , \8697 , \2094 );
and \U$15505 ( \15820 , \8378 , \2092 );
nor \U$15506 ( \15821 , \15819 , \15820 );
xnor \U$15507 ( \15822 , \15821 , \1942 );
and \U$15508 ( \15823 , \15817 , \15822 );
and \U$15509 ( \15824 , \15813 , \15822 );
or \U$15510 ( \15825 , \15818 , \15823 , \15824 );
and \U$15511 ( \15826 , \9550 , \1826 );
and \U$15512 ( \15827 , \8981 , \1824 );
nor \U$15513 ( \15828 , \15826 , \15827 );
xnor \U$15514 ( \15829 , \15828 , \1670 );
and \U$15515 ( \15830 , \10161 , \1554 );
and \U$15516 ( \15831 , \9558 , \1552 );
nor \U$15517 ( \15832 , \15830 , \15831 );
xnor \U$15518 ( \15833 , \15832 , \1441 );
and \U$15519 ( \15834 , \15829 , \15833 );
and \U$15520 ( \15835 , \10347 , \1360 );
and \U$15521 ( \15836 , \10166 , \1358 );
nor \U$15522 ( \15837 , \15835 , \15836 );
xnor \U$15523 ( \15838 , \15837 , \1224 );
and \U$15524 ( \15839 , \15833 , \15838 );
and \U$15525 ( \15840 , \15829 , \15838 );
or \U$15526 ( \15841 , \15834 , \15839 , \15840 );
and \U$15527 ( \15842 , \15825 , \15841 );
xor \U$15528 ( \15843 , \15512 , \15516 );
xor \U$15529 ( \15844 , \15843 , \15521 );
and \U$15530 ( \15845 , \15841 , \15844 );
and \U$15531 ( \15846 , \15825 , \15844 );
or \U$15532 ( \15847 , \15842 , \15845 , \15846 );
and \U$15533 ( \15848 , \15808 , \15847 );
and \U$15534 ( \15849 , \15760 , \15847 );
or \U$15535 ( \15850 , \15809 , \15848 , \15849 );
xor \U$15536 ( \15851 , \15496 , \15500 );
xor \U$15537 ( \15852 , \15851 , \15505 );
xor \U$15538 ( \15853 , \15589 , \15593 );
xor \U$15539 ( \15854 , \15853 , \15598 );
and \U$15540 ( \15855 , \15852 , \15854 );
xor \U$15541 ( \15856 , \15605 , \15609 );
xor \U$15542 ( \15857 , \15856 , \15614 );
and \U$15543 ( \15858 , \15854 , \15857 );
and \U$15544 ( \15859 , \15852 , \15857 );
or \U$15545 ( \15860 , \15855 , \15858 , \15859 );
xor \U$15546 ( \15861 , \15552 , \15556 );
xor \U$15547 ( \15862 , \15861 , \15561 );
xor \U$15548 ( \15863 , \15622 , \15626 );
xor \U$15549 ( \15864 , \15863 , \15631 );
and \U$15550 ( \15865 , \15862 , \15864 );
xor \U$15551 ( \15866 , \15569 , \15573 );
xor \U$15552 ( \15867 , \15866 , \15578 );
and \U$15553 ( \15868 , \15864 , \15867 );
and \U$15554 ( \15869 , \15862 , \15867 );
or \U$15555 ( \15870 , \15865 , \15868 , \15869 );
and \U$15556 ( \15871 , \15860 , \15870 );
xor \U$15557 ( \15872 , \15460 , \15462 );
xor \U$15558 ( \15873 , \15872 , \15465 );
and \U$15559 ( \15874 , \15870 , \15873 );
and \U$15560 ( \15875 , \15860 , \15873 );
or \U$15561 ( \15876 , \15871 , \15874 , \15875 );
and \U$15562 ( \15877 , \15850 , \15876 );
xor \U$15563 ( \15878 , \15508 , \15524 );
xor \U$15564 ( \15879 , \15878 , \15529 );
xor \U$15565 ( \15880 , \15470 , \15472 );
xor \U$15566 ( \15881 , \15880 , \15475 );
and \U$15567 ( \15882 , \15879 , \15881 );
xor \U$15568 ( \15883 , \15481 , \15483 );
xor \U$15569 ( \15884 , \15883 , \15486 );
and \U$15570 ( \15885 , \15881 , \15884 );
and \U$15571 ( \15886 , \15879 , \15884 );
or \U$15572 ( \15887 , \15882 , \15885 , \15886 );
and \U$15573 ( \15888 , \15876 , \15887 );
and \U$15574 ( \15889 , \15850 , \15887 );
or \U$15575 ( \15890 , \15877 , \15888 , \15889 );
xor \U$15576 ( \15891 , \15468 , \15478 );
xor \U$15577 ( \15892 , \15891 , \15489 );
xor \U$15578 ( \15893 , \15655 , \15657 );
xor \U$15579 ( \15894 , \15893 , \15660 );
and \U$15580 ( \15895 , \15892 , \15894 );
xor \U$15581 ( \15896 , \15643 , \15645 );
xor \U$15582 ( \15897 , \15896 , \15647 );
and \U$15583 ( \15898 , \15894 , \15897 );
and \U$15584 ( \15899 , \15892 , \15897 );
or \U$15585 ( \15900 , \15895 , \15898 , \15899 );
and \U$15586 ( \15901 , \15890 , \15900 );
xor \U$15587 ( \15902 , \15382 , \15392 );
xor \U$15588 ( \15903 , \15902 , \15398 );
and \U$15589 ( \15904 , \15900 , \15903 );
and \U$15590 ( \15905 , \15890 , \15903 );
or \U$15591 ( \15906 , \15901 , \15904 , \15905 );
xor \U$15592 ( \15907 , \15276 , \15316 );
xor \U$15593 ( \15908 , \15907 , \15369 );
xor \U$15594 ( \15909 , \15492 , \15640 );
xor \U$15595 ( \15910 , \15909 , \15650 );
and \U$15596 ( \15911 , \15908 , \15910 );
xor \U$15597 ( \15912 , \15663 , \15665 );
xor \U$15598 ( \15913 , \15912 , \15668 );
and \U$15599 ( \15914 , \15910 , \15913 );
and \U$15600 ( \15915 , \15908 , \15913 );
or \U$15601 ( \15916 , \15911 , \15914 , \15915 );
and \U$15602 ( \15917 , \15906 , \15916 );
xor \U$15603 ( \15918 , \15679 , \15681 );
xor \U$15604 ( \15919 , \15918 , \15684 );
and \U$15605 ( \15920 , \15916 , \15919 );
and \U$15606 ( \15921 , \15906 , \15919 );
or \U$15607 ( \15922 , \15917 , \15920 , \15921 );
xor \U$15608 ( \15923 , \15677 , \15687 );
xor \U$15609 ( \15924 , \15923 , \15690 );
and \U$15610 ( \15925 , \15922 , \15924 );
xor \U$15611 ( \15926 , \15695 , \15697 );
and \U$15612 ( \15927 , \15924 , \15926 );
and \U$15613 ( \15928 , \15922 , \15926 );
or \U$15614 ( \15929 , \15925 , \15927 , \15928 );
and \U$15615 ( \15930 , \15708 , \15929 );
xor \U$15616 ( \15931 , \15708 , \15929 );
xor \U$15617 ( \15932 , \15922 , \15924 );
xor \U$15618 ( \15933 , \15932 , \15926 );
and \U$15619 ( \15934 , \4016 , \5646 );
and \U$15620 ( \15935 , \4011 , \5644 );
nor \U$15621 ( \15936 , \15934 , \15935 );
xnor \U$15622 ( \15937 , \15936 , \5405 );
and \U$15623 ( \15938 , \4469 , \5180 );
and \U$15624 ( \15939 , \4272 , \5178 );
nor \U$15625 ( \15940 , \15938 , \15939 );
xnor \U$15626 ( \15941 , \15940 , \4992 );
and \U$15627 ( \15942 , \15937 , \15941 );
and \U$15628 ( \15943 , \4779 , \4806 );
and \U$15629 ( \15944 , \4771 , \4804 );
nor \U$15630 ( \15945 , \15943 , \15944 );
xnor \U$15631 ( \15946 , \15945 , \4574 );
and \U$15632 ( \15947 , \15941 , \15946 );
and \U$15633 ( \15948 , \15937 , \15946 );
or \U$15634 ( \15949 , \15942 , \15947 , \15948 );
and \U$15635 ( \15950 , \5253 , \4355 );
and \U$15636 ( \15951 , \5248 , \4353 );
nor \U$15637 ( \15952 , \15950 , \15951 );
xnor \U$15638 ( \15953 , \15952 , \4212 );
and \U$15639 ( \15954 , \5776 , \4032 );
and \U$15640 ( \15955 , \5517 , \4030 );
nor \U$15641 ( \15956 , \15954 , \15955 );
xnor \U$15642 ( \15957 , \15956 , \3786 );
and \U$15643 ( \15958 , \15953 , \15957 );
and \U$15644 ( \15959 , \6157 , \3637 );
and \U$15645 ( \15960 , \6148 , \3635 );
nor \U$15646 ( \15961 , \15959 , \15960 );
xnor \U$15647 ( \15962 , \15961 , \3450 );
and \U$15648 ( \15963 , \15957 , \15962 );
and \U$15649 ( \15964 , \15953 , \15962 );
or \U$15650 ( \15965 , \15958 , \15963 , \15964 );
and \U$15651 ( \15966 , \15949 , \15965 );
and \U$15652 ( \15967 , \6702 , \3324 );
and \U$15653 ( \15968 , \6500 , \3322 );
nor \U$15654 ( \15969 , \15967 , \15968 );
xnor \U$15655 ( \15970 , \15969 , \3119 );
and \U$15656 ( \15971 , \7177 , \2918 );
and \U$15657 ( \15972 , \7005 , \2916 );
nor \U$15658 ( \15973 , \15971 , \15972 );
xnor \U$15659 ( \15974 , \15973 , \2769 );
and \U$15660 ( \15975 , \15970 , \15974 );
and \U$15661 ( \15976 , \8127 , \2596 );
and \U$15662 ( \15977 , \7703 , \2594 );
nor \U$15663 ( \15978 , \15976 , \15977 );
xnor \U$15664 ( \15979 , \15978 , \2454 );
and \U$15665 ( \15980 , \15974 , \15979 );
and \U$15666 ( \15981 , \15970 , \15979 );
or \U$15667 ( \15982 , \15975 , \15980 , \15981 );
and \U$15668 ( \15983 , \15965 , \15982 );
and \U$15669 ( \15984 , \15949 , \15982 );
or \U$15670 ( \15985 , \15966 , \15983 , \15984 );
and \U$15671 ( \15986 , \2047 , \8896 );
and \U$15672 ( \15987 , \2042 , \8894 );
nor \U$15673 ( \15988 , \15986 , \15987 );
xnor \U$15674 ( \15989 , \15988 , \8525 );
and \U$15675 ( \15990 , \2377 , \8334 );
and \U$15676 ( \15991 , \2233 , \8332 );
nor \U$15677 ( \15992 , \15990 , \15991 );
xnor \U$15678 ( \15993 , \15992 , \8016 );
and \U$15679 ( \15994 , \15989 , \15993 );
and \U$15680 ( \15995 , \2666 , \7767 );
and \U$15681 ( \15996 , \2641 , \7765 );
nor \U$15682 ( \15997 , \15995 , \15996 );
xnor \U$15683 ( \15998 , \15997 , \7518 );
and \U$15684 ( \15999 , \15993 , \15998 );
and \U$15685 ( \16000 , \15989 , \15998 );
or \U$15686 ( \16001 , \15994 , \15999 , \16000 );
and \U$15687 ( \16002 , \3007 , \7238 );
and \U$15688 ( \16003 , \2840 , \7236 );
nor \U$15689 ( \16004 , \16002 , \16003 );
xnor \U$15690 ( \16005 , \16004 , \6978 );
and \U$15691 ( \16006 , \3264 , \6744 );
and \U$15692 ( \16007 , \3145 , \6742 );
nor \U$15693 ( \16008 , \16006 , \16007 );
xnor \U$15694 ( \16009 , \16008 , \6429 );
and \U$15695 ( \16010 , \16005 , \16009 );
and \U$15696 ( \16011 , \3889 , \6235 );
and \U$15697 ( \16012 , \3681 , \6233 );
nor \U$15698 ( \16013 , \16011 , \16012 );
xnor \U$15699 ( \16014 , \16013 , \5895 );
and \U$15700 ( \16015 , \16009 , \16014 );
and \U$15701 ( \16016 , \16005 , \16014 );
or \U$15702 ( \16017 , \16010 , \16015 , \16016 );
and \U$15703 ( \16018 , \16001 , \16017 );
and \U$15704 ( \16019 , \1384 , \10814 );
and \U$15705 ( \16020 , \1379 , \10811 );
nor \U$15706 ( \16021 , \16019 , \16020 );
xnor \U$15707 ( \16022 , \16021 , \9759 );
and \U$15708 ( \16023 , \1615 , \10001 );
and \U$15709 ( \16024 , \1500 , \9999 );
nor \U$15710 ( \16025 , \16023 , \16024 );
xnor \U$15711 ( \16026 , \16025 , \9762 );
and \U$15712 ( \16027 , \16022 , \16026 );
and \U$15713 ( \16028 , \1799 , \9433 );
and \U$15714 ( \16029 , \1791 , \9431 );
nor \U$15715 ( \16030 , \16028 , \16029 );
xnor \U$15716 ( \16031 , \16030 , \9123 );
and \U$15717 ( \16032 , \16026 , \16031 );
and \U$15718 ( \16033 , \16022 , \16031 );
or \U$15719 ( \16034 , \16027 , \16032 , \16033 );
and \U$15720 ( \16035 , \16017 , \16034 );
and \U$15721 ( \16036 , \16001 , \16034 );
or \U$15722 ( \16037 , \16018 , \16035 , \16036 );
and \U$15723 ( \16038 , \15985 , \16037 );
and \U$15724 ( \16039 , \8378 , \2300 );
and \U$15725 ( \16040 , \8373 , \2298 );
nor \U$15726 ( \16041 , \16039 , \16040 );
xnor \U$15727 ( \16042 , \16041 , \2163 );
and \U$15728 ( \16043 , \8981 , \2094 );
and \U$15729 ( \16044 , \8697 , \2092 );
nor \U$15730 ( \16045 , \16043 , \16044 );
xnor \U$15731 ( \16046 , \16045 , \1942 );
and \U$15732 ( \16047 , \16042 , \16046 );
and \U$15733 ( \16048 , \9558 , \1826 );
and \U$15734 ( \16049 , \9550 , \1824 );
nor \U$15735 ( \16050 , \16048 , \16049 );
xnor \U$15736 ( \16051 , \16050 , \1670 );
and \U$15737 ( \16052 , \16046 , \16051 );
and \U$15738 ( \16053 , \16042 , \16051 );
or \U$15739 ( \16054 , \16047 , \16052 , \16053 );
nand \U$15740 ( \16055 , \10967 , \1158 );
xnor \U$15741 ( \16056 , \16055 , \1082 );
and \U$15742 ( \16057 , \16054 , \16056 );
xor \U$15743 ( \16058 , \15829 , \15833 );
xor \U$15744 ( \16059 , \16058 , \15838 );
and \U$15745 ( \16060 , \16056 , \16059 );
and \U$15746 ( \16061 , \16054 , \16059 );
or \U$15747 ( \16062 , \16057 , \16060 , \16061 );
and \U$15748 ( \16063 , \16037 , \16062 );
and \U$15749 ( \16064 , \15985 , \16062 );
or \U$15750 ( \16065 , \16038 , \16063 , \16064 );
xor \U$15751 ( \16066 , \15712 , \15716 );
xor \U$15752 ( \16067 , \16066 , \15721 );
xor \U$15753 ( \16068 , \15813 , \15817 );
xor \U$15754 ( \16069 , \16068 , \15822 );
and \U$15755 ( \16070 , \16067 , \16069 );
xor \U$15756 ( \16071 , \15728 , \15732 );
xor \U$15757 ( \16072 , \16071 , \15737 );
and \U$15758 ( \16073 , \16069 , \16072 );
and \U$15759 ( \16074 , \16067 , \16072 );
or \U$15760 ( \16075 , \16070 , \16073 , \16074 );
xor \U$15761 ( \16076 , \15764 , \15768 );
xor \U$15762 ( \16077 , \16076 , \15773 );
xor \U$15763 ( \16078 , \15745 , \15749 );
xor \U$15764 ( \16079 , \16078 , \15754 );
and \U$15765 ( \16080 , \16077 , \16079 );
xor \U$15766 ( \16081 , \15793 , \15797 );
xor \U$15767 ( \16082 , \16081 , \15802 );
and \U$15768 ( \16083 , \16079 , \16082 );
and \U$15769 ( \16084 , \16077 , \16082 );
or \U$15770 ( \16085 , \16080 , \16083 , \16084 );
and \U$15771 ( \16086 , \16075 , \16085 );
xor \U$15772 ( \16087 , \15536 , \15540 );
xor \U$15773 ( \16088 , \16087 , \15545 );
and \U$15774 ( \16089 , \16085 , \16088 );
and \U$15775 ( \16090 , \16075 , \16088 );
or \U$15776 ( \16091 , \16086 , \16089 , \16090 );
and \U$15777 ( \16092 , \16065 , \16091 );
xor \U$15778 ( \16093 , \15852 , \15854 );
xor \U$15779 ( \16094 , \16093 , \15857 );
xor \U$15780 ( \16095 , \15862 , \15864 );
xor \U$15781 ( \16096 , \16095 , \15867 );
and \U$15782 ( \16097 , \16094 , \16096 );
xor \U$15783 ( \16098 , \15825 , \15841 );
xor \U$15784 ( \16099 , \16098 , \15844 );
and \U$15785 ( \16100 , \16096 , \16099 );
and \U$15786 ( \16101 , \16094 , \16099 );
or \U$15787 ( \16102 , \16097 , \16100 , \16101 );
and \U$15788 ( \16103 , \16091 , \16102 );
and \U$15789 ( \16104 , \16065 , \16102 );
or \U$15790 ( \16105 , \16092 , \16103 , \16104 );
xor \U$15791 ( \16106 , \15548 , \15564 );
xor \U$15792 ( \16107 , \16106 , \15581 );
xor \U$15793 ( \16108 , \15601 , \15617 );
xor \U$15794 ( \16109 , \16108 , \15634 );
and \U$15795 ( \16110 , \16107 , \16109 );
xor \U$15796 ( \16111 , \15879 , \15881 );
xor \U$15797 ( \16112 , \16111 , \15884 );
and \U$15798 ( \16113 , \16109 , \16112 );
and \U$15799 ( \16114 , \16107 , \16112 );
or \U$15800 ( \16115 , \16110 , \16113 , \16114 );
and \U$15801 ( \16116 , \16105 , \16115 );
xor \U$15802 ( \16117 , \15760 , \15808 );
xor \U$15803 ( \16118 , \16117 , \15847 );
xor \U$15804 ( \16119 , \15860 , \15870 );
xor \U$15805 ( \16120 , \16119 , \15873 );
and \U$15806 ( \16121 , \16118 , \16120 );
and \U$15807 ( \16122 , \16115 , \16121 );
and \U$15808 ( \16123 , \16105 , \16121 );
or \U$15809 ( \16124 , \16116 , \16122 , \16123 );
xor \U$15810 ( \16125 , \15532 , \15584 );
xor \U$15811 ( \16126 , \16125 , \15637 );
xor \U$15812 ( \16127 , \15850 , \15876 );
xor \U$15813 ( \16128 , \16127 , \15887 );
and \U$15814 ( \16129 , \16126 , \16128 );
xor \U$15815 ( \16130 , \15892 , \15894 );
xor \U$15816 ( \16131 , \16130 , \15897 );
and \U$15817 ( \16132 , \16128 , \16131 );
and \U$15818 ( \16133 , \16126 , \16131 );
or \U$15819 ( \16134 , \16129 , \16132 , \16133 );
and \U$15820 ( \16135 , \16124 , \16134 );
xor \U$15821 ( \16136 , \15908 , \15910 );
xor \U$15822 ( \16137 , \16136 , \15913 );
and \U$15823 ( \16138 , \16134 , \16137 );
and \U$15824 ( \16139 , \16124 , \16137 );
or \U$15825 ( \16140 , \16135 , \16138 , \16139 );
xor \U$15826 ( \16141 , \15653 , \15671 );
xor \U$15827 ( \16142 , \16141 , \15674 );
and \U$15828 ( \16143 , \16140 , \16142 );
xor \U$15829 ( \16144 , \15906 , \15916 );
xor \U$15830 ( \16145 , \16144 , \15919 );
and \U$15831 ( \16146 , \16142 , \16145 );
and \U$15832 ( \16147 , \16140 , \16145 );
or \U$15833 ( \16148 , \16143 , \16146 , \16147 );
and \U$15834 ( \16149 , \15933 , \16148 );
xor \U$15835 ( \16150 , \15933 , \16148 );
xor \U$15836 ( \16151 , \16140 , \16142 );
xor \U$15837 ( \16152 , \16151 , \16145 );
and \U$15838 ( \16153 , \1500 , \10814 );
and \U$15839 ( \16154 , \1384 , \10811 );
nor \U$15840 ( \16155 , \16153 , \16154 );
xnor \U$15841 ( \16156 , \16155 , \9759 );
and \U$15842 ( \16157 , \1791 , \10001 );
and \U$15843 ( \16158 , \1615 , \9999 );
nor \U$15844 ( \16159 , \16157 , \16158 );
xnor \U$15845 ( \16160 , \16159 , \9762 );
and \U$15846 ( \16161 , \16156 , \16160 );
and \U$15847 ( \16162 , \16160 , \1224 );
and \U$15848 ( \16163 , \16156 , \1224 );
or \U$15849 ( \16164 , \16161 , \16162 , \16163 );
and \U$15850 ( \16165 , \2840 , \7767 );
and \U$15851 ( \16166 , \2666 , \7765 );
nor \U$15852 ( \16167 , \16165 , \16166 );
xnor \U$15853 ( \16168 , \16167 , \7518 );
and \U$15854 ( \16169 , \3145 , \7238 );
and \U$15855 ( \16170 , \3007 , \7236 );
nor \U$15856 ( \16171 , \16169 , \16170 );
xnor \U$15857 ( \16172 , \16171 , \6978 );
and \U$15858 ( \16173 , \16168 , \16172 );
and \U$15859 ( \16174 , \3681 , \6744 );
and \U$15860 ( \16175 , \3264 , \6742 );
nor \U$15861 ( \16176 , \16174 , \16175 );
xnor \U$15862 ( \16177 , \16176 , \6429 );
and \U$15863 ( \16178 , \16172 , \16177 );
and \U$15864 ( \16179 , \16168 , \16177 );
or \U$15865 ( \16180 , \16173 , \16178 , \16179 );
and \U$15866 ( \16181 , \16164 , \16180 );
and \U$15867 ( \16182 , \2042 , \9433 );
and \U$15868 ( \16183 , \1799 , \9431 );
nor \U$15869 ( \16184 , \16182 , \16183 );
xnor \U$15870 ( \16185 , \16184 , \9123 );
and \U$15871 ( \16186 , \2233 , \8896 );
and \U$15872 ( \16187 , \2047 , \8894 );
nor \U$15873 ( \16188 , \16186 , \16187 );
xnor \U$15874 ( \16189 , \16188 , \8525 );
and \U$15875 ( \16190 , \16185 , \16189 );
and \U$15876 ( \16191 , \2641 , \8334 );
and \U$15877 ( \16192 , \2377 , \8332 );
nor \U$15878 ( \16193 , \16191 , \16192 );
xnor \U$15879 ( \16194 , \16193 , \8016 );
and \U$15880 ( \16195 , \16189 , \16194 );
and \U$15881 ( \16196 , \16185 , \16194 );
or \U$15882 ( \16197 , \16190 , \16195 , \16196 );
and \U$15883 ( \16198 , \16180 , \16197 );
and \U$15884 ( \16199 , \16164 , \16197 );
or \U$15885 ( \16200 , \16181 , \16198 , \16199 );
and \U$15886 ( \16201 , \4011 , \6235 );
and \U$15887 ( \16202 , \3889 , \6233 );
nor \U$15888 ( \16203 , \16201 , \16202 );
xnor \U$15889 ( \16204 , \16203 , \5895 );
and \U$15890 ( \16205 , \4272 , \5646 );
and \U$15891 ( \16206 , \4016 , \5644 );
nor \U$15892 ( \16207 , \16205 , \16206 );
xnor \U$15893 ( \16208 , \16207 , \5405 );
and \U$15894 ( \16209 , \16204 , \16208 );
and \U$15895 ( \16210 , \4771 , \5180 );
and \U$15896 ( \16211 , \4469 , \5178 );
nor \U$15897 ( \16212 , \16210 , \16211 );
xnor \U$15898 ( \16213 , \16212 , \4992 );
and \U$15899 ( \16214 , \16208 , \16213 );
and \U$15900 ( \16215 , \16204 , \16213 );
or \U$15901 ( \16216 , \16209 , \16214 , \16215 );
and \U$15902 ( \16217 , \5248 , \4806 );
and \U$15903 ( \16218 , \4779 , \4804 );
nor \U$15904 ( \16219 , \16217 , \16218 );
xnor \U$15905 ( \16220 , \16219 , \4574 );
and \U$15906 ( \16221 , \5517 , \4355 );
and \U$15907 ( \16222 , \5253 , \4353 );
nor \U$15908 ( \16223 , \16221 , \16222 );
xnor \U$15909 ( \16224 , \16223 , \4212 );
and \U$15910 ( \16225 , \16220 , \16224 );
and \U$15911 ( \16226 , \6148 , \4032 );
and \U$15912 ( \16227 , \5776 , \4030 );
nor \U$15913 ( \16228 , \16226 , \16227 );
xnor \U$15914 ( \16229 , \16228 , \3786 );
and \U$15915 ( \16230 , \16224 , \16229 );
and \U$15916 ( \16231 , \16220 , \16229 );
or \U$15917 ( \16232 , \16225 , \16230 , \16231 );
and \U$15918 ( \16233 , \16216 , \16232 );
and \U$15919 ( \16234 , \6500 , \3637 );
and \U$15920 ( \16235 , \6157 , \3635 );
nor \U$15921 ( \16236 , \16234 , \16235 );
xnor \U$15922 ( \16237 , \16236 , \3450 );
and \U$15923 ( \16238 , \7005 , \3324 );
and \U$15924 ( \16239 , \6702 , \3322 );
nor \U$15925 ( \16240 , \16238 , \16239 );
xnor \U$15926 ( \16241 , \16240 , \3119 );
and \U$15927 ( \16242 , \16237 , \16241 );
and \U$15928 ( \16243 , \7703 , \2918 );
and \U$15929 ( \16244 , \7177 , \2916 );
nor \U$15930 ( \16245 , \16243 , \16244 );
xnor \U$15931 ( \16246 , \16245 , \2769 );
and \U$15932 ( \16247 , \16241 , \16246 );
and \U$15933 ( \16248 , \16237 , \16246 );
or \U$15934 ( \16249 , \16242 , \16247 , \16248 );
and \U$15935 ( \16250 , \16232 , \16249 );
and \U$15936 ( \16251 , \16216 , \16249 );
or \U$15937 ( \16252 , \16233 , \16250 , \16251 );
and \U$15938 ( \16253 , \16200 , \16252 );
and \U$15939 ( \16254 , \10161 , \1826 );
and \U$15940 ( \16255 , \9558 , \1824 );
nor \U$15941 ( \16256 , \16254 , \16255 );
xnor \U$15942 ( \16257 , \16256 , \1670 );
and \U$15943 ( \16258 , \10347 , \1554 );
and \U$15944 ( \16259 , \10166 , \1552 );
nor \U$15945 ( \16260 , \16258 , \16259 );
xnor \U$15946 ( \16261 , \16260 , \1441 );
and \U$15947 ( \16262 , \16257 , \16261 );
nand \U$15948 ( \16263 , \10967 , \1358 );
xnor \U$15949 ( \16264 , \16263 , \1224 );
and \U$15950 ( \16265 , \16261 , \16264 );
and \U$15951 ( \16266 , \16257 , \16264 );
or \U$15952 ( \16267 , \16262 , \16265 , \16266 );
and \U$15953 ( \16268 , \8373 , \2596 );
and \U$15954 ( \16269 , \8127 , \2594 );
nor \U$15955 ( \16270 , \16268 , \16269 );
xnor \U$15956 ( \16271 , \16270 , \2454 );
and \U$15957 ( \16272 , \8697 , \2300 );
and \U$15958 ( \16273 , \8378 , \2298 );
nor \U$15959 ( \16274 , \16272 , \16273 );
xnor \U$15960 ( \16275 , \16274 , \2163 );
and \U$15961 ( \16276 , \16271 , \16275 );
and \U$15962 ( \16277 , \9550 , \2094 );
and \U$15963 ( \16278 , \8981 , \2092 );
nor \U$15964 ( \16279 , \16277 , \16278 );
xnor \U$15965 ( \16280 , \16279 , \1942 );
and \U$15966 ( \16281 , \16275 , \16280 );
and \U$15967 ( \16282 , \16271 , \16280 );
or \U$15968 ( \16283 , \16276 , \16281 , \16282 );
and \U$15969 ( \16284 , \16267 , \16283 );
and \U$15970 ( \16285 , \10166 , \1554 );
and \U$15971 ( \16286 , \10161 , \1552 );
nor \U$15972 ( \16287 , \16285 , \16286 );
xnor \U$15973 ( \16288 , \16287 , \1441 );
and \U$15974 ( \16289 , \16283 , \16288 );
and \U$15975 ( \16290 , \16267 , \16288 );
or \U$15976 ( \16291 , \16284 , \16289 , \16290 );
and \U$15977 ( \16292 , \16252 , \16291 );
and \U$15978 ( \16293 , \16200 , \16291 );
or \U$15979 ( \16294 , \16253 , \16292 , \16293 );
and \U$15980 ( \16295 , \10967 , \1360 );
and \U$15981 ( \16296 , \10347 , \1358 );
nor \U$15982 ( \16297 , \16295 , \16296 );
xnor \U$15983 ( \16298 , \16297 , \1224 );
xor \U$15984 ( \16299 , \15970 , \15974 );
xor \U$15985 ( \16300 , \16299 , \15979 );
and \U$15986 ( \16301 , \16298 , \16300 );
xor \U$15987 ( \16302 , \16042 , \16046 );
xor \U$15988 ( \16303 , \16302 , \16051 );
and \U$15989 ( \16304 , \16300 , \16303 );
and \U$15990 ( \16305 , \16298 , \16303 );
or \U$15991 ( \16306 , \16301 , \16304 , \16305 );
xor \U$15992 ( \16307 , \15937 , \15941 );
xor \U$15993 ( \16308 , \16307 , \15946 );
xor \U$15994 ( \16309 , \15953 , \15957 );
xor \U$15995 ( \16310 , \16309 , \15962 );
and \U$15996 ( \16311 , \16308 , \16310 );
xor \U$15997 ( \16312 , \16005 , \16009 );
xor \U$15998 ( \16313 , \16312 , \16014 );
and \U$15999 ( \16314 , \16310 , \16313 );
and \U$16000 ( \16315 , \16308 , \16313 );
or \U$16001 ( \16316 , \16311 , \16314 , \16315 );
and \U$16002 ( \16317 , \16306 , \16316 );
xor \U$16003 ( \16318 , \15780 , \15784 );
xor \U$16004 ( \16319 , \16318 , \1082 );
and \U$16005 ( \16320 , \16316 , \16319 );
and \U$16006 ( \16321 , \16306 , \16319 );
or \U$16007 ( \16322 , \16317 , \16320 , \16321 );
and \U$16008 ( \16323 , \16294 , \16322 );
xor \U$16009 ( \16324 , \16054 , \16056 );
xor \U$16010 ( \16325 , \16324 , \16059 );
xor \U$16011 ( \16326 , \16067 , \16069 );
xor \U$16012 ( \16327 , \16326 , \16072 );
and \U$16013 ( \16328 , \16325 , \16327 );
xor \U$16014 ( \16329 , \16077 , \16079 );
xor \U$16015 ( \16330 , \16329 , \16082 );
and \U$16016 ( \16331 , \16327 , \16330 );
and \U$16017 ( \16332 , \16325 , \16330 );
or \U$16018 ( \16333 , \16328 , \16331 , \16332 );
and \U$16019 ( \16334 , \16322 , \16333 );
and \U$16020 ( \16335 , \16294 , \16333 );
or \U$16021 ( \16336 , \16323 , \16334 , \16335 );
xor \U$16022 ( \16337 , \15724 , \15740 );
xor \U$16023 ( \16338 , \16337 , \15757 );
xor \U$16024 ( \16339 , \15776 , \15788 );
xor \U$16025 ( \16340 , \16339 , \15805 );
and \U$16026 ( \16341 , \16338 , \16340 );
xor \U$16027 ( \16342 , \16094 , \16096 );
xor \U$16028 ( \16343 , \16342 , \16099 );
and \U$16029 ( \16344 , \16340 , \16343 );
and \U$16030 ( \16345 , \16338 , \16343 );
or \U$16031 ( \16346 , \16341 , \16344 , \16345 );
and \U$16032 ( \16347 , \16336 , \16346 );
xor \U$16033 ( \16348 , \15985 , \16037 );
xor \U$16034 ( \16349 , \16348 , \16062 );
xor \U$16035 ( \16350 , \16075 , \16085 );
xor \U$16036 ( \16351 , \16350 , \16088 );
and \U$16037 ( \16352 , \16349 , \16351 );
and \U$16038 ( \16353 , \16346 , \16352 );
and \U$16039 ( \16354 , \16336 , \16352 );
or \U$16040 ( \16355 , \16347 , \16353 , \16354 );
xor \U$16041 ( \16356 , \16065 , \16091 );
xor \U$16042 ( \16357 , \16356 , \16102 );
xor \U$16043 ( \16358 , \16107 , \16109 );
xor \U$16044 ( \16359 , \16358 , \16112 );
and \U$16045 ( \16360 , \16357 , \16359 );
xor \U$16046 ( \16361 , \16118 , \16120 );
and \U$16047 ( \16362 , \16359 , \16361 );
and \U$16048 ( \16363 , \16357 , \16361 );
or \U$16049 ( \16364 , \16360 , \16362 , \16363 );
and \U$16050 ( \16365 , \16355 , \16364 );
xor \U$16051 ( \16366 , \16126 , \16128 );
xor \U$16052 ( \16367 , \16366 , \16131 );
and \U$16053 ( \16368 , \16364 , \16367 );
and \U$16054 ( \16369 , \16355 , \16367 );
or \U$16055 ( \16370 , \16365 , \16368 , \16369 );
xor \U$16056 ( \16371 , \15890 , \15900 );
xor \U$16057 ( \16372 , \16371 , \15903 );
and \U$16058 ( \16373 , \16370 , \16372 );
xor \U$16059 ( \16374 , \16124 , \16134 );
xor \U$16060 ( \16375 , \16374 , \16137 );
and \U$16061 ( \16376 , \16372 , \16375 );
and \U$16062 ( \16377 , \16370 , \16375 );
or \U$16063 ( \16378 , \16373 , \16376 , \16377 );
and \U$16064 ( \16379 , \16152 , \16378 );
xor \U$16065 ( \16380 , \16152 , \16378 );
xor \U$16066 ( \16381 , \16370 , \16372 );
xor \U$16067 ( \16382 , \16381 , \16375 );
and \U$16068 ( \16383 , \1615 , \10814 );
and \U$16069 ( \16384 , \1500 , \10811 );
nor \U$16070 ( \16385 , \16383 , \16384 );
xnor \U$16071 ( \16386 , \16385 , \9759 );
and \U$16072 ( \16387 , \1799 , \10001 );
and \U$16073 ( \16388 , \1791 , \9999 );
nor \U$16074 ( \16389 , \16387 , \16388 );
xnor \U$16075 ( \16390 , \16389 , \9762 );
and \U$16076 ( \16391 , \16386 , \16390 );
and \U$16077 ( \16392 , \2047 , \9433 );
and \U$16078 ( \16393 , \2042 , \9431 );
nor \U$16079 ( \16394 , \16392 , \16393 );
xnor \U$16080 ( \16395 , \16394 , \9123 );
and \U$16081 ( \16396 , \16390 , \16395 );
and \U$16082 ( \16397 , \16386 , \16395 );
or \U$16083 ( \16398 , \16391 , \16396 , \16397 );
and \U$16084 ( \16399 , \2377 , \8896 );
and \U$16085 ( \16400 , \2233 , \8894 );
nor \U$16086 ( \16401 , \16399 , \16400 );
xnor \U$16087 ( \16402 , \16401 , \8525 );
and \U$16088 ( \16403 , \2666 , \8334 );
and \U$16089 ( \16404 , \2641 , \8332 );
nor \U$16090 ( \16405 , \16403 , \16404 );
xnor \U$16091 ( \16406 , \16405 , \8016 );
and \U$16092 ( \16407 , \16402 , \16406 );
and \U$16093 ( \16408 , \3007 , \7767 );
and \U$16094 ( \16409 , \2840 , \7765 );
nor \U$16095 ( \16410 , \16408 , \16409 );
xnor \U$16096 ( \16411 , \16410 , \7518 );
and \U$16097 ( \16412 , \16406 , \16411 );
and \U$16098 ( \16413 , \16402 , \16411 );
or \U$16099 ( \16414 , \16407 , \16412 , \16413 );
and \U$16100 ( \16415 , \16398 , \16414 );
and \U$16101 ( \16416 , \3264 , \7238 );
and \U$16102 ( \16417 , \3145 , \7236 );
nor \U$16103 ( \16418 , \16416 , \16417 );
xnor \U$16104 ( \16419 , \16418 , \6978 );
and \U$16105 ( \16420 , \3889 , \6744 );
and \U$16106 ( \16421 , \3681 , \6742 );
nor \U$16107 ( \16422 , \16420 , \16421 );
xnor \U$16108 ( \16423 , \16422 , \6429 );
and \U$16109 ( \16424 , \16419 , \16423 );
and \U$16110 ( \16425 , \4016 , \6235 );
and \U$16111 ( \16426 , \4011 , \6233 );
nor \U$16112 ( \16427 , \16425 , \16426 );
xnor \U$16113 ( \16428 , \16427 , \5895 );
and \U$16114 ( \16429 , \16423 , \16428 );
and \U$16115 ( \16430 , \16419 , \16428 );
or \U$16116 ( \16431 , \16424 , \16429 , \16430 );
and \U$16117 ( \16432 , \16414 , \16431 );
and \U$16118 ( \16433 , \16398 , \16431 );
or \U$16119 ( \16434 , \16415 , \16432 , \16433 );
and \U$16120 ( \16435 , \5776 , \4355 );
and \U$16121 ( \16436 , \5517 , \4353 );
nor \U$16122 ( \16437 , \16435 , \16436 );
xnor \U$16123 ( \16438 , \16437 , \4212 );
and \U$16124 ( \16439 , \6157 , \4032 );
and \U$16125 ( \16440 , \6148 , \4030 );
nor \U$16126 ( \16441 , \16439 , \16440 );
xnor \U$16127 ( \16442 , \16441 , \3786 );
and \U$16128 ( \16443 , \16438 , \16442 );
and \U$16129 ( \16444 , \6702 , \3637 );
and \U$16130 ( \16445 , \6500 , \3635 );
nor \U$16131 ( \16446 , \16444 , \16445 );
xnor \U$16132 ( \16447 , \16446 , \3450 );
and \U$16133 ( \16448 , \16442 , \16447 );
and \U$16134 ( \16449 , \16438 , \16447 );
or \U$16135 ( \16450 , \16443 , \16448 , \16449 );
and \U$16136 ( \16451 , \7177 , \3324 );
and \U$16137 ( \16452 , \7005 , \3322 );
nor \U$16138 ( \16453 , \16451 , \16452 );
xnor \U$16139 ( \16454 , \16453 , \3119 );
and \U$16140 ( \16455 , \8127 , \2918 );
and \U$16141 ( \16456 , \7703 , \2916 );
nor \U$16142 ( \16457 , \16455 , \16456 );
xnor \U$16143 ( \16458 , \16457 , \2769 );
and \U$16144 ( \16459 , \16454 , \16458 );
and \U$16145 ( \16460 , \8378 , \2596 );
and \U$16146 ( \16461 , \8373 , \2594 );
nor \U$16147 ( \16462 , \16460 , \16461 );
xnor \U$16148 ( \16463 , \16462 , \2454 );
and \U$16149 ( \16464 , \16458 , \16463 );
and \U$16150 ( \16465 , \16454 , \16463 );
or \U$16151 ( \16466 , \16459 , \16464 , \16465 );
and \U$16152 ( \16467 , \16450 , \16466 );
and \U$16153 ( \16468 , \4469 , \5646 );
and \U$16154 ( \16469 , \4272 , \5644 );
nor \U$16155 ( \16470 , \16468 , \16469 );
xnor \U$16156 ( \16471 , \16470 , \5405 );
and \U$16157 ( \16472 , \4779 , \5180 );
and \U$16158 ( \16473 , \4771 , \5178 );
nor \U$16159 ( \16474 , \16472 , \16473 );
xnor \U$16160 ( \16475 , \16474 , \4992 );
and \U$16161 ( \16476 , \16471 , \16475 );
and \U$16162 ( \16477 , \5253 , \4806 );
and \U$16163 ( \16478 , \5248 , \4804 );
nor \U$16164 ( \16479 , \16477 , \16478 );
xnor \U$16165 ( \16480 , \16479 , \4574 );
and \U$16166 ( \16481 , \16475 , \16480 );
and \U$16167 ( \16482 , \16471 , \16480 );
or \U$16168 ( \16483 , \16476 , \16481 , \16482 );
and \U$16169 ( \16484 , \16466 , \16483 );
and \U$16170 ( \16485 , \16450 , \16483 );
or \U$16171 ( \16486 , \16467 , \16484 , \16485 );
and \U$16172 ( \16487 , \16434 , \16486 );
and \U$16173 ( \16488 , \8981 , \2300 );
and \U$16174 ( \16489 , \8697 , \2298 );
nor \U$16175 ( \16490 , \16488 , \16489 );
xnor \U$16176 ( \16491 , \16490 , \2163 );
and \U$16177 ( \16492 , \9558 , \2094 );
and \U$16178 ( \16493 , \9550 , \2092 );
nor \U$16179 ( \16494 , \16492 , \16493 );
xnor \U$16180 ( \16495 , \16494 , \1942 );
and \U$16181 ( \16496 , \16491 , \16495 );
and \U$16182 ( \16497 , \10166 , \1826 );
and \U$16183 ( \16498 , \10161 , \1824 );
nor \U$16184 ( \16499 , \16497 , \16498 );
xnor \U$16185 ( \16500 , \16499 , \1670 );
and \U$16186 ( \16501 , \16495 , \16500 );
and \U$16187 ( \16502 , \16491 , \16500 );
or \U$16188 ( \16503 , \16496 , \16501 , \16502 );
xor \U$16189 ( \16504 , \16257 , \16261 );
xor \U$16190 ( \16505 , \16504 , \16264 );
and \U$16191 ( \16506 , \16503 , \16505 );
xor \U$16192 ( \16507 , \16271 , \16275 );
xor \U$16193 ( \16508 , \16507 , \16280 );
and \U$16194 ( \16509 , \16505 , \16508 );
and \U$16195 ( \16510 , \16503 , \16508 );
or \U$16196 ( \16511 , \16506 , \16509 , \16510 );
and \U$16197 ( \16512 , \16486 , \16511 );
and \U$16198 ( \16513 , \16434 , \16511 );
or \U$16199 ( \16514 , \16487 , \16512 , \16513 );
xor \U$16200 ( \16515 , \16204 , \16208 );
xor \U$16201 ( \16516 , \16515 , \16213 );
xor \U$16202 ( \16517 , \16220 , \16224 );
xor \U$16203 ( \16518 , \16517 , \16229 );
and \U$16204 ( \16519 , \16516 , \16518 );
xor \U$16205 ( \16520 , \16237 , \16241 );
xor \U$16206 ( \16521 , \16520 , \16246 );
and \U$16207 ( \16522 , \16518 , \16521 );
and \U$16208 ( \16523 , \16516 , \16521 );
or \U$16209 ( \16524 , \16519 , \16522 , \16523 );
xor \U$16210 ( \16525 , \16156 , \16160 );
xor \U$16211 ( \16526 , \16525 , \1224 );
xor \U$16212 ( \16527 , \16168 , \16172 );
xor \U$16213 ( \16528 , \16527 , \16177 );
and \U$16214 ( \16529 , \16526 , \16528 );
xor \U$16215 ( \16530 , \16185 , \16189 );
xor \U$16216 ( \16531 , \16530 , \16194 );
and \U$16217 ( \16532 , \16528 , \16531 );
and \U$16218 ( \16533 , \16526 , \16531 );
or \U$16219 ( \16534 , \16529 , \16532 , \16533 );
and \U$16220 ( \16535 , \16524 , \16534 );
xor \U$16221 ( \16536 , \15989 , \15993 );
xor \U$16222 ( \16537 , \16536 , \15998 );
and \U$16223 ( \16538 , \16534 , \16537 );
and \U$16224 ( \16539 , \16524 , \16537 );
or \U$16225 ( \16540 , \16535 , \16538 , \16539 );
and \U$16226 ( \16541 , \16514 , \16540 );
xor \U$16227 ( \16542 , \16022 , \16026 );
xor \U$16228 ( \16543 , \16542 , \16031 );
xor \U$16229 ( \16544 , \16298 , \16300 );
xor \U$16230 ( \16545 , \16544 , \16303 );
and \U$16231 ( \16546 , \16543 , \16545 );
xor \U$16232 ( \16547 , \16308 , \16310 );
xor \U$16233 ( \16548 , \16547 , \16313 );
and \U$16234 ( \16549 , \16545 , \16548 );
and \U$16235 ( \16550 , \16543 , \16548 );
or \U$16236 ( \16551 , \16546 , \16549 , \16550 );
and \U$16237 ( \16552 , \16540 , \16551 );
and \U$16238 ( \16553 , \16514 , \16551 );
or \U$16239 ( \16554 , \16541 , \16552 , \16553 );
xor \U$16240 ( \16555 , \16164 , \16180 );
xor \U$16241 ( \16556 , \16555 , \16197 );
xor \U$16242 ( \16557 , \16216 , \16232 );
xor \U$16243 ( \16558 , \16557 , \16249 );
and \U$16244 ( \16559 , \16556 , \16558 );
xor \U$16245 ( \16560 , \16267 , \16283 );
xor \U$16246 ( \16561 , \16560 , \16288 );
and \U$16247 ( \16562 , \16558 , \16561 );
and \U$16248 ( \16563 , \16556 , \16561 );
or \U$16249 ( \16564 , \16559 , \16562 , \16563 );
xor \U$16250 ( \16565 , \15949 , \15965 );
xor \U$16251 ( \16566 , \16565 , \15982 );
and \U$16252 ( \16567 , \16564 , \16566 );
xor \U$16253 ( \16568 , \16001 , \16017 );
xor \U$16254 ( \16569 , \16568 , \16034 );
and \U$16255 ( \16570 , \16566 , \16569 );
and \U$16256 ( \16571 , \16564 , \16569 );
or \U$16257 ( \16572 , \16567 , \16570 , \16571 );
and \U$16258 ( \16573 , \16554 , \16572 );
xor \U$16259 ( \16574 , \16200 , \16252 );
xor \U$16260 ( \16575 , \16574 , \16291 );
xor \U$16261 ( \16576 , \16306 , \16316 );
xor \U$16262 ( \16577 , \16576 , \16319 );
and \U$16263 ( \16578 , \16575 , \16577 );
xor \U$16264 ( \16579 , \16325 , \16327 );
xor \U$16265 ( \16580 , \16579 , \16330 );
and \U$16266 ( \16581 , \16577 , \16580 );
and \U$16267 ( \16582 , \16575 , \16580 );
or \U$16268 ( \16583 , \16578 , \16581 , \16582 );
and \U$16269 ( \16584 , \16572 , \16583 );
and \U$16270 ( \16585 , \16554 , \16583 );
or \U$16271 ( \16586 , \16573 , \16584 , \16585 );
xor \U$16272 ( \16587 , \16294 , \16322 );
xor \U$16273 ( \16588 , \16587 , \16333 );
xor \U$16274 ( \16589 , \16338 , \16340 );
xor \U$16275 ( \16590 , \16589 , \16343 );
and \U$16276 ( \16591 , \16588 , \16590 );
xor \U$16277 ( \16592 , \16349 , \16351 );
and \U$16278 ( \16593 , \16590 , \16592 );
and \U$16279 ( \16594 , \16588 , \16592 );
or \U$16280 ( \16595 , \16591 , \16593 , \16594 );
and \U$16281 ( \16596 , \16586 , \16595 );
xor \U$16282 ( \16597 , \16357 , \16359 );
xor \U$16283 ( \16598 , \16597 , \16361 );
and \U$16284 ( \16599 , \16595 , \16598 );
and \U$16285 ( \16600 , \16586 , \16598 );
or \U$16286 ( \16601 , \16596 , \16599 , \16600 );
xor \U$16287 ( \16602 , \16105 , \16115 );
xor \U$16288 ( \16603 , \16602 , \16121 );
and \U$16289 ( \16604 , \16601 , \16603 );
xor \U$16290 ( \16605 , \16355 , \16364 );
xor \U$16291 ( \16606 , \16605 , \16367 );
and \U$16292 ( \16607 , \16603 , \16606 );
and \U$16293 ( \16608 , \16601 , \16606 );
or \U$16294 ( \16609 , \16604 , \16607 , \16608 );
and \U$16295 ( \16610 , \16382 , \16609 );
xor \U$16296 ( \16611 , \16382 , \16609 );
xor \U$16297 ( \16612 , \16601 , \16603 );
xor \U$16298 ( \16613 , \16612 , \16606 );
and \U$16299 ( \16614 , \7005 , \3637 );
and \U$16300 ( \16615 , \6702 , \3635 );
nor \U$16301 ( \16616 , \16614 , \16615 );
xnor \U$16302 ( \16617 , \16616 , \3450 );
and \U$16303 ( \16618 , \7703 , \3324 );
and \U$16304 ( \16619 , \7177 , \3322 );
nor \U$16305 ( \16620 , \16618 , \16619 );
xnor \U$16306 ( \16621 , \16620 , \3119 );
and \U$16307 ( \16622 , \16617 , \16621 );
and \U$16308 ( \16623 , \8373 , \2918 );
and \U$16309 ( \16624 , \8127 , \2916 );
nor \U$16310 ( \16625 , \16623 , \16624 );
xnor \U$16311 ( \16626 , \16625 , \2769 );
and \U$16312 ( \16627 , \16621 , \16626 );
and \U$16313 ( \16628 , \16617 , \16626 );
or \U$16314 ( \16629 , \16622 , \16627 , \16628 );
and \U$16315 ( \16630 , \4272 , \6235 );
and \U$16316 ( \16631 , \4016 , \6233 );
nor \U$16317 ( \16632 , \16630 , \16631 );
xnor \U$16318 ( \16633 , \16632 , \5895 );
and \U$16319 ( \16634 , \4771 , \5646 );
and \U$16320 ( \16635 , \4469 , \5644 );
nor \U$16321 ( \16636 , \16634 , \16635 );
xnor \U$16322 ( \16637 , \16636 , \5405 );
and \U$16323 ( \16638 , \16633 , \16637 );
and \U$16324 ( \16639 , \5248 , \5180 );
and \U$16325 ( \16640 , \4779 , \5178 );
nor \U$16326 ( \16641 , \16639 , \16640 );
xnor \U$16327 ( \16642 , \16641 , \4992 );
and \U$16328 ( \16643 , \16637 , \16642 );
and \U$16329 ( \16644 , \16633 , \16642 );
or \U$16330 ( \16645 , \16638 , \16643 , \16644 );
and \U$16331 ( \16646 , \16629 , \16645 );
and \U$16332 ( \16647 , \5517 , \4806 );
and \U$16333 ( \16648 , \5253 , \4804 );
nor \U$16334 ( \16649 , \16647 , \16648 );
xnor \U$16335 ( \16650 , \16649 , \4574 );
and \U$16336 ( \16651 , \6148 , \4355 );
and \U$16337 ( \16652 , \5776 , \4353 );
nor \U$16338 ( \16653 , \16651 , \16652 );
xnor \U$16339 ( \16654 , \16653 , \4212 );
and \U$16340 ( \16655 , \16650 , \16654 );
and \U$16341 ( \16656 , \6500 , \4032 );
and \U$16342 ( \16657 , \6157 , \4030 );
nor \U$16343 ( \16658 , \16656 , \16657 );
xnor \U$16344 ( \16659 , \16658 , \3786 );
and \U$16345 ( \16660 , \16654 , \16659 );
and \U$16346 ( \16661 , \16650 , \16659 );
or \U$16347 ( \16662 , \16655 , \16660 , \16661 );
and \U$16348 ( \16663 , \16645 , \16662 );
and \U$16349 ( \16664 , \16629 , \16662 );
or \U$16350 ( \16665 , \16646 , \16663 , \16664 );
and \U$16351 ( \16666 , \1791 , \10814 );
and \U$16352 ( \16667 , \1615 , \10811 );
nor \U$16353 ( \16668 , \16666 , \16667 );
xnor \U$16354 ( \16669 , \16668 , \9759 );
and \U$16355 ( \16670 , \2042 , \10001 );
and \U$16356 ( \16671 , \1799 , \9999 );
nor \U$16357 ( \16672 , \16670 , \16671 );
xnor \U$16358 ( \16673 , \16672 , \9762 );
and \U$16359 ( \16674 , \16669 , \16673 );
and \U$16360 ( \16675 , \16673 , \1441 );
and \U$16361 ( \16676 , \16669 , \1441 );
or \U$16362 ( \16677 , \16674 , \16675 , \16676 );
and \U$16363 ( \16678 , \3145 , \7767 );
and \U$16364 ( \16679 , \3007 , \7765 );
nor \U$16365 ( \16680 , \16678 , \16679 );
xnor \U$16366 ( \16681 , \16680 , \7518 );
and \U$16367 ( \16682 , \3681 , \7238 );
and \U$16368 ( \16683 , \3264 , \7236 );
nor \U$16369 ( \16684 , \16682 , \16683 );
xnor \U$16370 ( \16685 , \16684 , \6978 );
and \U$16371 ( \16686 , \16681 , \16685 );
and \U$16372 ( \16687 , \4011 , \6744 );
and \U$16373 ( \16688 , \3889 , \6742 );
nor \U$16374 ( \16689 , \16687 , \16688 );
xnor \U$16375 ( \16690 , \16689 , \6429 );
and \U$16376 ( \16691 , \16685 , \16690 );
and \U$16377 ( \16692 , \16681 , \16690 );
or \U$16378 ( \16693 , \16686 , \16691 , \16692 );
and \U$16379 ( \16694 , \16677 , \16693 );
and \U$16380 ( \16695 , \2233 , \9433 );
and \U$16381 ( \16696 , \2047 , \9431 );
nor \U$16382 ( \16697 , \16695 , \16696 );
xnor \U$16383 ( \16698 , \16697 , \9123 );
and \U$16384 ( \16699 , \2641 , \8896 );
and \U$16385 ( \16700 , \2377 , \8894 );
nor \U$16386 ( \16701 , \16699 , \16700 );
xnor \U$16387 ( \16702 , \16701 , \8525 );
and \U$16388 ( \16703 , \16698 , \16702 );
and \U$16389 ( \16704 , \2840 , \8334 );
and \U$16390 ( \16705 , \2666 , \8332 );
nor \U$16391 ( \16706 , \16704 , \16705 );
xnor \U$16392 ( \16707 , \16706 , \8016 );
and \U$16393 ( \16708 , \16702 , \16707 );
and \U$16394 ( \16709 , \16698 , \16707 );
or \U$16395 ( \16710 , \16703 , \16708 , \16709 );
and \U$16396 ( \16711 , \16693 , \16710 );
and \U$16397 ( \16712 , \16677 , \16710 );
or \U$16398 ( \16713 , \16694 , \16711 , \16712 );
and \U$16399 ( \16714 , \16665 , \16713 );
and \U$16400 ( \16715 , \8697 , \2596 );
and \U$16401 ( \16716 , \8378 , \2594 );
nor \U$16402 ( \16717 , \16715 , \16716 );
xnor \U$16403 ( \16718 , \16717 , \2454 );
and \U$16404 ( \16719 , \9550 , \2300 );
and \U$16405 ( \16720 , \8981 , \2298 );
nor \U$16406 ( \16721 , \16719 , \16720 );
xnor \U$16407 ( \16722 , \16721 , \2163 );
and \U$16408 ( \16723 , \16718 , \16722 );
and \U$16409 ( \16724 , \10161 , \2094 );
and \U$16410 ( \16725 , \9558 , \2092 );
nor \U$16411 ( \16726 , \16724 , \16725 );
xnor \U$16412 ( \16727 , \16726 , \1942 );
and \U$16413 ( \16728 , \16722 , \16727 );
and \U$16414 ( \16729 , \16718 , \16727 );
or \U$16415 ( \16730 , \16723 , \16728 , \16729 );
and \U$16416 ( \16731 , \10347 , \1826 );
and \U$16417 ( \16732 , \10166 , \1824 );
nor \U$16418 ( \16733 , \16731 , \16732 );
xnor \U$16419 ( \16734 , \16733 , \1670 );
nand \U$16420 ( \16735 , \10967 , \1552 );
xnor \U$16421 ( \16736 , \16735 , \1441 );
and \U$16422 ( \16737 , \16734 , \16736 );
and \U$16423 ( \16738 , \16730 , \16737 );
and \U$16424 ( \16739 , \10967 , \1554 );
and \U$16425 ( \16740 , \10347 , \1552 );
nor \U$16426 ( \16741 , \16739 , \16740 );
xnor \U$16427 ( \16742 , \16741 , \1441 );
and \U$16428 ( \16743 , \16737 , \16742 );
and \U$16429 ( \16744 , \16730 , \16742 );
or \U$16430 ( \16745 , \16738 , \16743 , \16744 );
and \U$16431 ( \16746 , \16713 , \16745 );
and \U$16432 ( \16747 , \16665 , \16745 );
or \U$16433 ( \16748 , \16714 , \16746 , \16747 );
xor \U$16434 ( \16749 , \16402 , \16406 );
xor \U$16435 ( \16750 , \16749 , \16411 );
xor \U$16436 ( \16751 , \16471 , \16475 );
xor \U$16437 ( \16752 , \16751 , \16480 );
and \U$16438 ( \16753 , \16750 , \16752 );
xor \U$16439 ( \16754 , \16419 , \16423 );
xor \U$16440 ( \16755 , \16754 , \16428 );
and \U$16441 ( \16756 , \16752 , \16755 );
and \U$16442 ( \16757 , \16750 , \16755 );
or \U$16443 ( \16758 , \16753 , \16756 , \16757 );
xor \U$16444 ( \16759 , \16438 , \16442 );
xor \U$16445 ( \16760 , \16759 , \16447 );
xor \U$16446 ( \16761 , \16491 , \16495 );
xor \U$16447 ( \16762 , \16761 , \16500 );
and \U$16448 ( \16763 , \16760 , \16762 );
xor \U$16449 ( \16764 , \16454 , \16458 );
xor \U$16450 ( \16765 , \16764 , \16463 );
and \U$16451 ( \16766 , \16762 , \16765 );
and \U$16452 ( \16767 , \16760 , \16765 );
or \U$16453 ( \16768 , \16763 , \16766 , \16767 );
and \U$16454 ( \16769 , \16758 , \16768 );
xor \U$16455 ( \16770 , \16526 , \16528 );
xor \U$16456 ( \16771 , \16770 , \16531 );
and \U$16457 ( \16772 , \16768 , \16771 );
and \U$16458 ( \16773 , \16758 , \16771 );
or \U$16459 ( \16774 , \16769 , \16772 , \16773 );
and \U$16460 ( \16775 , \16748 , \16774 );
xor \U$16461 ( \16776 , \16450 , \16466 );
xor \U$16462 ( \16777 , \16776 , \16483 );
xor \U$16463 ( \16778 , \16516 , \16518 );
xor \U$16464 ( \16779 , \16778 , \16521 );
and \U$16465 ( \16780 , \16777 , \16779 );
xor \U$16466 ( \16781 , \16503 , \16505 );
xor \U$16467 ( \16782 , \16781 , \16508 );
and \U$16468 ( \16783 , \16779 , \16782 );
and \U$16469 ( \16784 , \16777 , \16782 );
or \U$16470 ( \16785 , \16780 , \16783 , \16784 );
and \U$16471 ( \16786 , \16774 , \16785 );
and \U$16472 ( \16787 , \16748 , \16785 );
or \U$16473 ( \16788 , \16775 , \16786 , \16787 );
xor \U$16474 ( \16789 , \16556 , \16558 );
xor \U$16475 ( \16790 , \16789 , \16561 );
xor \U$16476 ( \16791 , \16524 , \16534 );
xor \U$16477 ( \16792 , \16791 , \16537 );
and \U$16478 ( \16793 , \16790 , \16792 );
xor \U$16479 ( \16794 , \16543 , \16545 );
xor \U$16480 ( \16795 , \16794 , \16548 );
and \U$16481 ( \16796 , \16792 , \16795 );
and \U$16482 ( \16797 , \16790 , \16795 );
or \U$16483 ( \16798 , \16793 , \16796 , \16797 );
and \U$16484 ( \16799 , \16788 , \16798 );
xor \U$16485 ( \16800 , \16575 , \16577 );
xor \U$16486 ( \16801 , \16800 , \16580 );
and \U$16487 ( \16802 , \16798 , \16801 );
and \U$16488 ( \16803 , \16788 , \16801 );
or \U$16489 ( \16804 , \16799 , \16802 , \16803 );
xor \U$16490 ( \16805 , \16554 , \16572 );
xor \U$16491 ( \16806 , \16805 , \16583 );
and \U$16492 ( \16807 , \16804 , \16806 );
xor \U$16493 ( \16808 , \16588 , \16590 );
xor \U$16494 ( \16809 , \16808 , \16592 );
and \U$16495 ( \16810 , \16806 , \16809 );
and \U$16496 ( \16811 , \16804 , \16809 );
or \U$16497 ( \16812 , \16807 , \16810 , \16811 );
xor \U$16498 ( \16813 , \16336 , \16346 );
xor \U$16499 ( \16814 , \16813 , \16352 );
and \U$16500 ( \16815 , \16812 , \16814 );
xor \U$16501 ( \16816 , \16586 , \16595 );
xor \U$16502 ( \16817 , \16816 , \16598 );
and \U$16503 ( \16818 , \16814 , \16817 );
and \U$16504 ( \16819 , \16812 , \16817 );
or \U$16505 ( \16820 , \16815 , \16818 , \16819 );
and \U$16506 ( \16821 , \16613 , \16820 );
xor \U$16507 ( \16822 , \16613 , \16820 );
xor \U$16508 ( \16823 , \16812 , \16814 );
xor \U$16509 ( \16824 , \16823 , \16817 );
and \U$16510 ( \16825 , \6157 , \4355 );
and \U$16511 ( \16826 , \6148 , \4353 );
nor \U$16512 ( \16827 , \16825 , \16826 );
xnor \U$16513 ( \16828 , \16827 , \4212 );
and \U$16514 ( \16829 , \6702 , \4032 );
and \U$16515 ( \16830 , \6500 , \4030 );
nor \U$16516 ( \16831 , \16829 , \16830 );
xnor \U$16517 ( \16832 , \16831 , \3786 );
and \U$16518 ( \16833 , \16828 , \16832 );
and \U$16519 ( \16834 , \7177 , \3637 );
and \U$16520 ( \16835 , \7005 , \3635 );
nor \U$16521 ( \16836 , \16834 , \16835 );
xnor \U$16522 ( \16837 , \16836 , \3450 );
and \U$16523 ( \16838 , \16832 , \16837 );
and \U$16524 ( \16839 , \16828 , \16837 );
or \U$16525 ( \16840 , \16833 , \16838 , \16839 );
and \U$16526 ( \16841 , \8127 , \3324 );
and \U$16527 ( \16842 , \7703 , \3322 );
nor \U$16528 ( \16843 , \16841 , \16842 );
xnor \U$16529 ( \16844 , \16843 , \3119 );
and \U$16530 ( \16845 , \8378 , \2918 );
and \U$16531 ( \16846 , \8373 , \2916 );
nor \U$16532 ( \16847 , \16845 , \16846 );
xnor \U$16533 ( \16848 , \16847 , \2769 );
and \U$16534 ( \16849 , \16844 , \16848 );
and \U$16535 ( \16850 , \8981 , \2596 );
and \U$16536 ( \16851 , \8697 , \2594 );
nor \U$16537 ( \16852 , \16850 , \16851 );
xnor \U$16538 ( \16853 , \16852 , \2454 );
and \U$16539 ( \16854 , \16848 , \16853 );
and \U$16540 ( \16855 , \16844 , \16853 );
or \U$16541 ( \16856 , \16849 , \16854 , \16855 );
and \U$16542 ( \16857 , \16840 , \16856 );
and \U$16543 ( \16858 , \4779 , \5646 );
and \U$16544 ( \16859 , \4771 , \5644 );
nor \U$16545 ( \16860 , \16858 , \16859 );
xnor \U$16546 ( \16861 , \16860 , \5405 );
and \U$16547 ( \16862 , \5253 , \5180 );
and \U$16548 ( \16863 , \5248 , \5178 );
nor \U$16549 ( \16864 , \16862 , \16863 );
xnor \U$16550 ( \16865 , \16864 , \4992 );
and \U$16551 ( \16866 , \16861 , \16865 );
and \U$16552 ( \16867 , \5776 , \4806 );
and \U$16553 ( \16868 , \5517 , \4804 );
nor \U$16554 ( \16869 , \16867 , \16868 );
xnor \U$16555 ( \16870 , \16869 , \4574 );
and \U$16556 ( \16871 , \16865 , \16870 );
and \U$16557 ( \16872 , \16861 , \16870 );
or \U$16558 ( \16873 , \16866 , \16871 , \16872 );
and \U$16559 ( \16874 , \16856 , \16873 );
and \U$16560 ( \16875 , \16840 , \16873 );
or \U$16561 ( \16876 , \16857 , \16874 , \16875 );
and \U$16562 ( \16877 , \3889 , \7238 );
and \U$16563 ( \16878 , \3681 , \7236 );
nor \U$16564 ( \16879 , \16877 , \16878 );
xnor \U$16565 ( \16880 , \16879 , \6978 );
and \U$16566 ( \16881 , \4016 , \6744 );
and \U$16567 ( \16882 , \4011 , \6742 );
nor \U$16568 ( \16883 , \16881 , \16882 );
xnor \U$16569 ( \16884 , \16883 , \6429 );
and \U$16570 ( \16885 , \16880 , \16884 );
and \U$16571 ( \16886 , \4469 , \6235 );
and \U$16572 ( \16887 , \4272 , \6233 );
nor \U$16573 ( \16888 , \16886 , \16887 );
xnor \U$16574 ( \16889 , \16888 , \5895 );
and \U$16575 ( \16890 , \16884 , \16889 );
and \U$16576 ( \16891 , \16880 , \16889 );
or \U$16577 ( \16892 , \16885 , \16890 , \16891 );
and \U$16578 ( \16893 , \2666 , \8896 );
and \U$16579 ( \16894 , \2641 , \8894 );
nor \U$16580 ( \16895 , \16893 , \16894 );
xnor \U$16581 ( \16896 , \16895 , \8525 );
and \U$16582 ( \16897 , \3007 , \8334 );
and \U$16583 ( \16898 , \2840 , \8332 );
nor \U$16584 ( \16899 , \16897 , \16898 );
xnor \U$16585 ( \16900 , \16899 , \8016 );
and \U$16586 ( \16901 , \16896 , \16900 );
and \U$16587 ( \16902 , \3264 , \7767 );
and \U$16588 ( \16903 , \3145 , \7765 );
nor \U$16589 ( \16904 , \16902 , \16903 );
xnor \U$16590 ( \16905 , \16904 , \7518 );
and \U$16591 ( \16906 , \16900 , \16905 );
and \U$16592 ( \16907 , \16896 , \16905 );
or \U$16593 ( \16908 , \16901 , \16906 , \16907 );
and \U$16594 ( \16909 , \16892 , \16908 );
and \U$16595 ( \16910 , \1799 , \10814 );
and \U$16596 ( \16911 , \1791 , \10811 );
nor \U$16597 ( \16912 , \16910 , \16911 );
xnor \U$16598 ( \16913 , \16912 , \9759 );
and \U$16599 ( \16914 , \2047 , \10001 );
and \U$16600 ( \16915 , \2042 , \9999 );
nor \U$16601 ( \16916 , \16914 , \16915 );
xnor \U$16602 ( \16917 , \16916 , \9762 );
and \U$16603 ( \16918 , \16913 , \16917 );
and \U$16604 ( \16919 , \2377 , \9433 );
and \U$16605 ( \16920 , \2233 , \9431 );
nor \U$16606 ( \16921 , \16919 , \16920 );
xnor \U$16607 ( \16922 , \16921 , \9123 );
and \U$16608 ( \16923 , \16917 , \16922 );
and \U$16609 ( \16924 , \16913 , \16922 );
or \U$16610 ( \16925 , \16918 , \16923 , \16924 );
and \U$16611 ( \16926 , \16908 , \16925 );
and \U$16612 ( \16927 , \16892 , \16925 );
or \U$16613 ( \16928 , \16909 , \16926 , \16927 );
and \U$16614 ( \16929 , \16876 , \16928 );
and \U$16615 ( \16930 , \9558 , \2300 );
and \U$16616 ( \16931 , \9550 , \2298 );
nor \U$16617 ( \16932 , \16930 , \16931 );
xnor \U$16618 ( \16933 , \16932 , \2163 );
and \U$16619 ( \16934 , \10166 , \2094 );
and \U$16620 ( \16935 , \10161 , \2092 );
nor \U$16621 ( \16936 , \16934 , \16935 );
xnor \U$16622 ( \16937 , \16936 , \1942 );
and \U$16623 ( \16938 , \16933 , \16937 );
and \U$16624 ( \16939 , \10967 , \1826 );
and \U$16625 ( \16940 , \10347 , \1824 );
nor \U$16626 ( \16941 , \16939 , \16940 );
xnor \U$16627 ( \16942 , \16941 , \1670 );
and \U$16628 ( \16943 , \16937 , \16942 );
and \U$16629 ( \16944 , \16933 , \16942 );
or \U$16630 ( \16945 , \16938 , \16943 , \16944 );
xor \U$16631 ( \16946 , \16718 , \16722 );
xor \U$16632 ( \16947 , \16946 , \16727 );
and \U$16633 ( \16948 , \16945 , \16947 );
xor \U$16634 ( \16949 , \16734 , \16736 );
and \U$16635 ( \16950 , \16947 , \16949 );
and \U$16636 ( \16951 , \16945 , \16949 );
or \U$16637 ( \16952 , \16948 , \16950 , \16951 );
and \U$16638 ( \16953 , \16928 , \16952 );
and \U$16639 ( \16954 , \16876 , \16952 );
or \U$16640 ( \16955 , \16929 , \16953 , \16954 );
xor \U$16641 ( \16956 , \16669 , \16673 );
xor \U$16642 ( \16957 , \16956 , \1441 );
xor \U$16643 ( \16958 , \16681 , \16685 );
xor \U$16644 ( \16959 , \16958 , \16690 );
and \U$16645 ( \16960 , \16957 , \16959 );
xor \U$16646 ( \16961 , \16698 , \16702 );
xor \U$16647 ( \16962 , \16961 , \16707 );
and \U$16648 ( \16963 , \16959 , \16962 );
and \U$16649 ( \16964 , \16957 , \16962 );
or \U$16650 ( \16965 , \16960 , \16963 , \16964 );
xor \U$16651 ( \16966 , \16617 , \16621 );
xor \U$16652 ( \16967 , \16966 , \16626 );
xor \U$16653 ( \16968 , \16633 , \16637 );
xor \U$16654 ( \16969 , \16968 , \16642 );
and \U$16655 ( \16970 , \16967 , \16969 );
xor \U$16656 ( \16971 , \16650 , \16654 );
xor \U$16657 ( \16972 , \16971 , \16659 );
and \U$16658 ( \16973 , \16969 , \16972 );
and \U$16659 ( \16974 , \16967 , \16972 );
or \U$16660 ( \16975 , \16970 , \16973 , \16974 );
and \U$16661 ( \16976 , \16965 , \16975 );
xor \U$16662 ( \16977 , \16386 , \16390 );
xor \U$16663 ( \16978 , \16977 , \16395 );
and \U$16664 ( \16979 , \16975 , \16978 );
and \U$16665 ( \16980 , \16965 , \16978 );
or \U$16666 ( \16981 , \16976 , \16979 , \16980 );
and \U$16667 ( \16982 , \16955 , \16981 );
xor \U$16668 ( \16983 , \16730 , \16737 );
xor \U$16669 ( \16984 , \16983 , \16742 );
xor \U$16670 ( \16985 , \16750 , \16752 );
xor \U$16671 ( \16986 , \16985 , \16755 );
and \U$16672 ( \16987 , \16984 , \16986 );
xor \U$16673 ( \16988 , \16760 , \16762 );
xor \U$16674 ( \16989 , \16988 , \16765 );
and \U$16675 ( \16990 , \16986 , \16989 );
and \U$16676 ( \16991 , \16984 , \16989 );
or \U$16677 ( \16992 , \16987 , \16990 , \16991 );
and \U$16678 ( \16993 , \16981 , \16992 );
and \U$16679 ( \16994 , \16955 , \16992 );
or \U$16680 ( \16995 , \16982 , \16993 , \16994 );
xor \U$16681 ( \16996 , \16398 , \16414 );
xor \U$16682 ( \16997 , \16996 , \16431 );
xor \U$16683 ( \16998 , \16758 , \16768 );
xor \U$16684 ( \16999 , \16998 , \16771 );
and \U$16685 ( \17000 , \16997 , \16999 );
xor \U$16686 ( \17001 , \16777 , \16779 );
xor \U$16687 ( \17002 , \17001 , \16782 );
and \U$16688 ( \17003 , \16999 , \17002 );
and \U$16689 ( \17004 , \16997 , \17002 );
or \U$16690 ( \17005 , \17000 , \17003 , \17004 );
and \U$16691 ( \17006 , \16995 , \17005 );
xor \U$16692 ( \17007 , \16434 , \16486 );
xor \U$16693 ( \17008 , \17007 , \16511 );
and \U$16694 ( \17009 , \17005 , \17008 );
and \U$16695 ( \17010 , \16995 , \17008 );
or \U$16696 ( \17011 , \17006 , \17009 , \17010 );
xor \U$16697 ( \17012 , \16748 , \16774 );
xor \U$16698 ( \17013 , \17012 , \16785 );
xor \U$16699 ( \17014 , \16790 , \16792 );
xor \U$16700 ( \17015 , \17014 , \16795 );
and \U$16701 ( \17016 , \17013 , \17015 );
and \U$16702 ( \17017 , \17011 , \17016 );
xor \U$16703 ( \17018 , \16564 , \16566 );
xor \U$16704 ( \17019 , \17018 , \16569 );
and \U$16705 ( \17020 , \17016 , \17019 );
and \U$16706 ( \17021 , \17011 , \17019 );
or \U$16707 ( \17022 , \17017 , \17020 , \17021 );
xor \U$16708 ( \17023 , \16514 , \16540 );
xor \U$16709 ( \17024 , \17023 , \16551 );
xor \U$16710 ( \17025 , \16788 , \16798 );
xor \U$16711 ( \17026 , \17025 , \16801 );
and \U$16712 ( \17027 , \17024 , \17026 );
and \U$16713 ( \17028 , \17022 , \17027 );
xor \U$16714 ( \17029 , \16804 , \16806 );
xor \U$16715 ( \17030 , \17029 , \16809 );
and \U$16716 ( \17031 , \17027 , \17030 );
and \U$16717 ( \17032 , \17022 , \17030 );
or \U$16718 ( \17033 , \17028 , \17031 , \17032 );
and \U$16719 ( \17034 , \16824 , \17033 );
xor \U$16720 ( \17035 , \16824 , \17033 );
xor \U$16721 ( \17036 , \17022 , \17027 );
xor \U$16722 ( \17037 , \17036 , \17030 );
and \U$16723 ( \17038 , \3681 , \7767 );
and \U$16724 ( \17039 , \3264 , \7765 );
nor \U$16725 ( \17040 , \17038 , \17039 );
xnor \U$16726 ( \17041 , \17040 , \7518 );
and \U$16727 ( \17042 , \4011 , \7238 );
and \U$16728 ( \17043 , \3889 , \7236 );
nor \U$16729 ( \17044 , \17042 , \17043 );
xnor \U$16730 ( \17045 , \17044 , \6978 );
and \U$16731 ( \17046 , \17041 , \17045 );
and \U$16732 ( \17047 , \4272 , \6744 );
and \U$16733 ( \17048 , \4016 , \6742 );
nor \U$16734 ( \17049 , \17047 , \17048 );
xnor \U$16735 ( \17050 , \17049 , \6429 );
and \U$16736 ( \17051 , \17045 , \17050 );
and \U$16737 ( \17052 , \17041 , \17050 );
or \U$16738 ( \17053 , \17046 , \17051 , \17052 );
and \U$16739 ( \17054 , \2641 , \9433 );
and \U$16740 ( \17055 , \2377 , \9431 );
nor \U$16741 ( \17056 , \17054 , \17055 );
xnor \U$16742 ( \17057 , \17056 , \9123 );
and \U$16743 ( \17058 , \2840 , \8896 );
and \U$16744 ( \17059 , \2666 , \8894 );
nor \U$16745 ( \17060 , \17058 , \17059 );
xnor \U$16746 ( \17061 , \17060 , \8525 );
and \U$16747 ( \17062 , \17057 , \17061 );
and \U$16748 ( \17063 , \3145 , \8334 );
and \U$16749 ( \17064 , \3007 , \8332 );
nor \U$16750 ( \17065 , \17063 , \17064 );
xnor \U$16751 ( \17066 , \17065 , \8016 );
and \U$16752 ( \17067 , \17061 , \17066 );
and \U$16753 ( \17068 , \17057 , \17066 );
or \U$16754 ( \17069 , \17062 , \17067 , \17068 );
and \U$16755 ( \17070 , \17053 , \17069 );
and \U$16756 ( \17071 , \2042 , \10814 );
and \U$16757 ( \17072 , \1799 , \10811 );
nor \U$16758 ( \17073 , \17071 , \17072 );
xnor \U$16759 ( \17074 , \17073 , \9759 );
and \U$16760 ( \17075 , \2233 , \10001 );
and \U$16761 ( \17076 , \2047 , \9999 );
nor \U$16762 ( \17077 , \17075 , \17076 );
xnor \U$16763 ( \17078 , \17077 , \9762 );
and \U$16764 ( \17079 , \17074 , \17078 );
and \U$16765 ( \17080 , \17078 , \1670 );
and \U$16766 ( \17081 , \17074 , \1670 );
or \U$16767 ( \17082 , \17079 , \17080 , \17081 );
and \U$16768 ( \17083 , \17069 , \17082 );
and \U$16769 ( \17084 , \17053 , \17082 );
or \U$16770 ( \17085 , \17070 , \17083 , \17084 );
and \U$16771 ( \17086 , \7703 , \3637 );
and \U$16772 ( \17087 , \7177 , \3635 );
nor \U$16773 ( \17088 , \17086 , \17087 );
xnor \U$16774 ( \17089 , \17088 , \3450 );
and \U$16775 ( \17090 , \8373 , \3324 );
and \U$16776 ( \17091 , \8127 , \3322 );
nor \U$16777 ( \17092 , \17090 , \17091 );
xnor \U$16778 ( \17093 , \17092 , \3119 );
and \U$16779 ( \17094 , \17089 , \17093 );
and \U$16780 ( \17095 , \8697 , \2918 );
and \U$16781 ( \17096 , \8378 , \2916 );
nor \U$16782 ( \17097 , \17095 , \17096 );
xnor \U$16783 ( \17098 , \17097 , \2769 );
and \U$16784 ( \17099 , \17093 , \17098 );
and \U$16785 ( \17100 , \17089 , \17098 );
or \U$16786 ( \17101 , \17094 , \17099 , \17100 );
and \U$16787 ( \17102 , \4771 , \6235 );
and \U$16788 ( \17103 , \4469 , \6233 );
nor \U$16789 ( \17104 , \17102 , \17103 );
xnor \U$16790 ( \17105 , \17104 , \5895 );
and \U$16791 ( \17106 , \5248 , \5646 );
and \U$16792 ( \17107 , \4779 , \5644 );
nor \U$16793 ( \17108 , \17106 , \17107 );
xnor \U$16794 ( \17109 , \17108 , \5405 );
and \U$16795 ( \17110 , \17105 , \17109 );
and \U$16796 ( \17111 , \5517 , \5180 );
and \U$16797 ( \17112 , \5253 , \5178 );
nor \U$16798 ( \17113 , \17111 , \17112 );
xnor \U$16799 ( \17114 , \17113 , \4992 );
and \U$16800 ( \17115 , \17109 , \17114 );
and \U$16801 ( \17116 , \17105 , \17114 );
or \U$16802 ( \17117 , \17110 , \17115 , \17116 );
and \U$16803 ( \17118 , \17101 , \17117 );
and \U$16804 ( \17119 , \6148 , \4806 );
and \U$16805 ( \17120 , \5776 , \4804 );
nor \U$16806 ( \17121 , \17119 , \17120 );
xnor \U$16807 ( \17122 , \17121 , \4574 );
and \U$16808 ( \17123 , \6500 , \4355 );
and \U$16809 ( \17124 , \6157 , \4353 );
nor \U$16810 ( \17125 , \17123 , \17124 );
xnor \U$16811 ( \17126 , \17125 , \4212 );
and \U$16812 ( \17127 , \17122 , \17126 );
and \U$16813 ( \17128 , \7005 , \4032 );
and \U$16814 ( \17129 , \6702 , \4030 );
nor \U$16815 ( \17130 , \17128 , \17129 );
xnor \U$16816 ( \17131 , \17130 , \3786 );
and \U$16817 ( \17132 , \17126 , \17131 );
and \U$16818 ( \17133 , \17122 , \17131 );
or \U$16819 ( \17134 , \17127 , \17132 , \17133 );
and \U$16820 ( \17135 , \17117 , \17134 );
and \U$16821 ( \17136 , \17101 , \17134 );
or \U$16822 ( \17137 , \17118 , \17135 , \17136 );
and \U$16823 ( \17138 , \17085 , \17137 );
and \U$16824 ( \17139 , \9550 , \2596 );
and \U$16825 ( \17140 , \8981 , \2594 );
nor \U$16826 ( \17141 , \17139 , \17140 );
xnor \U$16827 ( \17142 , \17141 , \2454 );
and \U$16828 ( \17143 , \10161 , \2300 );
and \U$16829 ( \17144 , \9558 , \2298 );
nor \U$16830 ( \17145 , \17143 , \17144 );
xnor \U$16831 ( \17146 , \17145 , \2163 );
and \U$16832 ( \17147 , \17142 , \17146 );
and \U$16833 ( \17148 , \10347 , \2094 );
and \U$16834 ( \17149 , \10166 , \2092 );
nor \U$16835 ( \17150 , \17148 , \17149 );
xnor \U$16836 ( \17151 , \17150 , \1942 );
and \U$16837 ( \17152 , \17146 , \17151 );
and \U$16838 ( \17153 , \17142 , \17151 );
or \U$16839 ( \17154 , \17147 , \17152 , \17153 );
xor \U$16840 ( \17155 , \16844 , \16848 );
xor \U$16841 ( \17156 , \17155 , \16853 );
and \U$16842 ( \17157 , \17154 , \17156 );
xor \U$16843 ( \17158 , \16933 , \16937 );
xor \U$16844 ( \17159 , \17158 , \16942 );
and \U$16845 ( \17160 , \17156 , \17159 );
and \U$16846 ( \17161 , \17154 , \17159 );
or \U$16847 ( \17162 , \17157 , \17160 , \17161 );
and \U$16848 ( \17163 , \17137 , \17162 );
and \U$16849 ( \17164 , \17085 , \17162 );
or \U$16850 ( \17165 , \17138 , \17163 , \17164 );
xor \U$16851 ( \17166 , \16828 , \16832 );
xor \U$16852 ( \17167 , \17166 , \16837 );
xor \U$16853 ( \17168 , \16880 , \16884 );
xor \U$16854 ( \17169 , \17168 , \16889 );
and \U$16855 ( \17170 , \17167 , \17169 );
xor \U$16856 ( \17171 , \16861 , \16865 );
xor \U$16857 ( \17172 , \17171 , \16870 );
and \U$16858 ( \17173 , \17169 , \17172 );
and \U$16859 ( \17174 , \17167 , \17172 );
or \U$16860 ( \17175 , \17170 , \17173 , \17174 );
xor \U$16861 ( \17176 , \16896 , \16900 );
xor \U$16862 ( \17177 , \17176 , \16905 );
xor \U$16863 ( \17178 , \16913 , \16917 );
xor \U$16864 ( \17179 , \17178 , \16922 );
and \U$16865 ( \17180 , \17177 , \17179 );
and \U$16866 ( \17181 , \17175 , \17180 );
xor \U$16867 ( \17182 , \16957 , \16959 );
xor \U$16868 ( \17183 , \17182 , \16962 );
and \U$16869 ( \17184 , \17180 , \17183 );
and \U$16870 ( \17185 , \17175 , \17183 );
or \U$16871 ( \17186 , \17181 , \17184 , \17185 );
and \U$16872 ( \17187 , \17165 , \17186 );
xor \U$16873 ( \17188 , \16840 , \16856 );
xor \U$16874 ( \17189 , \17188 , \16873 );
xor \U$16875 ( \17190 , \16967 , \16969 );
xor \U$16876 ( \17191 , \17190 , \16972 );
and \U$16877 ( \17192 , \17189 , \17191 );
xor \U$16878 ( \17193 , \16945 , \16947 );
xor \U$16879 ( \17194 , \17193 , \16949 );
and \U$16880 ( \17195 , \17191 , \17194 );
and \U$16881 ( \17196 , \17189 , \17194 );
or \U$16882 ( \17197 , \17192 , \17195 , \17196 );
and \U$16883 ( \17198 , \17186 , \17197 );
and \U$16884 ( \17199 , \17165 , \17197 );
or \U$16885 ( \17200 , \17187 , \17198 , \17199 );
xor \U$16886 ( \17201 , \16629 , \16645 );
xor \U$16887 ( \17202 , \17201 , \16662 );
xor \U$16888 ( \17203 , \16677 , \16693 );
xor \U$16889 ( \17204 , \17203 , \16710 );
and \U$16890 ( \17205 , \17202 , \17204 );
xor \U$16891 ( \17206 , \16984 , \16986 );
xor \U$16892 ( \17207 , \17206 , \16989 );
and \U$16893 ( \17208 , \17204 , \17207 );
and \U$16894 ( \17209 , \17202 , \17207 );
or \U$16895 ( \17210 , \17205 , \17208 , \17209 );
and \U$16896 ( \17211 , \17200 , \17210 );
xor \U$16897 ( \17212 , \16665 , \16713 );
xor \U$16898 ( \17213 , \17212 , \16745 );
and \U$16899 ( \17214 , \17210 , \17213 );
and \U$16900 ( \17215 , \17200 , \17213 );
or \U$16901 ( \17216 , \17211 , \17214 , \17215 );
xor \U$16902 ( \17217 , \16995 , \17005 );
xor \U$16903 ( \17218 , \17217 , \17008 );
and \U$16904 ( \17219 , \17216 , \17218 );
xor \U$16905 ( \17220 , \17013 , \17015 );
and \U$16906 ( \17221 , \17218 , \17220 );
and \U$16907 ( \17222 , \17216 , \17220 );
or \U$16908 ( \17223 , \17219 , \17221 , \17222 );
xor \U$16909 ( \17224 , \17011 , \17016 );
xor \U$16910 ( \17225 , \17224 , \17019 );
and \U$16911 ( \17226 , \17223 , \17225 );
xor \U$16912 ( \17227 , \17024 , \17026 );
and \U$16913 ( \17228 , \17225 , \17227 );
and \U$16914 ( \17229 , \17223 , \17227 );
or \U$16915 ( \17230 , \17226 , \17228 , \17229 );
and \U$16916 ( \17231 , \17037 , \17230 );
xor \U$16917 ( \17232 , \17037 , \17230 );
xor \U$16918 ( \17233 , \17223 , \17225 );
xor \U$16919 ( \17234 , \17233 , \17227 );
and \U$16920 ( \17235 , \2047 , \10814 );
and \U$16921 ( \17236 , \2042 , \10811 );
nor \U$16922 ( \17237 , \17235 , \17236 );
xnor \U$16923 ( \17238 , \17237 , \9759 );
and \U$16924 ( \17239 , \2377 , \10001 );
and \U$16925 ( \17240 , \2233 , \9999 );
nor \U$16926 ( \17241 , \17239 , \17240 );
xnor \U$16927 ( \17242 , \17241 , \9762 );
and \U$16928 ( \17243 , \17238 , \17242 );
and \U$16929 ( \17244 , \2666 , \9433 );
and \U$16930 ( \17245 , \2641 , \9431 );
nor \U$16931 ( \17246 , \17244 , \17245 );
xnor \U$16932 ( \17247 , \17246 , \9123 );
and \U$16933 ( \17248 , \17242 , \17247 );
and \U$16934 ( \17249 , \17238 , \17247 );
or \U$16935 ( \17250 , \17243 , \17248 , \17249 );
and \U$16936 ( \17251 , \3007 , \8896 );
and \U$16937 ( \17252 , \2840 , \8894 );
nor \U$16938 ( \17253 , \17251 , \17252 );
xnor \U$16939 ( \17254 , \17253 , \8525 );
and \U$16940 ( \17255 , \3264 , \8334 );
and \U$16941 ( \17256 , \3145 , \8332 );
nor \U$16942 ( \17257 , \17255 , \17256 );
xnor \U$16943 ( \17258 , \17257 , \8016 );
and \U$16944 ( \17259 , \17254 , \17258 );
and \U$16945 ( \17260 , \3889 , \7767 );
and \U$16946 ( \17261 , \3681 , \7765 );
nor \U$16947 ( \17262 , \17260 , \17261 );
xnor \U$16948 ( \17263 , \17262 , \7518 );
and \U$16949 ( \17264 , \17258 , \17263 );
and \U$16950 ( \17265 , \17254 , \17263 );
or \U$16951 ( \17266 , \17259 , \17264 , \17265 );
and \U$16952 ( \17267 , \17250 , \17266 );
and \U$16953 ( \17268 , \4016 , \7238 );
and \U$16954 ( \17269 , \4011 , \7236 );
nor \U$16955 ( \17270 , \17268 , \17269 );
xnor \U$16956 ( \17271 , \17270 , \6978 );
and \U$16957 ( \17272 , \4469 , \6744 );
and \U$16958 ( \17273 , \4272 , \6742 );
nor \U$16959 ( \17274 , \17272 , \17273 );
xnor \U$16960 ( \17275 , \17274 , \6429 );
and \U$16961 ( \17276 , \17271 , \17275 );
and \U$16962 ( \17277 , \4779 , \6235 );
and \U$16963 ( \17278 , \4771 , \6233 );
nor \U$16964 ( \17279 , \17277 , \17278 );
xnor \U$16965 ( \17280 , \17279 , \5895 );
and \U$16966 ( \17281 , \17275 , \17280 );
and \U$16967 ( \17282 , \17271 , \17280 );
or \U$16968 ( \17283 , \17276 , \17281 , \17282 );
and \U$16969 ( \17284 , \17266 , \17283 );
and \U$16970 ( \17285 , \17250 , \17283 );
or \U$16971 ( \17286 , \17267 , \17284 , \17285 );
and \U$16972 ( \17287 , \6702 , \4355 );
and \U$16973 ( \17288 , \6500 , \4353 );
nor \U$16974 ( \17289 , \17287 , \17288 );
xnor \U$16975 ( \17290 , \17289 , \4212 );
and \U$16976 ( \17291 , \7177 , \4032 );
and \U$16977 ( \17292 , \7005 , \4030 );
nor \U$16978 ( \17293 , \17291 , \17292 );
xnor \U$16979 ( \17294 , \17293 , \3786 );
and \U$16980 ( \17295 , \17290 , \17294 );
and \U$16981 ( \17296 , \8127 , \3637 );
and \U$16982 ( \17297 , \7703 , \3635 );
nor \U$16983 ( \17298 , \17296 , \17297 );
xnor \U$16984 ( \17299 , \17298 , \3450 );
and \U$16985 ( \17300 , \17294 , \17299 );
and \U$16986 ( \17301 , \17290 , \17299 );
or \U$16987 ( \17302 , \17295 , \17300 , \17301 );
and \U$16988 ( \17303 , \5253 , \5646 );
and \U$16989 ( \17304 , \5248 , \5644 );
nor \U$16990 ( \17305 , \17303 , \17304 );
xnor \U$16991 ( \17306 , \17305 , \5405 );
and \U$16992 ( \17307 , \5776 , \5180 );
and \U$16993 ( \17308 , \5517 , \5178 );
nor \U$16994 ( \17309 , \17307 , \17308 );
xnor \U$16995 ( \17310 , \17309 , \4992 );
and \U$16996 ( \17311 , \17306 , \17310 );
and \U$16997 ( \17312 , \6157 , \4806 );
and \U$16998 ( \17313 , \6148 , \4804 );
nor \U$16999 ( \17314 , \17312 , \17313 );
xnor \U$17000 ( \17315 , \17314 , \4574 );
and \U$17001 ( \17316 , \17310 , \17315 );
and \U$17002 ( \17317 , \17306 , \17315 );
or \U$17003 ( \17318 , \17311 , \17316 , \17317 );
and \U$17004 ( \17319 , \17302 , \17318 );
and \U$17005 ( \17320 , \8378 , \3324 );
and \U$17006 ( \17321 , \8373 , \3322 );
nor \U$17007 ( \17322 , \17320 , \17321 );
xnor \U$17008 ( \17323 , \17322 , \3119 );
and \U$17009 ( \17324 , \8981 , \2918 );
and \U$17010 ( \17325 , \8697 , \2916 );
nor \U$17011 ( \17326 , \17324 , \17325 );
xnor \U$17012 ( \17327 , \17326 , \2769 );
and \U$17013 ( \17328 , \17323 , \17327 );
and \U$17014 ( \17329 , \9558 , \2596 );
and \U$17015 ( \17330 , \9550 , \2594 );
nor \U$17016 ( \17331 , \17329 , \17330 );
xnor \U$17017 ( \17332 , \17331 , \2454 );
and \U$17018 ( \17333 , \17327 , \17332 );
and \U$17019 ( \17334 , \17323 , \17332 );
or \U$17020 ( \17335 , \17328 , \17333 , \17334 );
and \U$17021 ( \17336 , \17318 , \17335 );
and \U$17022 ( \17337 , \17302 , \17335 );
or \U$17023 ( \17338 , \17319 , \17336 , \17337 );
and \U$17024 ( \17339 , \17286 , \17338 );
nand \U$17025 ( \17340 , \10967 , \1824 );
xnor \U$17026 ( \17341 , \17340 , \1670 );
xor \U$17027 ( \17342 , \17089 , \17093 );
xor \U$17028 ( \17343 , \17342 , \17098 );
and \U$17029 ( \17344 , \17341 , \17343 );
xor \U$17030 ( \17345 , \17142 , \17146 );
xor \U$17031 ( \17346 , \17345 , \17151 );
and \U$17032 ( \17347 , \17343 , \17346 );
and \U$17033 ( \17348 , \17341 , \17346 );
or \U$17034 ( \17349 , \17344 , \17347 , \17348 );
and \U$17035 ( \17350 , \17338 , \17349 );
and \U$17036 ( \17351 , \17286 , \17349 );
or \U$17037 ( \17352 , \17339 , \17350 , \17351 );
xor \U$17038 ( \17353 , \17053 , \17069 );
xor \U$17039 ( \17354 , \17353 , \17082 );
xor \U$17040 ( \17355 , \17101 , \17117 );
xor \U$17041 ( \17356 , \17355 , \17134 );
and \U$17042 ( \17357 , \17354 , \17356 );
xor \U$17043 ( \17358 , \17154 , \17156 );
xor \U$17044 ( \17359 , \17358 , \17159 );
and \U$17045 ( \17360 , \17356 , \17359 );
and \U$17046 ( \17361 , \17354 , \17359 );
or \U$17047 ( \17362 , \17357 , \17360 , \17361 );
and \U$17048 ( \17363 , \17352 , \17362 );
xor \U$17049 ( \17364 , \17041 , \17045 );
xor \U$17050 ( \17365 , \17364 , \17050 );
xor \U$17051 ( \17366 , \17105 , \17109 );
xor \U$17052 ( \17367 , \17366 , \17114 );
and \U$17053 ( \17368 , \17365 , \17367 );
xor \U$17054 ( \17369 , \17122 , \17126 );
xor \U$17055 ( \17370 , \17369 , \17131 );
and \U$17056 ( \17371 , \17367 , \17370 );
and \U$17057 ( \17372 , \17365 , \17370 );
or \U$17058 ( \17373 , \17368 , \17371 , \17372 );
xor \U$17059 ( \17374 , \17167 , \17169 );
xor \U$17060 ( \17375 , \17374 , \17172 );
and \U$17061 ( \17376 , \17373 , \17375 );
xor \U$17062 ( \17377 , \17177 , \17179 );
and \U$17063 ( \17378 , \17375 , \17377 );
and \U$17064 ( \17379 , \17373 , \17377 );
or \U$17065 ( \17380 , \17376 , \17378 , \17379 );
and \U$17066 ( \17381 , \17362 , \17380 );
and \U$17067 ( \17382 , \17352 , \17380 );
or \U$17068 ( \17383 , \17363 , \17381 , \17382 );
xor \U$17069 ( \17384 , \16892 , \16908 );
xor \U$17070 ( \17385 , \17384 , \16925 );
xor \U$17071 ( \17386 , \17175 , \17180 );
xor \U$17072 ( \17387 , \17386 , \17183 );
and \U$17073 ( \17388 , \17385 , \17387 );
xor \U$17074 ( \17389 , \17189 , \17191 );
xor \U$17075 ( \17390 , \17389 , \17194 );
and \U$17076 ( \17391 , \17387 , \17390 );
and \U$17077 ( \17392 , \17385 , \17390 );
or \U$17078 ( \17393 , \17388 , \17391 , \17392 );
and \U$17079 ( \17394 , \17383 , \17393 );
xor \U$17080 ( \17395 , \16965 , \16975 );
xor \U$17081 ( \17396 , \17395 , \16978 );
and \U$17082 ( \17397 , \17393 , \17396 );
and \U$17083 ( \17398 , \17383 , \17396 );
or \U$17084 ( \17399 , \17394 , \17397 , \17398 );
xor \U$17085 ( \17400 , \16876 , \16928 );
xor \U$17086 ( \17401 , \17400 , \16952 );
xor \U$17087 ( \17402 , \17165 , \17186 );
xor \U$17088 ( \17403 , \17402 , \17197 );
and \U$17089 ( \17404 , \17401 , \17403 );
xor \U$17090 ( \17405 , \17202 , \17204 );
xor \U$17091 ( \17406 , \17405 , \17207 );
and \U$17092 ( \17407 , \17403 , \17406 );
and \U$17093 ( \17408 , \17401 , \17406 );
or \U$17094 ( \17409 , \17404 , \17407 , \17408 );
and \U$17095 ( \17410 , \17399 , \17409 );
xor \U$17096 ( \17411 , \16997 , \16999 );
xor \U$17097 ( \17412 , \17411 , \17002 );
and \U$17098 ( \17413 , \17409 , \17412 );
and \U$17099 ( \17414 , \17399 , \17412 );
or \U$17100 ( \17415 , \17410 , \17413 , \17414 );
xor \U$17101 ( \17416 , \16955 , \16981 );
xor \U$17102 ( \17417 , \17416 , \16992 );
xor \U$17103 ( \17418 , \17200 , \17210 );
xor \U$17104 ( \17419 , \17418 , \17213 );
and \U$17105 ( \17420 , \17417 , \17419 );
and \U$17106 ( \17421 , \17415 , \17420 );
xor \U$17107 ( \17422 , \17216 , \17218 );
xor \U$17108 ( \17423 , \17422 , \17220 );
and \U$17109 ( \17424 , \17420 , \17423 );
and \U$17110 ( \17425 , \17415 , \17423 );
or \U$17111 ( \17426 , \17421 , \17424 , \17425 );
and \U$17112 ( \17427 , \17234 , \17426 );
xor \U$17113 ( \17428 , \17234 , \17426 );
xor \U$17114 ( \17429 , \17415 , \17420 );
xor \U$17115 ( \17430 , \17429 , \17423 );
and \U$17116 ( \17431 , \2233 , \10814 );
and \U$17117 ( \17432 , \2047 , \10811 );
nor \U$17118 ( \17433 , \17431 , \17432 );
xnor \U$17119 ( \17434 , \17433 , \9759 );
and \U$17120 ( \17435 , \2641 , \10001 );
and \U$17121 ( \17436 , \2377 , \9999 );
nor \U$17122 ( \17437 , \17435 , \17436 );
xnor \U$17123 ( \17438 , \17437 , \9762 );
and \U$17124 ( \17439 , \17434 , \17438 );
and \U$17125 ( \17440 , \17438 , \1942 );
and \U$17126 ( \17441 , \17434 , \1942 );
or \U$17127 ( \17442 , \17439 , \17440 , \17441 );
and \U$17128 ( \17443 , \4011 , \7767 );
and \U$17129 ( \17444 , \3889 , \7765 );
nor \U$17130 ( \17445 , \17443 , \17444 );
xnor \U$17131 ( \17446 , \17445 , \7518 );
and \U$17132 ( \17447 , \4272 , \7238 );
and \U$17133 ( \17448 , \4016 , \7236 );
nor \U$17134 ( \17449 , \17447 , \17448 );
xnor \U$17135 ( \17450 , \17449 , \6978 );
and \U$17136 ( \17451 , \17446 , \17450 );
and \U$17137 ( \17452 , \4771 , \6744 );
and \U$17138 ( \17453 , \4469 , \6742 );
nor \U$17139 ( \17454 , \17452 , \17453 );
xnor \U$17140 ( \17455 , \17454 , \6429 );
and \U$17141 ( \17456 , \17450 , \17455 );
and \U$17142 ( \17457 , \17446 , \17455 );
or \U$17143 ( \17458 , \17451 , \17456 , \17457 );
and \U$17144 ( \17459 , \17442 , \17458 );
and \U$17145 ( \17460 , \2840 , \9433 );
and \U$17146 ( \17461 , \2666 , \9431 );
nor \U$17147 ( \17462 , \17460 , \17461 );
xnor \U$17148 ( \17463 , \17462 , \9123 );
and \U$17149 ( \17464 , \3145 , \8896 );
and \U$17150 ( \17465 , \3007 , \8894 );
nor \U$17151 ( \17466 , \17464 , \17465 );
xnor \U$17152 ( \17467 , \17466 , \8525 );
and \U$17153 ( \17468 , \17463 , \17467 );
and \U$17154 ( \17469 , \3681 , \8334 );
and \U$17155 ( \17470 , \3264 , \8332 );
nor \U$17156 ( \17471 , \17469 , \17470 );
xnor \U$17157 ( \17472 , \17471 , \8016 );
and \U$17158 ( \17473 , \17467 , \17472 );
and \U$17159 ( \17474 , \17463 , \17472 );
or \U$17160 ( \17475 , \17468 , \17473 , \17474 );
and \U$17161 ( \17476 , \17458 , \17475 );
and \U$17162 ( \17477 , \17442 , \17475 );
or \U$17163 ( \17478 , \17459 , \17476 , \17477 );
and \U$17164 ( \17479 , \10161 , \2596 );
and \U$17165 ( \17480 , \9558 , \2594 );
nor \U$17166 ( \17481 , \17479 , \17480 );
xnor \U$17167 ( \17482 , \17481 , \2454 );
and \U$17168 ( \17483 , \10347 , \2300 );
and \U$17169 ( \17484 , \10166 , \2298 );
nor \U$17170 ( \17485 , \17483 , \17484 );
xnor \U$17171 ( \17486 , \17485 , \2163 );
and \U$17172 ( \17487 , \17482 , \17486 );
nand \U$17173 ( \17488 , \10967 , \2092 );
xnor \U$17174 ( \17489 , \17488 , \1942 );
and \U$17175 ( \17490 , \17486 , \17489 );
and \U$17176 ( \17491 , \17482 , \17489 );
or \U$17177 ( \17492 , \17487 , \17490 , \17491 );
and \U$17178 ( \17493 , \10166 , \2300 );
and \U$17179 ( \17494 , \10161 , \2298 );
nor \U$17180 ( \17495 , \17493 , \17494 );
xnor \U$17181 ( \17496 , \17495 , \2163 );
and \U$17182 ( \17497 , \17492 , \17496 );
and \U$17183 ( \17498 , \10967 , \2094 );
and \U$17184 ( \17499 , \10347 , \2092 );
nor \U$17185 ( \17500 , \17498 , \17499 );
xnor \U$17186 ( \17501 , \17500 , \1942 );
and \U$17187 ( \17502 , \17496 , \17501 );
and \U$17188 ( \17503 , \17492 , \17501 );
or \U$17189 ( \17504 , \17497 , \17502 , \17503 );
and \U$17190 ( \17505 , \17478 , \17504 );
and \U$17191 ( \17506 , \5248 , \6235 );
and \U$17192 ( \17507 , \4779 , \6233 );
nor \U$17193 ( \17508 , \17506 , \17507 );
xnor \U$17194 ( \17509 , \17508 , \5895 );
and \U$17195 ( \17510 , \5517 , \5646 );
and \U$17196 ( \17511 , \5253 , \5644 );
nor \U$17197 ( \17512 , \17510 , \17511 );
xnor \U$17198 ( \17513 , \17512 , \5405 );
and \U$17199 ( \17514 , \17509 , \17513 );
and \U$17200 ( \17515 , \6148 , \5180 );
and \U$17201 ( \17516 , \5776 , \5178 );
nor \U$17202 ( \17517 , \17515 , \17516 );
xnor \U$17203 ( \17518 , \17517 , \4992 );
and \U$17204 ( \17519 , \17513 , \17518 );
and \U$17205 ( \17520 , \17509 , \17518 );
or \U$17206 ( \17521 , \17514 , \17519 , \17520 );
and \U$17207 ( \17522 , \8373 , \3637 );
and \U$17208 ( \17523 , \8127 , \3635 );
nor \U$17209 ( \17524 , \17522 , \17523 );
xnor \U$17210 ( \17525 , \17524 , \3450 );
and \U$17211 ( \17526 , \8697 , \3324 );
and \U$17212 ( \17527 , \8378 , \3322 );
nor \U$17213 ( \17528 , \17526 , \17527 );
xnor \U$17214 ( \17529 , \17528 , \3119 );
and \U$17215 ( \17530 , \17525 , \17529 );
and \U$17216 ( \17531 , \9550 , \2918 );
and \U$17217 ( \17532 , \8981 , \2916 );
nor \U$17218 ( \17533 , \17531 , \17532 );
xnor \U$17219 ( \17534 , \17533 , \2769 );
and \U$17220 ( \17535 , \17529 , \17534 );
and \U$17221 ( \17536 , \17525 , \17534 );
or \U$17222 ( \17537 , \17530 , \17535 , \17536 );
and \U$17223 ( \17538 , \17521 , \17537 );
and \U$17224 ( \17539 , \6500 , \4806 );
and \U$17225 ( \17540 , \6157 , \4804 );
nor \U$17226 ( \17541 , \17539 , \17540 );
xnor \U$17227 ( \17542 , \17541 , \4574 );
and \U$17228 ( \17543 , \7005 , \4355 );
and \U$17229 ( \17544 , \6702 , \4353 );
nor \U$17230 ( \17545 , \17543 , \17544 );
xnor \U$17231 ( \17546 , \17545 , \4212 );
and \U$17232 ( \17547 , \17542 , \17546 );
and \U$17233 ( \17548 , \7703 , \4032 );
and \U$17234 ( \17549 , \7177 , \4030 );
nor \U$17235 ( \17550 , \17548 , \17549 );
xnor \U$17236 ( \17551 , \17550 , \3786 );
and \U$17237 ( \17552 , \17546 , \17551 );
and \U$17238 ( \17553 , \17542 , \17551 );
or \U$17239 ( \17554 , \17547 , \17552 , \17553 );
and \U$17240 ( \17555 , \17537 , \17554 );
and \U$17241 ( \17556 , \17521 , \17554 );
or \U$17242 ( \17557 , \17538 , \17555 , \17556 );
and \U$17243 ( \17558 , \17504 , \17557 );
and \U$17244 ( \17559 , \17478 , \17557 );
or \U$17245 ( \17560 , \17505 , \17558 , \17559 );
xor \U$17246 ( \17561 , \17238 , \17242 );
xor \U$17247 ( \17562 , \17561 , \17247 );
xor \U$17248 ( \17563 , \17254 , \17258 );
xor \U$17249 ( \17564 , \17563 , \17263 );
and \U$17250 ( \17565 , \17562 , \17564 );
xor \U$17251 ( \17566 , \17271 , \17275 );
xor \U$17252 ( \17567 , \17566 , \17280 );
and \U$17253 ( \17568 , \17564 , \17567 );
and \U$17254 ( \17569 , \17562 , \17567 );
or \U$17255 ( \17570 , \17565 , \17568 , \17569 );
xor \U$17256 ( \17571 , \17290 , \17294 );
xor \U$17257 ( \17572 , \17571 , \17299 );
xor \U$17258 ( \17573 , \17306 , \17310 );
xor \U$17259 ( \17574 , \17573 , \17315 );
and \U$17260 ( \17575 , \17572 , \17574 );
xor \U$17261 ( \17576 , \17323 , \17327 );
xor \U$17262 ( \17577 , \17576 , \17332 );
and \U$17263 ( \17578 , \17574 , \17577 );
and \U$17264 ( \17579 , \17572 , \17577 );
or \U$17265 ( \17580 , \17575 , \17578 , \17579 );
and \U$17266 ( \17581 , \17570 , \17580 );
xor \U$17267 ( \17582 , \17057 , \17061 );
xor \U$17268 ( \17583 , \17582 , \17066 );
and \U$17269 ( \17584 , \17580 , \17583 );
and \U$17270 ( \17585 , \17570 , \17583 );
or \U$17271 ( \17586 , \17581 , \17584 , \17585 );
and \U$17272 ( \17587 , \17560 , \17586 );
xor \U$17273 ( \17588 , \17074 , \17078 );
xor \U$17274 ( \17589 , \17588 , \1670 );
xor \U$17275 ( \17590 , \17365 , \17367 );
xor \U$17276 ( \17591 , \17590 , \17370 );
and \U$17277 ( \17592 , \17589 , \17591 );
xor \U$17278 ( \17593 , \17341 , \17343 );
xor \U$17279 ( \17594 , \17593 , \17346 );
and \U$17280 ( \17595 , \17591 , \17594 );
and \U$17281 ( \17596 , \17589 , \17594 );
or \U$17282 ( \17597 , \17592 , \17595 , \17596 );
and \U$17283 ( \17598 , \17586 , \17597 );
and \U$17284 ( \17599 , \17560 , \17597 );
or \U$17285 ( \17600 , \17587 , \17598 , \17599 );
xor \U$17286 ( \17601 , \17286 , \17338 );
xor \U$17287 ( \17602 , \17601 , \17349 );
xor \U$17288 ( \17603 , \17354 , \17356 );
xor \U$17289 ( \17604 , \17603 , \17359 );
and \U$17290 ( \17605 , \17602 , \17604 );
xor \U$17291 ( \17606 , \17373 , \17375 );
xor \U$17292 ( \17607 , \17606 , \17377 );
and \U$17293 ( \17608 , \17604 , \17607 );
and \U$17294 ( \17609 , \17602 , \17607 );
or \U$17295 ( \17610 , \17605 , \17608 , \17609 );
and \U$17296 ( \17611 , \17600 , \17610 );
xor \U$17297 ( \17612 , \17085 , \17137 );
xor \U$17298 ( \17613 , \17612 , \17162 );
and \U$17299 ( \17614 , \17610 , \17613 );
and \U$17300 ( \17615 , \17600 , \17613 );
or \U$17301 ( \17616 , \17611 , \17614 , \17615 );
xor \U$17302 ( \17617 , \17352 , \17362 );
xor \U$17303 ( \17618 , \17617 , \17380 );
xor \U$17304 ( \17619 , \17385 , \17387 );
xor \U$17305 ( \17620 , \17619 , \17390 );
and \U$17306 ( \17621 , \17618 , \17620 );
and \U$17307 ( \17622 , \17616 , \17621 );
xor \U$17308 ( \17623 , \17401 , \17403 );
xor \U$17309 ( \17624 , \17623 , \17406 );
and \U$17310 ( \17625 , \17621 , \17624 );
and \U$17311 ( \17626 , \17616 , \17624 );
or \U$17312 ( \17627 , \17622 , \17625 , \17626 );
xor \U$17313 ( \17628 , \17399 , \17409 );
xor \U$17314 ( \17629 , \17628 , \17412 );
and \U$17315 ( \17630 , \17627 , \17629 );
xor \U$17316 ( \17631 , \17417 , \17419 );
and \U$17317 ( \17632 , \17629 , \17631 );
and \U$17318 ( \17633 , \17627 , \17631 );
or \U$17319 ( \17634 , \17630 , \17632 , \17633 );
and \U$17320 ( \17635 , \17430 , \17634 );
xor \U$17321 ( \17636 , \17430 , \17634 );
xor \U$17322 ( \17637 , \17627 , \17629 );
xor \U$17323 ( \17638 , \17637 , \17631 );
and \U$17324 ( \17639 , \8981 , \3324 );
and \U$17325 ( \17640 , \8697 , \3322 );
nor \U$17326 ( \17641 , \17639 , \17640 );
xnor \U$17327 ( \17642 , \17641 , \3119 );
and \U$17328 ( \17643 , \9558 , \2918 );
and \U$17329 ( \17644 , \9550 , \2916 );
nor \U$17330 ( \17645 , \17643 , \17644 );
xnor \U$17331 ( \17646 , \17645 , \2769 );
and \U$17332 ( \17647 , \17642 , \17646 );
and \U$17333 ( \17648 , \10166 , \2596 );
and \U$17334 ( \17649 , \10161 , \2594 );
nor \U$17335 ( \17650 , \17648 , \17649 );
xnor \U$17336 ( \17651 , \17650 , \2454 );
and \U$17337 ( \17652 , \17646 , \17651 );
and \U$17338 ( \17653 , \17642 , \17651 );
or \U$17339 ( \17654 , \17647 , \17652 , \17653 );
and \U$17340 ( \17655 , \5776 , \5646 );
and \U$17341 ( \17656 , \5517 , \5644 );
nor \U$17342 ( \17657 , \17655 , \17656 );
xnor \U$17343 ( \17658 , \17657 , \5405 );
and \U$17344 ( \17659 , \6157 , \5180 );
and \U$17345 ( \17660 , \6148 , \5178 );
nor \U$17346 ( \17661 , \17659 , \17660 );
xnor \U$17347 ( \17662 , \17661 , \4992 );
and \U$17348 ( \17663 , \17658 , \17662 );
and \U$17349 ( \17664 , \6702 , \4806 );
and \U$17350 ( \17665 , \6500 , \4804 );
nor \U$17351 ( \17666 , \17664 , \17665 );
xnor \U$17352 ( \17667 , \17666 , \4574 );
and \U$17353 ( \17668 , \17662 , \17667 );
and \U$17354 ( \17669 , \17658 , \17667 );
or \U$17355 ( \17670 , \17663 , \17668 , \17669 );
and \U$17356 ( \17671 , \17654 , \17670 );
and \U$17357 ( \17672 , \7177 , \4355 );
and \U$17358 ( \17673 , \7005 , \4353 );
nor \U$17359 ( \17674 , \17672 , \17673 );
xnor \U$17360 ( \17675 , \17674 , \4212 );
and \U$17361 ( \17676 , \8127 , \4032 );
and \U$17362 ( \17677 , \7703 , \4030 );
nor \U$17363 ( \17678 , \17676 , \17677 );
xnor \U$17364 ( \17679 , \17678 , \3786 );
and \U$17365 ( \17680 , \17675 , \17679 );
and \U$17366 ( \17681 , \8378 , \3637 );
and \U$17367 ( \17682 , \8373 , \3635 );
nor \U$17368 ( \17683 , \17681 , \17682 );
xnor \U$17369 ( \17684 , \17683 , \3450 );
and \U$17370 ( \17685 , \17679 , \17684 );
and \U$17371 ( \17686 , \17675 , \17684 );
or \U$17372 ( \17687 , \17680 , \17685 , \17686 );
and \U$17373 ( \17688 , \17670 , \17687 );
and \U$17374 ( \17689 , \17654 , \17687 );
or \U$17375 ( \17690 , \17671 , \17688 , \17689 );
and \U$17376 ( \17691 , \4469 , \7238 );
and \U$17377 ( \17692 , \4272 , \7236 );
nor \U$17378 ( \17693 , \17691 , \17692 );
xnor \U$17379 ( \17694 , \17693 , \6978 );
and \U$17380 ( \17695 , \4779 , \6744 );
and \U$17381 ( \17696 , \4771 , \6742 );
nor \U$17382 ( \17697 , \17695 , \17696 );
xnor \U$17383 ( \17698 , \17697 , \6429 );
and \U$17384 ( \17699 , \17694 , \17698 );
and \U$17385 ( \17700 , \5253 , \6235 );
and \U$17386 ( \17701 , \5248 , \6233 );
nor \U$17387 ( \17702 , \17700 , \17701 );
xnor \U$17388 ( \17703 , \17702 , \5895 );
and \U$17389 ( \17704 , \17698 , \17703 );
and \U$17390 ( \17705 , \17694 , \17703 );
or \U$17391 ( \17706 , \17699 , \17704 , \17705 );
and \U$17392 ( \17707 , \3264 , \8896 );
and \U$17393 ( \17708 , \3145 , \8894 );
nor \U$17394 ( \17709 , \17707 , \17708 );
xnor \U$17395 ( \17710 , \17709 , \8525 );
and \U$17396 ( \17711 , \3889 , \8334 );
and \U$17397 ( \17712 , \3681 , \8332 );
nor \U$17398 ( \17713 , \17711 , \17712 );
xnor \U$17399 ( \17714 , \17713 , \8016 );
and \U$17400 ( \17715 , \17710 , \17714 );
and \U$17401 ( \17716 , \4016 , \7767 );
and \U$17402 ( \17717 , \4011 , \7765 );
nor \U$17403 ( \17718 , \17716 , \17717 );
xnor \U$17404 ( \17719 , \17718 , \7518 );
and \U$17405 ( \17720 , \17714 , \17719 );
and \U$17406 ( \17721 , \17710 , \17719 );
or \U$17407 ( \17722 , \17715 , \17720 , \17721 );
and \U$17408 ( \17723 , \17706 , \17722 );
and \U$17409 ( \17724 , \2377 , \10814 );
and \U$17410 ( \17725 , \2233 , \10811 );
nor \U$17411 ( \17726 , \17724 , \17725 );
xnor \U$17412 ( \17727 , \17726 , \9759 );
and \U$17413 ( \17728 , \2666 , \10001 );
and \U$17414 ( \17729 , \2641 , \9999 );
nor \U$17415 ( \17730 , \17728 , \17729 );
xnor \U$17416 ( \17731 , \17730 , \9762 );
and \U$17417 ( \17732 , \17727 , \17731 );
and \U$17418 ( \17733 , \3007 , \9433 );
and \U$17419 ( \17734 , \2840 , \9431 );
nor \U$17420 ( \17735 , \17733 , \17734 );
xnor \U$17421 ( \17736 , \17735 , \9123 );
and \U$17422 ( \17737 , \17731 , \17736 );
and \U$17423 ( \17738 , \17727 , \17736 );
or \U$17424 ( \17739 , \17732 , \17737 , \17738 );
and \U$17425 ( \17740 , \17722 , \17739 );
and \U$17426 ( \17741 , \17706 , \17739 );
or \U$17427 ( \17742 , \17723 , \17740 , \17741 );
and \U$17428 ( \17743 , \17690 , \17742 );
xor \U$17429 ( \17744 , \17482 , \17486 );
xor \U$17430 ( \17745 , \17744 , \17489 );
xor \U$17431 ( \17746 , \17525 , \17529 );
xor \U$17432 ( \17747 , \17746 , \17534 );
and \U$17433 ( \17748 , \17745 , \17747 );
xor \U$17434 ( \17749 , \17542 , \17546 );
xor \U$17435 ( \17750 , \17749 , \17551 );
and \U$17436 ( \17751 , \17747 , \17750 );
and \U$17437 ( \17752 , \17745 , \17750 );
or \U$17438 ( \17753 , \17748 , \17751 , \17752 );
and \U$17439 ( \17754 , \17742 , \17753 );
and \U$17440 ( \17755 , \17690 , \17753 );
or \U$17441 ( \17756 , \17743 , \17754 , \17755 );
xor \U$17442 ( \17757 , \17442 , \17458 );
xor \U$17443 ( \17758 , \17757 , \17475 );
xor \U$17444 ( \17759 , \17492 , \17496 );
xor \U$17445 ( \17760 , \17759 , \17501 );
and \U$17446 ( \17761 , \17758 , \17760 );
xor \U$17447 ( \17762 , \17521 , \17537 );
xor \U$17448 ( \17763 , \17762 , \17554 );
and \U$17449 ( \17764 , \17760 , \17763 );
and \U$17450 ( \17765 , \17758 , \17763 );
or \U$17451 ( \17766 , \17761 , \17764 , \17765 );
and \U$17452 ( \17767 , \17756 , \17766 );
xor \U$17453 ( \17768 , \17509 , \17513 );
xor \U$17454 ( \17769 , \17768 , \17518 );
xor \U$17455 ( \17770 , \17446 , \17450 );
xor \U$17456 ( \17771 , \17770 , \17455 );
and \U$17457 ( \17772 , \17769 , \17771 );
xor \U$17458 ( \17773 , \17463 , \17467 );
xor \U$17459 ( \17774 , \17773 , \17472 );
and \U$17460 ( \17775 , \17771 , \17774 );
and \U$17461 ( \17776 , \17769 , \17774 );
or \U$17462 ( \17777 , \17772 , \17775 , \17776 );
xor \U$17463 ( \17778 , \17562 , \17564 );
xor \U$17464 ( \17779 , \17778 , \17567 );
and \U$17465 ( \17780 , \17777 , \17779 );
xor \U$17466 ( \17781 , \17572 , \17574 );
xor \U$17467 ( \17782 , \17781 , \17577 );
and \U$17468 ( \17783 , \17779 , \17782 );
and \U$17469 ( \17784 , \17777 , \17782 );
or \U$17470 ( \17785 , \17780 , \17783 , \17784 );
and \U$17471 ( \17786 , \17766 , \17785 );
and \U$17472 ( \17787 , \17756 , \17785 );
or \U$17473 ( \17788 , \17767 , \17786 , \17787 );
xor \U$17474 ( \17789 , \17250 , \17266 );
xor \U$17475 ( \17790 , \17789 , \17283 );
xor \U$17476 ( \17791 , \17302 , \17318 );
xor \U$17477 ( \17792 , \17791 , \17335 );
and \U$17478 ( \17793 , \17790 , \17792 );
xor \U$17479 ( \17794 , \17589 , \17591 );
xor \U$17480 ( \17795 , \17794 , \17594 );
and \U$17481 ( \17796 , \17792 , \17795 );
and \U$17482 ( \17797 , \17790 , \17795 );
or \U$17483 ( \17798 , \17793 , \17796 , \17797 );
and \U$17484 ( \17799 , \17788 , \17798 );
xor \U$17485 ( \17800 , \17602 , \17604 );
xor \U$17486 ( \17801 , \17800 , \17607 );
and \U$17487 ( \17802 , \17798 , \17801 );
and \U$17488 ( \17803 , \17788 , \17801 );
or \U$17489 ( \17804 , \17799 , \17802 , \17803 );
xor \U$17490 ( \17805 , \17600 , \17610 );
xor \U$17491 ( \17806 , \17805 , \17613 );
and \U$17492 ( \17807 , \17804 , \17806 );
xor \U$17493 ( \17808 , \17618 , \17620 );
and \U$17494 ( \17809 , \17806 , \17808 );
and \U$17495 ( \17810 , \17804 , \17808 );
or \U$17496 ( \17811 , \17807 , \17809 , \17810 );
xor \U$17497 ( \17812 , \17383 , \17393 );
xor \U$17498 ( \17813 , \17812 , \17396 );
and \U$17499 ( \17814 , \17811 , \17813 );
xor \U$17500 ( \17815 , \17616 , \17621 );
xor \U$17501 ( \17816 , \17815 , \17624 );
and \U$17502 ( \17817 , \17813 , \17816 );
and \U$17503 ( \17818 , \17811 , \17816 );
or \U$17504 ( \17819 , \17814 , \17817 , \17818 );
and \U$17505 ( \17820 , \17638 , \17819 );
xor \U$17506 ( \17821 , \17638 , \17819 );
xor \U$17507 ( \17822 , \17811 , \17813 );
xor \U$17508 ( \17823 , \17822 , \17816 );
and \U$17509 ( \17824 , \4272 , \7767 );
and \U$17510 ( \17825 , \4016 , \7765 );
nor \U$17511 ( \17826 , \17824 , \17825 );
xnor \U$17512 ( \17827 , \17826 , \7518 );
and \U$17513 ( \17828 , \4771 , \7238 );
and \U$17514 ( \17829 , \4469 , \7236 );
nor \U$17515 ( \17830 , \17828 , \17829 );
xnor \U$17516 ( \17831 , \17830 , \6978 );
and \U$17517 ( \17832 , \17827 , \17831 );
and \U$17518 ( \17833 , \5248 , \6744 );
and \U$17519 ( \17834 , \4779 , \6742 );
nor \U$17520 ( \17835 , \17833 , \17834 );
xnor \U$17521 ( \17836 , \17835 , \6429 );
and \U$17522 ( \17837 , \17831 , \17836 );
and \U$17523 ( \17838 , \17827 , \17836 );
or \U$17524 ( \17839 , \17832 , \17837 , \17838 );
and \U$17525 ( \17840 , \3145 , \9433 );
and \U$17526 ( \17841 , \3007 , \9431 );
nor \U$17527 ( \17842 , \17840 , \17841 );
xnor \U$17528 ( \17843 , \17842 , \9123 );
and \U$17529 ( \17844 , \3681 , \8896 );
and \U$17530 ( \17845 , \3264 , \8894 );
nor \U$17531 ( \17846 , \17844 , \17845 );
xnor \U$17532 ( \17847 , \17846 , \8525 );
and \U$17533 ( \17848 , \17843 , \17847 );
and \U$17534 ( \17849 , \4011 , \8334 );
and \U$17535 ( \17850 , \3889 , \8332 );
nor \U$17536 ( \17851 , \17849 , \17850 );
xnor \U$17537 ( \17852 , \17851 , \8016 );
and \U$17538 ( \17853 , \17847 , \17852 );
and \U$17539 ( \17854 , \17843 , \17852 );
or \U$17540 ( \17855 , \17848 , \17853 , \17854 );
and \U$17541 ( \17856 , \17839 , \17855 );
and \U$17542 ( \17857 , \2641 , \10814 );
and \U$17543 ( \17858 , \2377 , \10811 );
nor \U$17544 ( \17859 , \17857 , \17858 );
xnor \U$17545 ( \17860 , \17859 , \9759 );
and \U$17546 ( \17861 , \2840 , \10001 );
and \U$17547 ( \17862 , \2666 , \9999 );
nor \U$17548 ( \17863 , \17861 , \17862 );
xnor \U$17549 ( \17864 , \17863 , \9762 );
and \U$17550 ( \17865 , \17860 , \17864 );
and \U$17551 ( \17866 , \17864 , \2163 );
and \U$17552 ( \17867 , \17860 , \2163 );
or \U$17553 ( \17868 , \17865 , \17866 , \17867 );
and \U$17554 ( \17869 , \17855 , \17868 );
and \U$17555 ( \17870 , \17839 , \17868 );
or \U$17556 ( \17871 , \17856 , \17869 , \17870 );
and \U$17557 ( \17872 , \8697 , \3637 );
and \U$17558 ( \17873 , \8378 , \3635 );
nor \U$17559 ( \17874 , \17872 , \17873 );
xnor \U$17560 ( \17875 , \17874 , \3450 );
and \U$17561 ( \17876 , \9550 , \3324 );
and \U$17562 ( \17877 , \8981 , \3322 );
nor \U$17563 ( \17878 , \17876 , \17877 );
xnor \U$17564 ( \17879 , \17878 , \3119 );
and \U$17565 ( \17880 , \17875 , \17879 );
and \U$17566 ( \17881 , \10161 , \2918 );
and \U$17567 ( \17882 , \9558 , \2916 );
nor \U$17568 ( \17883 , \17881 , \17882 );
xnor \U$17569 ( \17884 , \17883 , \2769 );
and \U$17570 ( \17885 , \17879 , \17884 );
and \U$17571 ( \17886 , \17875 , \17884 );
or \U$17572 ( \17887 , \17880 , \17885 , \17886 );
and \U$17573 ( \17888 , \5517 , \6235 );
and \U$17574 ( \17889 , \5253 , \6233 );
nor \U$17575 ( \17890 , \17888 , \17889 );
xnor \U$17576 ( \17891 , \17890 , \5895 );
and \U$17577 ( \17892 , \6148 , \5646 );
and \U$17578 ( \17893 , \5776 , \5644 );
nor \U$17579 ( \17894 , \17892 , \17893 );
xnor \U$17580 ( \17895 , \17894 , \5405 );
and \U$17581 ( \17896 , \17891 , \17895 );
and \U$17582 ( \17897 , \6500 , \5180 );
and \U$17583 ( \17898 , \6157 , \5178 );
nor \U$17584 ( \17899 , \17897 , \17898 );
xnor \U$17585 ( \17900 , \17899 , \4992 );
and \U$17586 ( \17901 , \17895 , \17900 );
and \U$17587 ( \17902 , \17891 , \17900 );
or \U$17588 ( \17903 , \17896 , \17901 , \17902 );
and \U$17589 ( \17904 , \17887 , \17903 );
and \U$17590 ( \17905 , \7005 , \4806 );
and \U$17591 ( \17906 , \6702 , \4804 );
nor \U$17592 ( \17907 , \17905 , \17906 );
xnor \U$17593 ( \17908 , \17907 , \4574 );
and \U$17594 ( \17909 , \7703 , \4355 );
and \U$17595 ( \17910 , \7177 , \4353 );
nor \U$17596 ( \17911 , \17909 , \17910 );
xnor \U$17597 ( \17912 , \17911 , \4212 );
and \U$17598 ( \17913 , \17908 , \17912 );
and \U$17599 ( \17914 , \8373 , \4032 );
and \U$17600 ( \17915 , \8127 , \4030 );
nor \U$17601 ( \17916 , \17914 , \17915 );
xnor \U$17602 ( \17917 , \17916 , \3786 );
and \U$17603 ( \17918 , \17912 , \17917 );
and \U$17604 ( \17919 , \17908 , \17917 );
or \U$17605 ( \17920 , \17913 , \17918 , \17919 );
and \U$17606 ( \17921 , \17903 , \17920 );
and \U$17607 ( \17922 , \17887 , \17920 );
or \U$17608 ( \17923 , \17904 , \17921 , \17922 );
and \U$17609 ( \17924 , \17871 , \17923 );
and \U$17610 ( \17925 , \10967 , \2300 );
and \U$17611 ( \17926 , \10347 , \2298 );
nor \U$17612 ( \17927 , \17925 , \17926 );
xnor \U$17613 ( \17928 , \17927 , \2163 );
xor \U$17614 ( \17929 , \17642 , \17646 );
xor \U$17615 ( \17930 , \17929 , \17651 );
and \U$17616 ( \17931 , \17928 , \17930 );
xor \U$17617 ( \17932 , \17675 , \17679 );
xor \U$17618 ( \17933 , \17932 , \17684 );
and \U$17619 ( \17934 , \17930 , \17933 );
and \U$17620 ( \17935 , \17928 , \17933 );
or \U$17621 ( \17936 , \17931 , \17934 , \17935 );
and \U$17622 ( \17937 , \17923 , \17936 );
and \U$17623 ( \17938 , \17871 , \17936 );
or \U$17624 ( \17939 , \17924 , \17937 , \17938 );
xor \U$17625 ( \17940 , \17694 , \17698 );
xor \U$17626 ( \17941 , \17940 , \17703 );
xor \U$17627 ( \17942 , \17658 , \17662 );
xor \U$17628 ( \17943 , \17942 , \17667 );
and \U$17629 ( \17944 , \17941 , \17943 );
xor \U$17630 ( \17945 , \17710 , \17714 );
xor \U$17631 ( \17946 , \17945 , \17719 );
and \U$17632 ( \17947 , \17943 , \17946 );
and \U$17633 ( \17948 , \17941 , \17946 );
or \U$17634 ( \17949 , \17944 , \17947 , \17948 );
xor \U$17635 ( \17950 , \17434 , \17438 );
xor \U$17636 ( \17951 , \17950 , \1942 );
and \U$17637 ( \17952 , \17949 , \17951 );
xor \U$17638 ( \17953 , \17769 , \17771 );
xor \U$17639 ( \17954 , \17953 , \17774 );
and \U$17640 ( \17955 , \17951 , \17954 );
and \U$17641 ( \17956 , \17949 , \17954 );
or \U$17642 ( \17957 , \17952 , \17955 , \17956 );
and \U$17643 ( \17958 , \17939 , \17957 );
xor \U$17644 ( \17959 , \17654 , \17670 );
xor \U$17645 ( \17960 , \17959 , \17687 );
xor \U$17646 ( \17961 , \17706 , \17722 );
xor \U$17647 ( \17962 , \17961 , \17739 );
and \U$17648 ( \17963 , \17960 , \17962 );
xor \U$17649 ( \17964 , \17745 , \17747 );
xor \U$17650 ( \17965 , \17964 , \17750 );
and \U$17651 ( \17966 , \17962 , \17965 );
and \U$17652 ( \17967 , \17960 , \17965 );
or \U$17653 ( \17968 , \17963 , \17966 , \17967 );
and \U$17654 ( \17969 , \17957 , \17968 );
and \U$17655 ( \17970 , \17939 , \17968 );
or \U$17656 ( \17971 , \17958 , \17969 , \17970 );
xor \U$17657 ( \17972 , \17690 , \17742 );
xor \U$17658 ( \17973 , \17972 , \17753 );
xor \U$17659 ( \17974 , \17758 , \17760 );
xor \U$17660 ( \17975 , \17974 , \17763 );
and \U$17661 ( \17976 , \17973 , \17975 );
xor \U$17662 ( \17977 , \17777 , \17779 );
xor \U$17663 ( \17978 , \17977 , \17782 );
and \U$17664 ( \17979 , \17975 , \17978 );
and \U$17665 ( \17980 , \17973 , \17978 );
or \U$17666 ( \17981 , \17976 , \17979 , \17980 );
and \U$17667 ( \17982 , \17971 , \17981 );
xor \U$17668 ( \17983 , \17570 , \17580 );
xor \U$17669 ( \17984 , \17983 , \17583 );
and \U$17670 ( \17985 , \17981 , \17984 );
and \U$17671 ( \17986 , \17971 , \17984 );
or \U$17672 ( \17987 , \17982 , \17985 , \17986 );
xor \U$17673 ( \17988 , \17478 , \17504 );
xor \U$17674 ( \17989 , \17988 , \17557 );
xor \U$17675 ( \17990 , \17756 , \17766 );
xor \U$17676 ( \17991 , \17990 , \17785 );
and \U$17677 ( \17992 , \17989 , \17991 );
xor \U$17678 ( \17993 , \17790 , \17792 );
xor \U$17679 ( \17994 , \17993 , \17795 );
and \U$17680 ( \17995 , \17991 , \17994 );
and \U$17681 ( \17996 , \17989 , \17994 );
or \U$17682 ( \17997 , \17992 , \17995 , \17996 );
and \U$17683 ( \17998 , \17987 , \17997 );
xor \U$17684 ( \17999 , \17560 , \17586 );
xor \U$17685 ( \18000 , \17999 , \17597 );
and \U$17686 ( \18001 , \17997 , \18000 );
and \U$17687 ( \18002 , \17987 , \18000 );
or \U$17688 ( \18003 , \17998 , \18001 , \18002 );
xor \U$17689 ( \18004 , \17804 , \17806 );
xor \U$17690 ( \18005 , \18004 , \17808 );
and \U$17691 ( \18006 , \18003 , \18005 );
and \U$17692 ( \18007 , \17823 , \18006 );
xor \U$17693 ( \18008 , \17823 , \18006 );
xor \U$17694 ( \18009 , \18003 , \18005 );
and \U$17695 ( \18010 , \2666 , \10814 );
and \U$17696 ( \18011 , \2641 , \10811 );
nor \U$17697 ( \18012 , \18010 , \18011 );
xnor \U$17698 ( \18013 , \18012 , \9759 );
and \U$17699 ( \18014 , \3007 , \10001 );
and \U$17700 ( \18015 , \2840 , \9999 );
nor \U$17701 ( \18016 , \18014 , \18015 );
xnor \U$17702 ( \18017 , \18016 , \9762 );
and \U$17703 ( \18018 , \18013 , \18017 );
and \U$17704 ( \18019 , \3264 , \9433 );
and \U$17705 ( \18020 , \3145 , \9431 );
nor \U$17706 ( \18021 , \18019 , \18020 );
xnor \U$17707 ( \18022 , \18021 , \9123 );
and \U$17708 ( \18023 , \18017 , \18022 );
and \U$17709 ( \18024 , \18013 , \18022 );
or \U$17710 ( \18025 , \18018 , \18023 , \18024 );
and \U$17711 ( \18026 , \3889 , \8896 );
and \U$17712 ( \18027 , \3681 , \8894 );
nor \U$17713 ( \18028 , \18026 , \18027 );
xnor \U$17714 ( \18029 , \18028 , \8525 );
and \U$17715 ( \18030 , \4016 , \8334 );
and \U$17716 ( \18031 , \4011 , \8332 );
nor \U$17717 ( \18032 , \18030 , \18031 );
xnor \U$17718 ( \18033 , \18032 , \8016 );
and \U$17719 ( \18034 , \18029 , \18033 );
and \U$17720 ( \18035 , \4469 , \7767 );
and \U$17721 ( \18036 , \4272 , \7765 );
nor \U$17722 ( \18037 , \18035 , \18036 );
xnor \U$17723 ( \18038 , \18037 , \7518 );
and \U$17724 ( \18039 , \18033 , \18038 );
and \U$17725 ( \18040 , \18029 , \18038 );
or \U$17726 ( \18041 , \18034 , \18039 , \18040 );
and \U$17727 ( \18042 , \18025 , \18041 );
and \U$17728 ( \18043 , \4779 , \7238 );
and \U$17729 ( \18044 , \4771 , \7236 );
nor \U$17730 ( \18045 , \18043 , \18044 );
xnor \U$17731 ( \18046 , \18045 , \6978 );
and \U$17732 ( \18047 , \5253 , \6744 );
and \U$17733 ( \18048 , \5248 , \6742 );
nor \U$17734 ( \18049 , \18047 , \18048 );
xnor \U$17735 ( \18050 , \18049 , \6429 );
and \U$17736 ( \18051 , \18046 , \18050 );
and \U$17737 ( \18052 , \5776 , \6235 );
and \U$17738 ( \18053 , \5517 , \6233 );
nor \U$17739 ( \18054 , \18052 , \18053 );
xnor \U$17740 ( \18055 , \18054 , \5895 );
and \U$17741 ( \18056 , \18050 , \18055 );
and \U$17742 ( \18057 , \18046 , \18055 );
or \U$17743 ( \18058 , \18051 , \18056 , \18057 );
and \U$17744 ( \18059 , \18041 , \18058 );
and \U$17745 ( \18060 , \18025 , \18058 );
or \U$17746 ( \18061 , \18042 , \18059 , \18060 );
and \U$17747 ( \18062 , \9558 , \3324 );
and \U$17748 ( \18063 , \9550 , \3322 );
nor \U$17749 ( \18064 , \18062 , \18063 );
xnor \U$17750 ( \18065 , \18064 , \3119 );
and \U$17751 ( \18066 , \10166 , \2918 );
and \U$17752 ( \18067 , \10161 , \2916 );
nor \U$17753 ( \18068 , \18066 , \18067 );
xnor \U$17754 ( \18069 , \18068 , \2769 );
and \U$17755 ( \18070 , \18065 , \18069 );
and \U$17756 ( \18071 , \10967 , \2596 );
and \U$17757 ( \18072 , \10347 , \2594 );
nor \U$17758 ( \18073 , \18071 , \18072 );
xnor \U$17759 ( \18074 , \18073 , \2454 );
and \U$17760 ( \18075 , \18069 , \18074 );
and \U$17761 ( \18076 , \18065 , \18074 );
or \U$17762 ( \18077 , \18070 , \18075 , \18076 );
and \U$17763 ( \18078 , \8127 , \4355 );
and \U$17764 ( \18079 , \7703 , \4353 );
nor \U$17765 ( \18080 , \18078 , \18079 );
xnor \U$17766 ( \18081 , \18080 , \4212 );
and \U$17767 ( \18082 , \8378 , \4032 );
and \U$17768 ( \18083 , \8373 , \4030 );
nor \U$17769 ( \18084 , \18082 , \18083 );
xnor \U$17770 ( \18085 , \18084 , \3786 );
and \U$17771 ( \18086 , \18081 , \18085 );
and \U$17772 ( \18087 , \8981 , \3637 );
and \U$17773 ( \18088 , \8697 , \3635 );
nor \U$17774 ( \18089 , \18087 , \18088 );
xnor \U$17775 ( \18090 , \18089 , \3450 );
and \U$17776 ( \18091 , \18085 , \18090 );
and \U$17777 ( \18092 , \18081 , \18090 );
or \U$17778 ( \18093 , \18086 , \18091 , \18092 );
and \U$17779 ( \18094 , \18077 , \18093 );
and \U$17780 ( \18095 , \6157 , \5646 );
and \U$17781 ( \18096 , \6148 , \5644 );
nor \U$17782 ( \18097 , \18095 , \18096 );
xnor \U$17783 ( \18098 , \18097 , \5405 );
and \U$17784 ( \18099 , \6702 , \5180 );
and \U$17785 ( \18100 , \6500 , \5178 );
nor \U$17786 ( \18101 , \18099 , \18100 );
xnor \U$17787 ( \18102 , \18101 , \4992 );
and \U$17788 ( \18103 , \18098 , \18102 );
and \U$17789 ( \18104 , \7177 , \4806 );
and \U$17790 ( \18105 , \7005 , \4804 );
nor \U$17791 ( \18106 , \18104 , \18105 );
xnor \U$17792 ( \18107 , \18106 , \4574 );
and \U$17793 ( \18108 , \18102 , \18107 );
and \U$17794 ( \18109 , \18098 , \18107 );
or \U$17795 ( \18110 , \18103 , \18108 , \18109 );
and \U$17796 ( \18111 , \18093 , \18110 );
and \U$17797 ( \18112 , \18077 , \18110 );
or \U$17798 ( \18113 , \18094 , \18111 , \18112 );
and \U$17799 ( \18114 , \18061 , \18113 );
and \U$17800 ( \18115 , \10347 , \2596 );
and \U$17801 ( \18116 , \10166 , \2594 );
nor \U$17802 ( \18117 , \18115 , \18116 );
xnor \U$17803 ( \18118 , \18117 , \2454 );
nand \U$17804 ( \18119 , \10967 , \2298 );
xnor \U$17805 ( \18120 , \18119 , \2163 );
and \U$17806 ( \18121 , \18118 , \18120 );
xor \U$17807 ( \18122 , \17875 , \17879 );
xor \U$17808 ( \18123 , \18122 , \17884 );
and \U$17809 ( \18124 , \18120 , \18123 );
and \U$17810 ( \18125 , \18118 , \18123 );
or \U$17811 ( \18126 , \18121 , \18124 , \18125 );
and \U$17812 ( \18127 , \18113 , \18126 );
and \U$17813 ( \18128 , \18061 , \18126 );
or \U$17814 ( \18129 , \18114 , \18127 , \18128 );
xor \U$17815 ( \18130 , \17827 , \17831 );
xor \U$17816 ( \18131 , \18130 , \17836 );
xor \U$17817 ( \18132 , \17891 , \17895 );
xor \U$17818 ( \18133 , \18132 , \17900 );
and \U$17819 ( \18134 , \18131 , \18133 );
xor \U$17820 ( \18135 , \17908 , \17912 );
xor \U$17821 ( \18136 , \18135 , \17917 );
and \U$17822 ( \18137 , \18133 , \18136 );
and \U$17823 ( \18138 , \18131 , \18136 );
or \U$17824 ( \18139 , \18134 , \18137 , \18138 );
xor \U$17825 ( \18140 , \17843 , \17847 );
xor \U$17826 ( \18141 , \18140 , \17852 );
xor \U$17827 ( \18142 , \17860 , \17864 );
xor \U$17828 ( \18143 , \18142 , \2163 );
and \U$17829 ( \18144 , \18141 , \18143 );
and \U$17830 ( \18145 , \18139 , \18144 );
xor \U$17831 ( \18146 , \17727 , \17731 );
xor \U$17832 ( \18147 , \18146 , \17736 );
and \U$17833 ( \18148 , \18144 , \18147 );
and \U$17834 ( \18149 , \18139 , \18147 );
or \U$17835 ( \18150 , \18145 , \18148 , \18149 );
and \U$17836 ( \18151 , \18129 , \18150 );
xor \U$17837 ( \18152 , \17887 , \17903 );
xor \U$17838 ( \18153 , \18152 , \17920 );
xor \U$17839 ( \18154 , \17941 , \17943 );
xor \U$17840 ( \18155 , \18154 , \17946 );
and \U$17841 ( \18156 , \18153 , \18155 );
xor \U$17842 ( \18157 , \17928 , \17930 );
xor \U$17843 ( \18158 , \18157 , \17933 );
and \U$17844 ( \18159 , \18155 , \18158 );
and \U$17845 ( \18160 , \18153 , \18158 );
or \U$17846 ( \18161 , \18156 , \18159 , \18160 );
and \U$17847 ( \18162 , \18150 , \18161 );
and \U$17848 ( \18163 , \18129 , \18161 );
or \U$17849 ( \18164 , \18151 , \18162 , \18163 );
xor \U$17850 ( \18165 , \17871 , \17923 );
xor \U$17851 ( \18166 , \18165 , \17936 );
xor \U$17852 ( \18167 , \17949 , \17951 );
xor \U$17853 ( \18168 , \18167 , \17954 );
and \U$17854 ( \18169 , \18166 , \18168 );
xor \U$17855 ( \18170 , \17960 , \17962 );
xor \U$17856 ( \18171 , \18170 , \17965 );
and \U$17857 ( \18172 , \18168 , \18171 );
and \U$17858 ( \18173 , \18166 , \18171 );
or \U$17859 ( \18174 , \18169 , \18172 , \18173 );
and \U$17860 ( \18175 , \18164 , \18174 );
xor \U$17861 ( \18176 , \17973 , \17975 );
xor \U$17862 ( \18177 , \18176 , \17978 );
and \U$17863 ( \18178 , \18174 , \18177 );
and \U$17864 ( \18179 , \18164 , \18177 );
or \U$17865 ( \18180 , \18175 , \18178 , \18179 );
xor \U$17866 ( \18181 , \17971 , \17981 );
xor \U$17867 ( \18182 , \18181 , \17984 );
and \U$17868 ( \18183 , \18180 , \18182 );
xor \U$17869 ( \18184 , \17989 , \17991 );
xor \U$17870 ( \18185 , \18184 , \17994 );
and \U$17871 ( \18186 , \18182 , \18185 );
and \U$17872 ( \18187 , \18180 , \18185 );
or \U$17873 ( \18188 , \18183 , \18186 , \18187 );
xor \U$17874 ( \18189 , \17987 , \17997 );
xor \U$17875 ( \18190 , \18189 , \18000 );
and \U$17876 ( \18191 , \18188 , \18190 );
xor \U$17877 ( \18192 , \17788 , \17798 );
xor \U$17878 ( \18193 , \18192 , \17801 );
and \U$17879 ( \18194 , \18190 , \18193 );
and \U$17880 ( \18195 , \18188 , \18193 );
or \U$17881 ( \18196 , \18191 , \18194 , \18195 );
and \U$17882 ( \18197 , \18009 , \18196 );
xor \U$17883 ( \18198 , \18009 , \18196 );
xor \U$17884 ( \18199 , \18188 , \18190 );
xor \U$17885 ( \18200 , \18199 , \18193 );
and \U$17886 ( \18201 , \2840 , \10814 );
and \U$17887 ( \18202 , \2666 , \10811 );
nor \U$17888 ( \18203 , \18201 , \18202 );
xnor \U$17889 ( \18204 , \18203 , \9759 );
and \U$17890 ( \18205 , \3145 , \10001 );
and \U$17891 ( \18206 , \3007 , \9999 );
nor \U$17892 ( \18207 , \18205 , \18206 );
xnor \U$17893 ( \18208 , \18207 , \9762 );
and \U$17894 ( \18209 , \18204 , \18208 );
and \U$17895 ( \18210 , \18208 , \2454 );
and \U$17896 ( \18211 , \18204 , \2454 );
or \U$17897 ( \18212 , \18209 , \18210 , \18211 );
and \U$17898 ( \18213 , \3681 , \9433 );
and \U$17899 ( \18214 , \3264 , \9431 );
nor \U$17900 ( \18215 , \18213 , \18214 );
xnor \U$17901 ( \18216 , \18215 , \9123 );
and \U$17902 ( \18217 , \4011 , \8896 );
and \U$17903 ( \18218 , \3889 , \8894 );
nor \U$17904 ( \18219 , \18217 , \18218 );
xnor \U$17905 ( \18220 , \18219 , \8525 );
and \U$17906 ( \18221 , \18216 , \18220 );
and \U$17907 ( \18222 , \4272 , \8334 );
and \U$17908 ( \18223 , \4016 , \8332 );
nor \U$17909 ( \18224 , \18222 , \18223 );
xnor \U$17910 ( \18225 , \18224 , \8016 );
and \U$17911 ( \18226 , \18220 , \18225 );
and \U$17912 ( \18227 , \18216 , \18225 );
or \U$17913 ( \18228 , \18221 , \18226 , \18227 );
and \U$17914 ( \18229 , \18212 , \18228 );
and \U$17915 ( \18230 , \4771 , \7767 );
and \U$17916 ( \18231 , \4469 , \7765 );
nor \U$17917 ( \18232 , \18230 , \18231 );
xnor \U$17918 ( \18233 , \18232 , \7518 );
and \U$17919 ( \18234 , \5248 , \7238 );
and \U$17920 ( \18235 , \4779 , \7236 );
nor \U$17921 ( \18236 , \18234 , \18235 );
xnor \U$17922 ( \18237 , \18236 , \6978 );
and \U$17923 ( \18238 , \18233 , \18237 );
and \U$17924 ( \18239 , \5517 , \6744 );
and \U$17925 ( \18240 , \5253 , \6742 );
nor \U$17926 ( \18241 , \18239 , \18240 );
xnor \U$17927 ( \18242 , \18241 , \6429 );
and \U$17928 ( \18243 , \18237 , \18242 );
and \U$17929 ( \18244 , \18233 , \18242 );
or \U$17930 ( \18245 , \18238 , \18243 , \18244 );
and \U$17931 ( \18246 , \18228 , \18245 );
and \U$17932 ( \18247 , \18212 , \18245 );
or \U$17933 ( \18248 , \18229 , \18246 , \18247 );
and \U$17934 ( \18249 , \6148 , \6235 );
and \U$17935 ( \18250 , \5776 , \6233 );
nor \U$17936 ( \18251 , \18249 , \18250 );
xnor \U$17937 ( \18252 , \18251 , \5895 );
and \U$17938 ( \18253 , \6500 , \5646 );
and \U$17939 ( \18254 , \6157 , \5644 );
nor \U$17940 ( \18255 , \18253 , \18254 );
xnor \U$17941 ( \18256 , \18255 , \5405 );
and \U$17942 ( \18257 , \18252 , \18256 );
and \U$17943 ( \18258 , \7005 , \5180 );
and \U$17944 ( \18259 , \6702 , \5178 );
nor \U$17945 ( \18260 , \18258 , \18259 );
xnor \U$17946 ( \18261 , \18260 , \4992 );
and \U$17947 ( \18262 , \18256 , \18261 );
and \U$17948 ( \18263 , \18252 , \18261 );
or \U$17949 ( \18264 , \18257 , \18262 , \18263 );
and \U$17950 ( \18265 , \7703 , \4806 );
and \U$17951 ( \18266 , \7177 , \4804 );
nor \U$17952 ( \18267 , \18265 , \18266 );
xnor \U$17953 ( \18268 , \18267 , \4574 );
and \U$17954 ( \18269 , \8373 , \4355 );
and \U$17955 ( \18270 , \8127 , \4353 );
nor \U$17956 ( \18271 , \18269 , \18270 );
xnor \U$17957 ( \18272 , \18271 , \4212 );
and \U$17958 ( \18273 , \18268 , \18272 );
and \U$17959 ( \18274 , \8697 , \4032 );
and \U$17960 ( \18275 , \8378 , \4030 );
nor \U$17961 ( \18276 , \18274 , \18275 );
xnor \U$17962 ( \18277 , \18276 , \3786 );
and \U$17963 ( \18278 , \18272 , \18277 );
and \U$17964 ( \18279 , \18268 , \18277 );
or \U$17965 ( \18280 , \18273 , \18278 , \18279 );
and \U$17966 ( \18281 , \18264 , \18280 );
and \U$17967 ( \18282 , \9550 , \3637 );
and \U$17968 ( \18283 , \8981 , \3635 );
nor \U$17969 ( \18284 , \18282 , \18283 );
xnor \U$17970 ( \18285 , \18284 , \3450 );
and \U$17971 ( \18286 , \10161 , \3324 );
and \U$17972 ( \18287 , \9558 , \3322 );
nor \U$17973 ( \18288 , \18286 , \18287 );
xnor \U$17974 ( \18289 , \18288 , \3119 );
and \U$17975 ( \18290 , \18285 , \18289 );
and \U$17976 ( \18291 , \10347 , \2918 );
and \U$17977 ( \18292 , \10166 , \2916 );
nor \U$17978 ( \18293 , \18291 , \18292 );
xnor \U$17979 ( \18294 , \18293 , \2769 );
and \U$17980 ( \18295 , \18289 , \18294 );
and \U$17981 ( \18296 , \18285 , \18294 );
or \U$17982 ( \18297 , \18290 , \18295 , \18296 );
and \U$17983 ( \18298 , \18280 , \18297 );
and \U$17984 ( \18299 , \18264 , \18297 );
or \U$17985 ( \18300 , \18281 , \18298 , \18299 );
and \U$17986 ( \18301 , \18248 , \18300 );
xor \U$17987 ( \18302 , \18065 , \18069 );
xor \U$17988 ( \18303 , \18302 , \18074 );
xor \U$17989 ( \18304 , \18081 , \18085 );
xor \U$17990 ( \18305 , \18304 , \18090 );
and \U$17991 ( \18306 , \18303 , \18305 );
xor \U$17992 ( \18307 , \18098 , \18102 );
xor \U$17993 ( \18308 , \18307 , \18107 );
and \U$17994 ( \18309 , \18305 , \18308 );
and \U$17995 ( \18310 , \18303 , \18308 );
or \U$17996 ( \18311 , \18306 , \18309 , \18310 );
and \U$17997 ( \18312 , \18300 , \18311 );
and \U$17998 ( \18313 , \18248 , \18311 );
or \U$17999 ( \18314 , \18301 , \18312 , \18313 );
xor \U$18000 ( \18315 , \18025 , \18041 );
xor \U$18001 ( \18316 , \18315 , \18058 );
xor \U$18002 ( \18317 , \18077 , \18093 );
xor \U$18003 ( \18318 , \18317 , \18110 );
and \U$18004 ( \18319 , \18316 , \18318 );
xor \U$18005 ( \18320 , \18118 , \18120 );
xor \U$18006 ( \18321 , \18320 , \18123 );
and \U$18007 ( \18322 , \18318 , \18321 );
and \U$18008 ( \18323 , \18316 , \18321 );
or \U$18009 ( \18324 , \18319 , \18322 , \18323 );
and \U$18010 ( \18325 , \18314 , \18324 );
xor \U$18011 ( \18326 , \18013 , \18017 );
xor \U$18012 ( \18327 , \18326 , \18022 );
xor \U$18013 ( \18328 , \18029 , \18033 );
xor \U$18014 ( \18329 , \18328 , \18038 );
and \U$18015 ( \18330 , \18327 , \18329 );
xor \U$18016 ( \18331 , \18046 , \18050 );
xor \U$18017 ( \18332 , \18331 , \18055 );
and \U$18018 ( \18333 , \18329 , \18332 );
and \U$18019 ( \18334 , \18327 , \18332 );
or \U$18020 ( \18335 , \18330 , \18333 , \18334 );
xor \U$18021 ( \18336 , \18131 , \18133 );
xor \U$18022 ( \18337 , \18336 , \18136 );
and \U$18023 ( \18338 , \18335 , \18337 );
xor \U$18024 ( \18339 , \18141 , \18143 );
and \U$18025 ( \18340 , \18337 , \18339 );
and \U$18026 ( \18341 , \18335 , \18339 );
or \U$18027 ( \18342 , \18338 , \18340 , \18341 );
and \U$18028 ( \18343 , \18324 , \18342 );
and \U$18029 ( \18344 , \18314 , \18342 );
or \U$18030 ( \18345 , \18325 , \18343 , \18344 );
xor \U$18031 ( \18346 , \17839 , \17855 );
xor \U$18032 ( \18347 , \18346 , \17868 );
xor \U$18033 ( \18348 , \18139 , \18144 );
xor \U$18034 ( \18349 , \18348 , \18147 );
and \U$18035 ( \18350 , \18347 , \18349 );
xor \U$18036 ( \18351 , \18153 , \18155 );
xor \U$18037 ( \18352 , \18351 , \18158 );
and \U$18038 ( \18353 , \18349 , \18352 );
and \U$18039 ( \18354 , \18347 , \18352 );
or \U$18040 ( \18355 , \18350 , \18353 , \18354 );
and \U$18041 ( \18356 , \18345 , \18355 );
xor \U$18042 ( \18357 , \18166 , \18168 );
xor \U$18043 ( \18358 , \18357 , \18171 );
and \U$18044 ( \18359 , \18355 , \18358 );
and \U$18045 ( \18360 , \18345 , \18358 );
or \U$18046 ( \18361 , \18356 , \18359 , \18360 );
xor \U$18047 ( \18362 , \17939 , \17957 );
xor \U$18048 ( \18363 , \18362 , \17968 );
and \U$18049 ( \18364 , \18361 , \18363 );
xor \U$18050 ( \18365 , \18164 , \18174 );
xor \U$18051 ( \18366 , \18365 , \18177 );
and \U$18052 ( \18367 , \18363 , \18366 );
and \U$18053 ( \18368 , \18361 , \18366 );
or \U$18054 ( \18369 , \18364 , \18367 , \18368 );
xor \U$18055 ( \18370 , \18180 , \18182 );
xor \U$18056 ( \18371 , \18370 , \18185 );
and \U$18057 ( \18372 , \18369 , \18371 );
and \U$18058 ( \18373 , \18200 , \18372 );
xor \U$18059 ( \18374 , \18200 , \18372 );
xor \U$18060 ( \18375 , \18369 , \18371 );
and \U$18061 ( \18376 , \5253 , \7238 );
and \U$18062 ( \18377 , \5248 , \7236 );
nor \U$18063 ( \18378 , \18376 , \18377 );
xnor \U$18064 ( \18379 , \18378 , \6978 );
and \U$18065 ( \18380 , \5776 , \6744 );
and \U$18066 ( \18381 , \5517 , \6742 );
nor \U$18067 ( \18382 , \18380 , \18381 );
xnor \U$18068 ( \18383 , \18382 , \6429 );
and \U$18069 ( \18384 , \18379 , \18383 );
and \U$18070 ( \18385 , \6157 , \6235 );
and \U$18071 ( \18386 , \6148 , \6233 );
nor \U$18072 ( \18387 , \18385 , \18386 );
xnor \U$18073 ( \18388 , \18387 , \5895 );
and \U$18074 ( \18389 , \18383 , \18388 );
and \U$18075 ( \18390 , \18379 , \18388 );
or \U$18076 ( \18391 , \18384 , \18389 , \18390 );
and \U$18077 ( \18392 , \3007 , \10814 );
and \U$18078 ( \18393 , \2840 , \10811 );
nor \U$18079 ( \18394 , \18392 , \18393 );
xnor \U$18080 ( \18395 , \18394 , \9759 );
and \U$18081 ( \18396 , \3264 , \10001 );
and \U$18082 ( \18397 , \3145 , \9999 );
nor \U$18083 ( \18398 , \18396 , \18397 );
xnor \U$18084 ( \18399 , \18398 , \9762 );
and \U$18085 ( \18400 , \18395 , \18399 );
and \U$18086 ( \18401 , \3889 , \9433 );
and \U$18087 ( \18402 , \3681 , \9431 );
nor \U$18088 ( \18403 , \18401 , \18402 );
xnor \U$18089 ( \18404 , \18403 , \9123 );
and \U$18090 ( \18405 , \18399 , \18404 );
and \U$18091 ( \18406 , \18395 , \18404 );
or \U$18092 ( \18407 , \18400 , \18405 , \18406 );
and \U$18093 ( \18408 , \18391 , \18407 );
and \U$18094 ( \18409 , \4016 , \8896 );
and \U$18095 ( \18410 , \4011 , \8894 );
nor \U$18096 ( \18411 , \18409 , \18410 );
xnor \U$18097 ( \18412 , \18411 , \8525 );
and \U$18098 ( \18413 , \4469 , \8334 );
and \U$18099 ( \18414 , \4272 , \8332 );
nor \U$18100 ( \18415 , \18413 , \18414 );
xnor \U$18101 ( \18416 , \18415 , \8016 );
and \U$18102 ( \18417 , \18412 , \18416 );
and \U$18103 ( \18418 , \4779 , \7767 );
and \U$18104 ( \18419 , \4771 , \7765 );
nor \U$18105 ( \18420 , \18418 , \18419 );
xnor \U$18106 ( \18421 , \18420 , \7518 );
and \U$18107 ( \18422 , \18416 , \18421 );
and \U$18108 ( \18423 , \18412 , \18421 );
or \U$18109 ( \18424 , \18417 , \18422 , \18423 );
and \U$18110 ( \18425 , \18407 , \18424 );
and \U$18111 ( \18426 , \18391 , \18424 );
or \U$18112 ( \18427 , \18408 , \18425 , \18426 );
and \U$18113 ( \18428 , \8378 , \4355 );
and \U$18114 ( \18429 , \8373 , \4353 );
nor \U$18115 ( \18430 , \18428 , \18429 );
xnor \U$18116 ( \18431 , \18430 , \4212 );
and \U$18117 ( \18432 , \8981 , \4032 );
and \U$18118 ( \18433 , \8697 , \4030 );
nor \U$18119 ( \18434 , \18432 , \18433 );
xnor \U$18120 ( \18435 , \18434 , \3786 );
and \U$18121 ( \18436 , \18431 , \18435 );
and \U$18122 ( \18437 , \9558 , \3637 );
and \U$18123 ( \18438 , \9550 , \3635 );
nor \U$18124 ( \18439 , \18437 , \18438 );
xnor \U$18125 ( \18440 , \18439 , \3450 );
and \U$18126 ( \18441 , \18435 , \18440 );
and \U$18127 ( \18442 , \18431 , \18440 );
or \U$18128 ( \18443 , \18436 , \18441 , \18442 );
and \U$18129 ( \18444 , \6702 , \5646 );
and \U$18130 ( \18445 , \6500 , \5644 );
nor \U$18131 ( \18446 , \18444 , \18445 );
xnor \U$18132 ( \18447 , \18446 , \5405 );
and \U$18133 ( \18448 , \7177 , \5180 );
and \U$18134 ( \18449 , \7005 , \5178 );
nor \U$18135 ( \18450 , \18448 , \18449 );
xnor \U$18136 ( \18451 , \18450 , \4992 );
and \U$18137 ( \18452 , \18447 , \18451 );
and \U$18138 ( \18453 , \8127 , \4806 );
and \U$18139 ( \18454 , \7703 , \4804 );
nor \U$18140 ( \18455 , \18453 , \18454 );
xnor \U$18141 ( \18456 , \18455 , \4574 );
and \U$18142 ( \18457 , \18451 , \18456 );
and \U$18143 ( \18458 , \18447 , \18456 );
or \U$18144 ( \18459 , \18452 , \18457 , \18458 );
and \U$18145 ( \18460 , \18443 , \18459 );
and \U$18146 ( \18461 , \10166 , \3324 );
and \U$18147 ( \18462 , \10161 , \3322 );
nor \U$18148 ( \18463 , \18461 , \18462 );
xnor \U$18149 ( \18464 , \18463 , \3119 );
and \U$18150 ( \18465 , \10967 , \2918 );
and \U$18151 ( \18466 , \10347 , \2916 );
nor \U$18152 ( \18467 , \18465 , \18466 );
xnor \U$18153 ( \18468 , \18467 , \2769 );
and \U$18154 ( \18469 , \18464 , \18468 );
and \U$18155 ( \18470 , \18459 , \18469 );
and \U$18156 ( \18471 , \18443 , \18469 );
or \U$18157 ( \18472 , \18460 , \18470 , \18471 );
and \U$18158 ( \18473 , \18427 , \18472 );
nand \U$18159 ( \18474 , \10967 , \2594 );
xnor \U$18160 ( \18475 , \18474 , \2454 );
xor \U$18161 ( \18476 , \18268 , \18272 );
xor \U$18162 ( \18477 , \18476 , \18277 );
and \U$18163 ( \18478 , \18475 , \18477 );
xor \U$18164 ( \18479 , \18285 , \18289 );
xor \U$18165 ( \18480 , \18479 , \18294 );
and \U$18166 ( \18481 , \18477 , \18480 );
and \U$18167 ( \18482 , \18475 , \18480 );
or \U$18168 ( \18483 , \18478 , \18481 , \18482 );
and \U$18169 ( \18484 , \18472 , \18483 );
and \U$18170 ( \18485 , \18427 , \18483 );
or \U$18171 ( \18486 , \18473 , \18484 , \18485 );
xor \U$18172 ( \18487 , \18216 , \18220 );
xor \U$18173 ( \18488 , \18487 , \18225 );
xor \U$18174 ( \18489 , \18252 , \18256 );
xor \U$18175 ( \18490 , \18489 , \18261 );
and \U$18176 ( \18491 , \18488 , \18490 );
xor \U$18177 ( \18492 , \18233 , \18237 );
xor \U$18178 ( \18493 , \18492 , \18242 );
and \U$18179 ( \18494 , \18490 , \18493 );
and \U$18180 ( \18495 , \18488 , \18493 );
or \U$18181 ( \18496 , \18491 , \18494 , \18495 );
xor \U$18182 ( \18497 , \18303 , \18305 );
xor \U$18183 ( \18498 , \18497 , \18308 );
and \U$18184 ( \18499 , \18496 , \18498 );
xor \U$18185 ( \18500 , \18327 , \18329 );
xor \U$18186 ( \18501 , \18500 , \18332 );
and \U$18187 ( \18502 , \18498 , \18501 );
and \U$18188 ( \18503 , \18496 , \18501 );
or \U$18189 ( \18504 , \18499 , \18502 , \18503 );
and \U$18190 ( \18505 , \18486 , \18504 );
xor \U$18191 ( \18506 , \18212 , \18228 );
xor \U$18192 ( \18507 , \18506 , \18245 );
xor \U$18193 ( \18508 , \18264 , \18280 );
xor \U$18194 ( \18509 , \18508 , \18297 );
and \U$18195 ( \18510 , \18507 , \18509 );
and \U$18196 ( \18511 , \18504 , \18510 );
and \U$18197 ( \18512 , \18486 , \18510 );
or \U$18198 ( \18513 , \18505 , \18511 , \18512 );
xor \U$18199 ( \18514 , \18248 , \18300 );
xor \U$18200 ( \18515 , \18514 , \18311 );
xor \U$18201 ( \18516 , \18316 , \18318 );
xor \U$18202 ( \18517 , \18516 , \18321 );
and \U$18203 ( \18518 , \18515 , \18517 );
xor \U$18204 ( \18519 , \18335 , \18337 );
xor \U$18205 ( \18520 , \18519 , \18339 );
and \U$18206 ( \18521 , \18517 , \18520 );
and \U$18207 ( \18522 , \18515 , \18520 );
or \U$18208 ( \18523 , \18518 , \18521 , \18522 );
and \U$18209 ( \18524 , \18513 , \18523 );
xor \U$18210 ( \18525 , \18061 , \18113 );
xor \U$18211 ( \18526 , \18525 , \18126 );
and \U$18212 ( \18527 , \18523 , \18526 );
and \U$18213 ( \18528 , \18513 , \18526 );
or \U$18214 ( \18529 , \18524 , \18527 , \18528 );
xor \U$18215 ( \18530 , \18314 , \18324 );
xor \U$18216 ( \18531 , \18530 , \18342 );
xor \U$18217 ( \18532 , \18347 , \18349 );
xor \U$18218 ( \18533 , \18532 , \18352 );
and \U$18219 ( \18534 , \18531 , \18533 );
and \U$18220 ( \18535 , \18529 , \18534 );
xor \U$18221 ( \18536 , \18129 , \18150 );
xor \U$18222 ( \18537 , \18536 , \18161 );
and \U$18223 ( \18538 , \18534 , \18537 );
and \U$18224 ( \18539 , \18529 , \18537 );
or \U$18225 ( \18540 , \18535 , \18538 , \18539 );
xor \U$18226 ( \18541 , \18361 , \18363 );
xor \U$18227 ( \18542 , \18541 , \18366 );
and \U$18228 ( \18543 , \18540 , \18542 );
and \U$18229 ( \18544 , \18375 , \18543 );
xor \U$18230 ( \18545 , \18375 , \18543 );
xor \U$18231 ( \18546 , \18540 , \18542 );
xor \U$18232 ( \18547 , \18529 , \18534 );
xor \U$18233 ( \18548 , \18547 , \18537 );
xor \U$18234 ( \18549 , \18345 , \18355 );
xor \U$18235 ( \18550 , \18549 , \18358 );
and \U$18236 ( \18551 , \18548 , \18550 );
and \U$18237 ( \18552 , \18546 , \18551 );
xor \U$18238 ( \18553 , \18546 , \18551 );
xor \U$18239 ( \18554 , \18548 , \18550 );
and \U$18240 ( \18555 , \8373 , \4806 );
and \U$18241 ( \18556 , \8127 , \4804 );
nor \U$18242 ( \18557 , \18555 , \18556 );
xnor \U$18243 ( \18558 , \18557 , \4574 );
and \U$18244 ( \18559 , \8697 , \4355 );
and \U$18245 ( \18560 , \8378 , \4353 );
nor \U$18246 ( \18561 , \18559 , \18560 );
xnor \U$18247 ( \18562 , \18561 , \4212 );
and \U$18248 ( \18563 , \18558 , \18562 );
and \U$18249 ( \18564 , \9550 , \4032 );
and \U$18250 ( \18565 , \8981 , \4030 );
nor \U$18251 ( \18566 , \18564 , \18565 );
xnor \U$18252 ( \18567 , \18566 , \3786 );
and \U$18253 ( \18568 , \18562 , \18567 );
and \U$18254 ( \18569 , \18558 , \18567 );
or \U$18255 ( \18570 , \18563 , \18568 , \18569 );
and \U$18256 ( \18571 , \10161 , \3637 );
and \U$18257 ( \18572 , \9558 , \3635 );
nor \U$18258 ( \18573 , \18571 , \18572 );
xnor \U$18259 ( \18574 , \18573 , \3450 );
and \U$18260 ( \18575 , \10347 , \3324 );
and \U$18261 ( \18576 , \10166 , \3322 );
nor \U$18262 ( \18577 , \18575 , \18576 );
xnor \U$18263 ( \18578 , \18577 , \3119 );
and \U$18264 ( \18579 , \18574 , \18578 );
nand \U$18265 ( \18580 , \10967 , \2916 );
xnor \U$18266 ( \18581 , \18580 , \2769 );
and \U$18267 ( \18582 , \18578 , \18581 );
and \U$18268 ( \18583 , \18574 , \18581 );
or \U$18269 ( \18584 , \18579 , \18582 , \18583 );
and \U$18270 ( \18585 , \18570 , \18584 );
and \U$18271 ( \18586 , \6500 , \6235 );
and \U$18272 ( \18587 , \6157 , \6233 );
nor \U$18273 ( \18588 , \18586 , \18587 );
xnor \U$18274 ( \18589 , \18588 , \5895 );
and \U$18275 ( \18590 , \7005 , \5646 );
and \U$18276 ( \18591 , \6702 , \5644 );
nor \U$18277 ( \18592 , \18590 , \18591 );
xnor \U$18278 ( \18593 , \18592 , \5405 );
and \U$18279 ( \18594 , \18589 , \18593 );
and \U$18280 ( \18595 , \7703 , \5180 );
and \U$18281 ( \18596 , \7177 , \5178 );
nor \U$18282 ( \18597 , \18595 , \18596 );
xnor \U$18283 ( \18598 , \18597 , \4992 );
and \U$18284 ( \18599 , \18593 , \18598 );
and \U$18285 ( \18600 , \18589 , \18598 );
or \U$18286 ( \18601 , \18594 , \18599 , \18600 );
and \U$18287 ( \18602 , \18584 , \18601 );
and \U$18288 ( \18603 , \18570 , \18601 );
or \U$18289 ( \18604 , \18585 , \18602 , \18603 );
and \U$18290 ( \18605 , \5248 , \7767 );
and \U$18291 ( \18606 , \4779 , \7765 );
nor \U$18292 ( \18607 , \18605 , \18606 );
xnor \U$18293 ( \18608 , \18607 , \7518 );
and \U$18294 ( \18609 , \5517 , \7238 );
and \U$18295 ( \18610 , \5253 , \7236 );
nor \U$18296 ( \18611 , \18609 , \18610 );
xnor \U$18297 ( \18612 , \18611 , \6978 );
and \U$18298 ( \18613 , \18608 , \18612 );
and \U$18299 ( \18614 , \6148 , \6744 );
and \U$18300 ( \18615 , \5776 , \6742 );
nor \U$18301 ( \18616 , \18614 , \18615 );
xnor \U$18302 ( \18617 , \18616 , \6429 );
and \U$18303 ( \18618 , \18612 , \18617 );
and \U$18304 ( \18619 , \18608 , \18617 );
or \U$18305 ( \18620 , \18613 , \18618 , \18619 );
and \U$18306 ( \18621 , \3145 , \10814 );
and \U$18307 ( \18622 , \3007 , \10811 );
nor \U$18308 ( \18623 , \18621 , \18622 );
xnor \U$18309 ( \18624 , \18623 , \9759 );
and \U$18310 ( \18625 , \3681 , \10001 );
and \U$18311 ( \18626 , \3264 , \9999 );
nor \U$18312 ( \18627 , \18625 , \18626 );
xnor \U$18313 ( \18628 , \18627 , \9762 );
and \U$18314 ( \18629 , \18624 , \18628 );
and \U$18315 ( \18630 , \18628 , \2769 );
and \U$18316 ( \18631 , \18624 , \2769 );
or \U$18317 ( \18632 , \18629 , \18630 , \18631 );
and \U$18318 ( \18633 , \18620 , \18632 );
and \U$18319 ( \18634 , \4011 , \9433 );
and \U$18320 ( \18635 , \3889 , \9431 );
nor \U$18321 ( \18636 , \18634 , \18635 );
xnor \U$18322 ( \18637 , \18636 , \9123 );
and \U$18323 ( \18638 , \4272 , \8896 );
and \U$18324 ( \18639 , \4016 , \8894 );
nor \U$18325 ( \18640 , \18638 , \18639 );
xnor \U$18326 ( \18641 , \18640 , \8525 );
and \U$18327 ( \18642 , \18637 , \18641 );
and \U$18328 ( \18643 , \4771 , \8334 );
and \U$18329 ( \18644 , \4469 , \8332 );
nor \U$18330 ( \18645 , \18643 , \18644 );
xnor \U$18331 ( \18646 , \18645 , \8016 );
and \U$18332 ( \18647 , \18641 , \18646 );
and \U$18333 ( \18648 , \18637 , \18646 );
or \U$18334 ( \18649 , \18642 , \18647 , \18648 );
and \U$18335 ( \18650 , \18632 , \18649 );
and \U$18336 ( \18651 , \18620 , \18649 );
or \U$18337 ( \18652 , \18633 , \18650 , \18651 );
and \U$18338 ( \18653 , \18604 , \18652 );
xor \U$18339 ( \18654 , \18431 , \18435 );
xor \U$18340 ( \18655 , \18654 , \18440 );
xor \U$18341 ( \18656 , \18447 , \18451 );
xor \U$18342 ( \18657 , \18656 , \18456 );
and \U$18343 ( \18658 , \18655 , \18657 );
xor \U$18344 ( \18659 , \18464 , \18468 );
and \U$18345 ( \18660 , \18657 , \18659 );
and \U$18346 ( \18661 , \18655 , \18659 );
or \U$18347 ( \18662 , \18658 , \18660 , \18661 );
and \U$18348 ( \18663 , \18652 , \18662 );
and \U$18349 ( \18664 , \18604 , \18662 );
or \U$18350 ( \18665 , \18653 , \18663 , \18664 );
xor \U$18351 ( \18666 , \18379 , \18383 );
xor \U$18352 ( \18667 , \18666 , \18388 );
xor \U$18353 ( \18668 , \18395 , \18399 );
xor \U$18354 ( \18669 , \18668 , \18404 );
and \U$18355 ( \18670 , \18667 , \18669 );
xor \U$18356 ( \18671 , \18412 , \18416 );
xor \U$18357 ( \18672 , \18671 , \18421 );
and \U$18358 ( \18673 , \18669 , \18672 );
and \U$18359 ( \18674 , \18667 , \18672 );
or \U$18360 ( \18675 , \18670 , \18673 , \18674 );
xor \U$18361 ( \18676 , \18204 , \18208 );
xor \U$18362 ( \18677 , \18676 , \2454 );
and \U$18363 ( \18678 , \18675 , \18677 );
xor \U$18364 ( \18679 , \18488 , \18490 );
xor \U$18365 ( \18680 , \18679 , \18493 );
and \U$18366 ( \18681 , \18677 , \18680 );
and \U$18367 ( \18682 , \18675 , \18680 );
or \U$18368 ( \18683 , \18678 , \18681 , \18682 );
and \U$18369 ( \18684 , \18665 , \18683 );
xor \U$18370 ( \18685 , \18391 , \18407 );
xor \U$18371 ( \18686 , \18685 , \18424 );
xor \U$18372 ( \18687 , \18443 , \18459 );
xor \U$18373 ( \18688 , \18687 , \18469 );
and \U$18374 ( \18689 , \18686 , \18688 );
xor \U$18375 ( \18690 , \18475 , \18477 );
xor \U$18376 ( \18691 , \18690 , \18480 );
and \U$18377 ( \18692 , \18688 , \18691 );
and \U$18378 ( \18693 , \18686 , \18691 );
or \U$18379 ( \18694 , \18689 , \18692 , \18693 );
and \U$18380 ( \18695 , \18683 , \18694 );
and \U$18381 ( \18696 , \18665 , \18694 );
or \U$18382 ( \18697 , \18684 , \18695 , \18696 );
xor \U$18383 ( \18698 , \18427 , \18472 );
xor \U$18384 ( \18699 , \18698 , \18483 );
xor \U$18385 ( \18700 , \18496 , \18498 );
xor \U$18386 ( \18701 , \18700 , \18501 );
and \U$18387 ( \18702 , \18699 , \18701 );
xor \U$18388 ( \18703 , \18507 , \18509 );
and \U$18389 ( \18704 , \18701 , \18703 );
and \U$18390 ( \18705 , \18699 , \18703 );
or \U$18391 ( \18706 , \18702 , \18704 , \18705 );
and \U$18392 ( \18707 , \18697 , \18706 );
xor \U$18393 ( \18708 , \18515 , \18517 );
xor \U$18394 ( \18709 , \18708 , \18520 );
and \U$18395 ( \18710 , \18706 , \18709 );
and \U$18396 ( \18711 , \18697 , \18709 );
or \U$18397 ( \18712 , \18707 , \18710 , \18711 );
xor \U$18398 ( \18713 , \18513 , \18523 );
xor \U$18399 ( \18714 , \18713 , \18526 );
and \U$18400 ( \18715 , \18712 , \18714 );
xor \U$18401 ( \18716 , \18531 , \18533 );
and \U$18402 ( \18717 , \18714 , \18716 );
and \U$18403 ( \18718 , \18712 , \18716 );
or \U$18404 ( \18719 , \18715 , \18717 , \18718 );
and \U$18405 ( \18720 , \18554 , \18719 );
xor \U$18406 ( \18721 , \18554 , \18719 );
xor \U$18407 ( \18722 , \18712 , \18714 );
xor \U$18408 ( \18723 , \18722 , \18716 );
and \U$18409 ( \18724 , \4469 , \8896 );
and \U$18410 ( \18725 , \4272 , \8894 );
nor \U$18411 ( \18726 , \18724 , \18725 );
xnor \U$18412 ( \18727 , \18726 , \8525 );
and \U$18413 ( \18728 , \4779 , \8334 );
and \U$18414 ( \18729 , \4771 , \8332 );
nor \U$18415 ( \18730 , \18728 , \18729 );
xnor \U$18416 ( \18731 , \18730 , \8016 );
and \U$18417 ( \18732 , \18727 , \18731 );
and \U$18418 ( \18733 , \5253 , \7767 );
and \U$18419 ( \18734 , \5248 , \7765 );
nor \U$18420 ( \18735 , \18733 , \18734 );
xnor \U$18421 ( \18736 , \18735 , \7518 );
and \U$18422 ( \18737 , \18731 , \18736 );
and \U$18423 ( \18738 , \18727 , \18736 );
or \U$18424 ( \18739 , \18732 , \18737 , \18738 );
and \U$18425 ( \18740 , \3264 , \10814 );
and \U$18426 ( \18741 , \3145 , \10811 );
nor \U$18427 ( \18742 , \18740 , \18741 );
xnor \U$18428 ( \18743 , \18742 , \9759 );
and \U$18429 ( \18744 , \3889 , \10001 );
and \U$18430 ( \18745 , \3681 , \9999 );
nor \U$18431 ( \18746 , \18744 , \18745 );
xnor \U$18432 ( \18747 , \18746 , \9762 );
and \U$18433 ( \18748 , \18743 , \18747 );
and \U$18434 ( \18749 , \4016 , \9433 );
and \U$18435 ( \18750 , \4011 , \9431 );
nor \U$18436 ( \18751 , \18749 , \18750 );
xnor \U$18437 ( \18752 , \18751 , \9123 );
and \U$18438 ( \18753 , \18747 , \18752 );
and \U$18439 ( \18754 , \18743 , \18752 );
or \U$18440 ( \18755 , \18748 , \18753 , \18754 );
and \U$18441 ( \18756 , \18739 , \18755 );
and \U$18442 ( \18757 , \5776 , \7238 );
and \U$18443 ( \18758 , \5517 , \7236 );
nor \U$18444 ( \18759 , \18757 , \18758 );
xnor \U$18445 ( \18760 , \18759 , \6978 );
and \U$18446 ( \18761 , \6157 , \6744 );
and \U$18447 ( \18762 , \6148 , \6742 );
nor \U$18448 ( \18763 , \18761 , \18762 );
xnor \U$18449 ( \18764 , \18763 , \6429 );
and \U$18450 ( \18765 , \18760 , \18764 );
and \U$18451 ( \18766 , \6702 , \6235 );
and \U$18452 ( \18767 , \6500 , \6233 );
nor \U$18453 ( \18768 , \18766 , \18767 );
xnor \U$18454 ( \18769 , \18768 , \5895 );
and \U$18455 ( \18770 , \18764 , \18769 );
and \U$18456 ( \18771 , \18760 , \18769 );
or \U$18457 ( \18772 , \18765 , \18770 , \18771 );
and \U$18458 ( \18773 , \18755 , \18772 );
and \U$18459 ( \18774 , \18739 , \18772 );
or \U$18460 ( \18775 , \18756 , \18773 , \18774 );
xor \U$18461 ( \18776 , \18558 , \18562 );
xor \U$18462 ( \18777 , \18776 , \18567 );
xor \U$18463 ( \18778 , \18608 , \18612 );
xor \U$18464 ( \18779 , \18778 , \18617 );
and \U$18465 ( \18780 , \18777 , \18779 );
xor \U$18466 ( \18781 , \18589 , \18593 );
xor \U$18467 ( \18782 , \18781 , \18598 );
and \U$18468 ( \18783 , \18779 , \18782 );
and \U$18469 ( \18784 , \18777 , \18782 );
or \U$18470 ( \18785 , \18780 , \18783 , \18784 );
and \U$18471 ( \18786 , \18775 , \18785 );
and \U$18472 ( \18787 , \7177 , \5646 );
and \U$18473 ( \18788 , \7005 , \5644 );
nor \U$18474 ( \18789 , \18787 , \18788 );
xnor \U$18475 ( \18790 , \18789 , \5405 );
and \U$18476 ( \18791 , \8127 , \5180 );
and \U$18477 ( \18792 , \7703 , \5178 );
nor \U$18478 ( \18793 , \18791 , \18792 );
xnor \U$18479 ( \18794 , \18793 , \4992 );
and \U$18480 ( \18795 , \18790 , \18794 );
and \U$18481 ( \18796 , \8378 , \4806 );
and \U$18482 ( \18797 , \8373 , \4804 );
nor \U$18483 ( \18798 , \18796 , \18797 );
xnor \U$18484 ( \18799 , \18798 , \4574 );
and \U$18485 ( \18800 , \18794 , \18799 );
and \U$18486 ( \18801 , \18790 , \18799 );
or \U$18487 ( \18802 , \18795 , \18800 , \18801 );
and \U$18488 ( \18803 , \8981 , \4355 );
and \U$18489 ( \18804 , \8697 , \4353 );
nor \U$18490 ( \18805 , \18803 , \18804 );
xnor \U$18491 ( \18806 , \18805 , \4212 );
and \U$18492 ( \18807 , \9558 , \4032 );
and \U$18493 ( \18808 , \9550 , \4030 );
nor \U$18494 ( \18809 , \18807 , \18808 );
xnor \U$18495 ( \18810 , \18809 , \3786 );
and \U$18496 ( \18811 , \18806 , \18810 );
and \U$18497 ( \18812 , \10166 , \3637 );
and \U$18498 ( \18813 , \10161 , \3635 );
nor \U$18499 ( \18814 , \18812 , \18813 );
xnor \U$18500 ( \18815 , \18814 , \3450 );
and \U$18501 ( \18816 , \18810 , \18815 );
and \U$18502 ( \18817 , \18806 , \18815 );
or \U$18503 ( \18818 , \18811 , \18816 , \18817 );
and \U$18504 ( \18819 , \18802 , \18818 );
xor \U$18505 ( \18820 , \18574 , \18578 );
xor \U$18506 ( \18821 , \18820 , \18581 );
and \U$18507 ( \18822 , \18818 , \18821 );
and \U$18508 ( \18823 , \18802 , \18821 );
or \U$18509 ( \18824 , \18819 , \18822 , \18823 );
and \U$18510 ( \18825 , \18785 , \18824 );
and \U$18511 ( \18826 , \18775 , \18824 );
or \U$18512 ( \18827 , \18786 , \18825 , \18826 );
xor \U$18513 ( \18828 , \18570 , \18584 );
xor \U$18514 ( \18829 , \18828 , \18601 );
xor \U$18515 ( \18830 , \18667 , \18669 );
xor \U$18516 ( \18831 , \18830 , \18672 );
and \U$18517 ( \18832 , \18829 , \18831 );
xor \U$18518 ( \18833 , \18655 , \18657 );
xor \U$18519 ( \18834 , \18833 , \18659 );
and \U$18520 ( \18835 , \18831 , \18834 );
and \U$18521 ( \18836 , \18829 , \18834 );
or \U$18522 ( \18837 , \18832 , \18835 , \18836 );
and \U$18523 ( \18838 , \18827 , \18837 );
xor \U$18524 ( \18839 , \18686 , \18688 );
xor \U$18525 ( \18840 , \18839 , \18691 );
and \U$18526 ( \18841 , \18837 , \18840 );
and \U$18527 ( \18842 , \18827 , \18840 );
or \U$18528 ( \18843 , \18838 , \18841 , \18842 );
xor \U$18529 ( \18844 , \18665 , \18683 );
xor \U$18530 ( \18845 , \18844 , \18694 );
and \U$18531 ( \18846 , \18843 , \18845 );
xor \U$18532 ( \18847 , \18699 , \18701 );
xor \U$18533 ( \18848 , \18847 , \18703 );
and \U$18534 ( \18849 , \18845 , \18848 );
and \U$18535 ( \18850 , \18843 , \18848 );
or \U$18536 ( \18851 , \18846 , \18849 , \18850 );
xor \U$18537 ( \18852 , \18486 , \18504 );
xor \U$18538 ( \18853 , \18852 , \18510 );
and \U$18539 ( \18854 , \18851 , \18853 );
xor \U$18540 ( \18855 , \18697 , \18706 );
xor \U$18541 ( \18856 , \18855 , \18709 );
and \U$18542 ( \18857 , \18853 , \18856 );
and \U$18543 ( \18858 , \18851 , \18856 );
or \U$18544 ( \18859 , \18854 , \18857 , \18858 );
and \U$18545 ( \18860 , \18723 , \18859 );
xor \U$18546 ( \18861 , \18723 , \18859 );
xor \U$18547 ( \18862 , \18851 , \18853 );
xor \U$18548 ( \18863 , \18862 , \18856 );
and \U$18549 ( \18864 , \4272 , \9433 );
and \U$18550 ( \18865 , \4016 , \9431 );
nor \U$18551 ( \18866 , \18864 , \18865 );
xnor \U$18552 ( \18867 , \18866 , \9123 );
and \U$18553 ( \18868 , \4771 , \8896 );
and \U$18554 ( \18869 , \4469 , \8894 );
nor \U$18555 ( \18870 , \18868 , \18869 );
xnor \U$18556 ( \18871 , \18870 , \8525 );
and \U$18557 ( \18872 , \18867 , \18871 );
and \U$18558 ( \18873 , \5248 , \8334 );
and \U$18559 ( \18874 , \4779 , \8332 );
nor \U$18560 ( \18875 , \18873 , \18874 );
xnor \U$18561 ( \18876 , \18875 , \8016 );
and \U$18562 ( \18877 , \18871 , \18876 );
and \U$18563 ( \18878 , \18867 , \18876 );
or \U$18564 ( \18879 , \18872 , \18877 , \18878 );
and \U$18565 ( \18880 , \5517 , \7767 );
and \U$18566 ( \18881 , \5253 , \7765 );
nor \U$18567 ( \18882 , \18880 , \18881 );
xnor \U$18568 ( \18883 , \18882 , \7518 );
and \U$18569 ( \18884 , \6148 , \7238 );
and \U$18570 ( \18885 , \5776 , \7236 );
nor \U$18571 ( \18886 , \18884 , \18885 );
xnor \U$18572 ( \18887 , \18886 , \6978 );
and \U$18573 ( \18888 , \18883 , \18887 );
and \U$18574 ( \18889 , \6500 , \6744 );
and \U$18575 ( \18890 , \6157 , \6742 );
nor \U$18576 ( \18891 , \18889 , \18890 );
xnor \U$18577 ( \18892 , \18891 , \6429 );
and \U$18578 ( \18893 , \18887 , \18892 );
and \U$18579 ( \18894 , \18883 , \18892 );
or \U$18580 ( \18895 , \18888 , \18893 , \18894 );
and \U$18581 ( \18896 , \18879 , \18895 );
and \U$18582 ( \18897 , \3681 , \10814 );
and \U$18583 ( \18898 , \3264 , \10811 );
nor \U$18584 ( \18899 , \18897 , \18898 );
xnor \U$18585 ( \18900 , \18899 , \9759 );
and \U$18586 ( \18901 , \4011 , \10001 );
and \U$18587 ( \18902 , \3889 , \9999 );
nor \U$18588 ( \18903 , \18901 , \18902 );
xnor \U$18589 ( \18904 , \18903 , \9762 );
and \U$18590 ( \18905 , \18900 , \18904 );
and \U$18591 ( \18906 , \18904 , \3119 );
and \U$18592 ( \18907 , \18900 , \3119 );
or \U$18593 ( \18908 , \18905 , \18906 , \18907 );
and \U$18594 ( \18909 , \18895 , \18908 );
and \U$18595 ( \18910 , \18879 , \18908 );
or \U$18596 ( \18911 , \18896 , \18909 , \18910 );
and \U$18597 ( \18912 , \8697 , \4806 );
and \U$18598 ( \18913 , \8378 , \4804 );
nor \U$18599 ( \18914 , \18912 , \18913 );
xnor \U$18600 ( \18915 , \18914 , \4574 );
and \U$18601 ( \18916 , \9550 , \4355 );
and \U$18602 ( \18917 , \8981 , \4353 );
nor \U$18603 ( \18918 , \18916 , \18917 );
xnor \U$18604 ( \18919 , \18918 , \4212 );
and \U$18605 ( \18920 , \18915 , \18919 );
and \U$18606 ( \18921 , \10161 , \4032 );
and \U$18607 ( \18922 , \9558 , \4030 );
nor \U$18608 ( \18923 , \18921 , \18922 );
xnor \U$18609 ( \18924 , \18923 , \3786 );
and \U$18610 ( \18925 , \18919 , \18924 );
and \U$18611 ( \18926 , \18915 , \18924 );
or \U$18612 ( \18927 , \18920 , \18925 , \18926 );
and \U$18613 ( \18928 , \7005 , \6235 );
and \U$18614 ( \18929 , \6702 , \6233 );
nor \U$18615 ( \18930 , \18928 , \18929 );
xnor \U$18616 ( \18931 , \18930 , \5895 );
and \U$18617 ( \18932 , \7703 , \5646 );
and \U$18618 ( \18933 , \7177 , \5644 );
nor \U$18619 ( \18934 , \18932 , \18933 );
xnor \U$18620 ( \18935 , \18934 , \5405 );
and \U$18621 ( \18936 , \18931 , \18935 );
and \U$18622 ( \18937 , \8373 , \5180 );
and \U$18623 ( \18938 , \8127 , \5178 );
nor \U$18624 ( \18939 , \18937 , \18938 );
xnor \U$18625 ( \18940 , \18939 , \4992 );
and \U$18626 ( \18941 , \18935 , \18940 );
and \U$18627 ( \18942 , \18931 , \18940 );
or \U$18628 ( \18943 , \18936 , \18941 , \18942 );
and \U$18629 ( \18944 , \18927 , \18943 );
and \U$18630 ( \18945 , \10967 , \3324 );
and \U$18631 ( \18946 , \10347 , \3322 );
nor \U$18632 ( \18947 , \18945 , \18946 );
xnor \U$18633 ( \18948 , \18947 , \3119 );
and \U$18634 ( \18949 , \18943 , \18948 );
and \U$18635 ( \18950 , \18927 , \18948 );
or \U$18636 ( \18951 , \18944 , \18949 , \18950 );
and \U$18637 ( \18952 , \18911 , \18951 );
xor \U$18638 ( \18953 , \18790 , \18794 );
xor \U$18639 ( \18954 , \18953 , \18799 );
xor \U$18640 ( \18955 , \18806 , \18810 );
xor \U$18641 ( \18956 , \18955 , \18815 );
and \U$18642 ( \18957 , \18954 , \18956 );
xor \U$18643 ( \18958 , \18760 , \18764 );
xor \U$18644 ( \18959 , \18958 , \18769 );
and \U$18645 ( \18960 , \18956 , \18959 );
and \U$18646 ( \18961 , \18954 , \18959 );
or \U$18647 ( \18962 , \18957 , \18960 , \18961 );
and \U$18648 ( \18963 , \18951 , \18962 );
and \U$18649 ( \18964 , \18911 , \18962 );
or \U$18650 ( \18965 , \18952 , \18963 , \18964 );
xor \U$18651 ( \18966 , \18624 , \18628 );
xor \U$18652 ( \18967 , \18966 , \2769 );
xor \U$18653 ( \18968 , \18637 , \18641 );
xor \U$18654 ( \18969 , \18968 , \18646 );
and \U$18655 ( \18970 , \18967 , \18969 );
xor \U$18656 ( \18971 , \18777 , \18779 );
xor \U$18657 ( \18972 , \18971 , \18782 );
and \U$18658 ( \18973 , \18969 , \18972 );
and \U$18659 ( \18974 , \18967 , \18972 );
or \U$18660 ( \18975 , \18970 , \18973 , \18974 );
and \U$18661 ( \18976 , \18965 , \18975 );
xor \U$18662 ( \18977 , \18739 , \18755 );
xor \U$18663 ( \18978 , \18977 , \18772 );
xor \U$18664 ( \18979 , \18802 , \18818 );
xor \U$18665 ( \18980 , \18979 , \18821 );
and \U$18666 ( \18981 , \18978 , \18980 );
and \U$18667 ( \18982 , \18975 , \18981 );
and \U$18668 ( \18983 , \18965 , \18981 );
or \U$18669 ( \18984 , \18976 , \18982 , \18983 );
xor \U$18670 ( \18985 , \18620 , \18632 );
xor \U$18671 ( \18986 , \18985 , \18649 );
xor \U$18672 ( \18987 , \18775 , \18785 );
xor \U$18673 ( \18988 , \18987 , \18824 );
and \U$18674 ( \18989 , \18986 , \18988 );
xor \U$18675 ( \18990 , \18829 , \18831 );
xor \U$18676 ( \18991 , \18990 , \18834 );
and \U$18677 ( \18992 , \18988 , \18991 );
and \U$18678 ( \18993 , \18986 , \18991 );
or \U$18679 ( \18994 , \18989 , \18992 , \18993 );
and \U$18680 ( \18995 , \18984 , \18994 );
xor \U$18681 ( \18996 , \18675 , \18677 );
xor \U$18682 ( \18997 , \18996 , \18680 );
and \U$18683 ( \18998 , \18994 , \18997 );
and \U$18684 ( \18999 , \18984 , \18997 );
or \U$18685 ( \19000 , \18995 , \18998 , \18999 );
xor \U$18686 ( \19001 , \18604 , \18652 );
xor \U$18687 ( \19002 , \19001 , \18662 );
xor \U$18688 ( \19003 , \18827 , \18837 );
xor \U$18689 ( \19004 , \19003 , \18840 );
and \U$18690 ( \19005 , \19002 , \19004 );
and \U$18691 ( \19006 , \19000 , \19005 );
xor \U$18692 ( \19007 , \18843 , \18845 );
xor \U$18693 ( \19008 , \19007 , \18848 );
and \U$18694 ( \19009 , \19005 , \19008 );
and \U$18695 ( \19010 , \19000 , \19008 );
or \U$18696 ( \19011 , \19006 , \19009 , \19010 );
and \U$18697 ( \19012 , \18863 , \19011 );
xor \U$18698 ( \19013 , \18863 , \19011 );
xor \U$18699 ( \19014 , \19000 , \19005 );
xor \U$18700 ( \19015 , \19014 , \19008 );
and \U$18701 ( \19016 , \6157 , \7238 );
and \U$18702 ( \19017 , \6148 , \7236 );
nor \U$18703 ( \19018 , \19016 , \19017 );
xnor \U$18704 ( \19019 , \19018 , \6978 );
and \U$18705 ( \19020 , \6702 , \6744 );
and \U$18706 ( \19021 , \6500 , \6742 );
nor \U$18707 ( \19022 , \19020 , \19021 );
xnor \U$18708 ( \19023 , \19022 , \6429 );
and \U$18709 ( \19024 , \19019 , \19023 );
and \U$18710 ( \19025 , \7177 , \6235 );
and \U$18711 ( \19026 , \7005 , \6233 );
nor \U$18712 ( \19027 , \19025 , \19026 );
xnor \U$18713 ( \19028 , \19027 , \5895 );
and \U$18714 ( \19029 , \19023 , \19028 );
and \U$18715 ( \19030 , \19019 , \19028 );
or \U$18716 ( \19031 , \19024 , \19029 , \19030 );
and \U$18717 ( \19032 , \4779 , \8896 );
and \U$18718 ( \19033 , \4771 , \8894 );
nor \U$18719 ( \19034 , \19032 , \19033 );
xnor \U$18720 ( \19035 , \19034 , \8525 );
and \U$18721 ( \19036 , \5253 , \8334 );
and \U$18722 ( \19037 , \5248 , \8332 );
nor \U$18723 ( \19038 , \19036 , \19037 );
xnor \U$18724 ( \19039 , \19038 , \8016 );
and \U$18725 ( \19040 , \19035 , \19039 );
and \U$18726 ( \19041 , \5776 , \7767 );
and \U$18727 ( \19042 , \5517 , \7765 );
nor \U$18728 ( \19043 , \19041 , \19042 );
xnor \U$18729 ( \19044 , \19043 , \7518 );
and \U$18730 ( \19045 , \19039 , \19044 );
and \U$18731 ( \19046 , \19035 , \19044 );
or \U$18732 ( \19047 , \19040 , \19045 , \19046 );
and \U$18733 ( \19048 , \19031 , \19047 );
and \U$18734 ( \19049 , \3889 , \10814 );
and \U$18735 ( \19050 , \3681 , \10811 );
nor \U$18736 ( \19051 , \19049 , \19050 );
xnor \U$18737 ( \19052 , \19051 , \9759 );
and \U$18738 ( \19053 , \4016 , \10001 );
and \U$18739 ( \19054 , \4011 , \9999 );
nor \U$18740 ( \19055 , \19053 , \19054 );
xnor \U$18741 ( \19056 , \19055 , \9762 );
and \U$18742 ( \19057 , \19052 , \19056 );
and \U$18743 ( \19058 , \4469 , \9433 );
and \U$18744 ( \19059 , \4272 , \9431 );
nor \U$18745 ( \19060 , \19058 , \19059 );
xnor \U$18746 ( \19061 , \19060 , \9123 );
and \U$18747 ( \19062 , \19056 , \19061 );
and \U$18748 ( \19063 , \19052 , \19061 );
or \U$18749 ( \19064 , \19057 , \19062 , \19063 );
and \U$18750 ( \19065 , \19047 , \19064 );
and \U$18751 ( \19066 , \19031 , \19064 );
or \U$18752 ( \19067 , \19048 , \19065 , \19066 );
and \U$18753 ( \19068 , \9558 , \4355 );
and \U$18754 ( \19069 , \9550 , \4353 );
nor \U$18755 ( \19070 , \19068 , \19069 );
xnor \U$18756 ( \19071 , \19070 , \4212 );
and \U$18757 ( \19072 , \10166 , \4032 );
and \U$18758 ( \19073 , \10161 , \4030 );
nor \U$18759 ( \19074 , \19072 , \19073 );
xnor \U$18760 ( \19075 , \19074 , \3786 );
and \U$18761 ( \19076 , \19071 , \19075 );
and \U$18762 ( \19077 , \10967 , \3637 );
and \U$18763 ( \19078 , \10347 , \3635 );
nor \U$18764 ( \19079 , \19077 , \19078 );
xnor \U$18765 ( \19080 , \19079 , \3450 );
and \U$18766 ( \19081 , \19075 , \19080 );
and \U$18767 ( \19082 , \19071 , \19080 );
or \U$18768 ( \19083 , \19076 , \19081 , \19082 );
and \U$18769 ( \19084 , \8127 , \5646 );
and \U$18770 ( \19085 , \7703 , \5644 );
nor \U$18771 ( \19086 , \19084 , \19085 );
xnor \U$18772 ( \19087 , \19086 , \5405 );
and \U$18773 ( \19088 , \8378 , \5180 );
and \U$18774 ( \19089 , \8373 , \5178 );
nor \U$18775 ( \19090 , \19088 , \19089 );
xnor \U$18776 ( \19091 , \19090 , \4992 );
and \U$18777 ( \19092 , \19087 , \19091 );
and \U$18778 ( \19093 , \8981 , \4806 );
and \U$18779 ( \19094 , \8697 , \4804 );
nor \U$18780 ( \19095 , \19093 , \19094 );
xnor \U$18781 ( \19096 , \19095 , \4574 );
and \U$18782 ( \19097 , \19091 , \19096 );
and \U$18783 ( \19098 , \19087 , \19096 );
or \U$18784 ( \19099 , \19092 , \19097 , \19098 );
and \U$18785 ( \19100 , \19083 , \19099 );
and \U$18786 ( \19101 , \10347 , \3637 );
and \U$18787 ( \19102 , \10166 , \3635 );
nor \U$18788 ( \19103 , \19101 , \19102 );
xnor \U$18789 ( \19104 , \19103 , \3450 );
and \U$18790 ( \19105 , \19099 , \19104 );
and \U$18791 ( \19106 , \19083 , \19104 );
or \U$18792 ( \19107 , \19100 , \19105 , \19106 );
and \U$18793 ( \19108 , \19067 , \19107 );
nand \U$18794 ( \19109 , \10967 , \3322 );
xnor \U$18795 ( \19110 , \19109 , \3119 );
xor \U$18796 ( \19111 , \18915 , \18919 );
xor \U$18797 ( \19112 , \19111 , \18924 );
and \U$18798 ( \19113 , \19110 , \19112 );
xor \U$18799 ( \19114 , \18931 , \18935 );
xor \U$18800 ( \19115 , \19114 , \18940 );
and \U$18801 ( \19116 , \19112 , \19115 );
and \U$18802 ( \19117 , \19110 , \19115 );
or \U$18803 ( \19118 , \19113 , \19116 , \19117 );
and \U$18804 ( \19119 , \19107 , \19118 );
and \U$18805 ( \19120 , \19067 , \19118 );
or \U$18806 ( \19121 , \19108 , \19119 , \19120 );
xor \U$18807 ( \19122 , \18867 , \18871 );
xor \U$18808 ( \19123 , \19122 , \18876 );
xor \U$18809 ( \19124 , \18883 , \18887 );
xor \U$18810 ( \19125 , \19124 , \18892 );
and \U$18811 ( \19126 , \19123 , \19125 );
xor \U$18812 ( \19127 , \18900 , \18904 );
xor \U$18813 ( \19128 , \19127 , \3119 );
and \U$18814 ( \19129 , \19125 , \19128 );
and \U$18815 ( \19130 , \19123 , \19128 );
or \U$18816 ( \19131 , \19126 , \19129 , \19130 );
xor \U$18817 ( \19132 , \18727 , \18731 );
xor \U$18818 ( \19133 , \19132 , \18736 );
and \U$18819 ( \19134 , \19131 , \19133 );
xor \U$18820 ( \19135 , \18743 , \18747 );
xor \U$18821 ( \19136 , \19135 , \18752 );
and \U$18822 ( \19137 , \19133 , \19136 );
and \U$18823 ( \19138 , \19131 , \19136 );
or \U$18824 ( \19139 , \19134 , \19137 , \19138 );
and \U$18825 ( \19140 , \19121 , \19139 );
xor \U$18826 ( \19141 , \18879 , \18895 );
xor \U$18827 ( \19142 , \19141 , \18908 );
xor \U$18828 ( \19143 , \18927 , \18943 );
xor \U$18829 ( \19144 , \19143 , \18948 );
and \U$18830 ( \19145 , \19142 , \19144 );
xor \U$18831 ( \19146 , \18954 , \18956 );
xor \U$18832 ( \19147 , \19146 , \18959 );
and \U$18833 ( \19148 , \19144 , \19147 );
and \U$18834 ( \19149 , \19142 , \19147 );
or \U$18835 ( \19150 , \19145 , \19148 , \19149 );
and \U$18836 ( \19151 , \19139 , \19150 );
and \U$18837 ( \19152 , \19121 , \19150 );
or \U$18838 ( \19153 , \19140 , \19151 , \19152 );
xor \U$18839 ( \19154 , \18911 , \18951 );
xor \U$18840 ( \19155 , \19154 , \18962 );
xor \U$18841 ( \19156 , \18967 , \18969 );
xor \U$18842 ( \19157 , \19156 , \18972 );
and \U$18843 ( \19158 , \19155 , \19157 );
xor \U$18844 ( \19159 , \18978 , \18980 );
and \U$18845 ( \19160 , \19157 , \19159 );
and \U$18846 ( \19161 , \19155 , \19159 );
or \U$18847 ( \19162 , \19158 , \19160 , \19161 );
and \U$18848 ( \19163 , \19153 , \19162 );
xor \U$18849 ( \19164 , \18986 , \18988 );
xor \U$18850 ( \19165 , \19164 , \18991 );
and \U$18851 ( \19166 , \19162 , \19165 );
and \U$18852 ( \19167 , \19153 , \19165 );
or \U$18853 ( \19168 , \19163 , \19166 , \19167 );
xor \U$18854 ( \19169 , \18984 , \18994 );
xor \U$18855 ( \19170 , \19169 , \18997 );
and \U$18856 ( \19171 , \19168 , \19170 );
xor \U$18857 ( \19172 , \19002 , \19004 );
and \U$18858 ( \19173 , \19170 , \19172 );
and \U$18859 ( \19174 , \19168 , \19172 );
or \U$18860 ( \19175 , \19171 , \19173 , \19174 );
and \U$18861 ( \19176 , \19015 , \19175 );
xor \U$18862 ( \19177 , \19015 , \19175 );
xor \U$18863 ( \19178 , \19168 , \19170 );
xor \U$18864 ( \19179 , \19178 , \19172 );
and \U$18865 ( \19180 , \6148 , \7767 );
and \U$18866 ( \19181 , \5776 , \7765 );
nor \U$18867 ( \19182 , \19180 , \19181 );
xnor \U$18868 ( \19183 , \19182 , \7518 );
and \U$18869 ( \19184 , \6500 , \7238 );
and \U$18870 ( \19185 , \6157 , \7236 );
nor \U$18871 ( \19186 , \19184 , \19185 );
xnor \U$18872 ( \19187 , \19186 , \6978 );
and \U$18873 ( \19188 , \19183 , \19187 );
and \U$18874 ( \19189 , \7005 , \6744 );
and \U$18875 ( \19190 , \6702 , \6742 );
nor \U$18876 ( \19191 , \19189 , \19190 );
xnor \U$18877 ( \19192 , \19191 , \6429 );
and \U$18878 ( \19193 , \19187 , \19192 );
and \U$18879 ( \19194 , \19183 , \19192 );
or \U$18880 ( \19195 , \19188 , \19193 , \19194 );
and \U$18881 ( \19196 , \4771 , \9433 );
and \U$18882 ( \19197 , \4469 , \9431 );
nor \U$18883 ( \19198 , \19196 , \19197 );
xnor \U$18884 ( \19199 , \19198 , \9123 );
and \U$18885 ( \19200 , \5248 , \8896 );
and \U$18886 ( \19201 , \4779 , \8894 );
nor \U$18887 ( \19202 , \19200 , \19201 );
xnor \U$18888 ( \19203 , \19202 , \8525 );
and \U$18889 ( \19204 , \19199 , \19203 );
and \U$18890 ( \19205 , \5517 , \8334 );
and \U$18891 ( \19206 , \5253 , \8332 );
nor \U$18892 ( \19207 , \19205 , \19206 );
xnor \U$18893 ( \19208 , \19207 , \8016 );
and \U$18894 ( \19209 , \19203 , \19208 );
and \U$18895 ( \19210 , \19199 , \19208 );
or \U$18896 ( \19211 , \19204 , \19209 , \19210 );
and \U$18897 ( \19212 , \19195 , \19211 );
and \U$18898 ( \19213 , \4011 , \10814 );
and \U$18899 ( \19214 , \3889 , \10811 );
nor \U$18900 ( \19215 , \19213 , \19214 );
xnor \U$18901 ( \19216 , \19215 , \9759 );
and \U$18902 ( \19217 , \4272 , \10001 );
and \U$18903 ( \19218 , \4016 , \9999 );
nor \U$18904 ( \19219 , \19217 , \19218 );
xnor \U$18905 ( \19220 , \19219 , \9762 );
and \U$18906 ( \19221 , \19216 , \19220 );
and \U$18907 ( \19222 , \19220 , \3450 );
and \U$18908 ( \19223 , \19216 , \3450 );
or \U$18909 ( \19224 , \19221 , \19222 , \19223 );
and \U$18910 ( \19225 , \19211 , \19224 );
and \U$18911 ( \19226 , \19195 , \19224 );
or \U$18912 ( \19227 , \19212 , \19225 , \19226 );
and \U$18913 ( \19228 , \7703 , \6235 );
and \U$18914 ( \19229 , \7177 , \6233 );
nor \U$18915 ( \19230 , \19228 , \19229 );
xnor \U$18916 ( \19231 , \19230 , \5895 );
and \U$18917 ( \19232 , \8373 , \5646 );
and \U$18918 ( \19233 , \8127 , \5644 );
nor \U$18919 ( \19234 , \19232 , \19233 );
xnor \U$18920 ( \19235 , \19234 , \5405 );
and \U$18921 ( \19236 , \19231 , \19235 );
and \U$18922 ( \19237 , \8697 , \5180 );
and \U$18923 ( \19238 , \8378 , \5178 );
nor \U$18924 ( \19239 , \19237 , \19238 );
xnor \U$18925 ( \19240 , \19239 , \4992 );
and \U$18926 ( \19241 , \19235 , \19240 );
and \U$18927 ( \19242 , \19231 , \19240 );
or \U$18928 ( \19243 , \19236 , \19241 , \19242 );
and \U$18929 ( \19244 , \9550 , \4806 );
and \U$18930 ( \19245 , \8981 , \4804 );
nor \U$18931 ( \19246 , \19244 , \19245 );
xnor \U$18932 ( \19247 , \19246 , \4574 );
and \U$18933 ( \19248 , \10161 , \4355 );
and \U$18934 ( \19249 , \9558 , \4353 );
nor \U$18935 ( \19250 , \19248 , \19249 );
xnor \U$18936 ( \19251 , \19250 , \4212 );
and \U$18937 ( \19252 , \19247 , \19251 );
and \U$18938 ( \19253 , \10347 , \4032 );
and \U$18939 ( \19254 , \10166 , \4030 );
nor \U$18940 ( \19255 , \19253 , \19254 );
xnor \U$18941 ( \19256 , \19255 , \3786 );
and \U$18942 ( \19257 , \19251 , \19256 );
and \U$18943 ( \19258 , \19247 , \19256 );
or \U$18944 ( \19259 , \19252 , \19257 , \19258 );
and \U$18945 ( \19260 , \19243 , \19259 );
xor \U$18946 ( \19261 , \19071 , \19075 );
xor \U$18947 ( \19262 , \19261 , \19080 );
and \U$18948 ( \19263 , \19259 , \19262 );
and \U$18949 ( \19264 , \19243 , \19262 );
or \U$18950 ( \19265 , \19260 , \19263 , \19264 );
and \U$18951 ( \19266 , \19227 , \19265 );
xor \U$18952 ( \19267 , \19019 , \19023 );
xor \U$18953 ( \19268 , \19267 , \19028 );
xor \U$18954 ( \19269 , \19035 , \19039 );
xor \U$18955 ( \19270 , \19269 , \19044 );
and \U$18956 ( \19271 , \19268 , \19270 );
xor \U$18957 ( \19272 , \19087 , \19091 );
xor \U$18958 ( \19273 , \19272 , \19096 );
and \U$18959 ( \19274 , \19270 , \19273 );
and \U$18960 ( \19275 , \19268 , \19273 );
or \U$18961 ( \19276 , \19271 , \19274 , \19275 );
and \U$18962 ( \19277 , \19265 , \19276 );
and \U$18963 ( \19278 , \19227 , \19276 );
or \U$18964 ( \19279 , \19266 , \19277 , \19278 );
xor \U$18965 ( \19280 , \19083 , \19099 );
xor \U$18966 ( \19281 , \19280 , \19104 );
xor \U$18967 ( \19282 , \19123 , \19125 );
xor \U$18968 ( \19283 , \19282 , \19128 );
and \U$18969 ( \19284 , \19281 , \19283 );
xor \U$18970 ( \19285 , \19110 , \19112 );
xor \U$18971 ( \19286 , \19285 , \19115 );
and \U$18972 ( \19287 , \19283 , \19286 );
and \U$18973 ( \19288 , \19281 , \19286 );
or \U$18974 ( \19289 , \19284 , \19287 , \19288 );
and \U$18975 ( \19290 , \19279 , \19289 );
xor \U$18976 ( \19291 , \19142 , \19144 );
xor \U$18977 ( \19292 , \19291 , \19147 );
and \U$18978 ( \19293 , \19289 , \19292 );
and \U$18979 ( \19294 , \19279 , \19292 );
or \U$18980 ( \19295 , \19290 , \19293 , \19294 );
xor \U$18981 ( \19296 , \19067 , \19107 );
xor \U$18982 ( \19297 , \19296 , \19118 );
xor \U$18983 ( \19298 , \19131 , \19133 );
xor \U$18984 ( \19299 , \19298 , \19136 );
and \U$18985 ( \19300 , \19297 , \19299 );
and \U$18986 ( \19301 , \19295 , \19300 );
xor \U$18987 ( \19302 , \19155 , \19157 );
xor \U$18988 ( \19303 , \19302 , \19159 );
and \U$18989 ( \19304 , \19300 , \19303 );
and \U$18990 ( \19305 , \19295 , \19303 );
or \U$18991 ( \19306 , \19301 , \19304 , \19305 );
xor \U$18992 ( \19307 , \18965 , \18975 );
xor \U$18993 ( \19308 , \19307 , \18981 );
and \U$18994 ( \19309 , \19306 , \19308 );
xor \U$18995 ( \19310 , \19153 , \19162 );
xor \U$18996 ( \19311 , \19310 , \19165 );
and \U$18997 ( \19312 , \19308 , \19311 );
and \U$18998 ( \19313 , \19306 , \19311 );
or \U$18999 ( \19314 , \19309 , \19312 , \19313 );
and \U$19000 ( \19315 , \19179 , \19314 );
xor \U$19001 ( \19316 , \19179 , \19314 );
xor \U$19002 ( \19317 , \19306 , \19308 );
xor \U$19003 ( \19318 , \19317 , \19311 );
and \U$19004 ( \19319 , \4016 , \10814 );
and \U$19005 ( \19320 , \4011 , \10811 );
nor \U$19006 ( \19321 , \19319 , \19320 );
xnor \U$19007 ( \19322 , \19321 , \9759 );
and \U$19008 ( \19323 , \4469 , \10001 );
and \U$19009 ( \19324 , \4272 , \9999 );
nor \U$19010 ( \19325 , \19323 , \19324 );
xnor \U$19011 ( \19326 , \19325 , \9762 );
and \U$19012 ( \19327 , \19322 , \19326 );
and \U$19013 ( \19328 , \4779 , \9433 );
and \U$19014 ( \19329 , \4771 , \9431 );
nor \U$19015 ( \19330 , \19328 , \19329 );
xnor \U$19016 ( \19331 , \19330 , \9123 );
and \U$19017 ( \19332 , \19326 , \19331 );
and \U$19018 ( \19333 , \19322 , \19331 );
or \U$19019 ( \19334 , \19327 , \19332 , \19333 );
and \U$19020 ( \19335 , \6702 , \7238 );
and \U$19021 ( \19336 , \6500 , \7236 );
nor \U$19022 ( \19337 , \19335 , \19336 );
xnor \U$19023 ( \19338 , \19337 , \6978 );
and \U$19024 ( \19339 , \7177 , \6744 );
and \U$19025 ( \19340 , \7005 , \6742 );
nor \U$19026 ( \19341 , \19339 , \19340 );
xnor \U$19027 ( \19342 , \19341 , \6429 );
and \U$19028 ( \19343 , \19338 , \19342 );
and \U$19029 ( \19344 , \8127 , \6235 );
and \U$19030 ( \19345 , \7703 , \6233 );
nor \U$19031 ( \19346 , \19344 , \19345 );
xnor \U$19032 ( \19347 , \19346 , \5895 );
and \U$19033 ( \19348 , \19342 , \19347 );
and \U$19034 ( \19349 , \19338 , \19347 );
or \U$19035 ( \19350 , \19343 , \19348 , \19349 );
and \U$19036 ( \19351 , \19334 , \19350 );
and \U$19037 ( \19352 , \5253 , \8896 );
and \U$19038 ( \19353 , \5248 , \8894 );
nor \U$19039 ( \19354 , \19352 , \19353 );
xnor \U$19040 ( \19355 , \19354 , \8525 );
and \U$19041 ( \19356 , \5776 , \8334 );
and \U$19042 ( \19357 , \5517 , \8332 );
nor \U$19043 ( \19358 , \19356 , \19357 );
xnor \U$19044 ( \19359 , \19358 , \8016 );
and \U$19045 ( \19360 , \19355 , \19359 );
and \U$19046 ( \19361 , \6157 , \7767 );
and \U$19047 ( \19362 , \6148 , \7765 );
nor \U$19048 ( \19363 , \19361 , \19362 );
xnor \U$19049 ( \19364 , \19363 , \7518 );
and \U$19050 ( \19365 , \19359 , \19364 );
and \U$19051 ( \19366 , \19355 , \19364 );
or \U$19052 ( \19367 , \19360 , \19365 , \19366 );
and \U$19053 ( \19368 , \19350 , \19367 );
and \U$19054 ( \19369 , \19334 , \19367 );
or \U$19055 ( \19370 , \19351 , \19368 , \19369 );
xor \U$19056 ( \19371 , \19183 , \19187 );
xor \U$19057 ( \19372 , \19371 , \19192 );
xor \U$19058 ( \19373 , \19199 , \19203 );
xor \U$19059 ( \19374 , \19373 , \19208 );
and \U$19060 ( \19375 , \19372 , \19374 );
xor \U$19061 ( \19376 , \19231 , \19235 );
xor \U$19062 ( \19377 , \19376 , \19240 );
and \U$19063 ( \19378 , \19374 , \19377 );
and \U$19064 ( \19379 , \19372 , \19377 );
or \U$19065 ( \19380 , \19375 , \19378 , \19379 );
and \U$19066 ( \19381 , \19370 , \19380 );
and \U$19067 ( \19382 , \8378 , \5646 );
and \U$19068 ( \19383 , \8373 , \5644 );
nor \U$19069 ( \19384 , \19382 , \19383 );
xnor \U$19070 ( \19385 , \19384 , \5405 );
and \U$19071 ( \19386 , \8981 , \5180 );
and \U$19072 ( \19387 , \8697 , \5178 );
nor \U$19073 ( \19388 , \19386 , \19387 );
xnor \U$19074 ( \19389 , \19388 , \4992 );
and \U$19075 ( \19390 , \19385 , \19389 );
and \U$19076 ( \19391 , \9558 , \4806 );
and \U$19077 ( \19392 , \9550 , \4804 );
nor \U$19078 ( \19393 , \19391 , \19392 );
xnor \U$19079 ( \19394 , \19393 , \4574 );
and \U$19080 ( \19395 , \19389 , \19394 );
and \U$19081 ( \19396 , \19385 , \19394 );
or \U$19082 ( \19397 , \19390 , \19395 , \19396 );
nand \U$19083 ( \19398 , \10967 , \3635 );
xnor \U$19084 ( \19399 , \19398 , \3450 );
and \U$19085 ( \19400 , \19397 , \19399 );
xor \U$19086 ( \19401 , \19247 , \19251 );
xor \U$19087 ( \19402 , \19401 , \19256 );
and \U$19088 ( \19403 , \19399 , \19402 );
and \U$19089 ( \19404 , \19397 , \19402 );
or \U$19090 ( \19405 , \19400 , \19403 , \19404 );
and \U$19091 ( \19406 , \19380 , \19405 );
and \U$19092 ( \19407 , \19370 , \19405 );
or \U$19093 ( \19408 , \19381 , \19406 , \19407 );
xor \U$19094 ( \19409 , \19052 , \19056 );
xor \U$19095 ( \19410 , \19409 , \19061 );
xor \U$19096 ( \19411 , \19243 , \19259 );
xor \U$19097 ( \19412 , \19411 , \19262 );
and \U$19098 ( \19413 , \19410 , \19412 );
xor \U$19099 ( \19414 , \19268 , \19270 );
xor \U$19100 ( \19415 , \19414 , \19273 );
and \U$19101 ( \19416 , \19412 , \19415 );
and \U$19102 ( \19417 , \19410 , \19415 );
or \U$19103 ( \19418 , \19413 , \19416 , \19417 );
and \U$19104 ( \19419 , \19408 , \19418 );
xor \U$19105 ( \19420 , \19031 , \19047 );
xor \U$19106 ( \19421 , \19420 , \19064 );
and \U$19107 ( \19422 , \19418 , \19421 );
and \U$19108 ( \19423 , \19408 , \19421 );
or \U$19109 ( \19424 , \19419 , \19422 , \19423 );
xor \U$19110 ( \19425 , \19279 , \19289 );
xor \U$19111 ( \19426 , \19425 , \19292 );
and \U$19112 ( \19427 , \19424 , \19426 );
xor \U$19113 ( \19428 , \19297 , \19299 );
and \U$19114 ( \19429 , \19426 , \19428 );
and \U$19115 ( \19430 , \19424 , \19428 );
or \U$19116 ( \19431 , \19427 , \19429 , \19430 );
xor \U$19117 ( \19432 , \19121 , \19139 );
xor \U$19118 ( \19433 , \19432 , \19150 );
and \U$19119 ( \19434 , \19431 , \19433 );
xor \U$19120 ( \19435 , \19295 , \19300 );
xor \U$19121 ( \19436 , \19435 , \19303 );
and \U$19122 ( \19437 , \19433 , \19436 );
and \U$19123 ( \19438 , \19431 , \19436 );
or \U$19124 ( \19439 , \19434 , \19437 , \19438 );
and \U$19125 ( \19440 , \19318 , \19439 );
xor \U$19126 ( \19441 , \19318 , \19439 );
xor \U$19127 ( \19442 , \19431 , \19433 );
xor \U$19128 ( \19443 , \19442 , \19436 );
and \U$19129 ( \19444 , \8373 , \6235 );
and \U$19130 ( \19445 , \8127 , \6233 );
nor \U$19131 ( \19446 , \19444 , \19445 );
xnor \U$19132 ( \19447 , \19446 , \5895 );
and \U$19133 ( \19448 , \8697 , \5646 );
and \U$19134 ( \19449 , \8378 , \5644 );
nor \U$19135 ( \19450 , \19448 , \19449 );
xnor \U$19136 ( \19451 , \19450 , \5405 );
and \U$19137 ( \19452 , \19447 , \19451 );
and \U$19138 ( \19453 , \9550 , \5180 );
and \U$19139 ( \19454 , \8981 , \5178 );
nor \U$19140 ( \19455 , \19453 , \19454 );
xnor \U$19141 ( \19456 , \19455 , \4992 );
and \U$19142 ( \19457 , \19451 , \19456 );
and \U$19143 ( \19458 , \19447 , \19456 );
or \U$19144 ( \19459 , \19452 , \19457 , \19458 );
and \U$19145 ( \19460 , \10161 , \4806 );
and \U$19146 ( \19461 , \9558 , \4804 );
nor \U$19147 ( \19462 , \19460 , \19461 );
xnor \U$19148 ( \19463 , \19462 , \4574 );
and \U$19149 ( \19464 , \10347 , \4355 );
and \U$19150 ( \19465 , \10166 , \4353 );
nor \U$19151 ( \19466 , \19464 , \19465 );
xnor \U$19152 ( \19467 , \19466 , \4212 );
and \U$19153 ( \19468 , \19463 , \19467 );
nand \U$19154 ( \19469 , \10967 , \4030 );
xnor \U$19155 ( \19470 , \19469 , \3786 );
and \U$19156 ( \19471 , \19467 , \19470 );
and \U$19157 ( \19472 , \19463 , \19470 );
or \U$19158 ( \19473 , \19468 , \19471 , \19472 );
and \U$19159 ( \19474 , \19459 , \19473 );
and \U$19160 ( \19475 , \10166 , \4355 );
and \U$19161 ( \19476 , \10161 , \4353 );
nor \U$19162 ( \19477 , \19475 , \19476 );
xnor \U$19163 ( \19478 , \19477 , \4212 );
and \U$19164 ( \19479 , \19473 , \19478 );
and \U$19165 ( \19480 , \19459 , \19478 );
or \U$19166 ( \19481 , \19474 , \19479 , \19480 );
and \U$19167 ( \19482 , \6500 , \7767 );
and \U$19168 ( \19483 , \6157 , \7765 );
nor \U$19169 ( \19484 , \19482 , \19483 );
xnor \U$19170 ( \19485 , \19484 , \7518 );
and \U$19171 ( \19486 , \7005 , \7238 );
and \U$19172 ( \19487 , \6702 , \7236 );
nor \U$19173 ( \19488 , \19486 , \19487 );
xnor \U$19174 ( \19489 , \19488 , \6978 );
and \U$19175 ( \19490 , \19485 , \19489 );
and \U$19176 ( \19491 , \7703 , \6744 );
and \U$19177 ( \19492 , \7177 , \6742 );
nor \U$19178 ( \19493 , \19491 , \19492 );
xnor \U$19179 ( \19494 , \19493 , \6429 );
and \U$19180 ( \19495 , \19489 , \19494 );
and \U$19181 ( \19496 , \19485 , \19494 );
or \U$19182 ( \19497 , \19490 , \19495 , \19496 );
and \U$19183 ( \19498 , \4272 , \10814 );
and \U$19184 ( \19499 , \4016 , \10811 );
nor \U$19185 ( \19500 , \19498 , \19499 );
xnor \U$19186 ( \19501 , \19500 , \9759 );
and \U$19187 ( \19502 , \4771 , \10001 );
and \U$19188 ( \19503 , \4469 , \9999 );
nor \U$19189 ( \19504 , \19502 , \19503 );
xnor \U$19190 ( \19505 , \19504 , \9762 );
and \U$19191 ( \19506 , \19501 , \19505 );
and \U$19192 ( \19507 , \19505 , \3786 );
and \U$19193 ( \19508 , \19501 , \3786 );
or \U$19194 ( \19509 , \19506 , \19507 , \19508 );
and \U$19195 ( \19510 , \19497 , \19509 );
and \U$19196 ( \19511 , \5248 , \9433 );
and \U$19197 ( \19512 , \4779 , \9431 );
nor \U$19198 ( \19513 , \19511 , \19512 );
xnor \U$19199 ( \19514 , \19513 , \9123 );
and \U$19200 ( \19515 , \5517 , \8896 );
and \U$19201 ( \19516 , \5253 , \8894 );
nor \U$19202 ( \19517 , \19515 , \19516 );
xnor \U$19203 ( \19518 , \19517 , \8525 );
and \U$19204 ( \19519 , \19514 , \19518 );
and \U$19205 ( \19520 , \6148 , \8334 );
and \U$19206 ( \19521 , \5776 , \8332 );
nor \U$19207 ( \19522 , \19520 , \19521 );
xnor \U$19208 ( \19523 , \19522 , \8016 );
and \U$19209 ( \19524 , \19518 , \19523 );
and \U$19210 ( \19525 , \19514 , \19523 );
or \U$19211 ( \19526 , \19519 , \19524 , \19525 );
and \U$19212 ( \19527 , \19509 , \19526 );
and \U$19213 ( \19528 , \19497 , \19526 );
or \U$19214 ( \19529 , \19510 , \19527 , \19528 );
and \U$19215 ( \19530 , \19481 , \19529 );
and \U$19216 ( \19531 , \10967 , \4032 );
and \U$19217 ( \19532 , \10347 , \4030 );
nor \U$19218 ( \19533 , \19531 , \19532 );
xnor \U$19219 ( \19534 , \19533 , \3786 );
xor \U$19220 ( \19535 , \19385 , \19389 );
xor \U$19221 ( \19536 , \19535 , \19394 );
and \U$19222 ( \19537 , \19534 , \19536 );
xor \U$19223 ( \19538 , \19338 , \19342 );
xor \U$19224 ( \19539 , \19538 , \19347 );
and \U$19225 ( \19540 , \19536 , \19539 );
and \U$19226 ( \19541 , \19534 , \19539 );
or \U$19227 ( \19542 , \19537 , \19540 , \19541 );
and \U$19228 ( \19543 , \19529 , \19542 );
and \U$19229 ( \19544 , \19481 , \19542 );
or \U$19230 ( \19545 , \19530 , \19543 , \19544 );
xor \U$19231 ( \19546 , \19216 , \19220 );
xor \U$19232 ( \19547 , \19546 , \3450 );
xor \U$19233 ( \19548 , \19372 , \19374 );
xor \U$19234 ( \19549 , \19548 , \19377 );
and \U$19235 ( \19550 , \19547 , \19549 );
xor \U$19236 ( \19551 , \19397 , \19399 );
xor \U$19237 ( \19552 , \19551 , \19402 );
and \U$19238 ( \19553 , \19549 , \19552 );
and \U$19239 ( \19554 , \19547 , \19552 );
or \U$19240 ( \19555 , \19550 , \19553 , \19554 );
and \U$19241 ( \19556 , \19545 , \19555 );
xor \U$19242 ( \19557 , \19195 , \19211 );
xor \U$19243 ( \19558 , \19557 , \19224 );
and \U$19244 ( \19559 , \19555 , \19558 );
and \U$19245 ( \19560 , \19545 , \19558 );
or \U$19246 ( \19561 , \19556 , \19559 , \19560 );
xor \U$19247 ( \19562 , \19370 , \19380 );
xor \U$19248 ( \19563 , \19562 , \19405 );
xor \U$19249 ( \19564 , \19410 , \19412 );
xor \U$19250 ( \19565 , \19564 , \19415 );
and \U$19251 ( \19566 , \19563 , \19565 );
and \U$19252 ( \19567 , \19561 , \19566 );
xor \U$19253 ( \19568 , \19281 , \19283 );
xor \U$19254 ( \19569 , \19568 , \19286 );
and \U$19255 ( \19570 , \19566 , \19569 );
and \U$19256 ( \19571 , \19561 , \19569 );
or \U$19257 ( \19572 , \19567 , \19570 , \19571 );
xor \U$19258 ( \19573 , \19227 , \19265 );
xor \U$19259 ( \19574 , \19573 , \19276 );
xor \U$19260 ( \19575 , \19408 , \19418 );
xor \U$19261 ( \19576 , \19575 , \19421 );
and \U$19262 ( \19577 , \19574 , \19576 );
and \U$19263 ( \19578 , \19572 , \19577 );
xor \U$19264 ( \19579 , \19424 , \19426 );
xor \U$19265 ( \19580 , \19579 , \19428 );
and \U$19266 ( \19581 , \19577 , \19580 );
and \U$19267 ( \19582 , \19572 , \19580 );
or \U$19268 ( \19583 , \19578 , \19581 , \19582 );
and \U$19269 ( \19584 , \19443 , \19583 );
xor \U$19270 ( \19585 , \19443 , \19583 );
xor \U$19271 ( \19586 , \19572 , \19577 );
xor \U$19272 ( \19587 , \19586 , \19580 );
and \U$19273 ( \19588 , \5776 , \8896 );
and \U$19274 ( \19589 , \5517 , \8894 );
nor \U$19275 ( \19590 , \19588 , \19589 );
xnor \U$19276 ( \19591 , \19590 , \8525 );
and \U$19277 ( \19592 , \6157 , \8334 );
and \U$19278 ( \19593 , \6148 , \8332 );
nor \U$19279 ( \19594 , \19592 , \19593 );
xnor \U$19280 ( \19595 , \19594 , \8016 );
and \U$19281 ( \19596 , \19591 , \19595 );
and \U$19282 ( \19597 , \6702 , \7767 );
and \U$19283 ( \19598 , \6500 , \7765 );
nor \U$19284 ( \19599 , \19597 , \19598 );
xnor \U$19285 ( \19600 , \19599 , \7518 );
and \U$19286 ( \19601 , \19595 , \19600 );
and \U$19287 ( \19602 , \19591 , \19600 );
or \U$19288 ( \19603 , \19596 , \19601 , \19602 );
and \U$19289 ( \19604 , \4469 , \10814 );
and \U$19290 ( \19605 , \4272 , \10811 );
nor \U$19291 ( \19606 , \19604 , \19605 );
xnor \U$19292 ( \19607 , \19606 , \9759 );
and \U$19293 ( \19608 , \4779 , \10001 );
and \U$19294 ( \19609 , \4771 , \9999 );
nor \U$19295 ( \19610 , \19608 , \19609 );
xnor \U$19296 ( \19611 , \19610 , \9762 );
and \U$19297 ( \19612 , \19607 , \19611 );
and \U$19298 ( \19613 , \5253 , \9433 );
and \U$19299 ( \19614 , \5248 , \9431 );
nor \U$19300 ( \19615 , \19613 , \19614 );
xnor \U$19301 ( \19616 , \19615 , \9123 );
and \U$19302 ( \19617 , \19611 , \19616 );
and \U$19303 ( \19618 , \19607 , \19616 );
or \U$19304 ( \19619 , \19612 , \19617 , \19618 );
and \U$19305 ( \19620 , \19603 , \19619 );
and \U$19306 ( \19621 , \7177 , \7238 );
and \U$19307 ( \19622 , \7005 , \7236 );
nor \U$19308 ( \19623 , \19621 , \19622 );
xnor \U$19309 ( \19624 , \19623 , \6978 );
and \U$19310 ( \19625 , \8127 , \6744 );
and \U$19311 ( \19626 , \7703 , \6742 );
nor \U$19312 ( \19627 , \19625 , \19626 );
xnor \U$19313 ( \19628 , \19627 , \6429 );
and \U$19314 ( \19629 , \19624 , \19628 );
and \U$19315 ( \19630 , \8378 , \6235 );
and \U$19316 ( \19631 , \8373 , \6233 );
nor \U$19317 ( \19632 , \19630 , \19631 );
xnor \U$19318 ( \19633 , \19632 , \5895 );
and \U$19319 ( \19634 , \19628 , \19633 );
and \U$19320 ( \19635 , \19624 , \19633 );
or \U$19321 ( \19636 , \19629 , \19634 , \19635 );
and \U$19322 ( \19637 , \19619 , \19636 );
and \U$19323 ( \19638 , \19603 , \19636 );
or \U$19324 ( \19639 , \19620 , \19637 , \19638 );
xor \U$19325 ( \19640 , \19485 , \19489 );
xor \U$19326 ( \19641 , \19640 , \19494 );
xor \U$19327 ( \19642 , \19501 , \19505 );
xor \U$19328 ( \19643 , \19642 , \3786 );
and \U$19329 ( \19644 , \19641 , \19643 );
xor \U$19330 ( \19645 , \19514 , \19518 );
xor \U$19331 ( \19646 , \19645 , \19523 );
and \U$19332 ( \19647 , \19643 , \19646 );
and \U$19333 ( \19648 , \19641 , \19646 );
or \U$19334 ( \19649 , \19644 , \19647 , \19648 );
and \U$19335 ( \19650 , \19639 , \19649 );
and \U$19336 ( \19651 , \8981 , \5646 );
and \U$19337 ( \19652 , \8697 , \5644 );
nor \U$19338 ( \19653 , \19651 , \19652 );
xnor \U$19339 ( \19654 , \19653 , \5405 );
and \U$19340 ( \19655 , \9558 , \5180 );
and \U$19341 ( \19656 , \9550 , \5178 );
nor \U$19342 ( \19657 , \19655 , \19656 );
xnor \U$19343 ( \19658 , \19657 , \4992 );
and \U$19344 ( \19659 , \19654 , \19658 );
and \U$19345 ( \19660 , \10166 , \4806 );
and \U$19346 ( \19661 , \10161 , \4804 );
nor \U$19347 ( \19662 , \19660 , \19661 );
xnor \U$19348 ( \19663 , \19662 , \4574 );
and \U$19349 ( \19664 , \19658 , \19663 );
and \U$19350 ( \19665 , \19654 , \19663 );
or \U$19351 ( \19666 , \19659 , \19664 , \19665 );
xor \U$19352 ( \19667 , \19447 , \19451 );
xor \U$19353 ( \19668 , \19667 , \19456 );
and \U$19354 ( \19669 , \19666 , \19668 );
xor \U$19355 ( \19670 , \19463 , \19467 );
xor \U$19356 ( \19671 , \19670 , \19470 );
and \U$19357 ( \19672 , \19668 , \19671 );
and \U$19358 ( \19673 , \19666 , \19671 );
or \U$19359 ( \19674 , \19669 , \19672 , \19673 );
and \U$19360 ( \19675 , \19649 , \19674 );
and \U$19361 ( \19676 , \19639 , \19674 );
or \U$19362 ( \19677 , \19650 , \19675 , \19676 );
xor \U$19363 ( \19678 , \19322 , \19326 );
xor \U$19364 ( \19679 , \19678 , \19331 );
xor \U$19365 ( \19680 , \19355 , \19359 );
xor \U$19366 ( \19681 , \19680 , \19364 );
and \U$19367 ( \19682 , \19679 , \19681 );
xor \U$19368 ( \19683 , \19534 , \19536 );
xor \U$19369 ( \19684 , \19683 , \19539 );
and \U$19370 ( \19685 , \19681 , \19684 );
and \U$19371 ( \19686 , \19679 , \19684 );
or \U$19372 ( \19687 , \19682 , \19685 , \19686 );
and \U$19373 ( \19688 , \19677 , \19687 );
xor \U$19374 ( \19689 , \19334 , \19350 );
xor \U$19375 ( \19690 , \19689 , \19367 );
and \U$19376 ( \19691 , \19687 , \19690 );
and \U$19377 ( \19692 , \19677 , \19690 );
or \U$19378 ( \19693 , \19688 , \19691 , \19692 );
xor \U$19379 ( \19694 , \19545 , \19555 );
xor \U$19380 ( \19695 , \19694 , \19558 );
and \U$19381 ( \19696 , \19693 , \19695 );
xor \U$19382 ( \19697 , \19563 , \19565 );
and \U$19383 ( \19698 , \19695 , \19697 );
and \U$19384 ( \19699 , \19693 , \19697 );
or \U$19385 ( \19700 , \19696 , \19698 , \19699 );
xor \U$19386 ( \19701 , \19561 , \19566 );
xor \U$19387 ( \19702 , \19701 , \19569 );
and \U$19388 ( \19703 , \19700 , \19702 );
xor \U$19389 ( \19704 , \19574 , \19576 );
and \U$19390 ( \19705 , \19702 , \19704 );
and \U$19391 ( \19706 , \19700 , \19704 );
or \U$19392 ( \19707 , \19703 , \19705 , \19706 );
and \U$19393 ( \19708 , \19587 , \19707 );
xor \U$19394 ( \19709 , \19587 , \19707 );
xor \U$19395 ( \19710 , \19700 , \19702 );
xor \U$19396 ( \19711 , \19710 , \19704 );
and \U$19397 ( \19712 , \5517 , \9433 );
and \U$19398 ( \19713 , \5253 , \9431 );
nor \U$19399 ( \19714 , \19712 , \19713 );
xnor \U$19400 ( \19715 , \19714 , \9123 );
and \U$19401 ( \19716 , \6148 , \8896 );
and \U$19402 ( \19717 , \5776 , \8894 );
nor \U$19403 ( \19718 , \19716 , \19717 );
xnor \U$19404 ( \19719 , \19718 , \8525 );
and \U$19405 ( \19720 , \19715 , \19719 );
and \U$19406 ( \19721 , \6500 , \8334 );
and \U$19407 ( \19722 , \6157 , \8332 );
nor \U$19408 ( \19723 , \19721 , \19722 );
xnor \U$19409 ( \19724 , \19723 , \8016 );
and \U$19410 ( \19725 , \19719 , \19724 );
and \U$19411 ( \19726 , \19715 , \19724 );
or \U$19412 ( \19727 , \19720 , \19725 , \19726 );
and \U$19413 ( \19728 , \4771 , \10814 );
and \U$19414 ( \19729 , \4469 , \10811 );
nor \U$19415 ( \19730 , \19728 , \19729 );
xnor \U$19416 ( \19731 , \19730 , \9759 );
and \U$19417 ( \19732 , \5248 , \10001 );
and \U$19418 ( \19733 , \4779 , \9999 );
nor \U$19419 ( \19734 , \19732 , \19733 );
xnor \U$19420 ( \19735 , \19734 , \9762 );
and \U$19421 ( \19736 , \19731 , \19735 );
and \U$19422 ( \19737 , \19735 , \4212 );
and \U$19423 ( \19738 , \19731 , \4212 );
or \U$19424 ( \19739 , \19736 , \19737 , \19738 );
and \U$19425 ( \19740 , \19727 , \19739 );
and \U$19426 ( \19741 , \7005 , \7767 );
and \U$19427 ( \19742 , \6702 , \7765 );
nor \U$19428 ( \19743 , \19741 , \19742 );
xnor \U$19429 ( \19744 , \19743 , \7518 );
and \U$19430 ( \19745 , \7703 , \7238 );
and \U$19431 ( \19746 , \7177 , \7236 );
nor \U$19432 ( \19747 , \19745 , \19746 );
xnor \U$19433 ( \19748 , \19747 , \6978 );
and \U$19434 ( \19749 , \19744 , \19748 );
and \U$19435 ( \19750 , \8373 , \6744 );
and \U$19436 ( \19751 , \8127 , \6742 );
nor \U$19437 ( \19752 , \19750 , \19751 );
xnor \U$19438 ( \19753 , \19752 , \6429 );
and \U$19439 ( \19754 , \19748 , \19753 );
and \U$19440 ( \19755 , \19744 , \19753 );
or \U$19441 ( \19756 , \19749 , \19754 , \19755 );
and \U$19442 ( \19757 , \19739 , \19756 );
and \U$19443 ( \19758 , \19727 , \19756 );
or \U$19444 ( \19759 , \19740 , \19757 , \19758 );
and \U$19445 ( \19760 , \8697 , \6235 );
and \U$19446 ( \19761 , \8378 , \6233 );
nor \U$19447 ( \19762 , \19760 , \19761 );
xnor \U$19448 ( \19763 , \19762 , \5895 );
and \U$19449 ( \19764 , \9550 , \5646 );
and \U$19450 ( \19765 , \8981 , \5644 );
nor \U$19451 ( \19766 , \19764 , \19765 );
xnor \U$19452 ( \19767 , \19766 , \5405 );
and \U$19453 ( \19768 , \19763 , \19767 );
and \U$19454 ( \19769 , \10161 , \5180 );
and \U$19455 ( \19770 , \9558 , \5178 );
nor \U$19456 ( \19771 , \19769 , \19770 );
xnor \U$19457 ( \19772 , \19771 , \4992 );
and \U$19458 ( \19773 , \19767 , \19772 );
and \U$19459 ( \19774 , \19763 , \19772 );
or \U$19460 ( \19775 , \19768 , \19773 , \19774 );
and \U$19461 ( \19776 , \10347 , \4806 );
and \U$19462 ( \19777 , \10166 , \4804 );
nor \U$19463 ( \19778 , \19776 , \19777 );
xnor \U$19464 ( \19779 , \19778 , \4574 );
nand \U$19465 ( \19780 , \10967 , \4353 );
xnor \U$19466 ( \19781 , \19780 , \4212 );
and \U$19467 ( \19782 , \19779 , \19781 );
and \U$19468 ( \19783 , \19775 , \19782 );
and \U$19469 ( \19784 , \10967 , \4355 );
and \U$19470 ( \19785 , \10347 , \4353 );
nor \U$19471 ( \19786 , \19784 , \19785 );
xnor \U$19472 ( \19787 , \19786 , \4212 );
and \U$19473 ( \19788 , \19782 , \19787 );
and \U$19474 ( \19789 , \19775 , \19787 );
or \U$19475 ( \19790 , \19783 , \19788 , \19789 );
and \U$19476 ( \19791 , \19759 , \19790 );
xor \U$19477 ( \19792 , \19591 , \19595 );
xor \U$19478 ( \19793 , \19792 , \19600 );
xor \U$19479 ( \19794 , \19654 , \19658 );
xor \U$19480 ( \19795 , \19794 , \19663 );
and \U$19481 ( \19796 , \19793 , \19795 );
xor \U$19482 ( \19797 , \19624 , \19628 );
xor \U$19483 ( \19798 , \19797 , \19633 );
and \U$19484 ( \19799 , \19795 , \19798 );
and \U$19485 ( \19800 , \19793 , \19798 );
or \U$19486 ( \19801 , \19796 , \19799 , \19800 );
and \U$19487 ( \19802 , \19790 , \19801 );
and \U$19488 ( \19803 , \19759 , \19801 );
or \U$19489 ( \19804 , \19791 , \19802 , \19803 );
xor \U$19490 ( \19805 , \19603 , \19619 );
xor \U$19491 ( \19806 , \19805 , \19636 );
xor \U$19492 ( \19807 , \19641 , \19643 );
xor \U$19493 ( \19808 , \19807 , \19646 );
and \U$19494 ( \19809 , \19806 , \19808 );
xor \U$19495 ( \19810 , \19666 , \19668 );
xor \U$19496 ( \19811 , \19810 , \19671 );
and \U$19497 ( \19812 , \19808 , \19811 );
and \U$19498 ( \19813 , \19806 , \19811 );
or \U$19499 ( \19814 , \19809 , \19812 , \19813 );
and \U$19500 ( \19815 , \19804 , \19814 );
xor \U$19501 ( \19816 , \19459 , \19473 );
xor \U$19502 ( \19817 , \19816 , \19478 );
and \U$19503 ( \19818 , \19814 , \19817 );
and \U$19504 ( \19819 , \19804 , \19817 );
or \U$19505 ( \19820 , \19815 , \19818 , \19819 );
xor \U$19506 ( \19821 , \19497 , \19509 );
xor \U$19507 ( \19822 , \19821 , \19526 );
xor \U$19508 ( \19823 , \19639 , \19649 );
xor \U$19509 ( \19824 , \19823 , \19674 );
and \U$19510 ( \19825 , \19822 , \19824 );
xor \U$19511 ( \19826 , \19679 , \19681 );
xor \U$19512 ( \19827 , \19826 , \19684 );
and \U$19513 ( \19828 , \19824 , \19827 );
and \U$19514 ( \19829 , \19822 , \19827 );
or \U$19515 ( \19830 , \19825 , \19828 , \19829 );
and \U$19516 ( \19831 , \19820 , \19830 );
xor \U$19517 ( \19832 , \19547 , \19549 );
xor \U$19518 ( \19833 , \19832 , \19552 );
and \U$19519 ( \19834 , \19830 , \19833 );
and \U$19520 ( \19835 , \19820 , \19833 );
or \U$19521 ( \19836 , \19831 , \19834 , \19835 );
xor \U$19522 ( \19837 , \19481 , \19529 );
xor \U$19523 ( \19838 , \19837 , \19542 );
xor \U$19524 ( \19839 , \19677 , \19687 );
xor \U$19525 ( \19840 , \19839 , \19690 );
and \U$19526 ( \19841 , \19838 , \19840 );
and \U$19527 ( \19842 , \19836 , \19841 );
xor \U$19528 ( \19843 , \19693 , \19695 );
xor \U$19529 ( \19844 , \19843 , \19697 );
and \U$19530 ( \19845 , \19841 , \19844 );
and \U$19531 ( \19846 , \19836 , \19844 );
or \U$19532 ( \19847 , \19842 , \19845 , \19846 );
and \U$19533 ( \19848 , \19711 , \19847 );
xor \U$19534 ( \19849 , \19711 , \19847 );
xor \U$19535 ( \19850 , \19836 , \19841 );
xor \U$19536 ( \19851 , \19850 , \19844 );
and \U$19537 ( \19852 , \6157 , \8896 );
and \U$19538 ( \19853 , \6148 , \8894 );
nor \U$19539 ( \19854 , \19852 , \19853 );
xnor \U$19540 ( \19855 , \19854 , \8525 );
and \U$19541 ( \19856 , \6702 , \8334 );
and \U$19542 ( \19857 , \6500 , \8332 );
nor \U$19543 ( \19858 , \19856 , \19857 );
xnor \U$19544 ( \19859 , \19858 , \8016 );
and \U$19545 ( \19860 , \19855 , \19859 );
and \U$19546 ( \19861 , \7177 , \7767 );
and \U$19547 ( \19862 , \7005 , \7765 );
nor \U$19548 ( \19863 , \19861 , \19862 );
xnor \U$19549 ( \19864 , \19863 , \7518 );
and \U$19550 ( \19865 , \19859 , \19864 );
and \U$19551 ( \19866 , \19855 , \19864 );
or \U$19552 ( \19867 , \19860 , \19865 , \19866 );
and \U$19553 ( \19868 , \8127 , \7238 );
and \U$19554 ( \19869 , \7703 , \7236 );
nor \U$19555 ( \19870 , \19868 , \19869 );
xnor \U$19556 ( \19871 , \19870 , \6978 );
and \U$19557 ( \19872 , \8378 , \6744 );
and \U$19558 ( \19873 , \8373 , \6742 );
nor \U$19559 ( \19874 , \19872 , \19873 );
xnor \U$19560 ( \19875 , \19874 , \6429 );
and \U$19561 ( \19876 , \19871 , \19875 );
and \U$19562 ( \19877 , \8981 , \6235 );
and \U$19563 ( \19878 , \8697 , \6233 );
nor \U$19564 ( \19879 , \19877 , \19878 );
xnor \U$19565 ( \19880 , \19879 , \5895 );
and \U$19566 ( \19881 , \19875 , \19880 );
and \U$19567 ( \19882 , \19871 , \19880 );
or \U$19568 ( \19883 , \19876 , \19881 , \19882 );
and \U$19569 ( \19884 , \19867 , \19883 );
and \U$19570 ( \19885 , \4779 , \10814 );
and \U$19571 ( \19886 , \4771 , \10811 );
nor \U$19572 ( \19887 , \19885 , \19886 );
xnor \U$19573 ( \19888 , \19887 , \9759 );
and \U$19574 ( \19889 , \5253 , \10001 );
and \U$19575 ( \19890 , \5248 , \9999 );
nor \U$19576 ( \19891 , \19889 , \19890 );
xnor \U$19577 ( \19892 , \19891 , \9762 );
and \U$19578 ( \19893 , \19888 , \19892 );
and \U$19579 ( \19894 , \5776 , \9433 );
and \U$19580 ( \19895 , \5517 , \9431 );
nor \U$19581 ( \19896 , \19894 , \19895 );
xnor \U$19582 ( \19897 , \19896 , \9123 );
and \U$19583 ( \19898 , \19892 , \19897 );
and \U$19584 ( \19899 , \19888 , \19897 );
or \U$19585 ( \19900 , \19893 , \19898 , \19899 );
and \U$19586 ( \19901 , \19883 , \19900 );
and \U$19587 ( \19902 , \19867 , \19900 );
or \U$19588 ( \19903 , \19884 , \19901 , \19902 );
xor \U$19589 ( \19904 , \19715 , \19719 );
xor \U$19590 ( \19905 , \19904 , \19724 );
xor \U$19591 ( \19906 , \19731 , \19735 );
xor \U$19592 ( \19907 , \19906 , \4212 );
and \U$19593 ( \19908 , \19905 , \19907 );
xor \U$19594 ( \19909 , \19744 , \19748 );
xor \U$19595 ( \19910 , \19909 , \19753 );
and \U$19596 ( \19911 , \19907 , \19910 );
and \U$19597 ( \19912 , \19905 , \19910 );
or \U$19598 ( \19913 , \19908 , \19911 , \19912 );
and \U$19599 ( \19914 , \19903 , \19913 );
and \U$19600 ( \19915 , \9558 , \5646 );
and \U$19601 ( \19916 , \9550 , \5644 );
nor \U$19602 ( \19917 , \19915 , \19916 );
xnor \U$19603 ( \19918 , \19917 , \5405 );
and \U$19604 ( \19919 , \10166 , \5180 );
and \U$19605 ( \19920 , \10161 , \5178 );
nor \U$19606 ( \19921 , \19919 , \19920 );
xnor \U$19607 ( \19922 , \19921 , \4992 );
and \U$19608 ( \19923 , \19918 , \19922 );
and \U$19609 ( \19924 , \10967 , \4806 );
and \U$19610 ( \19925 , \10347 , \4804 );
nor \U$19611 ( \19926 , \19924 , \19925 );
xnor \U$19612 ( \19927 , \19926 , \4574 );
and \U$19613 ( \19928 , \19922 , \19927 );
and \U$19614 ( \19929 , \19918 , \19927 );
or \U$19615 ( \19930 , \19923 , \19928 , \19929 );
xor \U$19616 ( \19931 , \19763 , \19767 );
xor \U$19617 ( \19932 , \19931 , \19772 );
and \U$19618 ( \19933 , \19930 , \19932 );
xor \U$19619 ( \19934 , \19779 , \19781 );
and \U$19620 ( \19935 , \19932 , \19934 );
and \U$19621 ( \19936 , \19930 , \19934 );
or \U$19622 ( \19937 , \19933 , \19935 , \19936 );
and \U$19623 ( \19938 , \19913 , \19937 );
and \U$19624 ( \19939 , \19903 , \19937 );
or \U$19625 ( \19940 , \19914 , \19938 , \19939 );
xor \U$19626 ( \19941 , \19607 , \19611 );
xor \U$19627 ( \19942 , \19941 , \19616 );
xor \U$19628 ( \19943 , \19775 , \19782 );
xor \U$19629 ( \19944 , \19943 , \19787 );
and \U$19630 ( \19945 , \19942 , \19944 );
xor \U$19631 ( \19946 , \19793 , \19795 );
xor \U$19632 ( \19947 , \19946 , \19798 );
and \U$19633 ( \19948 , \19944 , \19947 );
and \U$19634 ( \19949 , \19942 , \19947 );
or \U$19635 ( \19950 , \19945 , \19948 , \19949 );
and \U$19636 ( \19951 , \19940 , \19950 );
xor \U$19637 ( \19952 , \19806 , \19808 );
xor \U$19638 ( \19953 , \19952 , \19811 );
and \U$19639 ( \19954 , \19950 , \19953 );
and \U$19640 ( \19955 , \19940 , \19953 );
or \U$19641 ( \19956 , \19951 , \19954 , \19955 );
xor \U$19642 ( \19957 , \19804 , \19814 );
xor \U$19643 ( \19958 , \19957 , \19817 );
and \U$19644 ( \19959 , \19956 , \19958 );
xor \U$19645 ( \19960 , \19822 , \19824 );
xor \U$19646 ( \19961 , \19960 , \19827 );
and \U$19647 ( \19962 , \19958 , \19961 );
and \U$19648 ( \19963 , \19956 , \19961 );
or \U$19649 ( \19964 , \19959 , \19962 , \19963 );
xor \U$19650 ( \19965 , \19820 , \19830 );
xor \U$19651 ( \19966 , \19965 , \19833 );
and \U$19652 ( \19967 , \19964 , \19966 );
xor \U$19653 ( \19968 , \19838 , \19840 );
and \U$19654 ( \19969 , \19966 , \19968 );
and \U$19655 ( \19970 , \19964 , \19968 );
or \U$19656 ( \19971 , \19967 , \19969 , \19970 );
and \U$19657 ( \19972 , \19851 , \19971 );
xor \U$19658 ( \19973 , \19851 , \19971 );
xor \U$19659 ( \19974 , \19964 , \19966 );
xor \U$19660 ( \19975 , \19974 , \19968 );
and \U$19661 ( \19976 , \6148 , \9433 );
and \U$19662 ( \19977 , \5776 , \9431 );
nor \U$19663 ( \19978 , \19976 , \19977 );
xnor \U$19664 ( \19979 , \19978 , \9123 );
and \U$19665 ( \19980 , \6500 , \8896 );
and \U$19666 ( \19981 , \6157 , \8894 );
nor \U$19667 ( \19982 , \19980 , \19981 );
xnor \U$19668 ( \19983 , \19982 , \8525 );
and \U$19669 ( \19984 , \19979 , \19983 );
and \U$19670 ( \19985 , \7005 , \8334 );
and \U$19671 ( \19986 , \6702 , \8332 );
nor \U$19672 ( \19987 , \19985 , \19986 );
xnor \U$19673 ( \19988 , \19987 , \8016 );
and \U$19674 ( \19989 , \19983 , \19988 );
and \U$19675 ( \19990 , \19979 , \19988 );
or \U$19676 ( \19991 , \19984 , \19989 , \19990 );
and \U$19677 ( \19992 , \7703 , \7767 );
and \U$19678 ( \19993 , \7177 , \7765 );
nor \U$19679 ( \19994 , \19992 , \19993 );
xnor \U$19680 ( \19995 , \19994 , \7518 );
and \U$19681 ( \19996 , \8373 , \7238 );
and \U$19682 ( \19997 , \8127 , \7236 );
nor \U$19683 ( \19998 , \19996 , \19997 );
xnor \U$19684 ( \19999 , \19998 , \6978 );
and \U$19685 ( \20000 , \19995 , \19999 );
and \U$19686 ( \20001 , \8697 , \6744 );
and \U$19687 ( \20002 , \8378 , \6742 );
nor \U$19688 ( \20003 , \20001 , \20002 );
xnor \U$19689 ( \20004 , \20003 , \6429 );
and \U$19690 ( \20005 , \19999 , \20004 );
and \U$19691 ( \20006 , \19995 , \20004 );
or \U$19692 ( \20007 , \20000 , \20005 , \20006 );
and \U$19693 ( \20008 , \19991 , \20007 );
and \U$19694 ( \20009 , \5248 , \10814 );
and \U$19695 ( \20010 , \4779 , \10811 );
nor \U$19696 ( \20011 , \20009 , \20010 );
xnor \U$19697 ( \20012 , \20011 , \9759 );
and \U$19698 ( \20013 , \5517 , \10001 );
and \U$19699 ( \20014 , \5253 , \9999 );
nor \U$19700 ( \20015 , \20013 , \20014 );
xnor \U$19701 ( \20016 , \20015 , \9762 );
and \U$19702 ( \20017 , \20012 , \20016 );
and \U$19703 ( \20018 , \20016 , \4574 );
and \U$19704 ( \20019 , \20012 , \4574 );
or \U$19705 ( \20020 , \20017 , \20018 , \20019 );
and \U$19706 ( \20021 , \20007 , \20020 );
and \U$19707 ( \20022 , \19991 , \20020 );
or \U$19708 ( \20023 , \20008 , \20021 , \20022 );
and \U$19709 ( \20024 , \9550 , \6235 );
and \U$19710 ( \20025 , \8981 , \6233 );
nor \U$19711 ( \20026 , \20024 , \20025 );
xnor \U$19712 ( \20027 , \20026 , \5895 );
and \U$19713 ( \20028 , \10161 , \5646 );
and \U$19714 ( \20029 , \9558 , \5644 );
nor \U$19715 ( \20030 , \20028 , \20029 );
xnor \U$19716 ( \20031 , \20030 , \5405 );
and \U$19717 ( \20032 , \20027 , \20031 );
and \U$19718 ( \20033 , \10347 , \5180 );
and \U$19719 ( \20034 , \10166 , \5178 );
nor \U$19720 ( \20035 , \20033 , \20034 );
xnor \U$19721 ( \20036 , \20035 , \4992 );
and \U$19722 ( \20037 , \20031 , \20036 );
and \U$19723 ( \20038 , \20027 , \20036 );
or \U$19724 ( \20039 , \20032 , \20037 , \20038 );
xor \U$19725 ( \20040 , \19871 , \19875 );
xor \U$19726 ( \20041 , \20040 , \19880 );
and \U$19727 ( \20042 , \20039 , \20041 );
xor \U$19728 ( \20043 , \19918 , \19922 );
xor \U$19729 ( \20044 , \20043 , \19927 );
and \U$19730 ( \20045 , \20041 , \20044 );
and \U$19731 ( \20046 , \20039 , \20044 );
or \U$19732 ( \20047 , \20042 , \20045 , \20046 );
and \U$19733 ( \20048 , \20023 , \20047 );
xor \U$19734 ( \20049 , \19855 , \19859 );
xor \U$19735 ( \20050 , \20049 , \19864 );
xor \U$19736 ( \20051 , \19888 , \19892 );
xor \U$19737 ( \20052 , \20051 , \19897 );
and \U$19738 ( \20053 , \20050 , \20052 );
and \U$19739 ( \20054 , \20047 , \20053 );
and \U$19740 ( \20055 , \20023 , \20053 );
or \U$19741 ( \20056 , \20048 , \20054 , \20055 );
xor \U$19742 ( \20057 , \19867 , \19883 );
xor \U$19743 ( \20058 , \20057 , \19900 );
xor \U$19744 ( \20059 , \19905 , \19907 );
xor \U$19745 ( \20060 , \20059 , \19910 );
and \U$19746 ( \20061 , \20058 , \20060 );
xor \U$19747 ( \20062 , \19930 , \19932 );
xor \U$19748 ( \20063 , \20062 , \19934 );
and \U$19749 ( \20064 , \20060 , \20063 );
and \U$19750 ( \20065 , \20058 , \20063 );
or \U$19751 ( \20066 , \20061 , \20064 , \20065 );
and \U$19752 ( \20067 , \20056 , \20066 );
xor \U$19753 ( \20068 , \19727 , \19739 );
xor \U$19754 ( \20069 , \20068 , \19756 );
and \U$19755 ( \20070 , \20066 , \20069 );
and \U$19756 ( \20071 , \20056 , \20069 );
or \U$19757 ( \20072 , \20067 , \20070 , \20071 );
xor \U$19758 ( \20073 , \19903 , \19913 );
xor \U$19759 ( \20074 , \20073 , \19937 );
xor \U$19760 ( \20075 , \19942 , \19944 );
xor \U$19761 ( \20076 , \20075 , \19947 );
and \U$19762 ( \20077 , \20074 , \20076 );
and \U$19763 ( \20078 , \20072 , \20077 );
xor \U$19764 ( \20079 , \19759 , \19790 );
xor \U$19765 ( \20080 , \20079 , \19801 );
and \U$19766 ( \20081 , \20077 , \20080 );
and \U$19767 ( \20082 , \20072 , \20080 );
or \U$19768 ( \20083 , \20078 , \20081 , \20082 );
xor \U$19769 ( \20084 , \19956 , \19958 );
xor \U$19770 ( \20085 , \20084 , \19961 );
and \U$19771 ( \20086 , \20083 , \20085 );
and \U$19772 ( \20087 , \19975 , \20086 );
xor \U$19773 ( \20088 , \19975 , \20086 );
xor \U$19774 ( \20089 , \20083 , \20085 );
xor \U$19775 ( \20090 , \20072 , \20077 );
xor \U$19776 ( \20091 , \20090 , \20080 );
xor \U$19777 ( \20092 , \19940 , \19950 );
xor \U$19778 ( \20093 , \20092 , \19953 );
and \U$19779 ( \20094 , \20091 , \20093 );
and \U$19780 ( \20095 , \20089 , \20094 );
xor \U$19781 ( \20096 , \20089 , \20094 );
xor \U$19782 ( \20097 , \20091 , \20093 );
and \U$19783 ( \20098 , \5253 , \10814 );
and \U$19784 ( \20099 , \5248 , \10811 );
nor \U$19785 ( \20100 , \20098 , \20099 );
xnor \U$19786 ( \20101 , \20100 , \9759 );
and \U$19787 ( \20102 , \5776 , \10001 );
and \U$19788 ( \20103 , \5517 , \9999 );
nor \U$19789 ( \20104 , \20102 , \20103 );
xnor \U$19790 ( \20105 , \20104 , \9762 );
and \U$19791 ( \20106 , \20101 , \20105 );
and \U$19792 ( \20107 , \6157 , \9433 );
and \U$19793 ( \20108 , \6148 , \9431 );
nor \U$19794 ( \20109 , \20107 , \20108 );
xnor \U$19795 ( \20110 , \20109 , \9123 );
and \U$19796 ( \20111 , \20105 , \20110 );
and \U$19797 ( \20112 , \20101 , \20110 );
or \U$19798 ( \20113 , \20106 , \20111 , \20112 );
and \U$19799 ( \20114 , \8378 , \7238 );
and \U$19800 ( \20115 , \8373 , \7236 );
nor \U$19801 ( \20116 , \20114 , \20115 );
xnor \U$19802 ( \20117 , \20116 , \6978 );
and \U$19803 ( \20118 , \8981 , \6744 );
and \U$19804 ( \20119 , \8697 , \6742 );
nor \U$19805 ( \20120 , \20118 , \20119 );
xnor \U$19806 ( \20121 , \20120 , \6429 );
and \U$19807 ( \20122 , \20117 , \20121 );
and \U$19808 ( \20123 , \9558 , \6235 );
and \U$19809 ( \20124 , \9550 , \6233 );
nor \U$19810 ( \20125 , \20123 , \20124 );
xnor \U$19811 ( \20126 , \20125 , \5895 );
and \U$19812 ( \20127 , \20121 , \20126 );
and \U$19813 ( \20128 , \20117 , \20126 );
or \U$19814 ( \20129 , \20122 , \20127 , \20128 );
and \U$19815 ( \20130 , \20113 , \20129 );
and \U$19816 ( \20131 , \6702 , \8896 );
and \U$19817 ( \20132 , \6500 , \8894 );
nor \U$19818 ( \20133 , \20131 , \20132 );
xnor \U$19819 ( \20134 , \20133 , \8525 );
and \U$19820 ( \20135 , \7177 , \8334 );
and \U$19821 ( \20136 , \7005 , \8332 );
nor \U$19822 ( \20137 , \20135 , \20136 );
xnor \U$19823 ( \20138 , \20137 , \8016 );
and \U$19824 ( \20139 , \20134 , \20138 );
and \U$19825 ( \20140 , \8127 , \7767 );
and \U$19826 ( \20141 , \7703 , \7765 );
nor \U$19827 ( \20142 , \20140 , \20141 );
xnor \U$19828 ( \20143 , \20142 , \7518 );
and \U$19829 ( \20144 , \20138 , \20143 );
and \U$19830 ( \20145 , \20134 , \20143 );
or \U$19831 ( \20146 , \20139 , \20144 , \20145 );
and \U$19832 ( \20147 , \20129 , \20146 );
and \U$19833 ( \20148 , \20113 , \20146 );
or \U$19834 ( \20149 , \20130 , \20147 , \20148 );
nand \U$19835 ( \20150 , \10967 , \4804 );
xnor \U$19836 ( \20151 , \20150 , \4574 );
xor \U$19837 ( \20152 , \19995 , \19999 );
xor \U$19838 ( \20153 , \20152 , \20004 );
and \U$19839 ( \20154 , \20151 , \20153 );
xor \U$19840 ( \20155 , \20027 , \20031 );
xor \U$19841 ( \20156 , \20155 , \20036 );
and \U$19842 ( \20157 , \20153 , \20156 );
and \U$19843 ( \20158 , \20151 , \20156 );
or \U$19844 ( \20159 , \20154 , \20157 , \20158 );
and \U$19845 ( \20160 , \20149 , \20159 );
xor \U$19846 ( \20161 , \19979 , \19983 );
xor \U$19847 ( \20162 , \20161 , \19988 );
xor \U$19848 ( \20163 , \20012 , \20016 );
xor \U$19849 ( \20164 , \20163 , \4574 );
and \U$19850 ( \20165 , \20162 , \20164 );
and \U$19851 ( \20166 , \20159 , \20165 );
and \U$19852 ( \20167 , \20149 , \20165 );
or \U$19853 ( \20168 , \20160 , \20166 , \20167 );
xor \U$19854 ( \20169 , \19991 , \20007 );
xor \U$19855 ( \20170 , \20169 , \20020 );
xor \U$19856 ( \20171 , \20039 , \20041 );
xor \U$19857 ( \20172 , \20171 , \20044 );
and \U$19858 ( \20173 , \20170 , \20172 );
xor \U$19859 ( \20174 , \20050 , \20052 );
and \U$19860 ( \20175 , \20172 , \20174 );
and \U$19861 ( \20176 , \20170 , \20174 );
or \U$19862 ( \20177 , \20173 , \20175 , \20176 );
and \U$19863 ( \20178 , \20168 , \20177 );
xor \U$19864 ( \20179 , \20058 , \20060 );
xor \U$19865 ( \20180 , \20179 , \20063 );
and \U$19866 ( \20181 , \20177 , \20180 );
and \U$19867 ( \20182 , \20168 , \20180 );
or \U$19868 ( \20183 , \20178 , \20181 , \20182 );
xor \U$19869 ( \20184 , \20056 , \20066 );
xor \U$19870 ( \20185 , \20184 , \20069 );
and \U$19871 ( \20186 , \20183 , \20185 );
xor \U$19872 ( \20187 , \20074 , \20076 );
and \U$19873 ( \20188 , \20185 , \20187 );
and \U$19874 ( \20189 , \20183 , \20187 );
or \U$19875 ( \20190 , \20186 , \20188 , \20189 );
and \U$19876 ( \20191 , \20097 , \20190 );
xor \U$19877 ( \20192 , \20097 , \20190 );
xor \U$19878 ( \20193 , \20183 , \20185 );
xor \U$19879 ( \20194 , \20193 , \20187 );
and \U$19880 ( \20195 , \10161 , \6235 );
and \U$19881 ( \20196 , \9558 , \6233 );
nor \U$19882 ( \20197 , \20195 , \20196 );
xnor \U$19883 ( \20198 , \20197 , \5895 );
and \U$19884 ( \20199 , \10347 , \5646 );
and \U$19885 ( \20200 , \10166 , \5644 );
nor \U$19886 ( \20201 , \20199 , \20200 );
xnor \U$19887 ( \20202 , \20201 , \5405 );
and \U$19888 ( \20203 , \20198 , \20202 );
nand \U$19889 ( \20204 , \10967 , \5178 );
xnor \U$19890 ( \20205 , \20204 , \4992 );
and \U$19891 ( \20206 , \20202 , \20205 );
and \U$19892 ( \20207 , \20198 , \20205 );
or \U$19893 ( \20208 , \20203 , \20206 , \20207 );
and \U$19894 ( \20209 , \10166 , \5646 );
and \U$19895 ( \20210 , \10161 , \5644 );
nor \U$19896 ( \20211 , \20209 , \20210 );
xnor \U$19897 ( \20212 , \20211 , \5405 );
and \U$19898 ( \20213 , \20208 , \20212 );
and \U$19899 ( \20214 , \10967 , \5180 );
and \U$19900 ( \20215 , \10347 , \5178 );
nor \U$19901 ( \20216 , \20214 , \20215 );
xnor \U$19902 ( \20217 , \20216 , \4992 );
and \U$19903 ( \20218 , \20212 , \20217 );
and \U$19904 ( \20219 , \20208 , \20217 );
or \U$19905 ( \20220 , \20213 , \20218 , \20219 );
and \U$19906 ( \20221 , \5517 , \10814 );
and \U$19907 ( \20222 , \5253 , \10811 );
nor \U$19908 ( \20223 , \20221 , \20222 );
xnor \U$19909 ( \20224 , \20223 , \9759 );
and \U$19910 ( \20225 , \6148 , \10001 );
and \U$19911 ( \20226 , \5776 , \9999 );
nor \U$19912 ( \20227 , \20225 , \20226 );
xnor \U$19913 ( \20228 , \20227 , \9762 );
and \U$19914 ( \20229 , \20224 , \20228 );
and \U$19915 ( \20230 , \20228 , \4992 );
and \U$19916 ( \20231 , \20224 , \4992 );
or \U$19917 ( \20232 , \20229 , \20230 , \20231 );
and \U$19918 ( \20233 , \6500 , \9433 );
and \U$19919 ( \20234 , \6157 , \9431 );
nor \U$19920 ( \20235 , \20233 , \20234 );
xnor \U$19921 ( \20236 , \20235 , \9123 );
and \U$19922 ( \20237 , \7005 , \8896 );
and \U$19923 ( \20238 , \6702 , \8894 );
nor \U$19924 ( \20239 , \20237 , \20238 );
xnor \U$19925 ( \20240 , \20239 , \8525 );
and \U$19926 ( \20241 , \20236 , \20240 );
and \U$19927 ( \20242 , \7703 , \8334 );
and \U$19928 ( \20243 , \7177 , \8332 );
nor \U$19929 ( \20244 , \20242 , \20243 );
xnor \U$19930 ( \20245 , \20244 , \8016 );
and \U$19931 ( \20246 , \20240 , \20245 );
and \U$19932 ( \20247 , \20236 , \20245 );
or \U$19933 ( \20248 , \20241 , \20246 , \20247 );
and \U$19934 ( \20249 , \20232 , \20248 );
and \U$19935 ( \20250 , \8373 , \7767 );
and \U$19936 ( \20251 , \8127 , \7765 );
nor \U$19937 ( \20252 , \20250 , \20251 );
xnor \U$19938 ( \20253 , \20252 , \7518 );
and \U$19939 ( \20254 , \8697 , \7238 );
and \U$19940 ( \20255 , \8378 , \7236 );
nor \U$19941 ( \20256 , \20254 , \20255 );
xnor \U$19942 ( \20257 , \20256 , \6978 );
and \U$19943 ( \20258 , \20253 , \20257 );
and \U$19944 ( \20259 , \9550 , \6744 );
and \U$19945 ( \20260 , \8981 , \6742 );
nor \U$19946 ( \20261 , \20259 , \20260 );
xnor \U$19947 ( \20262 , \20261 , \6429 );
and \U$19948 ( \20263 , \20257 , \20262 );
and \U$19949 ( \20264 , \20253 , \20262 );
or \U$19950 ( \20265 , \20258 , \20263 , \20264 );
and \U$19951 ( \20266 , \20248 , \20265 );
and \U$19952 ( \20267 , \20232 , \20265 );
or \U$19953 ( \20268 , \20249 , \20266 , \20267 );
and \U$19954 ( \20269 , \20220 , \20268 );
xor \U$19955 ( \20270 , \20101 , \20105 );
xor \U$19956 ( \20271 , \20270 , \20110 );
xor \U$19957 ( \20272 , \20117 , \20121 );
xor \U$19958 ( \20273 , \20272 , \20126 );
and \U$19959 ( \20274 , \20271 , \20273 );
xor \U$19960 ( \20275 , \20134 , \20138 );
xor \U$19961 ( \20276 , \20275 , \20143 );
and \U$19962 ( \20277 , \20273 , \20276 );
and \U$19963 ( \20278 , \20271 , \20276 );
or \U$19964 ( \20279 , \20274 , \20277 , \20278 );
and \U$19965 ( \20280 , \20268 , \20279 );
and \U$19966 ( \20281 , \20220 , \20279 );
or \U$19967 ( \20282 , \20269 , \20280 , \20281 );
xor \U$19968 ( \20283 , \20113 , \20129 );
xor \U$19969 ( \20284 , \20283 , \20146 );
xor \U$19970 ( \20285 , \20151 , \20153 );
xor \U$19971 ( \20286 , \20285 , \20156 );
and \U$19972 ( \20287 , \20284 , \20286 );
xor \U$19973 ( \20288 , \20162 , \20164 );
and \U$19974 ( \20289 , \20286 , \20288 );
and \U$19975 ( \20290 , \20284 , \20288 );
or \U$19976 ( \20291 , \20287 , \20289 , \20290 );
and \U$19977 ( \20292 , \20282 , \20291 );
xor \U$19978 ( \20293 , \20170 , \20172 );
xor \U$19979 ( \20294 , \20293 , \20174 );
and \U$19980 ( \20295 , \20291 , \20294 );
and \U$19981 ( \20296 , \20282 , \20294 );
or \U$19982 ( \20297 , \20292 , \20295 , \20296 );
xor \U$19983 ( \20298 , \20023 , \20047 );
xor \U$19984 ( \20299 , \20298 , \20053 );
and \U$19985 ( \20300 , \20297 , \20299 );
xor \U$19986 ( \20301 , \20168 , \20177 );
xor \U$19987 ( \20302 , \20301 , \20180 );
and \U$19988 ( \20303 , \20299 , \20302 );
and \U$19989 ( \20304 , \20297 , \20302 );
or \U$19990 ( \20305 , \20300 , \20303 , \20304 );
and \U$19991 ( \20306 , \20194 , \20305 );
xor \U$19992 ( \20307 , \20194 , \20305 );
xor \U$19993 ( \20308 , \20297 , \20299 );
xor \U$19994 ( \20309 , \20308 , \20302 );
and \U$19995 ( \20310 , \8981 , \7238 );
and \U$19996 ( \20311 , \8697 , \7236 );
nor \U$19997 ( \20312 , \20310 , \20311 );
xnor \U$19998 ( \20313 , \20312 , \6978 );
and \U$19999 ( \20314 , \9558 , \6744 );
and \U$20000 ( \20315 , \9550 , \6742 );
nor \U$20001 ( \20316 , \20314 , \20315 );
xnor \U$20002 ( \20317 , \20316 , \6429 );
and \U$20003 ( \20318 , \20313 , \20317 );
and \U$20004 ( \20319 , \10166 , \6235 );
and \U$20005 ( \20320 , \10161 , \6233 );
nor \U$20006 ( \20321 , \20319 , \20320 );
xnor \U$20007 ( \20322 , \20321 , \5895 );
and \U$20008 ( \20323 , \20317 , \20322 );
and \U$20009 ( \20324 , \20313 , \20322 );
or \U$20010 ( \20325 , \20318 , \20323 , \20324 );
and \U$20011 ( \20326 , \5776 , \10814 );
and \U$20012 ( \20327 , \5517 , \10811 );
nor \U$20013 ( \20328 , \20326 , \20327 );
xnor \U$20014 ( \20329 , \20328 , \9759 );
and \U$20015 ( \20330 , \6157 , \10001 );
and \U$20016 ( \20331 , \6148 , \9999 );
nor \U$20017 ( \20332 , \20330 , \20331 );
xnor \U$20018 ( \20333 , \20332 , \9762 );
and \U$20019 ( \20334 , \20329 , \20333 );
and \U$20020 ( \20335 , \6702 , \9433 );
and \U$20021 ( \20336 , \6500 , \9431 );
nor \U$20022 ( \20337 , \20335 , \20336 );
xnor \U$20023 ( \20338 , \20337 , \9123 );
and \U$20024 ( \20339 , \20333 , \20338 );
and \U$20025 ( \20340 , \20329 , \20338 );
or \U$20026 ( \20341 , \20334 , \20339 , \20340 );
and \U$20027 ( \20342 , \20325 , \20341 );
and \U$20028 ( \20343 , \7177 , \8896 );
and \U$20029 ( \20344 , \7005 , \8894 );
nor \U$20030 ( \20345 , \20343 , \20344 );
xnor \U$20031 ( \20346 , \20345 , \8525 );
and \U$20032 ( \20347 , \8127 , \8334 );
and \U$20033 ( \20348 , \7703 , \8332 );
nor \U$20034 ( \20349 , \20347 , \20348 );
xnor \U$20035 ( \20350 , \20349 , \8016 );
and \U$20036 ( \20351 , \20346 , \20350 );
and \U$20037 ( \20352 , \8378 , \7767 );
and \U$20038 ( \20353 , \8373 , \7765 );
nor \U$20039 ( \20354 , \20352 , \20353 );
xnor \U$20040 ( \20355 , \20354 , \7518 );
and \U$20041 ( \20356 , \20350 , \20355 );
and \U$20042 ( \20357 , \20346 , \20355 );
or \U$20043 ( \20358 , \20351 , \20356 , \20357 );
and \U$20044 ( \20359 , \20341 , \20358 );
and \U$20045 ( \20360 , \20325 , \20358 );
or \U$20046 ( \20361 , \20342 , \20359 , \20360 );
xor \U$20047 ( \20362 , \20236 , \20240 );
xor \U$20048 ( \20363 , \20362 , \20245 );
xor \U$20049 ( \20364 , \20198 , \20202 );
xor \U$20050 ( \20365 , \20364 , \20205 );
and \U$20051 ( \20366 , \20363 , \20365 );
xor \U$20052 ( \20367 , \20253 , \20257 );
xor \U$20053 ( \20368 , \20367 , \20262 );
and \U$20054 ( \20369 , \20365 , \20368 );
and \U$20055 ( \20370 , \20363 , \20368 );
or \U$20056 ( \20371 , \20366 , \20369 , \20370 );
and \U$20057 ( \20372 , \20361 , \20371 );
xor \U$20058 ( \20373 , \20271 , \20273 );
xor \U$20059 ( \20374 , \20373 , \20276 );
and \U$20060 ( \20375 , \20371 , \20374 );
and \U$20061 ( \20376 , \20361 , \20374 );
or \U$20062 ( \20377 , \20372 , \20375 , \20376 );
xor \U$20063 ( \20378 , \20220 , \20268 );
xor \U$20064 ( \20379 , \20378 , \20279 );
and \U$20065 ( \20380 , \20377 , \20379 );
xor \U$20066 ( \20381 , \20284 , \20286 );
xor \U$20067 ( \20382 , \20381 , \20288 );
and \U$20068 ( \20383 , \20379 , \20382 );
and \U$20069 ( \20384 , \20377 , \20382 );
or \U$20070 ( \20385 , \20380 , \20383 , \20384 );
xor \U$20071 ( \20386 , \20149 , \20159 );
xor \U$20072 ( \20387 , \20386 , \20165 );
and \U$20073 ( \20388 , \20385 , \20387 );
xor \U$20074 ( \20389 , \20282 , \20291 );
xor \U$20075 ( \20390 , \20389 , \20294 );
and \U$20076 ( \20391 , \20387 , \20390 );
and \U$20077 ( \20392 , \20385 , \20390 );
or \U$20078 ( \20393 , \20388 , \20391 , \20392 );
and \U$20079 ( \20394 , \20309 , \20393 );
xor \U$20080 ( \20395 , \20309 , \20393 );
xor \U$20081 ( \20396 , \20385 , \20387 );
xor \U$20082 ( \20397 , \20396 , \20390 );
and \U$20083 ( \20398 , \6148 , \10814 );
and \U$20084 ( \20399 , \5776 , \10811 );
nor \U$20085 ( \20400 , \20398 , \20399 );
xnor \U$20086 ( \20401 , \20400 , \9759 );
and \U$20087 ( \20402 , \6500 , \10001 );
and \U$20088 ( \20403 , \6157 , \9999 );
nor \U$20089 ( \20404 , \20402 , \20403 );
xnor \U$20090 ( \20405 , \20404 , \9762 );
and \U$20091 ( \20406 , \20401 , \20405 );
and \U$20092 ( \20407 , \20405 , \5405 );
and \U$20093 ( \20408 , \20401 , \5405 );
or \U$20094 ( \20409 , \20406 , \20407 , \20408 );
and \U$20095 ( \20410 , \8697 , \7767 );
and \U$20096 ( \20411 , \8378 , \7765 );
nor \U$20097 ( \20412 , \20410 , \20411 );
xnor \U$20098 ( \20413 , \20412 , \7518 );
and \U$20099 ( \20414 , \9550 , \7238 );
and \U$20100 ( \20415 , \8981 , \7236 );
nor \U$20101 ( \20416 , \20414 , \20415 );
xnor \U$20102 ( \20417 , \20416 , \6978 );
and \U$20103 ( \20418 , \20413 , \20417 );
and \U$20104 ( \20419 , \10161 , \6744 );
and \U$20105 ( \20420 , \9558 , \6742 );
nor \U$20106 ( \20421 , \20419 , \20420 );
xnor \U$20107 ( \20422 , \20421 , \6429 );
and \U$20108 ( \20423 , \20417 , \20422 );
and \U$20109 ( \20424 , \20413 , \20422 );
or \U$20110 ( \20425 , \20418 , \20423 , \20424 );
and \U$20111 ( \20426 , \20409 , \20425 );
and \U$20112 ( \20427 , \7005 , \9433 );
and \U$20113 ( \20428 , \6702 , \9431 );
nor \U$20114 ( \20429 , \20427 , \20428 );
xnor \U$20115 ( \20430 , \20429 , \9123 );
and \U$20116 ( \20431 , \7703 , \8896 );
and \U$20117 ( \20432 , \7177 , \8894 );
nor \U$20118 ( \20433 , \20431 , \20432 );
xnor \U$20119 ( \20434 , \20433 , \8525 );
and \U$20120 ( \20435 , \20430 , \20434 );
and \U$20121 ( \20436 , \8373 , \8334 );
and \U$20122 ( \20437 , \8127 , \8332 );
nor \U$20123 ( \20438 , \20436 , \20437 );
xnor \U$20124 ( \20439 , \20438 , \8016 );
and \U$20125 ( \20440 , \20434 , \20439 );
and \U$20126 ( \20441 , \20430 , \20439 );
or \U$20127 ( \20442 , \20435 , \20440 , \20441 );
and \U$20128 ( \20443 , \20425 , \20442 );
and \U$20129 ( \20444 , \20409 , \20442 );
or \U$20130 ( \20445 , \20426 , \20443 , \20444 );
and \U$20131 ( \20446 , \10967 , \5646 );
and \U$20132 ( \20447 , \10347 , \5644 );
nor \U$20133 ( \20448 , \20446 , \20447 );
xnor \U$20134 ( \20449 , \20448 , \5405 );
xor \U$20135 ( \20450 , \20313 , \20317 );
xor \U$20136 ( \20451 , \20450 , \20322 );
and \U$20137 ( \20452 , \20449 , \20451 );
xor \U$20138 ( \20453 , \20346 , \20350 );
xor \U$20139 ( \20454 , \20453 , \20355 );
and \U$20140 ( \20455 , \20451 , \20454 );
and \U$20141 ( \20456 , \20449 , \20454 );
or \U$20142 ( \20457 , \20452 , \20455 , \20456 );
and \U$20143 ( \20458 , \20445 , \20457 );
xor \U$20144 ( \20459 , \20224 , \20228 );
xor \U$20145 ( \20460 , \20459 , \4992 );
and \U$20146 ( \20461 , \20457 , \20460 );
and \U$20147 ( \20462 , \20445 , \20460 );
or \U$20148 ( \20463 , \20458 , \20461 , \20462 );
xor \U$20149 ( \20464 , \20325 , \20341 );
xor \U$20150 ( \20465 , \20464 , \20358 );
xor \U$20151 ( \20466 , \20363 , \20365 );
xor \U$20152 ( \20467 , \20466 , \20368 );
and \U$20153 ( \20468 , \20465 , \20467 );
and \U$20154 ( \20469 , \20463 , \20468 );
xor \U$20155 ( \20470 , \20208 , \20212 );
xor \U$20156 ( \20471 , \20470 , \20217 );
and \U$20157 ( \20472 , \20468 , \20471 );
and \U$20158 ( \20473 , \20463 , \20471 );
or \U$20159 ( \20474 , \20469 , \20472 , \20473 );
xor \U$20160 ( \20475 , \20232 , \20248 );
xor \U$20161 ( \20476 , \20475 , \20265 );
xor \U$20162 ( \20477 , \20361 , \20371 );
xor \U$20163 ( \20478 , \20477 , \20374 );
and \U$20164 ( \20479 , \20476 , \20478 );
and \U$20165 ( \20480 , \20474 , \20479 );
xor \U$20166 ( \20481 , \20377 , \20379 );
xor \U$20167 ( \20482 , \20481 , \20382 );
and \U$20168 ( \20483 , \20479 , \20482 );
and \U$20169 ( \20484 , \20474 , \20482 );
or \U$20170 ( \20485 , \20480 , \20483 , \20484 );
and \U$20171 ( \20486 , \20397 , \20485 );
xor \U$20172 ( \20487 , \20397 , \20485 );
xor \U$20173 ( \20488 , \20474 , \20479 );
xor \U$20174 ( \20489 , \20488 , \20482 );
and \U$20175 ( \20490 , \8127 , \8896 );
and \U$20176 ( \20491 , \7703 , \8894 );
nor \U$20177 ( \20492 , \20490 , \20491 );
xnor \U$20178 ( \20493 , \20492 , \8525 );
and \U$20179 ( \20494 , \8378 , \8334 );
and \U$20180 ( \20495 , \8373 , \8332 );
nor \U$20181 ( \20496 , \20494 , \20495 );
xnor \U$20182 ( \20497 , \20496 , \8016 );
and \U$20183 ( \20498 , \20493 , \20497 );
and \U$20184 ( \20499 , \8981 , \7767 );
and \U$20185 ( \20500 , \8697 , \7765 );
nor \U$20186 ( \20501 , \20499 , \20500 );
xnor \U$20187 ( \20502 , \20501 , \7518 );
and \U$20188 ( \20503 , \20497 , \20502 );
and \U$20189 ( \20504 , \20493 , \20502 );
or \U$20190 ( \20505 , \20498 , \20503 , \20504 );
and \U$20191 ( \20506 , \6157 , \10814 );
and \U$20192 ( \20507 , \6148 , \10811 );
nor \U$20193 ( \20508 , \20506 , \20507 );
xnor \U$20194 ( \20509 , \20508 , \9759 );
and \U$20195 ( \20510 , \6702 , \10001 );
and \U$20196 ( \20511 , \6500 , \9999 );
nor \U$20197 ( \20512 , \20510 , \20511 );
xnor \U$20198 ( \20513 , \20512 , \9762 );
and \U$20199 ( \20514 , \20509 , \20513 );
and \U$20200 ( \20515 , \7177 , \9433 );
and \U$20201 ( \20516 , \7005 , \9431 );
nor \U$20202 ( \20517 , \20515 , \20516 );
xnor \U$20203 ( \20518 , \20517 , \9123 );
and \U$20204 ( \20519 , \20513 , \20518 );
and \U$20205 ( \20520 , \20509 , \20518 );
or \U$20206 ( \20521 , \20514 , \20519 , \20520 );
and \U$20207 ( \20522 , \20505 , \20521 );
and \U$20208 ( \20523 , \9558 , \7238 );
and \U$20209 ( \20524 , \9550 , \7236 );
nor \U$20210 ( \20525 , \20523 , \20524 );
xnor \U$20211 ( \20526 , \20525 , \6978 );
and \U$20212 ( \20527 , \10166 , \6744 );
and \U$20213 ( \20528 , \10161 , \6742 );
nor \U$20214 ( \20529 , \20527 , \20528 );
xnor \U$20215 ( \20530 , \20529 , \6429 );
and \U$20216 ( \20531 , \20526 , \20530 );
and \U$20217 ( \20532 , \10967 , \6235 );
and \U$20218 ( \20533 , \10347 , \6233 );
nor \U$20219 ( \20534 , \20532 , \20533 );
xnor \U$20220 ( \20535 , \20534 , \5895 );
and \U$20221 ( \20536 , \20530 , \20535 );
and \U$20222 ( \20537 , \20526 , \20535 );
or \U$20223 ( \20538 , \20531 , \20536 , \20537 );
and \U$20224 ( \20539 , \20521 , \20538 );
and \U$20225 ( \20540 , \20505 , \20538 );
or \U$20226 ( \20541 , \20522 , \20539 , \20540 );
and \U$20227 ( \20542 , \10347 , \6235 );
and \U$20228 ( \20543 , \10166 , \6233 );
nor \U$20229 ( \20544 , \20542 , \20543 );
xnor \U$20230 ( \20545 , \20544 , \5895 );
nand \U$20231 ( \20546 , \10967 , \5644 );
xnor \U$20232 ( \20547 , \20546 , \5405 );
and \U$20233 ( \20548 , \20545 , \20547 );
xor \U$20234 ( \20549 , \20413 , \20417 );
xor \U$20235 ( \20550 , \20549 , \20422 );
and \U$20236 ( \20551 , \20547 , \20550 );
and \U$20237 ( \20552 , \20545 , \20550 );
or \U$20238 ( \20553 , \20548 , \20551 , \20552 );
and \U$20239 ( \20554 , \20541 , \20553 );
xor \U$20240 ( \20555 , \20329 , \20333 );
xor \U$20241 ( \20556 , \20555 , \20338 );
and \U$20242 ( \20557 , \20553 , \20556 );
and \U$20243 ( \20558 , \20541 , \20556 );
or \U$20244 ( \20559 , \20554 , \20557 , \20558 );
xor \U$20245 ( \20560 , \20445 , \20457 );
xor \U$20246 ( \20561 , \20560 , \20460 );
and \U$20247 ( \20562 , \20559 , \20561 );
xor \U$20248 ( \20563 , \20465 , \20467 );
and \U$20249 ( \20564 , \20561 , \20563 );
and \U$20250 ( \20565 , \20559 , \20563 );
or \U$20251 ( \20566 , \20562 , \20564 , \20565 );
xor \U$20252 ( \20567 , \20463 , \20468 );
xor \U$20253 ( \20568 , \20567 , \20471 );
and \U$20254 ( \20569 , \20566 , \20568 );
xor \U$20255 ( \20570 , \20476 , \20478 );
and \U$20256 ( \20571 , \20568 , \20570 );
and \U$20257 ( \20572 , \20566 , \20570 );
or \U$20258 ( \20573 , \20569 , \20571 , \20572 );
and \U$20259 ( \20574 , \20489 , \20573 );
xor \U$20260 ( \20575 , \20489 , \20573 );
xor \U$20261 ( \20576 , \20566 , \20568 );
xor \U$20262 ( \20577 , \20576 , \20570 );
and \U$20263 ( \20578 , \7703 , \9433 );
and \U$20264 ( \20579 , \7177 , \9431 );
nor \U$20265 ( \20580 , \20578 , \20579 );
xnor \U$20266 ( \20581 , \20580 , \9123 );
and \U$20267 ( \20582 , \8373 , \8896 );
and \U$20268 ( \20583 , \8127 , \8894 );
nor \U$20269 ( \20584 , \20582 , \20583 );
xnor \U$20270 ( \20585 , \20584 , \8525 );
and \U$20271 ( \20586 , \20581 , \20585 );
and \U$20272 ( \20587 , \8697 , \8334 );
and \U$20273 ( \20588 , \8378 , \8332 );
nor \U$20274 ( \20589 , \20587 , \20588 );
xnor \U$20275 ( \20590 , \20589 , \8016 );
and \U$20276 ( \20591 , \20585 , \20590 );
and \U$20277 ( \20592 , \20581 , \20590 );
or \U$20278 ( \20593 , \20586 , \20591 , \20592 );
and \U$20279 ( \20594 , \6500 , \10814 );
and \U$20280 ( \20595 , \6157 , \10811 );
nor \U$20281 ( \20596 , \20594 , \20595 );
xnor \U$20282 ( \20597 , \20596 , \9759 );
and \U$20283 ( \20598 , \7005 , \10001 );
and \U$20284 ( \20599 , \6702 , \9999 );
nor \U$20285 ( \20600 , \20598 , \20599 );
xnor \U$20286 ( \20601 , \20600 , \9762 );
and \U$20287 ( \20602 , \20597 , \20601 );
and \U$20288 ( \20603 , \20601 , \5895 );
and \U$20289 ( \20604 , \20597 , \5895 );
or \U$20290 ( \20605 , \20602 , \20603 , \20604 );
and \U$20291 ( \20606 , \20593 , \20605 );
and \U$20292 ( \20607 , \9550 , \7767 );
and \U$20293 ( \20608 , \8981 , \7765 );
nor \U$20294 ( \20609 , \20607 , \20608 );
xnor \U$20295 ( \20610 , \20609 , \7518 );
and \U$20296 ( \20611 , \10161 , \7238 );
and \U$20297 ( \20612 , \9558 , \7236 );
nor \U$20298 ( \20613 , \20611 , \20612 );
xnor \U$20299 ( \20614 , \20613 , \6978 );
and \U$20300 ( \20615 , \20610 , \20614 );
and \U$20301 ( \20616 , \10347 , \6744 );
and \U$20302 ( \20617 , \10166 , \6742 );
nor \U$20303 ( \20618 , \20616 , \20617 );
xnor \U$20304 ( \20619 , \20618 , \6429 );
and \U$20305 ( \20620 , \20614 , \20619 );
and \U$20306 ( \20621 , \20610 , \20619 );
or \U$20307 ( \20622 , \20615 , \20620 , \20621 );
and \U$20308 ( \20623 , \20605 , \20622 );
and \U$20309 ( \20624 , \20593 , \20622 );
or \U$20310 ( \20625 , \20606 , \20623 , \20624 );
xor \U$20311 ( \20626 , \20493 , \20497 );
xor \U$20312 ( \20627 , \20626 , \20502 );
xor \U$20313 ( \20628 , \20509 , \20513 );
xor \U$20314 ( \20629 , \20628 , \20518 );
and \U$20315 ( \20630 , \20627 , \20629 );
xor \U$20316 ( \20631 , \20526 , \20530 );
xor \U$20317 ( \20632 , \20631 , \20535 );
and \U$20318 ( \20633 , \20629 , \20632 );
and \U$20319 ( \20634 , \20627 , \20632 );
or \U$20320 ( \20635 , \20630 , \20633 , \20634 );
and \U$20321 ( \20636 , \20625 , \20635 );
xor \U$20322 ( \20637 , \20430 , \20434 );
xor \U$20323 ( \20638 , \20637 , \20439 );
and \U$20324 ( \20639 , \20635 , \20638 );
and \U$20325 ( \20640 , \20625 , \20638 );
or \U$20326 ( \20641 , \20636 , \20639 , \20640 );
xor \U$20327 ( \20642 , \20401 , \20405 );
xor \U$20328 ( \20643 , \20642 , \5405 );
xor \U$20329 ( \20644 , \20505 , \20521 );
xor \U$20330 ( \20645 , \20644 , \20538 );
and \U$20331 ( \20646 , \20643 , \20645 );
xor \U$20332 ( \20647 , \20545 , \20547 );
xor \U$20333 ( \20648 , \20647 , \20550 );
and \U$20334 ( \20649 , \20645 , \20648 );
and \U$20335 ( \20650 , \20643 , \20648 );
or \U$20336 ( \20651 , \20646 , \20649 , \20650 );
and \U$20337 ( \20652 , \20641 , \20651 );
xor \U$20338 ( \20653 , \20449 , \20451 );
xor \U$20339 ( \20654 , \20653 , \20454 );
and \U$20340 ( \20655 , \20651 , \20654 );
and \U$20341 ( \20656 , \20641 , \20654 );
or \U$20342 ( \20657 , \20652 , \20655 , \20656 );
xor \U$20343 ( \20658 , \20409 , \20425 );
xor \U$20344 ( \20659 , \20658 , \20442 );
xor \U$20345 ( \20660 , \20541 , \20553 );
xor \U$20346 ( \20661 , \20660 , \20556 );
and \U$20347 ( \20662 , \20659 , \20661 );
and \U$20348 ( \20663 , \20657 , \20662 );
xor \U$20349 ( \20664 , \20559 , \20561 );
xor \U$20350 ( \20665 , \20664 , \20563 );
and \U$20351 ( \20666 , \20662 , \20665 );
and \U$20352 ( \20667 , \20657 , \20665 );
or \U$20353 ( \20668 , \20663 , \20666 , \20667 );
and \U$20354 ( \20669 , \20577 , \20668 );
xor \U$20355 ( \20670 , \20577 , \20668 );
xor \U$20356 ( \20671 , \20657 , \20662 );
xor \U$20357 ( \20672 , \20671 , \20665 );
and \U$20358 ( \20673 , \6702 , \10814 );
and \U$20359 ( \20674 , \6500 , \10811 );
nor \U$20360 ( \20675 , \20673 , \20674 );
xnor \U$20361 ( \20676 , \20675 , \9759 );
and \U$20362 ( \20677 , \7177 , \10001 );
and \U$20363 ( \20678 , \7005 , \9999 );
nor \U$20364 ( \20679 , \20677 , \20678 );
xnor \U$20365 ( \20680 , \20679 , \9762 );
and \U$20366 ( \20681 , \20676 , \20680 );
and \U$20367 ( \20682 , \8127 , \9433 );
and \U$20368 ( \20683 , \7703 , \9431 );
nor \U$20369 ( \20684 , \20682 , \20683 );
xnor \U$20370 ( \20685 , \20684 , \9123 );
and \U$20371 ( \20686 , \20680 , \20685 );
and \U$20372 ( \20687 , \20676 , \20685 );
or \U$20373 ( \20688 , \20681 , \20686 , \20687 );
and \U$20374 ( \20689 , \8378 , \8896 );
and \U$20375 ( \20690 , \8373 , \8894 );
nor \U$20376 ( \20691 , \20689 , \20690 );
xnor \U$20377 ( \20692 , \20691 , \8525 );
and \U$20378 ( \20693 , \8981 , \8334 );
and \U$20379 ( \20694 , \8697 , \8332 );
nor \U$20380 ( \20695 , \20693 , \20694 );
xnor \U$20381 ( \20696 , \20695 , \8016 );
and \U$20382 ( \20697 , \20692 , \20696 );
and \U$20383 ( \20698 , \9558 , \7767 );
and \U$20384 ( \20699 , \9550 , \7765 );
nor \U$20385 ( \20700 , \20698 , \20699 );
xnor \U$20386 ( \20701 , \20700 , \7518 );
and \U$20387 ( \20702 , \20696 , \20701 );
and \U$20388 ( \20703 , \20692 , \20701 );
or \U$20389 ( \20704 , \20697 , \20702 , \20703 );
and \U$20390 ( \20705 , \20688 , \20704 );
and \U$20391 ( \20706 , \10166 , \7238 );
and \U$20392 ( \20707 , \10161 , \7236 );
nor \U$20393 ( \20708 , \20706 , \20707 );
xnor \U$20394 ( \20709 , \20708 , \6978 );
and \U$20395 ( \20710 , \10967 , \6744 );
and \U$20396 ( \20711 , \10347 , \6742 );
nor \U$20397 ( \20712 , \20710 , \20711 );
xnor \U$20398 ( \20713 , \20712 , \6429 );
and \U$20399 ( \20714 , \20709 , \20713 );
and \U$20400 ( \20715 , \20704 , \20714 );
and \U$20401 ( \20716 , \20688 , \20714 );
or \U$20402 ( \20717 , \20705 , \20715 , \20716 );
nand \U$20403 ( \20718 , \10967 , \6233 );
xnor \U$20404 ( \20719 , \20718 , \5895 );
xor \U$20405 ( \20720 , \20581 , \20585 );
xor \U$20406 ( \20721 , \20720 , \20590 );
and \U$20407 ( \20722 , \20719 , \20721 );
xor \U$20408 ( \20723 , \20610 , \20614 );
xor \U$20409 ( \20724 , \20723 , \20619 );
and \U$20410 ( \20725 , \20721 , \20724 );
and \U$20411 ( \20726 , \20719 , \20724 );
or \U$20412 ( \20727 , \20722 , \20725 , \20726 );
and \U$20413 ( \20728 , \20717 , \20727 );
xor \U$20414 ( \20729 , \20627 , \20629 );
xor \U$20415 ( \20730 , \20729 , \20632 );
and \U$20416 ( \20731 , \20727 , \20730 );
and \U$20417 ( \20732 , \20717 , \20730 );
or \U$20418 ( \20733 , \20728 , \20731 , \20732 );
xor \U$20419 ( \20734 , \20625 , \20635 );
xor \U$20420 ( \20735 , \20734 , \20638 );
and \U$20421 ( \20736 , \20733 , \20735 );
xor \U$20422 ( \20737 , \20643 , \20645 );
xor \U$20423 ( \20738 , \20737 , \20648 );
and \U$20424 ( \20739 , \20735 , \20738 );
and \U$20425 ( \20740 , \20733 , \20738 );
or \U$20426 ( \20741 , \20736 , \20739 , \20740 );
xor \U$20427 ( \20742 , \20641 , \20651 );
xor \U$20428 ( \20743 , \20742 , \20654 );
and \U$20429 ( \20744 , \20741 , \20743 );
xor \U$20430 ( \20745 , \20659 , \20661 );
and \U$20431 ( \20746 , \20743 , \20745 );
and \U$20432 ( \20747 , \20741 , \20745 );
or \U$20433 ( \20748 , \20744 , \20746 , \20747 );
and \U$20434 ( \20749 , \20672 , \20748 );
xor \U$20435 ( \20750 , \20672 , \20748 );
xor \U$20436 ( \20751 , \20741 , \20743 );
xor \U$20437 ( \20752 , \20751 , \20745 );
and \U$20438 ( \20753 , \10161 , \7767 );
and \U$20439 ( \20754 , \9558 , \7765 );
nor \U$20440 ( \20755 , \20753 , \20754 );
xnor \U$20441 ( \20756 , \20755 , \7518 );
and \U$20442 ( \20757 , \10347 , \7238 );
and \U$20443 ( \20758 , \10166 , \7236 );
nor \U$20444 ( \20759 , \20757 , \20758 );
xnor \U$20445 ( \20760 , \20759 , \6978 );
and \U$20446 ( \20761 , \20756 , \20760 );
nand \U$20447 ( \20762 , \10967 , \6742 );
xnor \U$20448 ( \20763 , \20762 , \6429 );
and \U$20449 ( \20764 , \20760 , \20763 );
and \U$20450 ( \20765 , \20756 , \20763 );
or \U$20451 ( \20766 , \20761 , \20764 , \20765 );
and \U$20452 ( \20767 , \7005 , \10814 );
and \U$20453 ( \20768 , \6702 , \10811 );
nor \U$20454 ( \20769 , \20767 , \20768 );
xnor \U$20455 ( \20770 , \20769 , \9759 );
and \U$20456 ( \20771 , \7703 , \10001 );
and \U$20457 ( \20772 , \7177 , \9999 );
nor \U$20458 ( \20773 , \20771 , \20772 );
xnor \U$20459 ( \20774 , \20773 , \9762 );
and \U$20460 ( \20775 , \20770 , \20774 );
and \U$20461 ( \20776 , \20774 , \6429 );
and \U$20462 ( \20777 , \20770 , \6429 );
or \U$20463 ( \20778 , \20775 , \20776 , \20777 );
and \U$20464 ( \20779 , \20766 , \20778 );
and \U$20465 ( \20780 , \8373 , \9433 );
and \U$20466 ( \20781 , \8127 , \9431 );
nor \U$20467 ( \20782 , \20780 , \20781 );
xnor \U$20468 ( \20783 , \20782 , \9123 );
and \U$20469 ( \20784 , \8697 , \8896 );
and \U$20470 ( \20785 , \8378 , \8894 );
nor \U$20471 ( \20786 , \20784 , \20785 );
xnor \U$20472 ( \20787 , \20786 , \8525 );
and \U$20473 ( \20788 , \20783 , \20787 );
and \U$20474 ( \20789 , \9550 , \8334 );
and \U$20475 ( \20790 , \8981 , \8332 );
nor \U$20476 ( \20791 , \20789 , \20790 );
xnor \U$20477 ( \20792 , \20791 , \8016 );
and \U$20478 ( \20793 , \20787 , \20792 );
and \U$20479 ( \20794 , \20783 , \20792 );
or \U$20480 ( \20795 , \20788 , \20793 , \20794 );
and \U$20481 ( \20796 , \20778 , \20795 );
and \U$20482 ( \20797 , \20766 , \20795 );
or \U$20483 ( \20798 , \20779 , \20796 , \20797 );
xor \U$20484 ( \20799 , \20676 , \20680 );
xor \U$20485 ( \20800 , \20799 , \20685 );
xor \U$20486 ( \20801 , \20692 , \20696 );
xor \U$20487 ( \20802 , \20801 , \20701 );
and \U$20488 ( \20803 , \20800 , \20802 );
xor \U$20489 ( \20804 , \20709 , \20713 );
and \U$20490 ( \20805 , \20802 , \20804 );
and \U$20491 ( \20806 , \20800 , \20804 );
or \U$20492 ( \20807 , \20803 , \20805 , \20806 );
and \U$20493 ( \20808 , \20798 , \20807 );
xor \U$20494 ( \20809 , \20597 , \20601 );
xor \U$20495 ( \20810 , \20809 , \5895 );
and \U$20496 ( \20811 , \20807 , \20810 );
and \U$20497 ( \20812 , \20798 , \20810 );
or \U$20498 ( \20813 , \20808 , \20811 , \20812 );
xor \U$20499 ( \20814 , \20688 , \20704 );
xor \U$20500 ( \20815 , \20814 , \20714 );
xor \U$20501 ( \20816 , \20719 , \20721 );
xor \U$20502 ( \20817 , \20816 , \20724 );
and \U$20503 ( \20818 , \20815 , \20817 );
and \U$20504 ( \20819 , \20813 , \20818 );
xor \U$20505 ( \20820 , \20593 , \20605 );
xor \U$20506 ( \20821 , \20820 , \20622 );
and \U$20507 ( \20822 , \20818 , \20821 );
and \U$20508 ( \20823 , \20813 , \20821 );
or \U$20509 ( \20824 , \20819 , \20822 , \20823 );
xor \U$20510 ( \20825 , \20733 , \20735 );
xor \U$20511 ( \20826 , \20825 , \20738 );
and \U$20512 ( \20827 , \20824 , \20826 );
and \U$20513 ( \20828 , \20752 , \20827 );
xor \U$20514 ( \20829 , \20752 , \20827 );
xor \U$20515 ( \20830 , \20824 , \20826 );
xor \U$20516 ( \20831 , \20813 , \20818 );
xor \U$20517 ( \20832 , \20831 , \20821 );
xor \U$20518 ( \20833 , \20717 , \20727 );
xor \U$20519 ( \20834 , \20833 , \20730 );
and \U$20520 ( \20835 , \20832 , \20834 );
and \U$20521 ( \20836 , \20830 , \20835 );
xor \U$20522 ( \20837 , \20830 , \20835 );
xor \U$20523 ( \20838 , \20832 , \20834 );
and \U$20524 ( \20839 , \7177 , \10814 );
and \U$20525 ( \20840 , \7005 , \10811 );
nor \U$20526 ( \20841 , \20839 , \20840 );
xnor \U$20527 ( \20842 , \20841 , \9759 );
and \U$20528 ( \20843 , \8127 , \10001 );
and \U$20529 ( \20844 , \7703 , \9999 );
nor \U$20530 ( \20845 , \20843 , \20844 );
xnor \U$20531 ( \20846 , \20845 , \9762 );
and \U$20532 ( \20847 , \20842 , \20846 );
and \U$20533 ( \20848 , \8378 , \9433 );
and \U$20534 ( \20849 , \8373 , \9431 );
nor \U$20535 ( \20850 , \20848 , \20849 );
xnor \U$20536 ( \20851 , \20850 , \9123 );
and \U$20537 ( \20852 , \20846 , \20851 );
and \U$20538 ( \20853 , \20842 , \20851 );
or \U$20539 ( \20854 , \20847 , \20852 , \20853 );
and \U$20540 ( \20855 , \8981 , \8896 );
and \U$20541 ( \20856 , \8697 , \8894 );
nor \U$20542 ( \20857 , \20855 , \20856 );
xnor \U$20543 ( \20858 , \20857 , \8525 );
and \U$20544 ( \20859 , \9558 , \8334 );
and \U$20545 ( \20860 , \9550 , \8332 );
nor \U$20546 ( \20861 , \20859 , \20860 );
xnor \U$20547 ( \20862 , \20861 , \8016 );
and \U$20548 ( \20863 , \20858 , \20862 );
and \U$20549 ( \20864 , \10166 , \7767 );
and \U$20550 ( \20865 , \10161 , \7765 );
nor \U$20551 ( \20866 , \20864 , \20865 );
xnor \U$20552 ( \20867 , \20866 , \7518 );
and \U$20553 ( \20868 , \20862 , \20867 );
and \U$20554 ( \20869 , \20858 , \20867 );
or \U$20555 ( \20870 , \20863 , \20868 , \20869 );
and \U$20556 ( \20871 , \20854 , \20870 );
xor \U$20557 ( \20872 , \20756 , \20760 );
xor \U$20558 ( \20873 , \20872 , \20763 );
and \U$20559 ( \20874 , \20870 , \20873 );
and \U$20560 ( \20875 , \20854 , \20873 );
or \U$20561 ( \20876 , \20871 , \20874 , \20875 );
xor \U$20562 ( \20877 , \20770 , \20774 );
xor \U$20563 ( \20878 , \20877 , \6429 );
xor \U$20564 ( \20879 , \20783 , \20787 );
xor \U$20565 ( \20880 , \20879 , \20792 );
and \U$20566 ( \20881 , \20878 , \20880 );
and \U$20567 ( \20882 , \20876 , \20881 );
xor \U$20568 ( \20883 , \20800 , \20802 );
xor \U$20569 ( \20884 , \20883 , \20804 );
and \U$20570 ( \20885 , \20881 , \20884 );
and \U$20571 ( \20886 , \20876 , \20884 );
or \U$20572 ( \20887 , \20882 , \20885 , \20886 );
xor \U$20573 ( \20888 , \20798 , \20807 );
xor \U$20574 ( \20889 , \20888 , \20810 );
and \U$20575 ( \20890 , \20887 , \20889 );
xor \U$20576 ( \20891 , \20815 , \20817 );
and \U$20577 ( \20892 , \20889 , \20891 );
and \U$20578 ( \20893 , \20887 , \20891 );
or \U$20579 ( \20894 , \20890 , \20892 , \20893 );
and \U$20580 ( \20895 , \20838 , \20894 );
xor \U$20581 ( \20896 , \20838 , \20894 );
xor \U$20582 ( \20897 , \20887 , \20889 );
xor \U$20583 ( \20898 , \20897 , \20891 );
and \U$20584 ( \20899 , \7703 , \10814 );
and \U$20585 ( \20900 , \7177 , \10811 );
nor \U$20586 ( \20901 , \20899 , \20900 );
xnor \U$20587 ( \20902 , \20901 , \9759 );
and \U$20588 ( \20903 , \8373 , \10001 );
and \U$20589 ( \20904 , \8127 , \9999 );
nor \U$20590 ( \20905 , \20903 , \20904 );
xnor \U$20591 ( \20906 , \20905 , \9762 );
and \U$20592 ( \20907 , \20902 , \20906 );
and \U$20593 ( \20908 , \20906 , \6978 );
and \U$20594 ( \20909 , \20902 , \6978 );
or \U$20595 ( \20910 , \20907 , \20908 , \20909 );
and \U$20596 ( \20911 , \8697 , \9433 );
and \U$20597 ( \20912 , \8378 , \9431 );
nor \U$20598 ( \20913 , \20911 , \20912 );
xnor \U$20599 ( \20914 , \20913 , \9123 );
and \U$20600 ( \20915 , \9550 , \8896 );
and \U$20601 ( \20916 , \8981 , \8894 );
nor \U$20602 ( \20917 , \20915 , \20916 );
xnor \U$20603 ( \20918 , \20917 , \8525 );
and \U$20604 ( \20919 , \20914 , \20918 );
and \U$20605 ( \20920 , \10161 , \8334 );
and \U$20606 ( \20921 , \9558 , \8332 );
nor \U$20607 ( \20922 , \20920 , \20921 );
xnor \U$20608 ( \20923 , \20922 , \8016 );
and \U$20609 ( \20924 , \20918 , \20923 );
and \U$20610 ( \20925 , \20914 , \20923 );
or \U$20611 ( \20926 , \20919 , \20924 , \20925 );
and \U$20612 ( \20927 , \20910 , \20926 );
and \U$20613 ( \20928 , \10967 , \7238 );
and \U$20614 ( \20929 , \10347 , \7236 );
nor \U$20615 ( \20930 , \20928 , \20929 );
xnor \U$20616 ( \20931 , \20930 , \6978 );
and \U$20617 ( \20932 , \20926 , \20931 );
and \U$20618 ( \20933 , \20910 , \20931 );
or \U$20619 ( \20934 , \20927 , \20932 , \20933 );
xor \U$20620 ( \20935 , \20854 , \20870 );
xor \U$20621 ( \20936 , \20935 , \20873 );
and \U$20622 ( \20937 , \20934 , \20936 );
xor \U$20623 ( \20938 , \20878 , \20880 );
and \U$20624 ( \20939 , \20936 , \20938 );
and \U$20625 ( \20940 , \20934 , \20938 );
or \U$20626 ( \20941 , \20937 , \20939 , \20940 );
xor \U$20627 ( \20942 , \20766 , \20778 );
xor \U$20628 ( \20943 , \20942 , \20795 );
and \U$20629 ( \20944 , \20941 , \20943 );
xor \U$20630 ( \20945 , \20876 , \20881 );
xor \U$20631 ( \20946 , \20945 , \20884 );
and \U$20632 ( \20947 , \20943 , \20946 );
and \U$20633 ( \20948 , \20941 , \20946 );
or \U$20634 ( \20949 , \20944 , \20947 , \20948 );
and \U$20635 ( \20950 , \20898 , \20949 );
xor \U$20636 ( \20951 , \20898 , \20949 );
xor \U$20637 ( \20952 , \20941 , \20943 );
xor \U$20638 ( \20953 , \20952 , \20946 );
and \U$20639 ( \20954 , \9558 , \8896 );
and \U$20640 ( \20955 , \9550 , \8894 );
nor \U$20641 ( \20956 , \20954 , \20955 );
xnor \U$20642 ( \20957 , \20956 , \8525 );
and \U$20643 ( \20958 , \10166 , \8334 );
and \U$20644 ( \20959 , \10161 , \8332 );
nor \U$20645 ( \20960 , \20958 , \20959 );
xnor \U$20646 ( \20961 , \20960 , \8016 );
and \U$20647 ( \20962 , \20957 , \20961 );
and \U$20648 ( \20963 , \10967 , \7767 );
and \U$20649 ( \20964 , \10347 , \7765 );
nor \U$20650 ( \20965 , \20963 , \20964 );
xnor \U$20651 ( \20966 , \20965 , \7518 );
and \U$20652 ( \20967 , \20961 , \20966 );
and \U$20653 ( \20968 , \20957 , \20966 );
or \U$20654 ( \20969 , \20962 , \20967 , \20968 );
and \U$20655 ( \20970 , \8127 , \10814 );
and \U$20656 ( \20971 , \7703 , \10811 );
nor \U$20657 ( \20972 , \20970 , \20971 );
xnor \U$20658 ( \20973 , \20972 , \9759 );
and \U$20659 ( \20974 , \8378 , \10001 );
and \U$20660 ( \20975 , \8373 , \9999 );
nor \U$20661 ( \20976 , \20974 , \20975 );
xnor \U$20662 ( \20977 , \20976 , \9762 );
and \U$20663 ( \20978 , \20973 , \20977 );
and \U$20664 ( \20979 , \8981 , \9433 );
and \U$20665 ( \20980 , \8697 , \9431 );
nor \U$20666 ( \20981 , \20979 , \20980 );
xnor \U$20667 ( \20982 , \20981 , \9123 );
and \U$20668 ( \20983 , \20977 , \20982 );
and \U$20669 ( \20984 , \20973 , \20982 );
or \U$20670 ( \20985 , \20978 , \20983 , \20984 );
and \U$20671 ( \20986 , \20969 , \20985 );
and \U$20672 ( \20987 , \10347 , \7767 );
and \U$20673 ( \20988 , \10166 , \7765 );
nor \U$20674 ( \20989 , \20987 , \20988 );
xnor \U$20675 ( \20990 , \20989 , \7518 );
and \U$20676 ( \20991 , \20985 , \20990 );
and \U$20677 ( \20992 , \20969 , \20990 );
or \U$20678 ( \20993 , \20986 , \20991 , \20992 );
nand \U$20679 ( \20994 , \10967 , \7236 );
xnor \U$20680 ( \20995 , \20994 , \6978 );
xor \U$20681 ( \20996 , \20902 , \20906 );
xor \U$20682 ( \20997 , \20996 , \6978 );
and \U$20683 ( \20998 , \20995 , \20997 );
xor \U$20684 ( \20999 , \20914 , \20918 );
xor \U$20685 ( \21000 , \20999 , \20923 );
and \U$20686 ( \21001 , \20997 , \21000 );
and \U$20687 ( \21002 , \20995 , \21000 );
or \U$20688 ( \21003 , \20998 , \21001 , \21002 );
and \U$20689 ( \21004 , \20993 , \21003 );
xor \U$20690 ( \21005 , \20858 , \20862 );
xor \U$20691 ( \21006 , \21005 , \20867 );
and \U$20692 ( \21007 , \21003 , \21006 );
and \U$20693 ( \21008 , \20993 , \21006 );
or \U$20694 ( \21009 , \21004 , \21007 , \21008 );
xor \U$20695 ( \21010 , \20842 , \20846 );
xor \U$20696 ( \21011 , \21010 , \20851 );
xor \U$20697 ( \21012 , \20910 , \20926 );
xor \U$20698 ( \21013 , \21012 , \20931 );
and \U$20699 ( \21014 , \21011 , \21013 );
and \U$20700 ( \21015 , \21009 , \21014 );
xor \U$20701 ( \21016 , \20934 , \20936 );
xor \U$20702 ( \21017 , \21016 , \20938 );
and \U$20703 ( \21018 , \21014 , \21017 );
and \U$20704 ( \21019 , \21009 , \21017 );
or \U$20705 ( \21020 , \21015 , \21018 , \21019 );
and \U$20706 ( \21021 , \20953 , \21020 );
xor \U$20707 ( \21022 , \20953 , \21020 );
xor \U$20708 ( \21023 , \21009 , \21014 );
xor \U$20709 ( \21024 , \21023 , \21017 );
and \U$20710 ( \21025 , \9550 , \9433 );
and \U$20711 ( \21026 , \8981 , \9431 );
nor \U$20712 ( \21027 , \21025 , \21026 );
xnor \U$20713 ( \21028 , \21027 , \9123 );
and \U$20714 ( \21029 , \10161 , \8896 );
and \U$20715 ( \21030 , \9558 , \8894 );
nor \U$20716 ( \21031 , \21029 , \21030 );
xnor \U$20717 ( \21032 , \21031 , \8525 );
and \U$20718 ( \21033 , \21028 , \21032 );
and \U$20719 ( \21034 , \10347 , \8334 );
and \U$20720 ( \21035 , \10166 , \8332 );
nor \U$20721 ( \21036 , \21034 , \21035 );
xnor \U$20722 ( \21037 , \21036 , \8016 );
and \U$20723 ( \21038 , \21032 , \21037 );
and \U$20724 ( \21039 , \21028 , \21037 );
or \U$20725 ( \21040 , \21033 , \21038 , \21039 );
and \U$20726 ( \21041 , \8373 , \10814 );
and \U$20727 ( \21042 , \8127 , \10811 );
nor \U$20728 ( \21043 , \21041 , \21042 );
xnor \U$20729 ( \21044 , \21043 , \9759 );
and \U$20730 ( \21045 , \8697 , \10001 );
and \U$20731 ( \21046 , \8378 , \9999 );
nor \U$20732 ( \21047 , \21045 , \21046 );
xnor \U$20733 ( \21048 , \21047 , \9762 );
and \U$20734 ( \21049 , \21044 , \21048 );
and \U$20735 ( \21050 , \21048 , \7518 );
and \U$20736 ( \21051 , \21044 , \7518 );
or \U$20737 ( \21052 , \21049 , \21050 , \21051 );
and \U$20738 ( \21053 , \21040 , \21052 );
xor \U$20739 ( \21054 , \20957 , \20961 );
xor \U$20740 ( \21055 , \21054 , \20966 );
and \U$20741 ( \21056 , \21052 , \21055 );
and \U$20742 ( \21057 , \21040 , \21055 );
or \U$20743 ( \21058 , \21053 , \21056 , \21057 );
xor \U$20744 ( \21059 , \20969 , \20985 );
xor \U$20745 ( \21060 , \21059 , \20990 );
and \U$20746 ( \21061 , \21058 , \21060 );
xor \U$20747 ( \21062 , \20995 , \20997 );
xor \U$20748 ( \21063 , \21062 , \21000 );
and \U$20749 ( \21064 , \21060 , \21063 );
and \U$20750 ( \21065 , \21058 , \21063 );
or \U$20751 ( \21066 , \21061 , \21064 , \21065 );
xor \U$20752 ( \21067 , \20993 , \21003 );
xor \U$20753 ( \21068 , \21067 , \21006 );
and \U$20754 ( \21069 , \21066 , \21068 );
xor \U$20755 ( \21070 , \21011 , \21013 );
and \U$20756 ( \21071 , \21068 , \21070 );
and \U$20757 ( \21072 , \21066 , \21070 );
or \U$20758 ( \21073 , \21069 , \21071 , \21072 );
and \U$20759 ( \21074 , \21024 , \21073 );
xor \U$20760 ( \21075 , \21024 , \21073 );
xor \U$20761 ( \21076 , \21066 , \21068 );
xor \U$20762 ( \21077 , \21076 , \21070 );
and \U$20763 ( \21078 , \8378 , \10814 );
and \U$20764 ( \21079 , \8373 , \10811 );
nor \U$20765 ( \21080 , \21078 , \21079 );
xnor \U$20766 ( \21081 , \21080 , \9759 );
and \U$20767 ( \21082 , \8981 , \10001 );
and \U$20768 ( \21083 , \8697 , \9999 );
nor \U$20769 ( \21084 , \21082 , \21083 );
xnor \U$20770 ( \21085 , \21084 , \9762 );
and \U$20771 ( \21086 , \21081 , \21085 );
and \U$20772 ( \21087 , \9558 , \9433 );
and \U$20773 ( \21088 , \9550 , \9431 );
nor \U$20774 ( \21089 , \21087 , \21088 );
xnor \U$20775 ( \21090 , \21089 , \9123 );
and \U$20776 ( \21091 , \21085 , \21090 );
and \U$20777 ( \21092 , \21081 , \21090 );
or \U$20778 ( \21093 , \21086 , \21091 , \21092 );
nand \U$20779 ( \21094 , \10967 , \7765 );
xnor \U$20780 ( \21095 , \21094 , \7518 );
and \U$20781 ( \21096 , \21093 , \21095 );
xor \U$20782 ( \21097 , \21028 , \21032 );
xor \U$20783 ( \21098 , \21097 , \21037 );
and \U$20784 ( \21099 , \21095 , \21098 );
and \U$20785 ( \21100 , \21093 , \21098 );
or \U$20786 ( \21101 , \21096 , \21099 , \21100 );
xor \U$20787 ( \21102 , \20973 , \20977 );
xor \U$20788 ( \21103 , \21102 , \20982 );
and \U$20789 ( \21104 , \21101 , \21103 );
xor \U$20790 ( \21105 , \21040 , \21052 );
xor \U$20791 ( \21106 , \21105 , \21055 );
and \U$20792 ( \21107 , \21103 , \21106 );
and \U$20793 ( \21108 , \21101 , \21106 );
or \U$20794 ( \21109 , \21104 , \21107 , \21108 );
xor \U$20795 ( \21110 , \21058 , \21060 );
xor \U$20796 ( \21111 , \21110 , \21063 );
and \U$20797 ( \21112 , \21109 , \21111 );
and \U$20798 ( \21113 , \21077 , \21112 );
xor \U$20799 ( \21114 , \21077 , \21112 );
xor \U$20800 ( \21115 , \21109 , \21111 );
and \U$20801 ( \21116 , \10161 , \9433 );
and \U$20802 ( \21117 , \9558 , \9431 );
nor \U$20803 ( \21118 , \21116 , \21117 );
xnor \U$20804 ( \21119 , \21118 , \9123 );
and \U$20805 ( \21120 , \10347 , \8896 );
and \U$20806 ( \21121 , \10166 , \8894 );
nor \U$20807 ( \21122 , \21120 , \21121 );
xnor \U$20808 ( \21123 , \21122 , \8525 );
and \U$20809 ( \21124 , \21119 , \21123 );
nand \U$20810 ( \21125 , \10967 , \8332 );
xnor \U$20811 ( \21126 , \21125 , \8016 );
and \U$20812 ( \21127 , \21123 , \21126 );
and \U$20813 ( \21128 , \21119 , \21126 );
or \U$20814 ( \21129 , \21124 , \21127 , \21128 );
and \U$20815 ( \21130 , \8697 , \10814 );
and \U$20816 ( \21131 , \8378 , \10811 );
nor \U$20817 ( \21132 , \21130 , \21131 );
xnor \U$20818 ( \21133 , \21132 , \9759 );
and \U$20819 ( \21134 , \9550 , \10001 );
and \U$20820 ( \21135 , \8981 , \9999 );
nor \U$20821 ( \21136 , \21134 , \21135 );
xnor \U$20822 ( \21137 , \21136 , \9762 );
and \U$20823 ( \21138 , \21133 , \21137 );
and \U$20824 ( \21139 , \21137 , \8016 );
and \U$20825 ( \21140 , \21133 , \8016 );
or \U$20826 ( \21141 , \21138 , \21139 , \21140 );
and \U$20827 ( \21142 , \21129 , \21141 );
and \U$20828 ( \21143 , \10166 , \8896 );
and \U$20829 ( \21144 , \10161 , \8894 );
nor \U$20830 ( \21145 , \21143 , \21144 );
xnor \U$20831 ( \21146 , \21145 , \8525 );
and \U$20832 ( \21147 , \21141 , \21146 );
and \U$20833 ( \21148 , \21129 , \21146 );
or \U$20834 ( \21149 , \21142 , \21147 , \21148 );
and \U$20835 ( \21150 , \10967 , \8334 );
and \U$20836 ( \21151 , \10347 , \8332 );
nor \U$20837 ( \21152 , \21150 , \21151 );
xnor \U$20838 ( \21153 , \21152 , \8016 );
xor \U$20839 ( \21154 , \21081 , \21085 );
xor \U$20840 ( \21155 , \21154 , \21090 );
and \U$20841 ( \21156 , \21153 , \21155 );
and \U$20842 ( \21157 , \21149 , \21156 );
xor \U$20843 ( \21158 , \21044 , \21048 );
xor \U$20844 ( \21159 , \21158 , \7518 );
and \U$20845 ( \21160 , \21156 , \21159 );
and \U$20846 ( \21161 , \21149 , \21159 );
or \U$20847 ( \21162 , \21157 , \21160 , \21161 );
xor \U$20848 ( \21163 , \21101 , \21103 );
xor \U$20849 ( \21164 , \21163 , \21106 );
and \U$20850 ( \21165 , \21162 , \21164 );
and \U$20851 ( \21166 , \21115 , \21165 );
xor \U$20852 ( \21167 , \21115 , \21165 );
xor \U$20853 ( \21168 , \21162 , \21164 );
xor \U$20854 ( \21169 , \21093 , \21095 );
xor \U$20855 ( \21170 , \21169 , \21098 );
xor \U$20856 ( \21171 , \21149 , \21156 );
xor \U$20857 ( \21172 , \21171 , \21159 );
and \U$20858 ( \21173 , \21170 , \21172 );
and \U$20859 ( \21174 , \21168 , \21173 );
xor \U$20860 ( \21175 , \21168 , \21173 );
xor \U$20861 ( \21176 , \21170 , \21172 );
and \U$20862 ( \21177 , \8981 , \10814 );
and \U$20863 ( \21178 , \8697 , \10811 );
nor \U$20864 ( \21179 , \21177 , \21178 );
xnor \U$20865 ( \21180 , \21179 , \9759 );
and \U$20866 ( \21181 , \9558 , \10001 );
and \U$20867 ( \21182 , \9550 , \9999 );
nor \U$20868 ( \21183 , \21181 , \21182 );
xnor \U$20869 ( \21184 , \21183 , \9762 );
and \U$20870 ( \21185 , \21180 , \21184 );
and \U$20871 ( \21186 , \10166 , \9433 );
and \U$20872 ( \21187 , \10161 , \9431 );
nor \U$20873 ( \21188 , \21186 , \21187 );
xnor \U$20874 ( \21189 , \21188 , \9123 );
and \U$20875 ( \21190 , \21184 , \21189 );
and \U$20876 ( \21191 , \21180 , \21189 );
or \U$20877 ( \21192 , \21185 , \21190 , \21191 );
xor \U$20878 ( \21193 , \21119 , \21123 );
xor \U$20879 ( \21194 , \21193 , \21126 );
and \U$20880 ( \21195 , \21192 , \21194 );
xor \U$20881 ( \21196 , \21133 , \21137 );
xor \U$20882 ( \21197 , \21196 , \8016 );
and \U$20883 ( \21198 , \21194 , \21197 );
and \U$20884 ( \21199 , \21192 , \21197 );
or \U$20885 ( \21200 , \21195 , \21198 , \21199 );
xor \U$20886 ( \21201 , \21129 , \21141 );
xor \U$20887 ( \21202 , \21201 , \21146 );
and \U$20888 ( \21203 , \21200 , \21202 );
xor \U$20889 ( \21204 , \21153 , \21155 );
and \U$20890 ( \21205 , \21202 , \21204 );
and \U$20891 ( \21206 , \21200 , \21204 );
or \U$20892 ( \21207 , \21203 , \21205 , \21206 );
and \U$20893 ( \21208 , \21176 , \21207 );
xor \U$20894 ( \21209 , \21176 , \21207 );
xor \U$20895 ( \21210 , \21200 , \21202 );
xor \U$20896 ( \21211 , \21210 , \21204 );
and \U$20897 ( \21212 , \9550 , \10814 );
and \U$20898 ( \21213 , \8981 , \10811 );
nor \U$20899 ( \21214 , \21212 , \21213 );
xnor \U$20900 ( \21215 , \21214 , \9759 );
and \U$20901 ( \21216 , \10161 , \10001 );
and \U$20902 ( \21217 , \9558 , \9999 );
nor \U$20903 ( \21218 , \21216 , \21217 );
xnor \U$20904 ( \21219 , \21218 , \9762 );
and \U$20905 ( \21220 , \21215 , \21219 );
and \U$20906 ( \21221 , \21219 , \8525 );
and \U$20907 ( \21222 , \21215 , \8525 );
or \U$20908 ( \21223 , \21220 , \21221 , \21222 );
and \U$20909 ( \21224 , \10347 , \9433 );
and \U$20910 ( \21225 , \10166 , \9431 );
nor \U$20911 ( \21226 , \21224 , \21225 );
xnor \U$20912 ( \21227 , \21226 , \9123 );
nand \U$20913 ( \21228 , \10967 , \8894 );
xnor \U$20914 ( \21229 , \21228 , \8525 );
and \U$20915 ( \21230 , \21227 , \21229 );
and \U$20916 ( \21231 , \21223 , \21230 );
and \U$20917 ( \21232 , \10967 , \8896 );
and \U$20918 ( \21233 , \10347 , \8894 );
nor \U$20919 ( \21234 , \21232 , \21233 );
xnor \U$20920 ( \21235 , \21234 , \8525 );
and \U$20921 ( \21236 , \21230 , \21235 );
and \U$20922 ( \21237 , \21223 , \21235 );
or \U$20923 ( \21238 , \21231 , \21236 , \21237 );
xor \U$20924 ( \21239 , \21192 , \21194 );
xor \U$20925 ( \21240 , \21239 , \21197 );
and \U$20926 ( \21241 , \21238 , \21240 );
and \U$20927 ( \21242 , \21211 , \21241 );
xor \U$20928 ( \21243 , \21211 , \21241 );
xor \U$20929 ( \21244 , \21238 , \21240 );
xor \U$20930 ( \21245 , \21180 , \21184 );
xor \U$20931 ( \21246 , \21245 , \21189 );
xor \U$20932 ( \21247 , \21223 , \21230 );
xor \U$20933 ( \21248 , \21247 , \21235 );
and \U$20934 ( \21249 , \21246 , \21248 );
and \U$20935 ( \21250 , \21244 , \21249 );
xor \U$20936 ( \21251 , \21244 , \21249 );
xor \U$20937 ( \21252 , \21246 , \21248 );
and \U$20938 ( \21253 , \9558 , \10814 );
and \U$20939 ( \21254 , \9550 , \10811 );
nor \U$20940 ( \21255 , \21253 , \21254 );
xnor \U$20941 ( \21256 , \21255 , \9759 );
and \U$20942 ( \21257 , \10166 , \10001 );
and \U$20943 ( \21258 , \10161 , \9999 );
nor \U$20944 ( \21259 , \21257 , \21258 );
xnor \U$20945 ( \21260 , \21259 , \9762 );
and \U$20946 ( \21261 , \21256 , \21260 );
and \U$20947 ( \21262 , \10967 , \9433 );
and \U$20948 ( \21263 , \10347 , \9431 );
nor \U$20949 ( \21264 , \21262 , \21263 );
xnor \U$20950 ( \21265 , \21264 , \9123 );
and \U$20951 ( \21266 , \21260 , \21265 );
and \U$20952 ( \21267 , \21256 , \21265 );
or \U$20953 ( \21268 , \21261 , \21266 , \21267 );
xor \U$20954 ( \21269 , \21215 , \21219 );
xor \U$20955 ( \21270 , \21269 , \8525 );
and \U$20956 ( \21271 , \21268 , \21270 );
xor \U$20957 ( \21272 , \21227 , \21229 );
and \U$20958 ( \21273 , \21270 , \21272 );
and \U$20959 ( \21274 , \21268 , \21272 );
or \U$20960 ( \21275 , \21271 , \21273 , \21274 );
and \U$20961 ( \21276 , \21252 , \21275 );
xor \U$20962 ( \21277 , \21252 , \21275 );
xor \U$20963 ( \21278 , \21268 , \21270 );
xor \U$20964 ( \21279 , \21278 , \21272 );
and \U$20965 ( \21280 , \10161 , \10814 );
and \U$20966 ( \21281 , \9558 , \10811 );
nor \U$20967 ( \21282 , \21280 , \21281 );
xnor \U$20968 ( \21283 , \21282 , \9759 );
and \U$20969 ( \21284 , \10347 , \10001 );
and \U$20970 ( \21285 , \10166 , \9999 );
nor \U$20971 ( \21286 , \21284 , \21285 );
xnor \U$20972 ( \21287 , \21286 , \9762 );
and \U$20973 ( \21288 , \21283 , \21287 );
and \U$20974 ( \21289 , \21287 , \9123 );
and \U$20975 ( \21290 , \21283 , \9123 );
or \U$20976 ( \21291 , \21288 , \21289 , \21290 );
xor \U$20977 ( \21292 , \21256 , \21260 );
xor \U$20978 ( \21293 , \21292 , \21265 );
and \U$20979 ( \21294 , \21291 , \21293 );
and \U$20980 ( \21295 , \21279 , \21294 );
xor \U$20981 ( \21296 , \21279 , \21294 );
xor \U$20982 ( \21297 , \21291 , \21293 );
nand \U$20983 ( \21298 , \10967 , \9431 );
xnor \U$20984 ( \21299 , \21298 , \9123 );
xor \U$20985 ( \21300 , \21283 , \21287 );
xor \U$20986 ( \21301 , \21300 , \9123 );
and \U$20987 ( \21302 , \21299 , \21301 );
and \U$20988 ( \21303 , \21297 , \21302 );
xor \U$20989 ( \21304 , \21297 , \21302 );
xor \U$20990 ( \21305 , \21299 , \21301 );
and \U$20991 ( \21306 , \10166 , \10814 );
and \U$20992 ( \21307 , \10161 , \10811 );
nor \U$20993 ( \21308 , \21306 , \21307 );
xnor \U$20994 ( \21309 , \21308 , \9759 );
and \U$20995 ( \21310 , \10967 , \10001 );
and \U$20996 ( \21311 , \10347 , \9999 );
nor \U$20997 ( \21312 , \21310 , \21311 );
xnor \U$20998 ( \21313 , \21312 , \9762 );
and \U$20999 ( \21314 , \21309 , \21313 );
and \U$21000 ( \21315 , \21305 , \21314 );
xor \U$21001 ( \21316 , \21305 , \21314 );
xor \U$21002 ( \21317 , \21309 , \21313 );
and \U$21003 ( \21318 , \10347 , \10814 );
and \U$21004 ( \21319 , \10166 , \10811 );
nor \U$21005 ( \21320 , \21318 , \21319 );
xnor \U$21006 ( \21321 , \21320 , \9759 );
and \U$21007 ( \21322 , \21321 , \9762 );
and \U$21008 ( \21323 , \21317 , \21322 );
xor \U$21009 ( \21324 , \21317 , \21322 );
nand \U$21010 ( \21325 , \10967 , \9999 );
xnor \U$21011 ( \21326 , \21325 , \9762 );
xor \U$21012 ( \21327 , \21321 , \9762 );
and \U$21013 ( \21328 , \21326 , \21327 );
xor \U$21014 ( \21329 , \21326 , \21327 );
and \U$21015 ( \21330 , \10967 , \10814 );
and \U$21016 ( \21331 , \10347 , \10811 );
nor \U$21017 ( \21332 , \21330 , \21331 );
xnor \U$21018 ( \21333 , \21332 , \9759 );
nand \U$21019 ( \21334 , \10967 , \10811 );
xnor \U$21020 ( \21335 , \21334 , \9759 );
and \U$21021 ( \21336 , \21335 , \9759 );
and \U$21022 ( \21337 , \21333 , \21336 );
and \U$21023 ( \21338 , \21329 , \21337 );
or \U$21024 ( \21339 , \21328 , \21338 );
and \U$21025 ( \21340 , \21324 , \21339 );
or \U$21026 ( \21341 , \21323 , \21340 );
and \U$21027 ( \21342 , \21316 , \21341 );
or \U$21028 ( \21343 , \21315 , \21342 );
and \U$21029 ( \21344 , \21304 , \21343 );
or \U$21030 ( \21345 , \21303 , \21344 );
and \U$21031 ( \21346 , \21296 , \21345 );
or \U$21032 ( \21347 , \21295 , \21346 );
and \U$21033 ( \21348 , \21277 , \21347 );
or \U$21034 ( \21349 , \21276 , \21348 );
and \U$21035 ( \21350 , \21251 , \21349 );
or \U$21036 ( \21351 , \21250 , \21350 );
and \U$21037 ( \21352 , \21243 , \21351 );
or \U$21038 ( \21353 , \21242 , \21352 );
and \U$21039 ( \21354 , \21209 , \21353 );
or \U$21040 ( \21355 , \21208 , \21354 );
and \U$21041 ( \21356 , \21175 , \21355 );
or \U$21042 ( \21357 , \21174 , \21356 );
and \U$21043 ( \21358 , \21167 , \21357 );
or \U$21044 ( \21359 , \21166 , \21358 );
and \U$21045 ( \21360 , \21114 , \21359 );
or \U$21046 ( \21361 , \21113 , \21360 );
and \U$21047 ( \21362 , \21075 , \21361 );
or \U$21048 ( \21363 , \21074 , \21362 );
and \U$21049 ( \21364 , \21022 , \21363 );
or \U$21050 ( \21365 , \21021 , \21364 );
and \U$21051 ( \21366 , \20951 , \21365 );
or \U$21052 ( \21367 , \20950 , \21366 );
and \U$21053 ( \21368 , \20896 , \21367 );
or \U$21054 ( \21369 , \20895 , \21368 );
and \U$21055 ( \21370 , \20837 , \21369 );
or \U$21056 ( \21371 , \20836 , \21370 );
and \U$21057 ( \21372 , \20829 , \21371 );
or \U$21058 ( \21373 , \20828 , \21372 );
and \U$21059 ( \21374 , \20750 , \21373 );
or \U$21060 ( \21375 , \20749 , \21374 );
and \U$21061 ( \21376 , \20670 , \21375 );
or \U$21062 ( \21377 , \20669 , \21376 );
and \U$21063 ( \21378 , \20575 , \21377 );
or \U$21064 ( \21379 , \20574 , \21378 );
and \U$21065 ( \21380 , \20487 , \21379 );
or \U$21066 ( \21381 , \20486 , \21380 );
and \U$21067 ( \21382 , \20395 , \21381 );
or \U$21068 ( \21383 , \20394 , \21382 );
and \U$21069 ( \21384 , \20307 , \21383 );
or \U$21070 ( \21385 , \20306 , \21384 );
and \U$21071 ( \21386 , \20192 , \21385 );
or \U$21072 ( \21387 , \20191 , \21386 );
and \U$21073 ( \21388 , \20096 , \21387 );
or \U$21074 ( \21389 , \20095 , \21388 );
and \U$21075 ( \21390 , \20088 , \21389 );
or \U$21076 ( \21391 , \20087 , \21390 );
and \U$21077 ( \21392 , \19973 , \21391 );
or \U$21078 ( \21393 , \19972 , \21392 );
and \U$21079 ( \21394 , \19849 , \21393 );
or \U$21080 ( \21395 , \19848 , \21394 );
and \U$21081 ( \21396 , \19709 , \21395 );
or \U$21082 ( \21397 , \19708 , \21396 );
and \U$21083 ( \21398 , \19585 , \21397 );
or \U$21084 ( \21399 , \19584 , \21398 );
and \U$21085 ( \21400 , \19441 , \21399 );
or \U$21086 ( \21401 , \19440 , \21400 );
and \U$21087 ( \21402 , \19316 , \21401 );
or \U$21088 ( \21403 , \19315 , \21402 );
and \U$21089 ( \21404 , \19177 , \21403 );
or \U$21090 ( \21405 , \19176 , \21404 );
and \U$21091 ( \21406 , \19013 , \21405 );
or \U$21092 ( \21407 , \19012 , \21406 );
and \U$21093 ( \21408 , \18861 , \21407 );
or \U$21094 ( \21409 , \18860 , \21408 );
and \U$21095 ( \21410 , \18721 , \21409 );
or \U$21096 ( \21411 , \18720 , \21410 );
and \U$21097 ( \21412 , \18553 , \21411 );
or \U$21098 ( \21413 , \18552 , \21412 );
and \U$21099 ( \21414 , \18545 , \21413 );
or \U$21100 ( \21415 , \18544 , \21414 );
and \U$21101 ( \21416 , \18374 , \21415 );
or \U$21102 ( \21417 , \18373 , \21416 );
and \U$21103 ( \21418 , \18198 , \21417 );
or \U$21104 ( \21419 , \18197 , \21418 );
and \U$21105 ( \21420 , \18008 , \21419 );
or \U$21106 ( \21421 , \18007 , \21420 );
and \U$21107 ( \21422 , \17821 , \21421 );
or \U$21108 ( \21423 , \17820 , \21422 );
and \U$21109 ( \21424 , \17636 , \21423 );
or \U$21110 ( \21425 , \17635 , \21424 );
and \U$21111 ( \21426 , \17428 , \21425 );
or \U$21112 ( \21427 , \17427 , \21426 );
and \U$21113 ( \21428 , \17232 , \21427 );
or \U$21114 ( \21429 , \17231 , \21428 );
and \U$21115 ( \21430 , \17035 , \21429 );
or \U$21116 ( \21431 , \17034 , \21430 );
and \U$21117 ( \21432 , \16822 , \21431 );
or \U$21118 ( \21433 , \16821 , \21432 );
and \U$21119 ( \21434 , \16611 , \21433 );
or \U$21120 ( \21435 , \16610 , \21434 );
and \U$21121 ( \21436 , \16380 , \21435 );
or \U$21122 ( \21437 , \16379 , \21436 );
and \U$21123 ( \21438 , \16150 , \21437 );
or \U$21124 ( \21439 , \16149 , \21438 );
and \U$21125 ( \21440 , \15931 , \21439 );
or \U$21126 ( \21441 , \15930 , \21440 );
and \U$21127 ( \21442 , \15706 , \21441 );
or \U$21128 ( \21443 , \15705 , \21442 );
and \U$21129 ( \21444 , \15456 , \21443 );
or \U$21130 ( \21445 , \15455 , \21444 );
and \U$21131 ( \21446 , \15226 , \21445 );
or \U$21132 ( \21447 , \15225 , \21446 );
and \U$21133 ( \21448 , \14980 , \21447 );
or \U$21134 ( \21449 , \14979 , \21448 );
and \U$21135 ( \21450 , \14972 , \21449 );
or \U$21136 ( \21451 , \14971 , \21450 );
and \U$21137 ( \21452 , \14711 , \21451 );
or \U$21138 ( \21453 , \14710 , \21452 );
and \U$21139 ( \21454 , \14449 , \21453 );
or \U$21140 ( \21455 , \14448 , \21454 );
and \U$21141 ( \21456 , \14179 , \21455 );
or \U$21142 ( \21457 , \14178 , \21456 );
and \U$21143 ( \21458 , \13902 , \21457 );
or \U$21144 ( \21459 , \13901 , \21458 );
and \U$21145 ( \21460 , \13626 , \21459 );
or \U$21146 ( \21461 , \13625 , \21460 );
and \U$21147 ( \21462 , \13355 , \21461 );
or \U$21148 ( \21463 , \13354 , \21462 );
and \U$21149 ( \21464 , \13052 , \21463 );
or \U$21150 ( \21465 , \13051 , \21464 );
and \U$21151 ( \21466 , \12773 , \21465 );
or \U$21152 ( \21467 , \12772 , \21466 );
and \U$21153 ( \21468 , \12488 , \21467 );
or \U$21154 ( \21469 , \12487 , \21468 );
and \U$21155 ( \21470 , \12172 , \21469 );
or \U$21156 ( \21471 , \12171 , \21470 );
and \U$21157 ( \21472 , \11872 , \21471 );
or \U$21158 ( \21473 , \11871 , \21472 );
and \U$21159 ( \21474 , \11556 , \21473 );
or \U$21160 ( \21475 , \11555 , \21474 );
and \U$21161 ( \21476 , \11238 , \21475 );
or \U$21162 ( \21477 , \11237 , \21476 );
and \U$21163 ( \21478 , \10927 , \21477 );
or \U$21164 ( \21479 , \10926 , \21478 );
and \U$21165 ( \21480 , \10614 , \21479 );
or \U$21166 ( \21481 , \10613 , \21480 );
and \U$21167 ( \21482 , \10298 , \21481 );
or \U$21168 ( \21483 , \10297 , \21482 );
and \U$21169 ( \21484 , \9980 , \21483 );
or \U$21170 ( \21485 , \9979 , \21484 );
and \U$21171 ( \21486 , \9671 , \21485 );
or \U$21172 ( \21487 , \9670 , \21486 );
and \U$21173 ( \21488 , \9375 , \21487 );
or \U$21174 ( \21489 , \9374 , \21488 );
and \U$21175 ( \21490 , \9074 , \21489 );
or \U$21176 ( \21491 , \9073 , \21490 );
and \U$21177 ( \21492 , \8786 , \21491 );
or \U$21178 ( \21493 , \8785 , \21492 );
and \U$21179 ( \21494 , \8503 , \21493 );
or \U$21180 ( \21495 , \8502 , \21494 );
and \U$21181 ( \21496 , \8208 , \21495 );
or \U$21182 ( \21497 , \8207 , \21496 );
and \U$21183 ( \21498 , \7942 , \21497 );
or \U$21184 ( \21499 , \7941 , \21498 );
and \U$21185 ( \21500 , \7676 , \21499 );
or \U$21186 ( \21501 , \7675 , \21500 );
and \U$21187 ( \21502 , \7415 , \21501 );
or \U$21188 ( \21503 , \7414 , \21502 );
and \U$21189 ( \21504 , \7150 , \21503 );
or \U$21190 ( \21505 , \7149 , \21504 );
and \U$21191 ( \21506 , \6887 , \21505 );
or \U$21192 ( \21507 , \6886 , \21506 );
and \U$21193 ( \21508 , \6630 , \21507 );
or \U$21194 ( \21509 , \6629 , \21508 );
and \U$21195 ( \21510 , \6374 , \21509 );
or \U$21196 ( \21511 , \6373 , \21510 );
and \U$21197 ( \21512 , \6121 , \21511 );
or \U$21198 ( \21513 , \6120 , \21512 );
and \U$21199 ( \21514 , \5873 , \21513 );
or \U$21200 ( \21515 , \5872 , \21514 );
and \U$21201 ( \21516 , \5641 , \21515 );
or \U$21202 ( \21517 , \5640 , \21516 );
and \U$21203 ( \21518 , \5398 , \21517 );
or \U$21204 ( \21519 , \5397 , \21518 );
and \U$21205 ( \21520 , \4969 , \21519 );
or \U$21206 ( \21521 , \4968 , \21520 );
and \U$21207 ( \21522 , \4759 , \21521 );
or \U$21208 ( \21523 , \4758 , \21522 );
and \U$21209 ( \21524 , \4552 , \21523 );
or \U$21210 ( \21525 , \4551 , \21524 );
and \U$21211 ( \21526 , \4350 , \21525 );
or \U$21212 ( \21527 , \4349 , \21526 );
and \U$21213 ( \21528 , \4154 , \21527 );
or \U$21214 ( \21529 , \4153 , \21528 );
and \U$21215 ( \21530 , \3957 , \21529 );
or \U$21216 ( \21531 , \3956 , \21530 );
and \U$21217 ( \21532 , \3780 , \21531 );
or \U$21218 ( \21533 , \3779 , \21532 );
and \U$21219 ( \21534 , \3599 , \21533 );
or \U$21220 ( \21535 , \3598 , \21534 );
and \U$21221 ( \21536 , \3428 , \21535 );
or \U$21222 ( \21537 , \3427 , \21536 );
and \U$21223 ( \21538 , \3253 , \21537 );
or \U$21224 ( \21539 , \3252 , \21538 );
and \U$21225 ( \21540 , \3080 , \21539 );
or \U$21226 ( \21541 , \3079 , \21540 );
and \U$21227 ( \21542 , \2913 , \21541 );
or \U$21228 ( \21543 , \2912 , \21542 );
and \U$21229 ( \21544 , \2747 , \21543 );
or \U$21230 ( \21545 , \2746 , \21544 );
and \U$21231 ( \21546 , \2574 , \21545 );
or \U$21232 ( \21547 , \2573 , \21546 );
and \U$21233 ( \21548 , \2294 , \21547 );
or \U$21234 ( \21549 , \2293 , \21548 );
and \U$21235 ( \21550 , \2157 , \21549 );
or \U$21236 ( \21551 , \2156 , \21550 );
and \U$21237 ( \21552 , \2024 , \21551 );
or \U$21238 ( \21553 , \2023 , \21552 );
and \U$21239 ( \21554 , \1903 , \21553 );
or \U$21240 ( \21555 , \1902 , \21554 );
and \U$21241 ( \21556 , \1780 , \21555 );
or \U$21242 ( \21557 , \1779 , \21556 );
and \U$21243 ( \21558 , \1664 , \21557 );
or \U$21244 ( \21559 , \1663 , \21558 );
and \U$21245 ( \21560 , \1549 , \21559 );
or \U$21246 ( \21561 , \1548 , \21560 );
and \U$21247 ( \21562 , \1435 , \21561 );
or \U$21248 ( \21563 , \1434 , \21562 );
and \U$21249 ( \21564 , \1321 , \21563 );
or \U$21250 ( \21565 , \1320 , \21564 );
and \U$21251 ( \21566 , \1139 , \21565 );
or \U$21252 ( \21567 , \1138 , \21566 );
and \U$21253 ( \21568 , \1060 , \21567 );
or \U$21254 ( \21569 , \1059 , \21568 );
and \U$21255 ( \21570 , \977 , \21569 );
or \U$21256 ( \21571 , \976 , \21570 );
and \U$21257 ( \21572 , \896 , \21571 );
or \U$21258 ( \21573 , \895 , \21572 );
and \U$21259 ( \21574 , \821 , \21573 );
or \U$21260 ( \21575 , \820 , \21574 );
and \U$21261 ( \21576 , \747 , \21575 );
or \U$21262 ( \21577 , \746 , \21576 );
and \U$21263 ( \21578 , \627 , \21577 );
or \U$21264 ( \21579 , \626 , \21578 );
and \U$21265 ( \21580 , \574 , \21579 );
or \U$21266 ( \21581 , \573 , \21580 );
and \U$21267 ( \21582 , \524 , \21581 );
or \U$21268 ( \21583 , \523 , \21582 );
and \U$21269 ( \21584 , \472 , \21583 );
or \U$21270 ( \21585 , \471 , \21584 );
and \U$21271 ( \21586 , \402 , \21585 );
or \U$21272 ( \21587 , \401 , \21586 );
xor \U$21273 ( \21588 , \355 , \21587 );
buf \U$21274 ( \21589 , \21588 );
buf \U$21275 ( \21590 , RIc0c9660_4);
buf \U$21276 ( \21591 , RIc0c95e8_5);
buf \U$21277 ( \21592 , RIc0c9570_6);
and \U$21278 ( \21593 , \21591 , \21592 );
not \U$21279 ( \21594 , \21593 );
and \U$21280 ( \21595 , \21590 , \21594 );
not \U$21281 ( \21596 , \21595 );
buf \U$21282 ( \21597 , RIc0c7950_66);
buf \U$21283 ( \21598 , RIc340698_130);
xor \U$21284 ( \21599 , \21597 , \21598 );
buf \U$21285 ( \21600 , RIc0c78d8_67);
buf \U$21286 ( \21601 , RIc340710_131);
and \U$21287 ( \21602 , \21600 , \21601 );
buf \U$21288 ( \21603 , RIc0c7860_68);
buf \U$21289 ( \21604 , RIc340788_132);
and \U$21290 ( \21605 , \21603 , \21604 );
buf \U$21291 ( \21606 , RIc0c77e8_69);
buf \U$21292 ( \21607 , RIc340800_133);
and \U$21293 ( \21608 , \21606 , \21607 );
buf \U$21294 ( \21609 , RIc0c7770_70);
buf \U$21295 ( \21610 , RIc340878_134);
and \U$21296 ( \21611 , \21609 , \21610 );
buf \U$21297 ( \21612 , RIc0c76f8_71);
buf \U$21298 ( \21613 , RIc3408f0_135);
and \U$21299 ( \21614 , \21612 , \21613 );
buf \U$21300 ( \21615 , RIc0c7680_72);
buf \U$21301 ( \21616 , RIc340968_136);
and \U$21302 ( \21617 , \21615 , \21616 );
buf \U$21303 ( \21618 , RIc0c7608_73);
buf \U$21304 ( \21619 , RIc3409e0_137);
and \U$21305 ( \21620 , \21618 , \21619 );
buf \U$21306 ( \21621 , RIc0c7590_74);
buf \U$21307 ( \21622 , RIc340a58_138);
and \U$21308 ( \21623 , \21621 , \21622 );
buf \U$21309 ( \21624 , RIc0c7518_75);
buf \U$21310 ( \21625 , RIc340ad0_139);
and \U$21311 ( \21626 , \21624 , \21625 );
buf \U$21312 ( \21627 , RIc0c74a0_76);
buf \U$21313 ( \21628 , RIc340b48_140);
and \U$21314 ( \21629 , \21627 , \21628 );
buf \U$21315 ( \21630 , RIc0c7428_77);
buf \U$21316 ( \21631 , RIc340bc0_141);
and \U$21317 ( \21632 , \21630 , \21631 );
buf \U$21318 ( \21633 , RIc0c73b0_78);
buf \U$21319 ( \21634 , RIc340c38_142);
and \U$21320 ( \21635 , \21633 , \21634 );
buf \U$21321 ( \21636 , RIc0c7338_79);
buf \U$21322 ( \21637 , RIc340cb0_143);
and \U$21323 ( \21638 , \21636 , \21637 );
buf \U$21324 ( \21639 , RIc0c72c0_80);
buf \U$21325 ( \21640 , RIc340d28_144);
and \U$21326 ( \21641 , \21639 , \21640 );
buf \U$21327 ( \21642 , RIc0c7248_81);
buf \U$21328 ( \21643 , RIc340da0_145);
and \U$21329 ( \21644 , \21642 , \21643 );
buf \U$21330 ( \21645 , RIc0c71d0_82);
buf \U$21331 ( \21646 , RIc340e18_146);
and \U$21332 ( \21647 , \21645 , \21646 );
buf \U$21333 ( \21648 , RIc0c7158_83);
buf \U$21334 ( \21649 , RIc340e90_147);
and \U$21335 ( \21650 , \21648 , \21649 );
buf \U$21336 ( \21651 , RIc0c70e0_84);
buf \U$21337 ( \21652 , RIc340f08_148);
and \U$21338 ( \21653 , \21651 , \21652 );
buf \U$21339 ( \21654 , RIc0c7068_85);
buf \U$21340 ( \21655 , RIc340f80_149);
and \U$21341 ( \21656 , \21654 , \21655 );
buf \U$21342 ( \21657 , RIc0c6ff0_86);
buf \U$21343 ( \21658 , RIc340ff8_150);
and \U$21344 ( \21659 , \21657 , \21658 );
buf \U$21345 ( \21660 , RIc0c6f78_87);
buf \U$21346 ( \21661 , RIc341070_151);
and \U$21347 ( \21662 , \21660 , \21661 );
buf \U$21348 ( \21663 , RIc0c6f00_88);
buf \U$21349 ( \21664 , RIc3410e8_152);
and \U$21350 ( \21665 , \21663 , \21664 );
buf \U$21351 ( \21666 , RIc0c6e88_89);
buf \U$21352 ( \21667 , RIc341160_153);
and \U$21353 ( \21668 , \21666 , \21667 );
buf \U$21354 ( \21669 , RIc0c6e10_90);
buf \U$21355 ( \21670 , RIc3411d8_154);
and \U$21356 ( \21671 , \21669 , \21670 );
buf \U$21357 ( \21672 , RIc0c6d98_91);
buf \U$21358 ( \21673 , RIc341250_155);
and \U$21359 ( \21674 , \21672 , \21673 );
buf \U$21360 ( \21675 , RIc0c6d20_92);
buf \U$21361 ( \21676 , RIc3412c8_156);
and \U$21362 ( \21677 , \21675 , \21676 );
buf \U$21363 ( \21678 , RIc0c6ca8_93);
buf \U$21364 ( \21679 , RIc341340_157);
and \U$21365 ( \21680 , \21678 , \21679 );
buf \U$21366 ( \21681 , RIc0c6c30_94);
buf \U$21367 ( \21682 , RIc3413b8_158);
and \U$21368 ( \21683 , \21681 , \21682 );
buf \U$21369 ( \21684 , RIc0c6bb8_95);
buf \U$21370 ( \21685 , RIc341430_159);
and \U$21371 ( \21686 , \21684 , \21685 );
buf \U$21372 ( \21687 , RIc0c6b40_96);
buf \U$21373 ( \21688 , RIc3414a8_160);
and \U$21374 ( \21689 , \21687 , \21688 );
buf \U$21375 ( \21690 , RIc0c6ac8_97);
buf \U$21376 ( \21691 , RIc341520_161);
and \U$21377 ( \21692 , \21690 , \21691 );
buf \U$21378 ( \21693 , RIc0c6a50_98);
buf \U$21379 ( \21694 , RIc341598_162);
and \U$21380 ( \21695 , \21693 , \21694 );
buf \U$21381 ( \21696 , RIc0c69d8_99);
buf \U$21382 ( \21697 , RIc341610_163);
and \U$21383 ( \21698 , \21696 , \21697 );
buf \U$21384 ( \21699 , RIc0c6960_100);
buf \U$21385 ( \21700 , RIc341688_164);
and \U$21386 ( \21701 , \21699 , \21700 );
buf \U$21387 ( \21702 , RIc0c68e8_101);
buf \U$21388 ( \21703 , RIc341700_165);
and \U$21389 ( \21704 , \21702 , \21703 );
buf \U$21390 ( \21705 , RIc0c6870_102);
buf \U$21391 ( \21706 , RIc341778_166);
and \U$21392 ( \21707 , \21705 , \21706 );
buf \U$21393 ( \21708 , RIc0c67f8_103);
buf \U$21394 ( \21709 , RIc3417f0_167);
and \U$21395 ( \21710 , \21708 , \21709 );
buf \U$21396 ( \21711 , RIc0c6780_104);
buf \U$21397 ( \21712 , RIc341868_168);
and \U$21398 ( \21713 , \21711 , \21712 );
buf \U$21399 ( \21714 , RIc0c6708_105);
buf \U$21400 ( \21715 , RIc3418e0_169);
and \U$21401 ( \21716 , \21714 , \21715 );
buf \U$21402 ( \21717 , RIc0c6690_106);
buf \U$21403 ( \21718 , RIc341958_170);
and \U$21404 ( \21719 , \21717 , \21718 );
buf \U$21405 ( \21720 , RIc0c6618_107);
buf \U$21406 ( \21721 , RIc3419d0_171);
and \U$21407 ( \21722 , \21720 , \21721 );
buf \U$21408 ( \21723 , RIc0c65a0_108);
buf \U$21409 ( \21724 , RIc341a48_172);
and \U$21410 ( \21725 , \21723 , \21724 );
buf \U$21411 ( \21726 , RIc0c6528_109);
buf \U$21412 ( \21727 , RIc341ac0_173);
and \U$21413 ( \21728 , \21726 , \21727 );
buf \U$21414 ( \21729 , RIc0c64b0_110);
buf \U$21415 ( \21730 , RIc341b38_174);
and \U$21416 ( \21731 , \21729 , \21730 );
buf \U$21417 ( \21732 , RIc0c6438_111);
buf \U$21418 ( \21733 , RIc341bb0_175);
and \U$21419 ( \21734 , \21732 , \21733 );
buf \U$21420 ( \21735 , RIc0c63c0_112);
buf \U$21421 ( \21736 , RIc341c28_176);
and \U$21422 ( \21737 , \21735 , \21736 );
buf \U$21423 ( \21738 , RIc0c6348_113);
buf \U$21424 ( \21739 , RIc341ca0_177);
and \U$21425 ( \21740 , \21738 , \21739 );
buf \U$21426 ( \21741 , RIc0c62d0_114);
buf \U$21427 ( \21742 , RIc341d18_178);
and \U$21428 ( \21743 , \21741 , \21742 );
buf \U$21429 ( \21744 , RIc0c6258_115);
buf \U$21430 ( \21745 , RIc341d90_179);
and \U$21431 ( \21746 , \21744 , \21745 );
buf \U$21432 ( \21747 , RIc0c61e0_116);
buf \U$21433 ( \21748 , RIc341e08_180);
and \U$21434 ( \21749 , \21747 , \21748 );
buf \U$21435 ( \21750 , RIc0c6168_117);
buf \U$21436 ( \21751 , RIc341e80_181);
and \U$21437 ( \21752 , \21750 , \21751 );
buf \U$21438 ( \21753 , RIc0c60f0_118);
buf \U$21439 ( \21754 , RIc341ef8_182);
and \U$21440 ( \21755 , \21753 , \21754 );
buf \U$21441 ( \21756 , RIc0c6078_119);
buf \U$21442 ( \21757 , RIc341f70_183);
and \U$21443 ( \21758 , \21756 , \21757 );
buf \U$21444 ( \21759 , RIc0c6000_120);
buf \U$21445 ( \21760 , RIc341fe8_184);
and \U$21446 ( \21761 , \21759 , \21760 );
buf \U$21447 ( \21762 , RIc0c5f88_121);
buf \U$21448 ( \21763 , RIc342060_185);
and \U$21449 ( \21764 , \21762 , \21763 );
buf \U$21450 ( \21765 , RIc0c5f10_122);
buf \U$21451 ( \21766 , RIc3420d8_186);
and \U$21452 ( \21767 , \21765 , \21766 );
buf \U$21453 ( \21768 , RIc0c5e98_123);
buf \U$21454 ( \21769 , RIc342150_187);
and \U$21455 ( \21770 , \21768 , \21769 );
buf \U$21456 ( \21771 , RIc0c5e20_124);
buf \U$21457 ( \21772 , RIc3421c8_188);
and \U$21458 ( \21773 , \21771 , \21772 );
buf \U$21459 ( \21774 , RIc0c5da8_125);
buf \U$21460 ( \21775 , RIc342240_189);
and \U$21461 ( \21776 , \21774 , \21775 );
buf \U$21462 ( \21777 , RIc0c5d30_126);
buf \U$21463 ( \21778 , RIc3422b8_190);
and \U$21464 ( \21779 , \21777 , \21778 );
buf \U$21465 ( \21780 , RIc340530_127);
buf \U$21466 ( \21781 , RIc342330_191);
and \U$21467 ( \21782 , \21780 , \21781 );
buf \U$21468 ( \21783 , RIc3405a8_128);
buf \U$21469 ( \21784 , RIc3423a8_192);
and \U$21470 ( \21785 , \21783 , \21784 );
buf \U$21471 ( \21786 , RIc340620_129);
buf \U$21472 ( \21787 , RIc342420_193);
and \U$21473 ( \21788 , \21786 , \21787 );
and \U$21474 ( \21789 , \21784 , \21788 );
and \U$21475 ( \21790 , \21783 , \21788 );
or \U$21476 ( \21791 , \21785 , \21789 , \21790 );
and \U$21477 ( \21792 , \21781 , \21791 );
and \U$21478 ( \21793 , \21780 , \21791 );
or \U$21479 ( \21794 , \21782 , \21792 , \21793 );
and \U$21480 ( \21795 , \21778 , \21794 );
and \U$21481 ( \21796 , \21777 , \21794 );
or \U$21482 ( \21797 , \21779 , \21795 , \21796 );
and \U$21483 ( \21798 , \21775 , \21797 );
and \U$21484 ( \21799 , \21774 , \21797 );
or \U$21485 ( \21800 , \21776 , \21798 , \21799 );
and \U$21486 ( \21801 , \21772 , \21800 );
and \U$21487 ( \21802 , \21771 , \21800 );
or \U$21488 ( \21803 , \21773 , \21801 , \21802 );
and \U$21489 ( \21804 , \21769 , \21803 );
and \U$21490 ( \21805 , \21768 , \21803 );
or \U$21491 ( \21806 , \21770 , \21804 , \21805 );
and \U$21492 ( \21807 , \21766 , \21806 );
and \U$21493 ( \21808 , \21765 , \21806 );
or \U$21494 ( \21809 , \21767 , \21807 , \21808 );
and \U$21495 ( \21810 , \21763 , \21809 );
and \U$21496 ( \21811 , \21762 , \21809 );
or \U$21497 ( \21812 , \21764 , \21810 , \21811 );
and \U$21498 ( \21813 , \21760 , \21812 );
and \U$21499 ( \21814 , \21759 , \21812 );
or \U$21500 ( \21815 , \21761 , \21813 , \21814 );
and \U$21501 ( \21816 , \21757 , \21815 );
and \U$21502 ( \21817 , \21756 , \21815 );
or \U$21503 ( \21818 , \21758 , \21816 , \21817 );
and \U$21504 ( \21819 , \21754 , \21818 );
and \U$21505 ( \21820 , \21753 , \21818 );
or \U$21506 ( \21821 , \21755 , \21819 , \21820 );
and \U$21507 ( \21822 , \21751 , \21821 );
and \U$21508 ( \21823 , \21750 , \21821 );
or \U$21509 ( \21824 , \21752 , \21822 , \21823 );
and \U$21510 ( \21825 , \21748 , \21824 );
and \U$21511 ( \21826 , \21747 , \21824 );
or \U$21512 ( \21827 , \21749 , \21825 , \21826 );
and \U$21513 ( \21828 , \21745 , \21827 );
and \U$21514 ( \21829 , \21744 , \21827 );
or \U$21515 ( \21830 , \21746 , \21828 , \21829 );
and \U$21516 ( \21831 , \21742 , \21830 );
and \U$21517 ( \21832 , \21741 , \21830 );
or \U$21518 ( \21833 , \21743 , \21831 , \21832 );
and \U$21519 ( \21834 , \21739 , \21833 );
and \U$21520 ( \21835 , \21738 , \21833 );
or \U$21521 ( \21836 , \21740 , \21834 , \21835 );
and \U$21522 ( \21837 , \21736 , \21836 );
and \U$21523 ( \21838 , \21735 , \21836 );
or \U$21524 ( \21839 , \21737 , \21837 , \21838 );
and \U$21525 ( \21840 , \21733 , \21839 );
and \U$21526 ( \21841 , \21732 , \21839 );
or \U$21527 ( \21842 , \21734 , \21840 , \21841 );
and \U$21528 ( \21843 , \21730 , \21842 );
and \U$21529 ( \21844 , \21729 , \21842 );
or \U$21530 ( \21845 , \21731 , \21843 , \21844 );
and \U$21531 ( \21846 , \21727 , \21845 );
and \U$21532 ( \21847 , \21726 , \21845 );
or \U$21533 ( \21848 , \21728 , \21846 , \21847 );
and \U$21534 ( \21849 , \21724 , \21848 );
and \U$21535 ( \21850 , \21723 , \21848 );
or \U$21536 ( \21851 , \21725 , \21849 , \21850 );
and \U$21537 ( \21852 , \21721 , \21851 );
and \U$21538 ( \21853 , \21720 , \21851 );
or \U$21539 ( \21854 , \21722 , \21852 , \21853 );
and \U$21540 ( \21855 , \21718 , \21854 );
and \U$21541 ( \21856 , \21717 , \21854 );
or \U$21542 ( \21857 , \21719 , \21855 , \21856 );
and \U$21543 ( \21858 , \21715 , \21857 );
and \U$21544 ( \21859 , \21714 , \21857 );
or \U$21545 ( \21860 , \21716 , \21858 , \21859 );
and \U$21546 ( \21861 , \21712 , \21860 );
and \U$21547 ( \21862 , \21711 , \21860 );
or \U$21548 ( \21863 , \21713 , \21861 , \21862 );
and \U$21549 ( \21864 , \21709 , \21863 );
and \U$21550 ( \21865 , \21708 , \21863 );
or \U$21551 ( \21866 , \21710 , \21864 , \21865 );
and \U$21552 ( \21867 , \21706 , \21866 );
and \U$21553 ( \21868 , \21705 , \21866 );
or \U$21554 ( \21869 , \21707 , \21867 , \21868 );
and \U$21555 ( \21870 , \21703 , \21869 );
and \U$21556 ( \21871 , \21702 , \21869 );
or \U$21557 ( \21872 , \21704 , \21870 , \21871 );
and \U$21558 ( \21873 , \21700 , \21872 );
and \U$21559 ( \21874 , \21699 , \21872 );
or \U$21560 ( \21875 , \21701 , \21873 , \21874 );
and \U$21561 ( \21876 , \21697 , \21875 );
and \U$21562 ( \21877 , \21696 , \21875 );
or \U$21563 ( \21878 , \21698 , \21876 , \21877 );
and \U$21564 ( \21879 , \21694 , \21878 );
and \U$21565 ( \21880 , \21693 , \21878 );
or \U$21566 ( \21881 , \21695 , \21879 , \21880 );
and \U$21567 ( \21882 , \21691 , \21881 );
and \U$21568 ( \21883 , \21690 , \21881 );
or \U$21569 ( \21884 , \21692 , \21882 , \21883 );
and \U$21570 ( \21885 , \21688 , \21884 );
and \U$21571 ( \21886 , \21687 , \21884 );
or \U$21572 ( \21887 , \21689 , \21885 , \21886 );
and \U$21573 ( \21888 , \21685 , \21887 );
and \U$21574 ( \21889 , \21684 , \21887 );
or \U$21575 ( \21890 , \21686 , \21888 , \21889 );
and \U$21576 ( \21891 , \21682 , \21890 );
and \U$21577 ( \21892 , \21681 , \21890 );
or \U$21578 ( \21893 , \21683 , \21891 , \21892 );
and \U$21579 ( \21894 , \21679 , \21893 );
and \U$21580 ( \21895 , \21678 , \21893 );
or \U$21581 ( \21896 , \21680 , \21894 , \21895 );
and \U$21582 ( \21897 , \21676 , \21896 );
and \U$21583 ( \21898 , \21675 , \21896 );
or \U$21584 ( \21899 , \21677 , \21897 , \21898 );
and \U$21585 ( \21900 , \21673 , \21899 );
and \U$21586 ( \21901 , \21672 , \21899 );
or \U$21587 ( \21902 , \21674 , \21900 , \21901 );
and \U$21588 ( \21903 , \21670 , \21902 );
and \U$21589 ( \21904 , \21669 , \21902 );
or \U$21590 ( \21905 , \21671 , \21903 , \21904 );
and \U$21591 ( \21906 , \21667 , \21905 );
and \U$21592 ( \21907 , \21666 , \21905 );
or \U$21593 ( \21908 , \21668 , \21906 , \21907 );
and \U$21594 ( \21909 , \21664 , \21908 );
and \U$21595 ( \21910 , \21663 , \21908 );
or \U$21596 ( \21911 , \21665 , \21909 , \21910 );
and \U$21597 ( \21912 , \21661 , \21911 );
and \U$21598 ( \21913 , \21660 , \21911 );
or \U$21599 ( \21914 , \21662 , \21912 , \21913 );
and \U$21600 ( \21915 , \21658 , \21914 );
and \U$21601 ( \21916 , \21657 , \21914 );
or \U$21602 ( \21917 , \21659 , \21915 , \21916 );
and \U$21603 ( \21918 , \21655 , \21917 );
and \U$21604 ( \21919 , \21654 , \21917 );
or \U$21605 ( \21920 , \21656 , \21918 , \21919 );
and \U$21606 ( \21921 , \21652 , \21920 );
and \U$21607 ( \21922 , \21651 , \21920 );
or \U$21608 ( \21923 , \21653 , \21921 , \21922 );
and \U$21609 ( \21924 , \21649 , \21923 );
and \U$21610 ( \21925 , \21648 , \21923 );
or \U$21611 ( \21926 , \21650 , \21924 , \21925 );
and \U$21612 ( \21927 , \21646 , \21926 );
and \U$21613 ( \21928 , \21645 , \21926 );
or \U$21614 ( \21929 , \21647 , \21927 , \21928 );
and \U$21615 ( \21930 , \21643 , \21929 );
and \U$21616 ( \21931 , \21642 , \21929 );
or \U$21617 ( \21932 , \21644 , \21930 , \21931 );
and \U$21618 ( \21933 , \21640 , \21932 );
and \U$21619 ( \21934 , \21639 , \21932 );
or \U$21620 ( \21935 , \21641 , \21933 , \21934 );
and \U$21621 ( \21936 , \21637 , \21935 );
and \U$21622 ( \21937 , \21636 , \21935 );
or \U$21623 ( \21938 , \21638 , \21936 , \21937 );
and \U$21624 ( \21939 , \21634 , \21938 );
and \U$21625 ( \21940 , \21633 , \21938 );
or \U$21626 ( \21941 , \21635 , \21939 , \21940 );
and \U$21627 ( \21942 , \21631 , \21941 );
and \U$21628 ( \21943 , \21630 , \21941 );
or \U$21629 ( \21944 , \21632 , \21942 , \21943 );
and \U$21630 ( \21945 , \21628 , \21944 );
and \U$21631 ( \21946 , \21627 , \21944 );
or \U$21632 ( \21947 , \21629 , \21945 , \21946 );
and \U$21633 ( \21948 , \21625 , \21947 );
and \U$21634 ( \21949 , \21624 , \21947 );
or \U$21635 ( \21950 , \21626 , \21948 , \21949 );
and \U$21636 ( \21951 , \21622 , \21950 );
and \U$21637 ( \21952 , \21621 , \21950 );
or \U$21638 ( \21953 , \21623 , \21951 , \21952 );
and \U$21639 ( \21954 , \21619 , \21953 );
and \U$21640 ( \21955 , \21618 , \21953 );
or \U$21641 ( \21956 , \21620 , \21954 , \21955 );
and \U$21642 ( \21957 , \21616 , \21956 );
and \U$21643 ( \21958 , \21615 , \21956 );
or \U$21644 ( \21959 , \21617 , \21957 , \21958 );
and \U$21645 ( \21960 , \21613 , \21959 );
and \U$21646 ( \21961 , \21612 , \21959 );
or \U$21647 ( \21962 , \21614 , \21960 , \21961 );
and \U$21648 ( \21963 , \21610 , \21962 );
and \U$21649 ( \21964 , \21609 , \21962 );
or \U$21650 ( \21965 , \21611 , \21963 , \21964 );
and \U$21651 ( \21966 , \21607 , \21965 );
and \U$21652 ( \21967 , \21606 , \21965 );
or \U$21653 ( \21968 , \21608 , \21966 , \21967 );
and \U$21654 ( \21969 , \21604 , \21968 );
and \U$21655 ( \21970 , \21603 , \21968 );
or \U$21656 ( \21971 , \21605 , \21969 , \21970 );
and \U$21657 ( \21972 , \21601 , \21971 );
and \U$21658 ( \21973 , \21600 , \21971 );
or \U$21659 ( \21974 , \21602 , \21972 , \21973 );
xor \U$21660 ( \21975 , \21599 , \21974 );
buf \U$21661 ( \21976 , \21975 );
buf \U$21662 ( \21977 , \21976 );
buf \U$21663 ( \21978 , RIc0c9750_2);
buf \U$21664 ( \21979 , RIc0c96d8_3);
xor \U$21665 ( \21980 , \21978 , \21979 );
xor \U$21666 ( \21981 , \21979 , \21590 );
not \U$21667 ( \21982 , \21981 );
and \U$21668 ( \21983 , \21980 , \21982 );
and \U$21669 ( \21984 , \21977 , \21983 );
and \U$21670 ( \21985 , \21597 , \21598 );
and \U$21671 ( \21986 , \21598 , \21974 );
and \U$21672 ( \21987 , \21597 , \21974 );
or \U$21673 ( \21988 , \21985 , \21986 , \21987 );
buf \U$21674 ( \21989 , \21988 );
buf \U$21675 ( \21990 , \21989 );
and \U$21676 ( \21991 , \21990 , \21981 );
nor \U$21677 ( \21992 , \21984 , \21991 );
and \U$21678 ( \21993 , \21979 , \21590 );
not \U$21679 ( \21994 , \21993 );
and \U$21680 ( \21995 , \21978 , \21994 );
xnor \U$21681 ( \21996 , \21992 , \21995 );
and \U$21682 ( \21997 , \21596 , \21996 );
xor \U$21683 ( \21998 , \21600 , \21601 );
xor \U$21684 ( \21999 , \21998 , \21971 );
buf \U$21685 ( \22000 , \21999 );
buf \U$21686 ( \22001 , \22000 );
and \U$21687 ( \22002 , \22001 , \21978 );
and \U$21688 ( \22003 , \21996 , \22002 );
and \U$21689 ( \22004 , \21596 , \22002 );
or \U$21690 ( \22005 , \21997 , \22003 , \22004 );
and \U$21691 ( \22006 , \21990 , \21983 );
not \U$21692 ( \22007 , \22006 );
xnor \U$21693 ( \22008 , \22007 , \21995 );
and \U$21694 ( \22009 , \21977 , \21978 );
xnor \U$21695 ( \22010 , \22008 , \22009 );
xor \U$21696 ( \22011 , \22005 , \22010 );
buf \U$21697 ( \22012 , RIc0c94f8_7);
buf \U$21698 ( \22013 , RIc0c9480_8);
and \U$21699 ( \22014 , \22012 , \22013 );
not \U$21700 ( \22015 , \22014 );
and \U$21701 ( \22016 , \21592 , \22015 );
not \U$21702 ( \22017 , \22016 );
xor \U$21703 ( \22018 , \21590 , \21591 );
xor \U$21704 ( \22019 , \21591 , \21592 );
not \U$21705 ( \22020 , \22019 );
and \U$21706 ( \22021 , \22018 , \22020 );
and \U$21707 ( \22022 , \21977 , \22021 );
and \U$21708 ( \22023 , \21990 , \22019 );
nor \U$21709 ( \22024 , \22022 , \22023 );
xnor \U$21710 ( \22025 , \22024 , \21595 );
and \U$21711 ( \22026 , \22017 , \22025 );
xor \U$21712 ( \22027 , \21603 , \21604 );
xor \U$21713 ( \22028 , \22027 , \21968 );
buf \U$21714 ( \22029 , \22028 );
buf \U$21715 ( \22030 , \22029 );
and \U$21716 ( \22031 , \22030 , \21983 );
and \U$21717 ( \22032 , \22001 , \21981 );
nor \U$21718 ( \22033 , \22031 , \22032 );
xnor \U$21719 ( \22034 , \22033 , \21995 );
and \U$21720 ( \22035 , \22025 , \22034 );
and \U$21721 ( \22036 , \22017 , \22034 );
or \U$21722 ( \22037 , \22026 , \22035 , \22036 );
and \U$21723 ( \22038 , \21990 , \22021 );
not \U$21724 ( \22039 , \22038 );
xnor \U$21725 ( \22040 , \22039 , \21595 );
and \U$21726 ( \22041 , \22001 , \21983 );
and \U$21727 ( \22042 , \21977 , \21981 );
nor \U$21728 ( \22043 , \22041 , \22042 );
xnor \U$21729 ( \22044 , \22043 , \21995 );
xor \U$21730 ( \22045 , \22040 , \22044 );
and \U$21731 ( \22046 , \22030 , \21978 );
xor \U$21732 ( \22047 , \22045 , \22046 );
or \U$21733 ( \22048 , \22037 , \22047 );
and \U$21734 ( \22049 , \22040 , \22044 );
and \U$21735 ( \22050 , \22044 , \22046 );
and \U$21736 ( \22051 , \22040 , \22046 );
or \U$21737 ( \22052 , \22049 , \22050 , \22051 );
and \U$21738 ( \22053 , \22048 , \22052 );
xor \U$21739 ( \22054 , \21596 , \21996 );
xor \U$21740 ( \22055 , \22054 , \22002 );
and \U$21741 ( \22056 , \22052 , \22055 );
and \U$21742 ( \22057 , \22048 , \22055 );
or \U$21743 ( \22058 , \22053 , \22056 , \22057 );
nand \U$21744 ( \22059 , \22011 , \22058 );
nor \U$21745 ( \22060 , \22011 , \22058 );
not \U$21746 ( \22061 , \22060 );
nand \U$21747 ( \22062 , \22059 , \22061 );
buf \U$21748 ( \22063 , RIc0c9408_9);
buf \U$21749 ( \22064 , RIc0c9390_10);
and \U$21750 ( \22065 , \22063 , \22064 );
not \U$21751 ( \22066 , \22065 );
and \U$21752 ( \22067 , \22013 , \22066 );
xor \U$21753 ( \22068 , \21621 , \21622 );
xor \U$21754 ( \22069 , \22068 , \21950 );
buf \U$21755 ( \22070 , \22069 );
buf \U$21756 ( \22071 , \22070 );
buf \U$21757 ( \22072 , RIc0c7a40_64);
buf \U$21758 ( \22073 , RIc0c79c8_65);
xor \U$21759 ( \22074 , \22072 , \22073 );
not \U$21760 ( \22075 , \22073 );
and \U$21761 ( \22076 , \22074 , \22075 );
and \U$21762 ( \22077 , \22071 , \22076 );
xor \U$21763 ( \22078 , \21618 , \21619 );
xor \U$21764 ( \22079 , \22078 , \21953 );
buf \U$21765 ( \22080 , \22079 );
buf \U$21766 ( \22081 , \22080 );
and \U$21767 ( \22082 , \22081 , \22073 );
nor \U$21768 ( \22083 , \22077 , \22082 );
xnor \U$21769 ( \22084 , \22083 , \22072 );
and \U$21770 ( \22085 , \22067 , \22084 );
xor \U$21771 ( \22086 , \21627 , \21628 );
xor \U$21772 ( \22087 , \22086 , \21944 );
buf \U$21773 ( \22088 , \22087 );
buf \U$21774 ( \22089 , \22088 );
buf \U$21775 ( \22090 , RIc0c7b30_62);
buf \U$21776 ( \22091 , RIc0c7ab8_63);
xor \U$21777 ( \22092 , \22090 , \22091 );
xor \U$21778 ( \22093 , \22091 , \22072 );
not \U$21779 ( \22094 , \22093 );
and \U$21780 ( \22095 , \22092 , \22094 );
and \U$21781 ( \22096 , \22089 , \22095 );
xor \U$21782 ( \22097 , \21624 , \21625 );
xor \U$21783 ( \22098 , \22097 , \21947 );
buf \U$21784 ( \22099 , \22098 );
buf \U$21785 ( \22100 , \22099 );
and \U$21786 ( \22101 , \22100 , \22093 );
nor \U$21787 ( \22102 , \22096 , \22101 );
and \U$21788 ( \22103 , \22091 , \22072 );
not \U$21789 ( \22104 , \22103 );
and \U$21790 ( \22105 , \22090 , \22104 );
xnor \U$21791 ( \22106 , \22102 , \22105 );
and \U$21792 ( \22107 , \22084 , \22106 );
and \U$21793 ( \22108 , \22067 , \22106 );
or \U$21794 ( \22109 , \22085 , \22107 , \22108 );
xor \U$21795 ( \22110 , \21633 , \21634 );
xor \U$21796 ( \22111 , \22110 , \21938 );
buf \U$21797 ( \22112 , \22111 );
buf \U$21798 ( \22113 , \22112 );
buf \U$21799 ( \22114 , RIc0c7c20_60);
buf \U$21800 ( \22115 , RIc0c7ba8_61);
xor \U$21801 ( \22116 , \22114 , \22115 );
xor \U$21802 ( \22117 , \22115 , \22090 );
not \U$21803 ( \22118 , \22117 );
and \U$21804 ( \22119 , \22116 , \22118 );
and \U$21805 ( \22120 , \22113 , \22119 );
xor \U$21806 ( \22121 , \21630 , \21631 );
xor \U$21807 ( \22122 , \22121 , \21941 );
buf \U$21808 ( \22123 , \22122 );
buf \U$21809 ( \22124 , \22123 );
and \U$21810 ( \22125 , \22124 , \22117 );
nor \U$21811 ( \22126 , \22120 , \22125 );
and \U$21812 ( \22127 , \22115 , \22090 );
not \U$21813 ( \22128 , \22127 );
and \U$21814 ( \22129 , \22114 , \22128 );
xnor \U$21815 ( \22130 , \22126 , \22129 );
xor \U$21816 ( \22131 , \21639 , \21640 );
xor \U$21817 ( \22132 , \22131 , \21932 );
buf \U$21818 ( \22133 , \22132 );
buf \U$21819 ( \22134 , \22133 );
buf \U$21820 ( \22135 , RIc0c7d10_58);
buf \U$21821 ( \22136 , RIc0c7c98_59);
xor \U$21822 ( \22137 , \22135 , \22136 );
xor \U$21823 ( \22138 , \22136 , \22114 );
not \U$21824 ( \22139 , \22138 );
and \U$21825 ( \22140 , \22137 , \22139 );
and \U$21826 ( \22141 , \22134 , \22140 );
xor \U$21827 ( \22142 , \21636 , \21637 );
xor \U$21828 ( \22143 , \22142 , \21935 );
buf \U$21829 ( \22144 , \22143 );
buf \U$21830 ( \22145 , \22144 );
and \U$21831 ( \22146 , \22145 , \22138 );
nor \U$21832 ( \22147 , \22141 , \22146 );
and \U$21833 ( \22148 , \22136 , \22114 );
not \U$21834 ( \22149 , \22148 );
and \U$21835 ( \22150 , \22135 , \22149 );
xnor \U$21836 ( \22151 , \22147 , \22150 );
and \U$21837 ( \22152 , \22130 , \22151 );
xor \U$21838 ( \22153 , \21645 , \21646 );
xor \U$21839 ( \22154 , \22153 , \21926 );
buf \U$21840 ( \22155 , \22154 );
buf \U$21841 ( \22156 , \22155 );
buf \U$21842 ( \22157 , RIc0c7e00_56);
buf \U$21843 ( \22158 , RIc0c7d88_57);
xor \U$21844 ( \22159 , \22157 , \22158 );
xor \U$21845 ( \22160 , \22158 , \22135 );
not \U$21846 ( \22161 , \22160 );
and \U$21847 ( \22162 , \22159 , \22161 );
and \U$21848 ( \22163 , \22156 , \22162 );
xor \U$21849 ( \22164 , \21642 , \21643 );
xor \U$21850 ( \22165 , \22164 , \21929 );
buf \U$21851 ( \22166 , \22165 );
buf \U$21852 ( \22167 , \22166 );
and \U$21853 ( \22168 , \22167 , \22160 );
nor \U$21854 ( \22169 , \22163 , \22168 );
and \U$21855 ( \22170 , \22158 , \22135 );
not \U$21856 ( \22171 , \22170 );
and \U$21857 ( \22172 , \22157 , \22171 );
xnor \U$21858 ( \22173 , \22169 , \22172 );
and \U$21859 ( \22174 , \22151 , \22173 );
and \U$21860 ( \22175 , \22130 , \22173 );
or \U$21861 ( \22176 , \22152 , \22174 , \22175 );
and \U$21862 ( \22177 , \22109 , \22176 );
xor \U$21863 ( \22178 , \21651 , \21652 );
xor \U$21864 ( \22179 , \22178 , \21920 );
buf \U$21865 ( \22180 , \22179 );
buf \U$21866 ( \22181 , \22180 );
buf \U$21867 ( \22182 , RIc0c7ef0_54);
buf \U$21868 ( \22183 , RIc0c7e78_55);
xor \U$21869 ( \22184 , \22182 , \22183 );
xor \U$21870 ( \22185 , \22183 , \22157 );
not \U$21871 ( \22186 , \22185 );
and \U$21872 ( \22187 , \22184 , \22186 );
and \U$21873 ( \22188 , \22181 , \22187 );
xor \U$21874 ( \22189 , \21648 , \21649 );
xor \U$21875 ( \22190 , \22189 , \21923 );
buf \U$21876 ( \22191 , \22190 );
buf \U$21877 ( \22192 , \22191 );
and \U$21878 ( \22193 , \22192 , \22185 );
nor \U$21879 ( \22194 , \22188 , \22193 );
and \U$21880 ( \22195 , \22183 , \22157 );
not \U$21881 ( \22196 , \22195 );
and \U$21882 ( \22197 , \22182 , \22196 );
xnor \U$21883 ( \22198 , \22194 , \22197 );
xor \U$21884 ( \22199 , \21657 , \21658 );
xor \U$21885 ( \22200 , \22199 , \21914 );
buf \U$21886 ( \22201 , \22200 );
buf \U$21887 ( \22202 , \22201 );
buf \U$21888 ( \22203 , RIc0c7fe0_52);
buf \U$21889 ( \22204 , RIc0c7f68_53);
xor \U$21890 ( \22205 , \22203 , \22204 );
xor \U$21891 ( \22206 , \22204 , \22182 );
not \U$21892 ( \22207 , \22206 );
and \U$21893 ( \22208 , \22205 , \22207 );
and \U$21894 ( \22209 , \22202 , \22208 );
xor \U$21895 ( \22210 , \21654 , \21655 );
xor \U$21896 ( \22211 , \22210 , \21917 );
buf \U$21897 ( \22212 , \22211 );
buf \U$21898 ( \22213 , \22212 );
and \U$21899 ( \22214 , \22213 , \22206 );
nor \U$21900 ( \22215 , \22209 , \22214 );
and \U$21901 ( \22216 , \22204 , \22182 );
not \U$21902 ( \22217 , \22216 );
and \U$21903 ( \22218 , \22203 , \22217 );
xnor \U$21904 ( \22219 , \22215 , \22218 );
and \U$21905 ( \22220 , \22198 , \22219 );
xor \U$21906 ( \22221 , \21663 , \21664 );
xor \U$21907 ( \22222 , \22221 , \21908 );
buf \U$21908 ( \22223 , \22222 );
buf \U$21909 ( \22224 , \22223 );
buf \U$21910 ( \22225 , RIc0c80d0_50);
buf \U$21911 ( \22226 , RIc0c8058_51);
xor \U$21912 ( \22227 , \22225 , \22226 );
xor \U$21913 ( \22228 , \22226 , \22203 );
not \U$21914 ( \22229 , \22228 );
and \U$21915 ( \22230 , \22227 , \22229 );
and \U$21916 ( \22231 , \22224 , \22230 );
xor \U$21917 ( \22232 , \21660 , \21661 );
xor \U$21918 ( \22233 , \22232 , \21911 );
buf \U$21919 ( \22234 , \22233 );
buf \U$21920 ( \22235 , \22234 );
and \U$21921 ( \22236 , \22235 , \22228 );
nor \U$21922 ( \22237 , \22231 , \22236 );
and \U$21923 ( \22238 , \22226 , \22203 );
not \U$21924 ( \22239 , \22238 );
and \U$21925 ( \22240 , \22225 , \22239 );
xnor \U$21926 ( \22241 , \22237 , \22240 );
and \U$21927 ( \22242 , \22219 , \22241 );
and \U$21928 ( \22243 , \22198 , \22241 );
or \U$21929 ( \22244 , \22220 , \22242 , \22243 );
and \U$21930 ( \22245 , \22176 , \22244 );
and \U$21931 ( \22246 , \22109 , \22244 );
or \U$21932 ( \22247 , \22177 , \22245 , \22246 );
xor \U$21933 ( \22248 , \21669 , \21670 );
xor \U$21934 ( \22249 , \22248 , \21902 );
buf \U$21935 ( \22250 , \22249 );
buf \U$21936 ( \22251 , \22250 );
buf \U$21937 ( \22252 , RIc0c81c0_48);
buf \U$21938 ( \22253 , RIc0c8148_49);
xor \U$21939 ( \22254 , \22252 , \22253 );
xor \U$21940 ( \22255 , \22253 , \22225 );
not \U$21941 ( \22256 , \22255 );
and \U$21942 ( \22257 , \22254 , \22256 );
and \U$21943 ( \22258 , \22251 , \22257 );
xor \U$21944 ( \22259 , \21666 , \21667 );
xor \U$21945 ( \22260 , \22259 , \21905 );
buf \U$21946 ( \22261 , \22260 );
buf \U$21947 ( \22262 , \22261 );
and \U$21948 ( \22263 , \22262 , \22255 );
nor \U$21949 ( \22264 , \22258 , \22263 );
and \U$21950 ( \22265 , \22253 , \22225 );
not \U$21951 ( \22266 , \22265 );
and \U$21952 ( \22267 , \22252 , \22266 );
xnor \U$21953 ( \22268 , \22264 , \22267 );
xor \U$21954 ( \22269 , \21675 , \21676 );
xor \U$21955 ( \22270 , \22269 , \21896 );
buf \U$21956 ( \22271 , \22270 );
buf \U$21957 ( \22272 , \22271 );
buf \U$21958 ( \22273 , RIc0c82b0_46);
buf \U$21959 ( \22274 , RIc0c8238_47);
xor \U$21960 ( \22275 , \22273 , \22274 );
xor \U$21961 ( \22276 , \22274 , \22252 );
not \U$21962 ( \22277 , \22276 );
and \U$21963 ( \22278 , \22275 , \22277 );
and \U$21964 ( \22279 , \22272 , \22278 );
xor \U$21965 ( \22280 , \21672 , \21673 );
xor \U$21966 ( \22281 , \22280 , \21899 );
buf \U$21967 ( \22282 , \22281 );
buf \U$21968 ( \22283 , \22282 );
and \U$21969 ( \22284 , \22283 , \22276 );
nor \U$21970 ( \22285 , \22279 , \22284 );
and \U$21971 ( \22286 , \22274 , \22252 );
not \U$21972 ( \22287 , \22286 );
and \U$21973 ( \22288 , \22273 , \22287 );
xnor \U$21974 ( \22289 , \22285 , \22288 );
and \U$21975 ( \22290 , \22268 , \22289 );
xor \U$21976 ( \22291 , \21681 , \21682 );
xor \U$21977 ( \22292 , \22291 , \21890 );
buf \U$21978 ( \22293 , \22292 );
buf \U$21979 ( \22294 , \22293 );
buf \U$21980 ( \22295 , RIc0c83a0_44);
buf \U$21981 ( \22296 , RIc0c8328_45);
xor \U$21982 ( \22297 , \22295 , \22296 );
xor \U$21983 ( \22298 , \22296 , \22273 );
not \U$21984 ( \22299 , \22298 );
and \U$21985 ( \22300 , \22297 , \22299 );
and \U$21986 ( \22301 , \22294 , \22300 );
xor \U$21987 ( \22302 , \21678 , \21679 );
xor \U$21988 ( \22303 , \22302 , \21893 );
buf \U$21989 ( \22304 , \22303 );
buf \U$21990 ( \22305 , \22304 );
and \U$21991 ( \22306 , \22305 , \22298 );
nor \U$21992 ( \22307 , \22301 , \22306 );
and \U$21993 ( \22308 , \22296 , \22273 );
not \U$21994 ( \22309 , \22308 );
and \U$21995 ( \22310 , \22295 , \22309 );
xnor \U$21996 ( \22311 , \22307 , \22310 );
and \U$21997 ( \22312 , \22289 , \22311 );
and \U$21998 ( \22313 , \22268 , \22311 );
or \U$21999 ( \22314 , \22290 , \22312 , \22313 );
xor \U$22000 ( \22315 , \21687 , \21688 );
xor \U$22001 ( \22316 , \22315 , \21884 );
buf \U$22002 ( \22317 , \22316 );
buf \U$22003 ( \22318 , \22317 );
buf \U$22004 ( \22319 , RIc0c8490_42);
buf \U$22005 ( \22320 , RIc0c8418_43);
xor \U$22006 ( \22321 , \22319 , \22320 );
xor \U$22007 ( \22322 , \22320 , \22295 );
not \U$22008 ( \22323 , \22322 );
and \U$22009 ( \22324 , \22321 , \22323 );
and \U$22010 ( \22325 , \22318 , \22324 );
xor \U$22011 ( \22326 , \21684 , \21685 );
xor \U$22012 ( \22327 , \22326 , \21887 );
buf \U$22013 ( \22328 , \22327 );
buf \U$22014 ( \22329 , \22328 );
and \U$22015 ( \22330 , \22329 , \22322 );
nor \U$22016 ( \22331 , \22325 , \22330 );
and \U$22017 ( \22332 , \22320 , \22295 );
not \U$22018 ( \22333 , \22332 );
and \U$22019 ( \22334 , \22319 , \22333 );
xnor \U$22020 ( \22335 , \22331 , \22334 );
xor \U$22021 ( \22336 , \21693 , \21694 );
xor \U$22022 ( \22337 , \22336 , \21878 );
buf \U$22023 ( \22338 , \22337 );
buf \U$22024 ( \22339 , \22338 );
buf \U$22025 ( \22340 , RIc0c8580_40);
buf \U$22026 ( \22341 , RIc0c8508_41);
xor \U$22027 ( \22342 , \22340 , \22341 );
xor \U$22028 ( \22343 , \22341 , \22319 );
not \U$22029 ( \22344 , \22343 );
and \U$22030 ( \22345 , \22342 , \22344 );
and \U$22031 ( \22346 , \22339 , \22345 );
xor \U$22032 ( \22347 , \21690 , \21691 );
xor \U$22033 ( \22348 , \22347 , \21881 );
buf \U$22034 ( \22349 , \22348 );
buf \U$22035 ( \22350 , \22349 );
and \U$22036 ( \22351 , \22350 , \22343 );
nor \U$22037 ( \22352 , \22346 , \22351 );
and \U$22038 ( \22353 , \22341 , \22319 );
not \U$22039 ( \22354 , \22353 );
and \U$22040 ( \22355 , \22340 , \22354 );
xnor \U$22041 ( \22356 , \22352 , \22355 );
and \U$22042 ( \22357 , \22335 , \22356 );
xor \U$22043 ( \22358 , \21699 , \21700 );
xor \U$22044 ( \22359 , \22358 , \21872 );
buf \U$22045 ( \22360 , \22359 );
buf \U$22046 ( \22361 , \22360 );
buf \U$22047 ( \22362 , RIc0c8670_38);
buf \U$22048 ( \22363 , RIc0c85f8_39);
xor \U$22049 ( \22364 , \22362 , \22363 );
xor \U$22050 ( \22365 , \22363 , \22340 );
not \U$22051 ( \22366 , \22365 );
and \U$22052 ( \22367 , \22364 , \22366 );
and \U$22053 ( \22368 , \22361 , \22367 );
xor \U$22054 ( \22369 , \21696 , \21697 );
xor \U$22055 ( \22370 , \22369 , \21875 );
buf \U$22056 ( \22371 , \22370 );
buf \U$22057 ( \22372 , \22371 );
and \U$22058 ( \22373 , \22372 , \22365 );
nor \U$22059 ( \22374 , \22368 , \22373 );
and \U$22060 ( \22375 , \22363 , \22340 );
not \U$22061 ( \22376 , \22375 );
and \U$22062 ( \22377 , \22362 , \22376 );
xnor \U$22063 ( \22378 , \22374 , \22377 );
and \U$22064 ( \22379 , \22356 , \22378 );
and \U$22065 ( \22380 , \22335 , \22378 );
or \U$22066 ( \22381 , \22357 , \22379 , \22380 );
and \U$22067 ( \22382 , \22314 , \22381 );
xor \U$22068 ( \22383 , \21705 , \21706 );
xor \U$22069 ( \22384 , \22383 , \21866 );
buf \U$22070 ( \22385 , \22384 );
buf \U$22071 ( \22386 , \22385 );
buf \U$22072 ( \22387 , RIc0c8760_36);
buf \U$22073 ( \22388 , RIc0c86e8_37);
xor \U$22074 ( \22389 , \22387 , \22388 );
xor \U$22075 ( \22390 , \22388 , \22362 );
not \U$22076 ( \22391 , \22390 );
and \U$22077 ( \22392 , \22389 , \22391 );
and \U$22078 ( \22393 , \22386 , \22392 );
xor \U$22079 ( \22394 , \21702 , \21703 );
xor \U$22080 ( \22395 , \22394 , \21869 );
buf \U$22081 ( \22396 , \22395 );
buf \U$22082 ( \22397 , \22396 );
and \U$22083 ( \22398 , \22397 , \22390 );
nor \U$22084 ( \22399 , \22393 , \22398 );
and \U$22085 ( \22400 , \22388 , \22362 );
not \U$22086 ( \22401 , \22400 );
and \U$22087 ( \22402 , \22387 , \22401 );
xnor \U$22088 ( \22403 , \22399 , \22402 );
xor \U$22089 ( \22404 , \21711 , \21712 );
xor \U$22090 ( \22405 , \22404 , \21860 );
buf \U$22091 ( \22406 , \22405 );
buf \U$22092 ( \22407 , \22406 );
buf \U$22093 ( \22408 , RIc0c8850_34);
buf \U$22094 ( \22409 , RIc0c87d8_35);
xor \U$22095 ( \22410 , \22408 , \22409 );
xor \U$22096 ( \22411 , \22409 , \22387 );
not \U$22097 ( \22412 , \22411 );
and \U$22098 ( \22413 , \22410 , \22412 );
and \U$22099 ( \22414 , \22407 , \22413 );
xor \U$22100 ( \22415 , \21708 , \21709 );
xor \U$22101 ( \22416 , \22415 , \21863 );
buf \U$22102 ( \22417 , \22416 );
buf \U$22103 ( \22418 , \22417 );
and \U$22104 ( \22419 , \22418 , \22411 );
nor \U$22105 ( \22420 , \22414 , \22419 );
and \U$22106 ( \22421 , \22409 , \22387 );
not \U$22107 ( \22422 , \22421 );
and \U$22108 ( \22423 , \22408 , \22422 );
xnor \U$22109 ( \22424 , \22420 , \22423 );
and \U$22110 ( \22425 , \22403 , \22424 );
xor \U$22111 ( \22426 , \21717 , \21718 );
xor \U$22112 ( \22427 , \22426 , \21854 );
buf \U$22113 ( \22428 , \22427 );
buf \U$22114 ( \22429 , \22428 );
buf \U$22115 ( \22430 , RIc0c8940_32);
buf \U$22116 ( \22431 , RIc0c88c8_33);
xor \U$22117 ( \22432 , \22430 , \22431 );
xor \U$22118 ( \22433 , \22431 , \22408 );
not \U$22119 ( \22434 , \22433 );
and \U$22120 ( \22435 , \22432 , \22434 );
and \U$22121 ( \22436 , \22429 , \22435 );
xor \U$22122 ( \22437 , \21714 , \21715 );
xor \U$22123 ( \22438 , \22437 , \21857 );
buf \U$22124 ( \22439 , \22438 );
buf \U$22125 ( \22440 , \22439 );
and \U$22126 ( \22441 , \22440 , \22433 );
nor \U$22127 ( \22442 , \22436 , \22441 );
and \U$22128 ( \22443 , \22431 , \22408 );
not \U$22129 ( \22444 , \22443 );
and \U$22130 ( \22445 , \22430 , \22444 );
xnor \U$22131 ( \22446 , \22442 , \22445 );
and \U$22132 ( \22447 , \22424 , \22446 );
and \U$22133 ( \22448 , \22403 , \22446 );
or \U$22134 ( \22449 , \22425 , \22447 , \22448 );
and \U$22135 ( \22450 , \22381 , \22449 );
and \U$22136 ( \22451 , \22314 , \22449 );
or \U$22137 ( \22452 , \22382 , \22450 , \22451 );
and \U$22138 ( \22453 , \22247 , \22452 );
xor \U$22139 ( \22454 , \21723 , \21724 );
xor \U$22140 ( \22455 , \22454 , \21848 );
buf \U$22141 ( \22456 , \22455 );
buf \U$22142 ( \22457 , \22456 );
buf \U$22143 ( \22458 , RIc0c8a30_30);
buf \U$22144 ( \22459 , RIc0c89b8_31);
xor \U$22145 ( \22460 , \22458 , \22459 );
xor \U$22146 ( \22461 , \22459 , \22430 );
not \U$22147 ( \22462 , \22461 );
and \U$22148 ( \22463 , \22460 , \22462 );
and \U$22149 ( \22464 , \22457 , \22463 );
xor \U$22150 ( \22465 , \21720 , \21721 );
xor \U$22151 ( \22466 , \22465 , \21851 );
buf \U$22152 ( \22467 , \22466 );
buf \U$22153 ( \22468 , \22467 );
and \U$22154 ( \22469 , \22468 , \22461 );
nor \U$22155 ( \22470 , \22464 , \22469 );
and \U$22156 ( \22471 , \22459 , \22430 );
not \U$22157 ( \22472 , \22471 );
and \U$22158 ( \22473 , \22458 , \22472 );
xnor \U$22159 ( \22474 , \22470 , \22473 );
xor \U$22160 ( \22475 , \21729 , \21730 );
xor \U$22161 ( \22476 , \22475 , \21842 );
buf \U$22162 ( \22477 , \22476 );
buf \U$22163 ( \22478 , \22477 );
buf \U$22164 ( \22479 , RIc0c8b20_28);
buf \U$22165 ( \22480 , RIc0c8aa8_29);
xor \U$22166 ( \22481 , \22479 , \22480 );
xor \U$22167 ( \22482 , \22480 , \22458 );
not \U$22168 ( \22483 , \22482 );
and \U$22169 ( \22484 , \22481 , \22483 );
and \U$22170 ( \22485 , \22478 , \22484 );
xor \U$22171 ( \22486 , \21726 , \21727 );
xor \U$22172 ( \22487 , \22486 , \21845 );
buf \U$22173 ( \22488 , \22487 );
buf \U$22174 ( \22489 , \22488 );
and \U$22175 ( \22490 , \22489 , \22482 );
nor \U$22176 ( \22491 , \22485 , \22490 );
and \U$22177 ( \22492 , \22480 , \22458 );
not \U$22178 ( \22493 , \22492 );
and \U$22179 ( \22494 , \22479 , \22493 );
xnor \U$22180 ( \22495 , \22491 , \22494 );
and \U$22181 ( \22496 , \22474 , \22495 );
xor \U$22182 ( \22497 , \21735 , \21736 );
xor \U$22183 ( \22498 , \22497 , \21836 );
buf \U$22184 ( \22499 , \22498 );
buf \U$22185 ( \22500 , \22499 );
buf \U$22186 ( \22501 , RIc0c8c10_26);
buf \U$22187 ( \22502 , RIc0c8b98_27);
xor \U$22188 ( \22503 , \22501 , \22502 );
xor \U$22189 ( \22504 , \22502 , \22479 );
not \U$22190 ( \22505 , \22504 );
and \U$22191 ( \22506 , \22503 , \22505 );
and \U$22192 ( \22507 , \22500 , \22506 );
xor \U$22193 ( \22508 , \21732 , \21733 );
xor \U$22194 ( \22509 , \22508 , \21839 );
buf \U$22195 ( \22510 , \22509 );
buf \U$22196 ( \22511 , \22510 );
and \U$22197 ( \22512 , \22511 , \22504 );
nor \U$22198 ( \22513 , \22507 , \22512 );
and \U$22199 ( \22514 , \22502 , \22479 );
not \U$22200 ( \22515 , \22514 );
and \U$22201 ( \22516 , \22501 , \22515 );
xnor \U$22202 ( \22517 , \22513 , \22516 );
and \U$22203 ( \22518 , \22495 , \22517 );
and \U$22204 ( \22519 , \22474 , \22517 );
or \U$22205 ( \22520 , \22496 , \22518 , \22519 );
xor \U$22206 ( \22521 , \21741 , \21742 );
xor \U$22207 ( \22522 , \22521 , \21830 );
buf \U$22208 ( \22523 , \22522 );
buf \U$22209 ( \22524 , \22523 );
buf \U$22210 ( \22525 , RIc0c8d00_24);
buf \U$22211 ( \22526 , RIc0c8c88_25);
xor \U$22212 ( \22527 , \22525 , \22526 );
xor \U$22213 ( \22528 , \22526 , \22501 );
not \U$22214 ( \22529 , \22528 );
and \U$22215 ( \22530 , \22527 , \22529 );
and \U$22216 ( \22531 , \22524 , \22530 );
xor \U$22217 ( \22532 , \21738 , \21739 );
xor \U$22218 ( \22533 , \22532 , \21833 );
buf \U$22219 ( \22534 , \22533 );
buf \U$22220 ( \22535 , \22534 );
and \U$22221 ( \22536 , \22535 , \22528 );
nor \U$22222 ( \22537 , \22531 , \22536 );
and \U$22223 ( \22538 , \22526 , \22501 );
not \U$22224 ( \22539 , \22538 );
and \U$22225 ( \22540 , \22525 , \22539 );
xnor \U$22226 ( \22541 , \22537 , \22540 );
xor \U$22227 ( \22542 , \21747 , \21748 );
xor \U$22228 ( \22543 , \22542 , \21824 );
buf \U$22229 ( \22544 , \22543 );
buf \U$22230 ( \22545 , \22544 );
buf \U$22231 ( \22546 , RIc0c8df0_22);
buf \U$22232 ( \22547 , RIc0c8d78_23);
xor \U$22233 ( \22548 , \22546 , \22547 );
xor \U$22234 ( \22549 , \22547 , \22525 );
not \U$22235 ( \22550 , \22549 );
and \U$22236 ( \22551 , \22548 , \22550 );
and \U$22237 ( \22552 , \22545 , \22551 );
xor \U$22238 ( \22553 , \21744 , \21745 );
xor \U$22239 ( \22554 , \22553 , \21827 );
buf \U$22240 ( \22555 , \22554 );
buf \U$22241 ( \22556 , \22555 );
and \U$22242 ( \22557 , \22556 , \22549 );
nor \U$22243 ( \22558 , \22552 , \22557 );
and \U$22244 ( \22559 , \22547 , \22525 );
not \U$22245 ( \22560 , \22559 );
and \U$22246 ( \22561 , \22546 , \22560 );
xnor \U$22247 ( \22562 , \22558 , \22561 );
and \U$22248 ( \22563 , \22541 , \22562 );
xor \U$22249 ( \22564 , \21753 , \21754 );
xor \U$22250 ( \22565 , \22564 , \21818 );
buf \U$22251 ( \22566 , \22565 );
buf \U$22252 ( \22567 , \22566 );
buf \U$22253 ( \22568 , RIc0c8ee0_20);
buf \U$22254 ( \22569 , RIc0c8e68_21);
xor \U$22255 ( \22570 , \22568 , \22569 );
xor \U$22256 ( \22571 , \22569 , \22546 );
not \U$22257 ( \22572 , \22571 );
and \U$22258 ( \22573 , \22570 , \22572 );
and \U$22259 ( \22574 , \22567 , \22573 );
xor \U$22260 ( \22575 , \21750 , \21751 );
xor \U$22261 ( \22576 , \22575 , \21821 );
buf \U$22262 ( \22577 , \22576 );
buf \U$22263 ( \22578 , \22577 );
and \U$22264 ( \22579 , \22578 , \22571 );
nor \U$22265 ( \22580 , \22574 , \22579 );
and \U$22266 ( \22581 , \22569 , \22546 );
not \U$22267 ( \22582 , \22581 );
and \U$22268 ( \22583 , \22568 , \22582 );
xnor \U$22269 ( \22584 , \22580 , \22583 );
and \U$22270 ( \22585 , \22562 , \22584 );
and \U$22271 ( \22586 , \22541 , \22584 );
or \U$22272 ( \22587 , \22563 , \22585 , \22586 );
and \U$22273 ( \22588 , \22520 , \22587 );
xor \U$22274 ( \22589 , \21759 , \21760 );
xor \U$22275 ( \22590 , \22589 , \21812 );
buf \U$22276 ( \22591 , \22590 );
buf \U$22277 ( \22592 , \22591 );
buf \U$22278 ( \22593 , RIc0c8fd0_18);
buf \U$22279 ( \22594 , RIc0c8f58_19);
xor \U$22280 ( \22595 , \22593 , \22594 );
xor \U$22281 ( \22596 , \22594 , \22568 );
not \U$22282 ( \22597 , \22596 );
and \U$22283 ( \22598 , \22595 , \22597 );
and \U$22284 ( \22599 , \22592 , \22598 );
xor \U$22285 ( \22600 , \21756 , \21757 );
xor \U$22286 ( \22601 , \22600 , \21815 );
buf \U$22287 ( \22602 , \22601 );
buf \U$22288 ( \22603 , \22602 );
and \U$22289 ( \22604 , \22603 , \22596 );
nor \U$22290 ( \22605 , \22599 , \22604 );
and \U$22291 ( \22606 , \22594 , \22568 );
not \U$22292 ( \22607 , \22606 );
and \U$22293 ( \22608 , \22593 , \22607 );
xnor \U$22294 ( \22609 , \22605 , \22608 );
xor \U$22295 ( \22610 , \21765 , \21766 );
xor \U$22296 ( \22611 , \22610 , \21806 );
buf \U$22297 ( \22612 , \22611 );
buf \U$22298 ( \22613 , \22612 );
buf \U$22299 ( \22614 , RIc0c90c0_16);
buf \U$22300 ( \22615 , RIc0c9048_17);
xor \U$22301 ( \22616 , \22614 , \22615 );
xor \U$22302 ( \22617 , \22615 , \22593 );
not \U$22303 ( \22618 , \22617 );
and \U$22304 ( \22619 , \22616 , \22618 );
and \U$22305 ( \22620 , \22613 , \22619 );
xor \U$22306 ( \22621 , \21762 , \21763 );
xor \U$22307 ( \22622 , \22621 , \21809 );
buf \U$22308 ( \22623 , \22622 );
buf \U$22309 ( \22624 , \22623 );
and \U$22310 ( \22625 , \22624 , \22617 );
nor \U$22311 ( \22626 , \22620 , \22625 );
and \U$22312 ( \22627 , \22615 , \22593 );
not \U$22313 ( \22628 , \22627 );
and \U$22314 ( \22629 , \22614 , \22628 );
xnor \U$22315 ( \22630 , \22626 , \22629 );
and \U$22316 ( \22631 , \22609 , \22630 );
xor \U$22317 ( \22632 , \21771 , \21772 );
xor \U$22318 ( \22633 , \22632 , \21800 );
buf \U$22319 ( \22634 , \22633 );
buf \U$22320 ( \22635 , \22634 );
buf \U$22321 ( \22636 , RIc0c91b0_14);
buf \U$22322 ( \22637 , RIc0c9138_15);
xor \U$22323 ( \22638 , \22636 , \22637 );
xor \U$22324 ( \22639 , \22637 , \22614 );
not \U$22325 ( \22640 , \22639 );
and \U$22326 ( \22641 , \22638 , \22640 );
and \U$22327 ( \22642 , \22635 , \22641 );
xor \U$22328 ( \22643 , \21768 , \21769 );
xor \U$22329 ( \22644 , \22643 , \21803 );
buf \U$22330 ( \22645 , \22644 );
buf \U$22331 ( \22646 , \22645 );
and \U$22332 ( \22647 , \22646 , \22639 );
nor \U$22333 ( \22648 , \22642 , \22647 );
and \U$22334 ( \22649 , \22637 , \22614 );
not \U$22335 ( \22650 , \22649 );
and \U$22336 ( \22651 , \22636 , \22650 );
xnor \U$22337 ( \22652 , \22648 , \22651 );
and \U$22338 ( \22653 , \22630 , \22652 );
and \U$22339 ( \22654 , \22609 , \22652 );
or \U$22340 ( \22655 , \22631 , \22653 , \22654 );
and \U$22341 ( \22656 , \22587 , \22655 );
and \U$22342 ( \22657 , \22520 , \22655 );
or \U$22343 ( \22658 , \22588 , \22656 , \22657 );
and \U$22344 ( \22659 , \22452 , \22658 );
and \U$22345 ( \22660 , \22247 , \22658 );
or \U$22346 ( \22661 , \22453 , \22659 , \22660 );
xor \U$22347 ( \22662 , \21777 , \21778 );
xor \U$22348 ( \22663 , \22662 , \21794 );
buf \U$22349 ( \22664 , \22663 );
buf \U$22350 ( \22665 , \22664 );
buf \U$22351 ( \22666 , RIc0c92a0_12);
buf \U$22352 ( \22667 , RIc0c9228_13);
xor \U$22353 ( \22668 , \22666 , \22667 );
xor \U$22354 ( \22669 , \22667 , \22636 );
not \U$22355 ( \22670 , \22669 );
and \U$22356 ( \22671 , \22668 , \22670 );
and \U$22357 ( \22672 , \22665 , \22671 );
xor \U$22358 ( \22673 , \21774 , \21775 );
xor \U$22359 ( \22674 , \22673 , \21797 );
buf \U$22360 ( \22675 , \22674 );
buf \U$22361 ( \22676 , \22675 );
and \U$22362 ( \22677 , \22676 , \22669 );
nor \U$22363 ( \22678 , \22672 , \22677 );
and \U$22364 ( \22679 , \22667 , \22636 );
not \U$22365 ( \22680 , \22679 );
and \U$22366 ( \22681 , \22666 , \22680 );
xnor \U$22367 ( \22682 , \22678 , \22681 );
xor \U$22368 ( \22683 , \21783 , \21784 );
xor \U$22369 ( \22684 , \22683 , \21788 );
buf \U$22370 ( \22685 , \22684 );
buf \U$22371 ( \22686 , \22685 );
buf \U$22372 ( \22687 , RIc0c9318_11);
xor \U$22373 ( \22688 , \22064 , \22687 );
xor \U$22374 ( \22689 , \22687 , \22666 );
not \U$22375 ( \22690 , \22689 );
and \U$22376 ( \22691 , \22688 , \22690 );
and \U$22377 ( \22692 , \22686 , \22691 );
xor \U$22378 ( \22693 , \21780 , \21781 );
xor \U$22379 ( \22694 , \22693 , \21791 );
buf \U$22380 ( \22695 , \22694 );
buf \U$22381 ( \22696 , \22695 );
and \U$22382 ( \22697 , \22696 , \22689 );
nor \U$22383 ( \22698 , \22692 , \22697 );
and \U$22384 ( \22699 , \22687 , \22666 );
not \U$22385 ( \22700 , \22699 );
and \U$22386 ( \22701 , \22064 , \22700 );
xnor \U$22387 ( \22702 , \22698 , \22701 );
and \U$22388 ( \22703 , \22682 , \22702 );
xor \U$22389 ( \22704 , \21786 , \21787 );
buf \U$22390 ( \22705 , \22704 );
buf \U$22391 ( \22706 , \22705 );
xor \U$22392 ( \22707 , \22063 , \22064 );
nand \U$22393 ( \22708 , \22706 , \22707 );
xnor \U$22394 ( \22709 , \22708 , \22067 );
and \U$22395 ( \22710 , \22702 , \22709 );
and \U$22396 ( \22711 , \22682 , \22709 );
or \U$22397 ( \22712 , \22703 , \22710 , \22711 );
and \U$22398 ( \22713 , \22696 , \22691 );
and \U$22399 ( \22714 , \22665 , \22689 );
nor \U$22400 ( \22715 , \22713 , \22714 );
xnor \U$22401 ( \22716 , \22715 , \22701 );
and \U$22402 ( \22717 , \22712 , \22716 );
xor \U$22403 ( \22718 , \22013 , \22063 );
not \U$22404 ( \22719 , \22707 );
and \U$22405 ( \22720 , \22718 , \22719 );
and \U$22406 ( \22721 , \22706 , \22720 );
and \U$22407 ( \22722 , \22686 , \22707 );
nor \U$22408 ( \22723 , \22721 , \22722 );
xnor \U$22409 ( \22724 , \22723 , \22067 );
and \U$22410 ( \22725 , \22716 , \22724 );
and \U$22411 ( \22726 , \22712 , \22724 );
or \U$22412 ( \22727 , \22717 , \22725 , \22726 );
and \U$22413 ( \22728 , \22624 , \22619 );
and \U$22414 ( \22729 , \22592 , \22617 );
nor \U$22415 ( \22730 , \22728 , \22729 );
xnor \U$22416 ( \22731 , \22730 , \22629 );
and \U$22417 ( \22732 , \22646 , \22641 );
and \U$22418 ( \22733 , \22613 , \22639 );
nor \U$22419 ( \22734 , \22732 , \22733 );
xnor \U$22420 ( \22735 , \22734 , \22651 );
xor \U$22421 ( \22736 , \22731 , \22735 );
and \U$22422 ( \22737 , \22676 , \22671 );
and \U$22423 ( \22738 , \22635 , \22669 );
nor \U$22424 ( \22739 , \22737 , \22738 );
xnor \U$22425 ( \22740 , \22739 , \22681 );
xor \U$22426 ( \22741 , \22736 , \22740 );
and \U$22427 ( \22742 , \22556 , \22551 );
and \U$22428 ( \22743 , \22524 , \22549 );
nor \U$22429 ( \22744 , \22742 , \22743 );
xnor \U$22430 ( \22745 , \22744 , \22561 );
and \U$22431 ( \22746 , \22578 , \22573 );
and \U$22432 ( \22747 , \22545 , \22571 );
nor \U$22433 ( \22748 , \22746 , \22747 );
xnor \U$22434 ( \22749 , \22748 , \22583 );
xor \U$22435 ( \22750 , \22745 , \22749 );
and \U$22436 ( \22751 , \22603 , \22598 );
and \U$22437 ( \22752 , \22567 , \22596 );
nor \U$22438 ( \22753 , \22751 , \22752 );
xnor \U$22439 ( \22754 , \22753 , \22608 );
xor \U$22440 ( \22755 , \22750 , \22754 );
and \U$22441 ( \22756 , \22741 , \22755 );
and \U$22442 ( \22757 , \22489 , \22484 );
and \U$22443 ( \22758 , \22457 , \22482 );
nor \U$22444 ( \22759 , \22757 , \22758 );
xnor \U$22445 ( \22760 , \22759 , \22494 );
and \U$22446 ( \22761 , \22511 , \22506 );
and \U$22447 ( \22762 , \22478 , \22504 );
nor \U$22448 ( \22763 , \22761 , \22762 );
xnor \U$22449 ( \22764 , \22763 , \22516 );
xor \U$22450 ( \22765 , \22760 , \22764 );
and \U$22451 ( \22766 , \22535 , \22530 );
and \U$22452 ( \22767 , \22500 , \22528 );
nor \U$22453 ( \22768 , \22766 , \22767 );
xnor \U$22454 ( \22769 , \22768 , \22540 );
xor \U$22455 ( \22770 , \22765 , \22769 );
and \U$22456 ( \22771 , \22755 , \22770 );
and \U$22457 ( \22772 , \22741 , \22770 );
or \U$22458 ( \22773 , \22756 , \22771 , \22772 );
and \U$22459 ( \22774 , \22727 , \22773 );
and \U$22460 ( \22775 , \22418 , \22413 );
and \U$22461 ( \22776 , \22386 , \22411 );
nor \U$22462 ( \22777 , \22775 , \22776 );
xnor \U$22463 ( \22778 , \22777 , \22423 );
and \U$22464 ( \22779 , \22440 , \22435 );
and \U$22465 ( \22780 , \22407 , \22433 );
nor \U$22466 ( \22781 , \22779 , \22780 );
xnor \U$22467 ( \22782 , \22781 , \22445 );
xor \U$22468 ( \22783 , \22778 , \22782 );
and \U$22469 ( \22784 , \22468 , \22463 );
and \U$22470 ( \22785 , \22429 , \22461 );
nor \U$22471 ( \22786 , \22784 , \22785 );
xnor \U$22472 ( \22787 , \22786 , \22473 );
xor \U$22473 ( \22788 , \22783 , \22787 );
and \U$22474 ( \22789 , \22350 , \22345 );
and \U$22475 ( \22790 , \22318 , \22343 );
nor \U$22476 ( \22791 , \22789 , \22790 );
xnor \U$22477 ( \22792 , \22791 , \22355 );
and \U$22478 ( \22793 , \22372 , \22367 );
and \U$22479 ( \22794 , \22339 , \22365 );
nor \U$22480 ( \22795 , \22793 , \22794 );
xnor \U$22481 ( \22796 , \22795 , \22377 );
xor \U$22482 ( \22797 , \22792 , \22796 );
and \U$22483 ( \22798 , \22397 , \22392 );
and \U$22484 ( \22799 , \22361 , \22390 );
nor \U$22485 ( \22800 , \22798 , \22799 );
xnor \U$22486 ( \22801 , \22800 , \22402 );
xor \U$22487 ( \22802 , \22797 , \22801 );
and \U$22488 ( \22803 , \22788 , \22802 );
and \U$22489 ( \22804 , \22283 , \22278 );
and \U$22490 ( \22805 , \22251 , \22276 );
nor \U$22491 ( \22806 , \22804 , \22805 );
xnor \U$22492 ( \22807 , \22806 , \22288 );
and \U$22493 ( \22808 , \22305 , \22300 );
and \U$22494 ( \22809 , \22272 , \22298 );
nor \U$22495 ( \22810 , \22808 , \22809 );
xnor \U$22496 ( \22811 , \22810 , \22310 );
xor \U$22497 ( \22812 , \22807 , \22811 );
and \U$22498 ( \22813 , \22329 , \22324 );
and \U$22499 ( \22814 , \22294 , \22322 );
nor \U$22500 ( \22815 , \22813 , \22814 );
xnor \U$22501 ( \22816 , \22815 , \22334 );
xor \U$22502 ( \22817 , \22812 , \22816 );
and \U$22503 ( \22818 , \22802 , \22817 );
and \U$22504 ( \22819 , \22788 , \22817 );
or \U$22505 ( \22820 , \22803 , \22818 , \22819 );
and \U$22506 ( \22821 , \22773 , \22820 );
and \U$22507 ( \22822 , \22727 , \22820 );
or \U$22508 ( \22823 , \22774 , \22821 , \22822 );
and \U$22509 ( \22824 , \22661 , \22823 );
and \U$22510 ( \22825 , \22213 , \22208 );
and \U$22511 ( \22826 , \22181 , \22206 );
nor \U$22512 ( \22827 , \22825 , \22826 );
xnor \U$22513 ( \22828 , \22827 , \22218 );
and \U$22514 ( \22829 , \22235 , \22230 );
and \U$22515 ( \22830 , \22202 , \22228 );
nor \U$22516 ( \22831 , \22829 , \22830 );
xnor \U$22517 ( \22832 , \22831 , \22240 );
xor \U$22518 ( \22833 , \22828 , \22832 );
and \U$22519 ( \22834 , \22262 , \22257 );
and \U$22520 ( \22835 , \22224 , \22255 );
nor \U$22521 ( \22836 , \22834 , \22835 );
xnor \U$22522 ( \22837 , \22836 , \22267 );
xor \U$22523 ( \22838 , \22833 , \22837 );
and \U$22524 ( \22839 , \22145 , \22140 );
and \U$22525 ( \22840 , \22113 , \22138 );
nor \U$22526 ( \22841 , \22839 , \22840 );
xnor \U$22527 ( \22842 , \22841 , \22150 );
and \U$22528 ( \22843 , \22167 , \22162 );
and \U$22529 ( \22844 , \22134 , \22160 );
nor \U$22530 ( \22845 , \22843 , \22844 );
xnor \U$22531 ( \22846 , \22845 , \22172 );
xor \U$22532 ( \22847 , \22842 , \22846 );
and \U$22533 ( \22848 , \22192 , \22187 );
and \U$22534 ( \22849 , \22156 , \22185 );
nor \U$22535 ( \22850 , \22848 , \22849 );
xnor \U$22536 ( \22851 , \22850 , \22197 );
xor \U$22537 ( \22852 , \22847 , \22851 );
and \U$22538 ( \22853 , \22838 , \22852 );
and \U$22539 ( \22854 , \22081 , \22076 );
xor \U$22540 ( \22855 , \21615 , \21616 );
xor \U$22541 ( \22856 , \22855 , \21956 );
buf \U$22542 ( \22857 , \22856 );
buf \U$22543 ( \22858 , \22857 );
and \U$22544 ( \22859 , \22858 , \22073 );
nor \U$22545 ( \22860 , \22854 , \22859 );
xnor \U$22546 ( \22861 , \22860 , \22072 );
and \U$22547 ( \22862 , \22100 , \22095 );
and \U$22548 ( \22863 , \22071 , \22093 );
nor \U$22549 ( \22864 , \22862 , \22863 );
xnor \U$22550 ( \22865 , \22864 , \22105 );
xor \U$22551 ( \22866 , \22861 , \22865 );
and \U$22552 ( \22867 , \22124 , \22119 );
and \U$22553 ( \22868 , \22089 , \22117 );
nor \U$22554 ( \22869 , \22867 , \22868 );
xnor \U$22555 ( \22870 , \22869 , \22129 );
xor \U$22556 ( \22871 , \22866 , \22870 );
and \U$22557 ( \22872 , \22852 , \22871 );
and \U$22558 ( \22873 , \22838 , \22871 );
or \U$22559 ( \22874 , \22853 , \22872 , \22873 );
and \U$22560 ( \22875 , \22089 , \22119 );
and \U$22561 ( \22876 , \22100 , \22117 );
nor \U$22562 ( \22877 , \22875 , \22876 );
xnor \U$22563 ( \22878 , \22877 , \22129 );
and \U$22564 ( \22879 , \22113 , \22140 );
and \U$22565 ( \22880 , \22124 , \22138 );
nor \U$22566 ( \22881 , \22879 , \22880 );
xnor \U$22567 ( \22882 , \22881 , \22150 );
xor \U$22568 ( \22883 , \22878 , \22882 );
and \U$22569 ( \22884 , \22134 , \22162 );
and \U$22570 ( \22885 , \22145 , \22160 );
nor \U$22571 ( \22886 , \22884 , \22885 );
xnor \U$22572 ( \22887 , \22886 , \22172 );
xor \U$22573 ( \22888 , \22883 , \22887 );
and \U$22574 ( \22889 , \22874 , \22888 );
and \U$22575 ( \22890 , \22858 , \22076 );
xor \U$22576 ( \22891 , \21612 , \21613 );
xor \U$22577 ( \22892 , \22891 , \21959 );
buf \U$22578 ( \22893 , \22892 );
buf \U$22579 ( \22894 , \22893 );
and \U$22580 ( \22895 , \22894 , \22073 );
nor \U$22581 ( \22896 , \22890 , \22895 );
xnor \U$22582 ( \22897 , \22896 , \22072 );
xor \U$22583 ( \22898 , \22016 , \22897 );
and \U$22584 ( \22899 , \22071 , \22095 );
and \U$22585 ( \22900 , \22081 , \22093 );
nor \U$22586 ( \22901 , \22899 , \22900 );
xnor \U$22587 ( \22902 , \22901 , \22105 );
xor \U$22588 ( \22903 , \22898 , \22902 );
and \U$22589 ( \22904 , \22888 , \22903 );
and \U$22590 ( \22905 , \22874 , \22903 );
or \U$22591 ( \22906 , \22889 , \22904 , \22905 );
and \U$22592 ( \22907 , \22823 , \22906 );
and \U$22593 ( \22908 , \22661 , \22906 );
or \U$22594 ( \22909 , \22824 , \22907 , \22908 );
and \U$22595 ( \22910 , \22294 , \22324 );
and \U$22596 ( \22911 , \22305 , \22322 );
nor \U$22597 ( \22912 , \22910 , \22911 );
xnor \U$22598 ( \22913 , \22912 , \22334 );
and \U$22599 ( \22914 , \22318 , \22345 );
and \U$22600 ( \22915 , \22329 , \22343 );
nor \U$22601 ( \22916 , \22914 , \22915 );
xnor \U$22602 ( \22917 , \22916 , \22355 );
xor \U$22603 ( \22918 , \22913 , \22917 );
and \U$22604 ( \22919 , \22339 , \22367 );
and \U$22605 ( \22920 , \22350 , \22365 );
nor \U$22606 ( \22921 , \22919 , \22920 );
xnor \U$22607 ( \22922 , \22921 , \22377 );
xor \U$22608 ( \22923 , \22918 , \22922 );
and \U$22609 ( \22924 , \22224 , \22257 );
and \U$22610 ( \22925 , \22235 , \22255 );
nor \U$22611 ( \22926 , \22924 , \22925 );
xnor \U$22612 ( \22927 , \22926 , \22267 );
and \U$22613 ( \22928 , \22251 , \22278 );
and \U$22614 ( \22929 , \22262 , \22276 );
nor \U$22615 ( \22930 , \22928 , \22929 );
xnor \U$22616 ( \22931 , \22930 , \22288 );
xor \U$22617 ( \22932 , \22927 , \22931 );
and \U$22618 ( \22933 , \22272 , \22300 );
and \U$22619 ( \22934 , \22283 , \22298 );
nor \U$22620 ( \22935 , \22933 , \22934 );
xnor \U$22621 ( \22936 , \22935 , \22310 );
xor \U$22622 ( \22937 , \22932 , \22936 );
xor \U$22623 ( \22938 , \22923 , \22937 );
and \U$22624 ( \22939 , \22156 , \22187 );
and \U$22625 ( \22940 , \22167 , \22185 );
nor \U$22626 ( \22941 , \22939 , \22940 );
xnor \U$22627 ( \22942 , \22941 , \22197 );
and \U$22628 ( \22943 , \22181 , \22208 );
and \U$22629 ( \22944 , \22192 , \22206 );
nor \U$22630 ( \22945 , \22943 , \22944 );
xnor \U$22631 ( \22946 , \22945 , \22218 );
xor \U$22632 ( \22947 , \22942 , \22946 );
and \U$22633 ( \22948 , \22202 , \22230 );
and \U$22634 ( \22949 , \22213 , \22228 );
nor \U$22635 ( \22950 , \22948 , \22949 );
xnor \U$22636 ( \22951 , \22950 , \22240 );
xor \U$22637 ( \22952 , \22947 , \22951 );
xor \U$22638 ( \22953 , \22938 , \22952 );
and \U$22639 ( \22954 , \22500 , \22530 );
and \U$22640 ( \22955 , \22511 , \22528 );
nor \U$22641 ( \22956 , \22954 , \22955 );
xnor \U$22642 ( \22957 , \22956 , \22540 );
and \U$22643 ( \22958 , \22524 , \22551 );
and \U$22644 ( \22959 , \22535 , \22549 );
nor \U$22645 ( \22960 , \22958 , \22959 );
xnor \U$22646 ( \22961 , \22960 , \22561 );
xor \U$22647 ( \22962 , \22957 , \22961 );
and \U$22648 ( \22963 , \22545 , \22573 );
and \U$22649 ( \22964 , \22556 , \22571 );
nor \U$22650 ( \22965 , \22963 , \22964 );
xnor \U$22651 ( \22966 , \22965 , \22583 );
xor \U$22652 ( \22967 , \22962 , \22966 );
and \U$22653 ( \22968 , \22429 , \22463 );
and \U$22654 ( \22969 , \22440 , \22461 );
nor \U$22655 ( \22970 , \22968 , \22969 );
xnor \U$22656 ( \22971 , \22970 , \22473 );
and \U$22657 ( \22972 , \22457 , \22484 );
and \U$22658 ( \22973 , \22468 , \22482 );
nor \U$22659 ( \22974 , \22972 , \22973 );
xnor \U$22660 ( \22975 , \22974 , \22494 );
xor \U$22661 ( \22976 , \22971 , \22975 );
and \U$22662 ( \22977 , \22478 , \22506 );
and \U$22663 ( \22978 , \22489 , \22504 );
nor \U$22664 ( \22979 , \22977 , \22978 );
xnor \U$22665 ( \22980 , \22979 , \22516 );
xor \U$22666 ( \22981 , \22976 , \22980 );
xor \U$22667 ( \22982 , \22967 , \22981 );
and \U$22668 ( \22983 , \22361 , \22392 );
and \U$22669 ( \22984 , \22372 , \22390 );
nor \U$22670 ( \22985 , \22983 , \22984 );
xnor \U$22671 ( \22986 , \22985 , \22402 );
and \U$22672 ( \22987 , \22386 , \22413 );
and \U$22673 ( \22988 , \22397 , \22411 );
nor \U$22674 ( \22989 , \22987 , \22988 );
xnor \U$22675 ( \22990 , \22989 , \22423 );
xor \U$22676 ( \22991 , \22986 , \22990 );
and \U$22677 ( \22992 , \22407 , \22435 );
and \U$22678 ( \22993 , \22418 , \22433 );
nor \U$22679 ( \22994 , \22992 , \22993 );
xnor \U$22680 ( \22995 , \22994 , \22445 );
xor \U$22681 ( \22996 , \22991 , \22995 );
xor \U$22682 ( \22997 , \22982 , \22996 );
and \U$22683 ( \22998 , \22953 , \22997 );
xor \U$22684 ( \22999 , \22012 , \22013 );
nand \U$22685 ( \23000 , \22706 , \22999 );
xnor \U$22686 ( \23001 , \23000 , \22016 );
and \U$22687 ( \23002 , \22635 , \22671 );
and \U$22688 ( \23003 , \22646 , \22669 );
nor \U$22689 ( \23004 , \23002 , \23003 );
xnor \U$22690 ( \23005 , \23004 , \22681 );
and \U$22691 ( \23006 , \22665 , \22691 );
and \U$22692 ( \23007 , \22676 , \22689 );
nor \U$22693 ( \23008 , \23006 , \23007 );
xnor \U$22694 ( \23009 , \23008 , \22701 );
xor \U$22695 ( \23010 , \23005 , \23009 );
and \U$22696 ( \23011 , \22686 , \22720 );
and \U$22697 ( \23012 , \22696 , \22707 );
nor \U$22698 ( \23013 , \23011 , \23012 );
xnor \U$22699 ( \23014 , \23013 , \22067 );
xor \U$22700 ( \23015 , \23010 , \23014 );
xor \U$22701 ( \23016 , \23001 , \23015 );
and \U$22702 ( \23017 , \22567 , \22598 );
and \U$22703 ( \23018 , \22578 , \22596 );
nor \U$22704 ( \23019 , \23017 , \23018 );
xnor \U$22705 ( \23020 , \23019 , \22608 );
and \U$22706 ( \23021 , \22592 , \22619 );
and \U$22707 ( \23022 , \22603 , \22617 );
nor \U$22708 ( \23023 , \23021 , \23022 );
xnor \U$22709 ( \23024 , \23023 , \22629 );
xor \U$22710 ( \23025 , \23020 , \23024 );
and \U$22711 ( \23026 , \22613 , \22641 );
and \U$22712 ( \23027 , \22624 , \22639 );
nor \U$22713 ( \23028 , \23026 , \23027 );
xnor \U$22714 ( \23029 , \23028 , \22651 );
xor \U$22715 ( \23030 , \23025 , \23029 );
xor \U$22716 ( \23031 , \23016 , \23030 );
and \U$22717 ( \23032 , \22997 , \23031 );
and \U$22718 ( \23033 , \22953 , \23031 );
or \U$22719 ( \23034 , \22998 , \23032 , \23033 );
and \U$22720 ( \23035 , \22760 , \22764 );
and \U$22721 ( \23036 , \22764 , \22769 );
and \U$22722 ( \23037 , \22760 , \22769 );
or \U$22723 ( \23038 , \23035 , \23036 , \23037 );
and \U$22724 ( \23039 , \22745 , \22749 );
and \U$22725 ( \23040 , \22749 , \22754 );
and \U$22726 ( \23041 , \22745 , \22754 );
or \U$22727 ( \23042 , \23039 , \23040 , \23041 );
xor \U$22728 ( \23043 , \23038 , \23042 );
and \U$22729 ( \23044 , \22731 , \22735 );
and \U$22730 ( \23045 , \22735 , \22740 );
and \U$22731 ( \23046 , \22731 , \22740 );
or \U$22732 ( \23047 , \23044 , \23045 , \23046 );
xor \U$22733 ( \23048 , \23043 , \23047 );
and \U$22734 ( \23049 , \22807 , \22811 );
and \U$22735 ( \23050 , \22811 , \22816 );
and \U$22736 ( \23051 , \22807 , \22816 );
or \U$22737 ( \23052 , \23049 , \23050 , \23051 );
and \U$22738 ( \23053 , \22792 , \22796 );
and \U$22739 ( \23054 , \22796 , \22801 );
and \U$22740 ( \23055 , \22792 , \22801 );
or \U$22741 ( \23056 , \23053 , \23054 , \23055 );
xor \U$22742 ( \23057 , \23052 , \23056 );
and \U$22743 ( \23058 , \22778 , \22782 );
and \U$22744 ( \23059 , \22782 , \22787 );
and \U$22745 ( \23060 , \22778 , \22787 );
or \U$22746 ( \23061 , \23058 , \23059 , \23060 );
xor \U$22747 ( \23062 , \23057 , \23061 );
and \U$22748 ( \23063 , \23048 , \23062 );
and \U$22749 ( \23064 , \22861 , \22865 );
and \U$22750 ( \23065 , \22865 , \22870 );
and \U$22751 ( \23066 , \22861 , \22870 );
or \U$22752 ( \23067 , \23064 , \23065 , \23066 );
and \U$22753 ( \23068 , \22842 , \22846 );
and \U$22754 ( \23069 , \22846 , \22851 );
and \U$22755 ( \23070 , \22842 , \22851 );
or \U$22756 ( \23071 , \23068 , \23069 , \23070 );
xor \U$22757 ( \23072 , \23067 , \23071 );
and \U$22758 ( \23073 , \22828 , \22832 );
and \U$22759 ( \23074 , \22832 , \22837 );
and \U$22760 ( \23075 , \22828 , \22837 );
or \U$22761 ( \23076 , \23073 , \23074 , \23075 );
xor \U$22762 ( \23077 , \23072 , \23076 );
and \U$22763 ( \23078 , \23062 , \23077 );
and \U$22764 ( \23079 , \23048 , \23077 );
or \U$22765 ( \23080 , \23063 , \23078 , \23079 );
and \U$22766 ( \23081 , \23034 , \23080 );
and \U$22767 ( \23082 , \22927 , \22931 );
and \U$22768 ( \23083 , \22931 , \22936 );
and \U$22769 ( \23084 , \22927 , \22936 );
or \U$22770 ( \23085 , \23082 , \23083 , \23084 );
and \U$22771 ( \23086 , \22913 , \22917 );
and \U$22772 ( \23087 , \22917 , \22922 );
and \U$22773 ( \23088 , \22913 , \22922 );
or \U$22774 ( \23089 , \23086 , \23087 , \23088 );
xor \U$22775 ( \23090 , \23085 , \23089 );
and \U$22776 ( \23091 , \22986 , \22990 );
and \U$22777 ( \23092 , \22990 , \22995 );
and \U$22778 ( \23093 , \22986 , \22995 );
or \U$22779 ( \23094 , \23091 , \23092 , \23093 );
xor \U$22780 ( \23095 , \23090 , \23094 );
and \U$22781 ( \23096 , \23080 , \23095 );
and \U$22782 ( \23097 , \23034 , \23095 );
or \U$22783 ( \23098 , \23081 , \23096 , \23097 );
and \U$22784 ( \23099 , \22909 , \23098 );
and \U$22785 ( \23100 , \22016 , \22897 );
and \U$22786 ( \23101 , \22897 , \22902 );
and \U$22787 ( \23102 , \22016 , \22902 );
or \U$22788 ( \23103 , \23100 , \23101 , \23102 );
and \U$22789 ( \23104 , \22878 , \22882 );
and \U$22790 ( \23105 , \22882 , \22887 );
and \U$22791 ( \23106 , \22878 , \22887 );
or \U$22792 ( \23107 , \23104 , \23105 , \23106 );
xor \U$22793 ( \23108 , \23103 , \23107 );
and \U$22794 ( \23109 , \22942 , \22946 );
and \U$22795 ( \23110 , \22946 , \22951 );
and \U$22796 ( \23111 , \22942 , \22951 );
or \U$22797 ( \23112 , \23109 , \23110 , \23111 );
xor \U$22798 ( \23113 , \23108 , \23112 );
and \U$22799 ( \23114 , \22535 , \22551 );
and \U$22800 ( \23115 , \22500 , \22549 );
nor \U$22801 ( \23116 , \23114 , \23115 );
xnor \U$22802 ( \23117 , \23116 , \22561 );
and \U$22803 ( \23118 , \22556 , \22573 );
and \U$22804 ( \23119 , \22524 , \22571 );
nor \U$22805 ( \23120 , \23118 , \23119 );
xnor \U$22806 ( \23121 , \23120 , \22583 );
xor \U$22807 ( \23122 , \23117 , \23121 );
and \U$22808 ( \23123 , \22578 , \22598 );
and \U$22809 ( \23124 , \22545 , \22596 );
nor \U$22810 ( \23125 , \23123 , \23124 );
xnor \U$22811 ( \23126 , \23125 , \22608 );
xor \U$22812 ( \23127 , \23122 , \23126 );
and \U$22813 ( \23128 , \22468 , \22484 );
and \U$22814 ( \23129 , \22429 , \22482 );
nor \U$22815 ( \23130 , \23128 , \23129 );
xnor \U$22816 ( \23131 , \23130 , \22494 );
and \U$22817 ( \23132 , \22489 , \22506 );
and \U$22818 ( \23133 , \22457 , \22504 );
nor \U$22819 ( \23134 , \23132 , \23133 );
xnor \U$22820 ( \23135 , \23134 , \22516 );
xor \U$22821 ( \23136 , \23131 , \23135 );
and \U$22822 ( \23137 , \22511 , \22530 );
and \U$22823 ( \23138 , \22478 , \22528 );
nor \U$22824 ( \23139 , \23137 , \23138 );
xnor \U$22825 ( \23140 , \23139 , \22540 );
xor \U$22826 ( \23141 , \23136 , \23140 );
xor \U$22827 ( \23142 , \23127 , \23141 );
and \U$22828 ( \23143 , \22397 , \22413 );
and \U$22829 ( \23144 , \22361 , \22411 );
nor \U$22830 ( \23145 , \23143 , \23144 );
xnor \U$22831 ( \23146 , \23145 , \22423 );
and \U$22832 ( \23147 , \22418 , \22435 );
and \U$22833 ( \23148 , \22386 , \22433 );
nor \U$22834 ( \23149 , \23147 , \23148 );
xnor \U$22835 ( \23150 , \23149 , \22445 );
xor \U$22836 ( \23151 , \23146 , \23150 );
and \U$22837 ( \23152 , \22440 , \22463 );
and \U$22838 ( \23153 , \22407 , \22461 );
nor \U$22839 ( \23154 , \23152 , \23153 );
xnor \U$22840 ( \23155 , \23154 , \22473 );
xor \U$22841 ( \23156 , \23151 , \23155 );
xor \U$22842 ( \23157 , \23142 , \23156 );
and \U$22843 ( \23158 , \23005 , \23009 );
and \U$22844 ( \23159 , \23009 , \23014 );
and \U$22845 ( \23160 , \23005 , \23014 );
or \U$22846 ( \23161 , \23158 , \23159 , \23160 );
and \U$22847 ( \23162 , \22676 , \22691 );
and \U$22848 ( \23163 , \22635 , \22689 );
nor \U$22849 ( \23164 , \23162 , \23163 );
xnor \U$22850 ( \23165 , \23164 , \22701 );
and \U$22851 ( \23166 , \22696 , \22720 );
and \U$22852 ( \23167 , \22665 , \22707 );
nor \U$22853 ( \23168 , \23166 , \23167 );
xnor \U$22854 ( \23169 , \23168 , \22067 );
xor \U$22855 ( \23170 , \23165 , \23169 );
xor \U$22856 ( \23171 , \21592 , \22012 );
not \U$22857 ( \23172 , \22999 );
and \U$22858 ( \23173 , \23171 , \23172 );
and \U$22859 ( \23174 , \22706 , \23173 );
and \U$22860 ( \23175 , \22686 , \22999 );
nor \U$22861 ( \23176 , \23174 , \23175 );
xnor \U$22862 ( \23177 , \23176 , \22016 );
xor \U$22863 ( \23178 , \23170 , \23177 );
xor \U$22864 ( \23179 , \23161 , \23178 );
and \U$22865 ( \23180 , \22603 , \22619 );
and \U$22866 ( \23181 , \22567 , \22617 );
nor \U$22867 ( \23182 , \23180 , \23181 );
xnor \U$22868 ( \23183 , \23182 , \22629 );
and \U$22869 ( \23184 , \22624 , \22641 );
and \U$22870 ( \23185 , \22592 , \22639 );
nor \U$22871 ( \23186 , \23184 , \23185 );
xnor \U$22872 ( \23187 , \23186 , \22651 );
xor \U$22873 ( \23188 , \23183 , \23187 );
and \U$22874 ( \23189 , \22646 , \22671 );
and \U$22875 ( \23190 , \22613 , \22669 );
nor \U$22876 ( \23191 , \23189 , \23190 );
xnor \U$22877 ( \23192 , \23191 , \22681 );
xor \U$22878 ( \23193 , \23188 , \23192 );
xor \U$22879 ( \23194 , \23179 , \23193 );
xor \U$22880 ( \23195 , \23157 , \23194 );
and \U$22881 ( \23196 , \22971 , \22975 );
and \U$22882 ( \23197 , \22975 , \22980 );
and \U$22883 ( \23198 , \22971 , \22980 );
or \U$22884 ( \23199 , \23196 , \23197 , \23198 );
and \U$22885 ( \23200 , \22957 , \22961 );
and \U$22886 ( \23201 , \22961 , \22966 );
and \U$22887 ( \23202 , \22957 , \22966 );
or \U$22888 ( \23203 , \23200 , \23201 , \23202 );
xor \U$22889 ( \23204 , \23199 , \23203 );
and \U$22890 ( \23205 , \23020 , \23024 );
and \U$22891 ( \23206 , \23024 , \23029 );
and \U$22892 ( \23207 , \23020 , \23029 );
or \U$22893 ( \23208 , \23205 , \23206 , \23207 );
xor \U$22894 ( \23209 , \23204 , \23208 );
xor \U$22895 ( \23210 , \23195 , \23209 );
and \U$22896 ( \23211 , \23113 , \23210 );
and \U$22897 ( \23212 , \22124 , \22140 );
and \U$22898 ( \23213 , \22089 , \22138 );
nor \U$22899 ( \23214 , \23212 , \23213 );
xnor \U$22900 ( \23215 , \23214 , \22150 );
and \U$22901 ( \23216 , \22145 , \22162 );
and \U$22902 ( \23217 , \22113 , \22160 );
nor \U$22903 ( \23218 , \23216 , \23217 );
xnor \U$22904 ( \23219 , \23218 , \22172 );
xor \U$22905 ( \23220 , \23215 , \23219 );
and \U$22906 ( \23221 , \22167 , \22187 );
and \U$22907 ( \23222 , \22134 , \22185 );
nor \U$22908 ( \23223 , \23221 , \23222 );
xnor \U$22909 ( \23224 , \23223 , \22197 );
xor \U$22910 ( \23225 , \23220 , \23224 );
and \U$22911 ( \23226 , \22894 , \22076 );
xor \U$22912 ( \23227 , \21609 , \21610 );
xor \U$22913 ( \23228 , \23227 , \21962 );
buf \U$22914 ( \23229 , \23228 );
buf \U$22915 ( \23230 , \23229 );
and \U$22916 ( \23231 , \23230 , \22073 );
nor \U$22917 ( \23232 , \23226 , \23231 );
xnor \U$22918 ( \23233 , \23232 , \22072 );
and \U$22919 ( \23234 , \22081 , \22095 );
and \U$22920 ( \23235 , \22858 , \22093 );
nor \U$22921 ( \23236 , \23234 , \23235 );
xnor \U$22922 ( \23237 , \23236 , \22105 );
xor \U$22923 ( \23238 , \23233 , \23237 );
and \U$22924 ( \23239 , \22100 , \22119 );
and \U$22925 ( \23240 , \22071 , \22117 );
nor \U$22926 ( \23241 , \23239 , \23240 );
xnor \U$22927 ( \23242 , \23241 , \22129 );
xor \U$22928 ( \23243 , \23238 , \23242 );
xor \U$22929 ( \23244 , \23225 , \23243 );
and \U$22930 ( \23245 , \22329 , \22345 );
and \U$22931 ( \23246 , \22294 , \22343 );
nor \U$22932 ( \23247 , \23245 , \23246 );
xnor \U$22933 ( \23248 , \23247 , \22355 );
and \U$22934 ( \23249 , \22350 , \22367 );
and \U$22935 ( \23250 , \22318 , \22365 );
nor \U$22936 ( \23251 , \23249 , \23250 );
xnor \U$22937 ( \23252 , \23251 , \22377 );
xor \U$22938 ( \23253 , \23248 , \23252 );
and \U$22939 ( \23254 , \22372 , \22392 );
and \U$22940 ( \23255 , \22339 , \22390 );
nor \U$22941 ( \23256 , \23254 , \23255 );
xnor \U$22942 ( \23257 , \23256 , \22402 );
xor \U$22943 ( \23258 , \23253 , \23257 );
and \U$22944 ( \23259 , \22262 , \22278 );
and \U$22945 ( \23260 , \22224 , \22276 );
nor \U$22946 ( \23261 , \23259 , \23260 );
xnor \U$22947 ( \23262 , \23261 , \22288 );
and \U$22948 ( \23263 , \22283 , \22300 );
and \U$22949 ( \23264 , \22251 , \22298 );
nor \U$22950 ( \23265 , \23263 , \23264 );
xnor \U$22951 ( \23266 , \23265 , \22310 );
xor \U$22952 ( \23267 , \23262 , \23266 );
and \U$22953 ( \23268 , \22305 , \22324 );
and \U$22954 ( \23269 , \22272 , \22322 );
nor \U$22955 ( \23270 , \23268 , \23269 );
xnor \U$22956 ( \23271 , \23270 , \22334 );
xor \U$22957 ( \23272 , \23267 , \23271 );
xor \U$22958 ( \23273 , \23258 , \23272 );
and \U$22959 ( \23274 , \22192 , \22208 );
and \U$22960 ( \23275 , \22156 , \22206 );
nor \U$22961 ( \23276 , \23274 , \23275 );
xnor \U$22962 ( \23277 , \23276 , \22218 );
and \U$22963 ( \23278 , \22213 , \22230 );
and \U$22964 ( \23279 , \22181 , \22228 );
nor \U$22965 ( \23280 , \23278 , \23279 );
xnor \U$22966 ( \23281 , \23280 , \22240 );
xor \U$22967 ( \23282 , \23277 , \23281 );
and \U$22968 ( \23283 , \22235 , \22257 );
and \U$22969 ( \23284 , \22202 , \22255 );
nor \U$22970 ( \23285 , \23283 , \23284 );
xnor \U$22971 ( \23286 , \23285 , \22267 );
xor \U$22972 ( \23287 , \23282 , \23286 );
xor \U$22973 ( \23288 , \23273 , \23287 );
xor \U$22974 ( \23289 , \23244 , \23288 );
and \U$22975 ( \23290 , \23210 , \23289 );
and \U$22976 ( \23291 , \23113 , \23289 );
or \U$22977 ( \23292 , \23211 , \23290 , \23291 );
and \U$22978 ( \23293 , \23098 , \23292 );
and \U$22979 ( \23294 , \22909 , \23292 );
or \U$22980 ( \23295 , \23099 , \23293 , \23294 );
and \U$22981 ( \23296 , \22134 , \22187 );
and \U$22982 ( \23297 , \22145 , \22185 );
nor \U$22983 ( \23298 , \23296 , \23297 );
xnor \U$22984 ( \23299 , \23298 , \22197 );
and \U$22985 ( \23300 , \22156 , \22208 );
and \U$22986 ( \23301 , \22167 , \22206 );
nor \U$22987 ( \23302 , \23300 , \23301 );
xnor \U$22988 ( \23303 , \23302 , \22218 );
xor \U$22989 ( \23304 , \23299 , \23303 );
and \U$22990 ( \23305 , \22181 , \22230 );
and \U$22991 ( \23306 , \22192 , \22228 );
nor \U$22992 ( \23307 , \23305 , \23306 );
xnor \U$22993 ( \23308 , \23307 , \22240 );
xor \U$22994 ( \23309 , \23304 , \23308 );
and \U$22995 ( \23310 , \22071 , \22119 );
and \U$22996 ( \23311 , \22081 , \22117 );
nor \U$22997 ( \23312 , \23310 , \23311 );
xnor \U$22998 ( \23313 , \23312 , \22129 );
and \U$22999 ( \23314 , \22089 , \22140 );
and \U$23000 ( \23315 , \22100 , \22138 );
nor \U$23001 ( \23316 , \23314 , \23315 );
xnor \U$23002 ( \23317 , \23316 , \22150 );
xor \U$23003 ( \23318 , \23313 , \23317 );
and \U$23004 ( \23319 , \22113 , \22162 );
and \U$23005 ( \23320 , \22124 , \22160 );
nor \U$23006 ( \23321 , \23319 , \23320 );
xnor \U$23007 ( \23322 , \23321 , \22172 );
xor \U$23008 ( \23323 , \23318 , \23322 );
xor \U$23009 ( \23324 , \23309 , \23323 );
and \U$23010 ( \23325 , \23230 , \22076 );
xor \U$23011 ( \23326 , \21606 , \21607 );
xor \U$23012 ( \23327 , \23326 , \21965 );
buf \U$23013 ( \23328 , \23327 );
buf \U$23014 ( \23329 , \23328 );
and \U$23015 ( \23330 , \23329 , \22073 );
nor \U$23016 ( \23331 , \23325 , \23330 );
xnor \U$23017 ( \23332 , \23331 , \22072 );
xor \U$23018 ( \23333 , \21595 , \23332 );
and \U$23019 ( \23334 , \22858 , \22095 );
and \U$23020 ( \23335 , \22894 , \22093 );
nor \U$23021 ( \23336 , \23334 , \23335 );
xnor \U$23022 ( \23337 , \23336 , \22105 );
xor \U$23023 ( \23338 , \23333 , \23337 );
xor \U$23024 ( \23339 , \23324 , \23338 );
and \U$23025 ( \23340 , \22339 , \22392 );
and \U$23026 ( \23341 , \22350 , \22390 );
nor \U$23027 ( \23342 , \23340 , \23341 );
xnor \U$23028 ( \23343 , \23342 , \22402 );
and \U$23029 ( \23344 , \22361 , \22413 );
and \U$23030 ( \23345 , \22372 , \22411 );
nor \U$23031 ( \23346 , \23344 , \23345 );
xnor \U$23032 ( \23347 , \23346 , \22423 );
xor \U$23033 ( \23348 , \23343 , \23347 );
and \U$23034 ( \23349 , \22386 , \22435 );
and \U$23035 ( \23350 , \22397 , \22433 );
nor \U$23036 ( \23351 , \23349 , \23350 );
xnor \U$23037 ( \23352 , \23351 , \22445 );
xor \U$23038 ( \23353 , \23348 , \23352 );
and \U$23039 ( \23354 , \22272 , \22324 );
and \U$23040 ( \23355 , \22283 , \22322 );
nor \U$23041 ( \23356 , \23354 , \23355 );
xnor \U$23042 ( \23357 , \23356 , \22334 );
and \U$23043 ( \23358 , \22294 , \22345 );
and \U$23044 ( \23359 , \22305 , \22343 );
nor \U$23045 ( \23360 , \23358 , \23359 );
xnor \U$23046 ( \23361 , \23360 , \22355 );
xor \U$23047 ( \23362 , \23357 , \23361 );
and \U$23048 ( \23363 , \22318 , \22367 );
and \U$23049 ( \23364 , \22329 , \22365 );
nor \U$23050 ( \23365 , \23363 , \23364 );
xnor \U$23051 ( \23366 , \23365 , \22377 );
xor \U$23052 ( \23367 , \23362 , \23366 );
xor \U$23053 ( \23368 , \23353 , \23367 );
and \U$23054 ( \23369 , \22202 , \22257 );
and \U$23055 ( \23370 , \22213 , \22255 );
nor \U$23056 ( \23371 , \23369 , \23370 );
xnor \U$23057 ( \23372 , \23371 , \22267 );
and \U$23058 ( \23373 , \22224 , \22278 );
and \U$23059 ( \23374 , \22235 , \22276 );
nor \U$23060 ( \23375 , \23373 , \23374 );
xnor \U$23061 ( \23376 , \23375 , \22288 );
xor \U$23062 ( \23377 , \23372 , \23376 );
and \U$23063 ( \23378 , \22251 , \22300 );
and \U$23064 ( \23379 , \22262 , \22298 );
nor \U$23065 ( \23380 , \23378 , \23379 );
xnor \U$23066 ( \23381 , \23380 , \22310 );
xor \U$23067 ( \23382 , \23377 , \23381 );
xor \U$23068 ( \23383 , \23368 , \23382 );
xor \U$23069 ( \23384 , \23339 , \23383 );
and \U$23070 ( \23385 , \22545 , \22598 );
and \U$23071 ( \23386 , \22556 , \22596 );
nor \U$23072 ( \23387 , \23385 , \23386 );
xnor \U$23073 ( \23388 , \23387 , \22608 );
and \U$23074 ( \23389 , \22567 , \22619 );
and \U$23075 ( \23390 , \22578 , \22617 );
nor \U$23076 ( \23391 , \23389 , \23390 );
xnor \U$23077 ( \23392 , \23391 , \22629 );
xor \U$23078 ( \23393 , \23388 , \23392 );
and \U$23079 ( \23394 , \22592 , \22641 );
and \U$23080 ( \23395 , \22603 , \22639 );
nor \U$23081 ( \23396 , \23394 , \23395 );
xnor \U$23082 ( \23397 , \23396 , \22651 );
xor \U$23083 ( \23398 , \23393 , \23397 );
and \U$23084 ( \23399 , \22478 , \22530 );
and \U$23085 ( \23400 , \22489 , \22528 );
nor \U$23086 ( \23401 , \23399 , \23400 );
xnor \U$23087 ( \23402 , \23401 , \22540 );
and \U$23088 ( \23403 , \22500 , \22551 );
and \U$23089 ( \23404 , \22511 , \22549 );
nor \U$23090 ( \23405 , \23403 , \23404 );
xnor \U$23091 ( \23406 , \23405 , \22561 );
xor \U$23092 ( \23407 , \23402 , \23406 );
and \U$23093 ( \23408 , \22524 , \22573 );
and \U$23094 ( \23409 , \22535 , \22571 );
nor \U$23095 ( \23410 , \23408 , \23409 );
xnor \U$23096 ( \23411 , \23410 , \22583 );
xor \U$23097 ( \23412 , \23407 , \23411 );
xor \U$23098 ( \23413 , \23398 , \23412 );
and \U$23099 ( \23414 , \22407 , \22463 );
and \U$23100 ( \23415 , \22418 , \22461 );
nor \U$23101 ( \23416 , \23414 , \23415 );
xnor \U$23102 ( \23417 , \23416 , \22473 );
and \U$23103 ( \23418 , \22429 , \22484 );
and \U$23104 ( \23419 , \22440 , \22482 );
nor \U$23105 ( \23420 , \23418 , \23419 );
xnor \U$23106 ( \23421 , \23420 , \22494 );
xor \U$23107 ( \23422 , \23417 , \23421 );
and \U$23108 ( \23423 , \22457 , \22506 );
and \U$23109 ( \23424 , \22468 , \22504 );
nor \U$23110 ( \23425 , \23423 , \23424 );
xnor \U$23111 ( \23426 , \23425 , \22516 );
xor \U$23112 ( \23427 , \23422 , \23426 );
xor \U$23113 ( \23428 , \23413 , \23427 );
xor \U$23114 ( \23429 , \23384 , \23428 );
and \U$23115 ( \23430 , \23161 , \23178 );
and \U$23116 ( \23431 , \23178 , \23193 );
and \U$23117 ( \23432 , \23161 , \23193 );
or \U$23118 ( \23433 , \23430 , \23431 , \23432 );
and \U$23119 ( \23434 , \23127 , \23141 );
and \U$23120 ( \23435 , \23141 , \23156 );
and \U$23121 ( \23436 , \23127 , \23156 );
or \U$23122 ( \23437 , \23434 , \23435 , \23436 );
xor \U$23123 ( \23438 , \23433 , \23437 );
and \U$23124 ( \23439 , \23258 , \23272 );
and \U$23125 ( \23440 , \23272 , \23287 );
and \U$23126 ( \23441 , \23258 , \23287 );
or \U$23127 ( \23442 , \23439 , \23440 , \23441 );
xor \U$23128 ( \23443 , \23438 , \23442 );
xor \U$23129 ( \23444 , \23429 , \23443 );
and \U$23130 ( \23445 , \23103 , \23107 );
and \U$23131 ( \23446 , \23107 , \23112 );
and \U$23132 ( \23447 , \23103 , \23112 );
or \U$23133 ( \23448 , \23445 , \23446 , \23447 );
and \U$23134 ( \23449 , \23085 , \23089 );
and \U$23135 ( \23450 , \23089 , \23094 );
and \U$23136 ( \23451 , \23085 , \23094 );
or \U$23137 ( \23452 , \23449 , \23450 , \23451 );
xor \U$23138 ( \23453 , \23448 , \23452 );
and \U$23139 ( \23454 , \23199 , \23203 );
and \U$23140 ( \23455 , \23203 , \23208 );
and \U$23141 ( \23456 , \23199 , \23208 );
or \U$23142 ( \23457 , \23454 , \23455 , \23456 );
xor \U$23143 ( \23458 , \23453 , \23457 );
xor \U$23144 ( \23459 , \23444 , \23458 );
and \U$23145 ( \23460 , \23157 , \23194 );
and \U$23146 ( \23461 , \23194 , \23209 );
and \U$23147 ( \23462 , \23157 , \23209 );
or \U$23148 ( \23463 , \23460 , \23461 , \23462 );
and \U$23149 ( \23464 , \23233 , \23237 );
and \U$23150 ( \23465 , \23237 , \23242 );
and \U$23151 ( \23466 , \23233 , \23242 );
or \U$23152 ( \23467 , \23464 , \23465 , \23466 );
and \U$23153 ( \23468 , \23215 , \23219 );
and \U$23154 ( \23469 , \23219 , \23224 );
and \U$23155 ( \23470 , \23215 , \23224 );
or \U$23156 ( \23471 , \23468 , \23469 , \23470 );
xor \U$23157 ( \23472 , \23467 , \23471 );
and \U$23158 ( \23473 , \23277 , \23281 );
and \U$23159 ( \23474 , \23281 , \23286 );
and \U$23160 ( \23475 , \23277 , \23286 );
or \U$23161 ( \23476 , \23473 , \23474 , \23475 );
xor \U$23162 ( \23477 , \23472 , \23476 );
xor \U$23163 ( \23478 , \23463 , \23477 );
and \U$23164 ( \23479 , \23165 , \23169 );
and \U$23165 ( \23480 , \23169 , \23177 );
and \U$23166 ( \23481 , \23165 , \23177 );
or \U$23167 ( \23482 , \23479 , \23480 , \23481 );
and \U$23168 ( \23483 , \22686 , \23173 );
and \U$23169 ( \23484 , \22696 , \22999 );
nor \U$23170 ( \23485 , \23483 , \23484 );
xnor \U$23171 ( \23486 , \23485 , \22016 );
nand \U$23172 ( \23487 , \22706 , \22019 );
xnor \U$23173 ( \23488 , \23487 , \21595 );
xor \U$23174 ( \23489 , \23486 , \23488 );
xor \U$23175 ( \23490 , \23482 , \23489 );
and \U$23176 ( \23491 , \22613 , \22671 );
and \U$23177 ( \23492 , \22624 , \22669 );
nor \U$23178 ( \23493 , \23491 , \23492 );
xnor \U$23179 ( \23494 , \23493 , \22681 );
and \U$23180 ( \23495 , \22635 , \22691 );
and \U$23181 ( \23496 , \22646 , \22689 );
nor \U$23182 ( \23497 , \23495 , \23496 );
xnor \U$23183 ( \23498 , \23497 , \22701 );
xor \U$23184 ( \23499 , \23494 , \23498 );
and \U$23185 ( \23500 , \22665 , \22720 );
and \U$23186 ( \23501 , \22676 , \22707 );
nor \U$23187 ( \23502 , \23500 , \23501 );
xnor \U$23188 ( \23503 , \23502 , \22067 );
xor \U$23189 ( \23504 , \23499 , \23503 );
xor \U$23190 ( \23505 , \23490 , \23504 );
and \U$23191 ( \23506 , \23131 , \23135 );
and \U$23192 ( \23507 , \23135 , \23140 );
and \U$23193 ( \23508 , \23131 , \23140 );
or \U$23194 ( \23509 , \23506 , \23507 , \23508 );
and \U$23195 ( \23510 , \23117 , \23121 );
and \U$23196 ( \23511 , \23121 , \23126 );
and \U$23197 ( \23512 , \23117 , \23126 );
or \U$23198 ( \23513 , \23510 , \23511 , \23512 );
xor \U$23199 ( \23514 , \23509 , \23513 );
and \U$23200 ( \23515 , \23183 , \23187 );
and \U$23201 ( \23516 , \23187 , \23192 );
and \U$23202 ( \23517 , \23183 , \23192 );
or \U$23203 ( \23518 , \23515 , \23516 , \23517 );
xor \U$23204 ( \23519 , \23514 , \23518 );
xor \U$23205 ( \23520 , \23505 , \23519 );
and \U$23206 ( \23521 , \23262 , \23266 );
and \U$23207 ( \23522 , \23266 , \23271 );
and \U$23208 ( \23523 , \23262 , \23271 );
or \U$23209 ( \23524 , \23521 , \23522 , \23523 );
and \U$23210 ( \23525 , \23248 , \23252 );
and \U$23211 ( \23526 , \23252 , \23257 );
and \U$23212 ( \23527 , \23248 , \23257 );
or \U$23213 ( \23528 , \23525 , \23526 , \23527 );
xor \U$23214 ( \23529 , \23524 , \23528 );
and \U$23215 ( \23530 , \23146 , \23150 );
and \U$23216 ( \23531 , \23150 , \23155 );
and \U$23217 ( \23532 , \23146 , \23155 );
or \U$23218 ( \23533 , \23530 , \23531 , \23532 );
xor \U$23219 ( \23534 , \23529 , \23533 );
xor \U$23220 ( \23535 , \23520 , \23534 );
xor \U$23221 ( \23536 , \23478 , \23535 );
and \U$23222 ( \23537 , \23459 , \23536 );
and \U$23223 ( \23538 , \23067 , \23071 );
and \U$23224 ( \23539 , \23071 , \23076 );
and \U$23225 ( \23540 , \23067 , \23076 );
or \U$23226 ( \23541 , \23538 , \23539 , \23540 );
and \U$23227 ( \23542 , \23052 , \23056 );
and \U$23228 ( \23543 , \23056 , \23061 );
and \U$23229 ( \23544 , \23052 , \23061 );
or \U$23230 ( \23545 , \23542 , \23543 , \23544 );
and \U$23231 ( \23546 , \23541 , \23545 );
and \U$23232 ( \23547 , \23038 , \23042 );
and \U$23233 ( \23548 , \23042 , \23047 );
and \U$23234 ( \23549 , \23038 , \23047 );
or \U$23235 ( \23550 , \23547 , \23548 , \23549 );
and \U$23236 ( \23551 , \23545 , \23550 );
and \U$23237 ( \23552 , \23541 , \23550 );
or \U$23238 ( \23553 , \23546 , \23551 , \23552 );
and \U$23239 ( \23554 , \23001 , \23015 );
and \U$23240 ( \23555 , \23015 , \23030 );
and \U$23241 ( \23556 , \23001 , \23030 );
or \U$23242 ( \23557 , \23554 , \23555 , \23556 );
and \U$23243 ( \23558 , \22967 , \22981 );
and \U$23244 ( \23559 , \22981 , \22996 );
and \U$23245 ( \23560 , \22967 , \22996 );
or \U$23246 ( \23561 , \23558 , \23559 , \23560 );
and \U$23247 ( \23562 , \23557 , \23561 );
and \U$23248 ( \23563 , \22923 , \22937 );
and \U$23249 ( \23564 , \22937 , \22952 );
and \U$23250 ( \23565 , \22923 , \22952 );
or \U$23251 ( \23566 , \23563 , \23564 , \23565 );
and \U$23252 ( \23567 , \23561 , \23566 );
and \U$23253 ( \23568 , \23557 , \23566 );
or \U$23254 ( \23569 , \23562 , \23567 , \23568 );
xor \U$23255 ( \23570 , \23553 , \23569 );
and \U$23256 ( \23571 , \23225 , \23243 );
and \U$23257 ( \23572 , \23243 , \23288 );
and \U$23258 ( \23573 , \23225 , \23288 );
or \U$23259 ( \23574 , \23571 , \23572 , \23573 );
xor \U$23260 ( \23575 , \23570 , \23574 );
and \U$23261 ( \23576 , \23536 , \23575 );
and \U$23262 ( \23577 , \23459 , \23575 );
or \U$23263 ( \23578 , \23537 , \23576 , \23577 );
and \U$23264 ( \23579 , \23295 , \23578 );
and \U$23265 ( \23580 , \23309 , \23323 );
and \U$23266 ( \23581 , \23323 , \23338 );
and \U$23267 ( \23582 , \23309 , \23338 );
or \U$23268 ( \23583 , \23580 , \23581 , \23582 );
and \U$23269 ( \23584 , \23329 , \22076 );
and \U$23270 ( \23585 , \22030 , \22073 );
nor \U$23271 ( \23586 , \23584 , \23585 );
xnor \U$23272 ( \23587 , \23586 , \22072 );
and \U$23273 ( \23588 , \22894 , \22095 );
and \U$23274 ( \23589 , \23230 , \22093 );
nor \U$23275 ( \23590 , \23588 , \23589 );
xnor \U$23276 ( \23591 , \23590 , \22105 );
xor \U$23277 ( \23592 , \23587 , \23591 );
and \U$23278 ( \23593 , \22081 , \22119 );
and \U$23279 ( \23594 , \22858 , \22117 );
nor \U$23280 ( \23595 , \23593 , \23594 );
xnor \U$23281 ( \23596 , \23595 , \22129 );
xor \U$23282 ( \23597 , \23592 , \23596 );
xor \U$23283 ( \23598 , \23583 , \23597 );
and \U$23284 ( \23599 , \22235 , \22278 );
and \U$23285 ( \23600 , \22202 , \22276 );
nor \U$23286 ( \23601 , \23599 , \23600 );
xnor \U$23287 ( \23602 , \23601 , \22288 );
and \U$23288 ( \23603 , \22262 , \22300 );
and \U$23289 ( \23604 , \22224 , \22298 );
nor \U$23290 ( \23605 , \23603 , \23604 );
xnor \U$23291 ( \23606 , \23605 , \22310 );
xor \U$23292 ( \23607 , \23602 , \23606 );
and \U$23293 ( \23608 , \22283 , \22324 );
and \U$23294 ( \23609 , \22251 , \22322 );
nor \U$23295 ( \23610 , \23608 , \23609 );
xnor \U$23296 ( \23611 , \23610 , \22334 );
xor \U$23297 ( \23612 , \23607 , \23611 );
and \U$23298 ( \23613 , \22167 , \22208 );
and \U$23299 ( \23614 , \22134 , \22206 );
nor \U$23300 ( \23615 , \23613 , \23614 );
xnor \U$23301 ( \23616 , \23615 , \22218 );
and \U$23302 ( \23617 , \22192 , \22230 );
and \U$23303 ( \23618 , \22156 , \22228 );
nor \U$23304 ( \23619 , \23617 , \23618 );
xnor \U$23305 ( \23620 , \23619 , \22240 );
xor \U$23306 ( \23621 , \23616 , \23620 );
and \U$23307 ( \23622 , \22213 , \22257 );
and \U$23308 ( \23623 , \22181 , \22255 );
nor \U$23309 ( \23624 , \23622 , \23623 );
xnor \U$23310 ( \23625 , \23624 , \22267 );
xor \U$23311 ( \23626 , \23621 , \23625 );
xor \U$23312 ( \23627 , \23612 , \23626 );
and \U$23313 ( \23628 , \22100 , \22140 );
and \U$23314 ( \23629 , \22071 , \22138 );
nor \U$23315 ( \23630 , \23628 , \23629 );
xnor \U$23316 ( \23631 , \23630 , \22150 );
and \U$23317 ( \23632 , \22124 , \22162 );
and \U$23318 ( \23633 , \22089 , \22160 );
nor \U$23319 ( \23634 , \23632 , \23633 );
xnor \U$23320 ( \23635 , \23634 , \22172 );
xor \U$23321 ( \23636 , \23631 , \23635 );
and \U$23322 ( \23637 , \22145 , \22187 );
and \U$23323 ( \23638 , \22113 , \22185 );
nor \U$23324 ( \23639 , \23637 , \23638 );
xnor \U$23325 ( \23640 , \23639 , \22197 );
xor \U$23326 ( \23641 , \23636 , \23640 );
xor \U$23327 ( \23642 , \23627 , \23641 );
xor \U$23328 ( \23643 , \23598 , \23642 );
and \U$23329 ( \23644 , \23482 , \23489 );
and \U$23330 ( \23645 , \23489 , \23504 );
and \U$23331 ( \23646 , \23482 , \23504 );
or \U$23332 ( \23647 , \23644 , \23645 , \23646 );
and \U$23333 ( \23648 , \23398 , \23412 );
and \U$23334 ( \23649 , \23412 , \23427 );
and \U$23335 ( \23650 , \23398 , \23427 );
or \U$23336 ( \23651 , \23648 , \23649 , \23650 );
xor \U$23337 ( \23652 , \23647 , \23651 );
and \U$23338 ( \23653 , \23353 , \23367 );
and \U$23339 ( \23654 , \23367 , \23382 );
and \U$23340 ( \23655 , \23353 , \23382 );
or \U$23341 ( \23656 , \23653 , \23654 , \23655 );
xor \U$23342 ( \23657 , \23652 , \23656 );
xor \U$23343 ( \23658 , \23643 , \23657 );
and \U$23344 ( \23659 , \23467 , \23471 );
and \U$23345 ( \23660 , \23471 , \23476 );
and \U$23346 ( \23661 , \23467 , \23476 );
or \U$23347 ( \23662 , \23659 , \23660 , \23661 );
and \U$23348 ( \23663 , \23524 , \23528 );
and \U$23349 ( \23664 , \23528 , \23533 );
and \U$23350 ( \23665 , \23524 , \23533 );
or \U$23351 ( \23666 , \23663 , \23664 , \23665 );
xor \U$23352 ( \23667 , \23662 , \23666 );
and \U$23353 ( \23668 , \23509 , \23513 );
and \U$23354 ( \23669 , \23513 , \23518 );
and \U$23355 ( \23670 , \23509 , \23518 );
or \U$23356 ( \23671 , \23668 , \23669 , \23670 );
xor \U$23357 ( \23672 , \23667 , \23671 );
xor \U$23358 ( \23673 , \23658 , \23672 );
and \U$23359 ( \23674 , \23505 , \23519 );
and \U$23360 ( \23675 , \23519 , \23534 );
and \U$23361 ( \23676 , \23505 , \23534 );
or \U$23362 ( \23677 , \23674 , \23675 , \23676 );
and \U$23363 ( \23678 , \23417 , \23421 );
and \U$23364 ( \23679 , \23421 , \23426 );
and \U$23365 ( \23680 , \23417 , \23426 );
or \U$23366 ( \23681 , \23678 , \23679 , \23680 );
and \U$23367 ( \23682 , \23402 , \23406 );
and \U$23368 ( \23683 , \23406 , \23411 );
and \U$23369 ( \23684 , \23402 , \23411 );
or \U$23370 ( \23685 , \23682 , \23683 , \23684 );
xor \U$23371 ( \23686 , \23681 , \23685 );
and \U$23372 ( \23687 , \23388 , \23392 );
and \U$23373 ( \23688 , \23392 , \23397 );
and \U$23374 ( \23689 , \23388 , \23397 );
or \U$23375 ( \23690 , \23687 , \23688 , \23689 );
xor \U$23376 ( \23691 , \23686 , \23690 );
and \U$23377 ( \23692 , \23372 , \23376 );
and \U$23378 ( \23693 , \23376 , \23381 );
and \U$23379 ( \23694 , \23372 , \23381 );
or \U$23380 ( \23695 , \23692 , \23693 , \23694 );
and \U$23381 ( \23696 , \23357 , \23361 );
and \U$23382 ( \23697 , \23361 , \23366 );
and \U$23383 ( \23698 , \23357 , \23366 );
or \U$23384 ( \23699 , \23696 , \23697 , \23698 );
xor \U$23385 ( \23700 , \23695 , \23699 );
and \U$23386 ( \23701 , \23343 , \23347 );
and \U$23387 ( \23702 , \23347 , \23352 );
and \U$23388 ( \23703 , \23343 , \23352 );
or \U$23389 ( \23704 , \23701 , \23702 , \23703 );
xor \U$23390 ( \23705 , \23700 , \23704 );
xor \U$23391 ( \23706 , \23691 , \23705 );
and \U$23392 ( \23707 , \21595 , \23332 );
and \U$23393 ( \23708 , \23332 , \23337 );
and \U$23394 ( \23709 , \21595 , \23337 );
or \U$23395 ( \23710 , \23707 , \23708 , \23709 );
and \U$23396 ( \23711 , \23313 , \23317 );
and \U$23397 ( \23712 , \23317 , \23322 );
and \U$23398 ( \23713 , \23313 , \23322 );
or \U$23399 ( \23714 , \23711 , \23712 , \23713 );
xor \U$23400 ( \23715 , \23710 , \23714 );
and \U$23401 ( \23716 , \23299 , \23303 );
and \U$23402 ( \23717 , \23303 , \23308 );
and \U$23403 ( \23718 , \23299 , \23308 );
or \U$23404 ( \23719 , \23716 , \23717 , \23718 );
xor \U$23405 ( \23720 , \23715 , \23719 );
xor \U$23406 ( \23721 , \23706 , \23720 );
xor \U$23407 ( \23722 , \23677 , \23721 );
and \U$23408 ( \23723 , \22440 , \22484 );
and \U$23409 ( \23724 , \22407 , \22482 );
nor \U$23410 ( \23725 , \23723 , \23724 );
xnor \U$23411 ( \23726 , \23725 , \22494 );
and \U$23412 ( \23727 , \22468 , \22506 );
and \U$23413 ( \23728 , \22429 , \22504 );
nor \U$23414 ( \23729 , \23727 , \23728 );
xnor \U$23415 ( \23730 , \23729 , \22516 );
xor \U$23416 ( \23731 , \23726 , \23730 );
and \U$23417 ( \23732 , \22489 , \22530 );
and \U$23418 ( \23733 , \22457 , \22528 );
nor \U$23419 ( \23734 , \23732 , \23733 );
xnor \U$23420 ( \23735 , \23734 , \22540 );
xor \U$23421 ( \23736 , \23731 , \23735 );
and \U$23422 ( \23737 , \22372 , \22413 );
and \U$23423 ( \23738 , \22339 , \22411 );
nor \U$23424 ( \23739 , \23737 , \23738 );
xnor \U$23425 ( \23740 , \23739 , \22423 );
and \U$23426 ( \23741 , \22397 , \22435 );
and \U$23427 ( \23742 , \22361 , \22433 );
nor \U$23428 ( \23743 , \23741 , \23742 );
xnor \U$23429 ( \23744 , \23743 , \22445 );
xor \U$23430 ( \23745 , \23740 , \23744 );
and \U$23431 ( \23746 , \22418 , \22463 );
and \U$23432 ( \23747 , \22386 , \22461 );
nor \U$23433 ( \23748 , \23746 , \23747 );
xnor \U$23434 ( \23749 , \23748 , \22473 );
xor \U$23435 ( \23750 , \23745 , \23749 );
xor \U$23436 ( \23751 , \23736 , \23750 );
and \U$23437 ( \23752 , \22305 , \22345 );
and \U$23438 ( \23753 , \22272 , \22343 );
nor \U$23439 ( \23754 , \23752 , \23753 );
xnor \U$23440 ( \23755 , \23754 , \22355 );
and \U$23441 ( \23756 , \22329 , \22367 );
and \U$23442 ( \23757 , \22294 , \22365 );
nor \U$23443 ( \23758 , \23756 , \23757 );
xnor \U$23444 ( \23759 , \23758 , \22377 );
xor \U$23445 ( \23760 , \23755 , \23759 );
and \U$23446 ( \23761 , \22350 , \22392 );
and \U$23447 ( \23762 , \22318 , \22390 );
nor \U$23448 ( \23763 , \23761 , \23762 );
xnor \U$23449 ( \23764 , \23763 , \22402 );
xor \U$23450 ( \23765 , \23760 , \23764 );
xor \U$23451 ( \23766 , \23751 , \23765 );
and \U$23452 ( \23767 , \22646 , \22691 );
and \U$23453 ( \23768 , \22613 , \22689 );
nor \U$23454 ( \23769 , \23767 , \23768 );
xnor \U$23455 ( \23770 , \23769 , \22701 );
and \U$23456 ( \23771 , \22676 , \22720 );
and \U$23457 ( \23772 , \22635 , \22707 );
nor \U$23458 ( \23773 , \23771 , \23772 );
xnor \U$23459 ( \23774 , \23773 , \22067 );
xor \U$23460 ( \23775 , \23770 , \23774 );
and \U$23461 ( \23776 , \22696 , \23173 );
and \U$23462 ( \23777 , \22665 , \22999 );
nor \U$23463 ( \23778 , \23776 , \23777 );
xnor \U$23464 ( \23779 , \23778 , \22016 );
xor \U$23465 ( \23780 , \23775 , \23779 );
and \U$23466 ( \23781 , \22578 , \22619 );
and \U$23467 ( \23782 , \22545 , \22617 );
nor \U$23468 ( \23783 , \23781 , \23782 );
xnor \U$23469 ( \23784 , \23783 , \22629 );
and \U$23470 ( \23785 , \22603 , \22641 );
and \U$23471 ( \23786 , \22567 , \22639 );
nor \U$23472 ( \23787 , \23785 , \23786 );
xnor \U$23473 ( \23788 , \23787 , \22651 );
xor \U$23474 ( \23789 , \23784 , \23788 );
and \U$23475 ( \23790 , \22624 , \22671 );
and \U$23476 ( \23791 , \22592 , \22669 );
nor \U$23477 ( \23792 , \23790 , \23791 );
xnor \U$23478 ( \23793 , \23792 , \22681 );
xor \U$23479 ( \23794 , \23789 , \23793 );
xor \U$23480 ( \23795 , \23780 , \23794 );
and \U$23481 ( \23796 , \22511 , \22551 );
and \U$23482 ( \23797 , \22478 , \22549 );
nor \U$23483 ( \23798 , \23796 , \23797 );
xnor \U$23484 ( \23799 , \23798 , \22561 );
and \U$23485 ( \23800 , \22535 , \22573 );
and \U$23486 ( \23801 , \22500 , \22571 );
nor \U$23487 ( \23802 , \23800 , \23801 );
xnor \U$23488 ( \23803 , \23802 , \22583 );
xor \U$23489 ( \23804 , \23799 , \23803 );
and \U$23490 ( \23805 , \22556 , \22598 );
and \U$23491 ( \23806 , \22524 , \22596 );
nor \U$23492 ( \23807 , \23805 , \23806 );
xnor \U$23493 ( \23808 , \23807 , \22608 );
xor \U$23494 ( \23809 , \23804 , \23808 );
xor \U$23495 ( \23810 , \23795 , \23809 );
xor \U$23496 ( \23811 , \23766 , \23810 );
and \U$23497 ( \23812 , \23494 , \23498 );
and \U$23498 ( \23813 , \23498 , \23503 );
and \U$23499 ( \23814 , \23494 , \23503 );
or \U$23500 ( \23815 , \23812 , \23813 , \23814 );
and \U$23501 ( \23816 , \23486 , \23488 );
xor \U$23502 ( \23817 , \23815 , \23816 );
and \U$23503 ( \23818 , \22706 , \22021 );
and \U$23504 ( \23819 , \22686 , \22019 );
nor \U$23505 ( \23820 , \23818 , \23819 );
xnor \U$23506 ( \23821 , \23820 , \21595 );
xor \U$23507 ( \23822 , \23817 , \23821 );
xor \U$23508 ( \23823 , \23811 , \23822 );
xor \U$23509 ( \23824 , \23722 , \23823 );
xor \U$23510 ( \23825 , \23673 , \23824 );
and \U$23511 ( \23826 , \23448 , \23452 );
and \U$23512 ( \23827 , \23452 , \23457 );
and \U$23513 ( \23828 , \23448 , \23457 );
or \U$23514 ( \23829 , \23826 , \23827 , \23828 );
and \U$23515 ( \23830 , \23433 , \23437 );
and \U$23516 ( \23831 , \23437 , \23442 );
and \U$23517 ( \23832 , \23433 , \23442 );
or \U$23518 ( \23833 , \23830 , \23831 , \23832 );
xor \U$23519 ( \23834 , \23829 , \23833 );
and \U$23520 ( \23835 , \23339 , \23383 );
and \U$23521 ( \23836 , \23383 , \23428 );
and \U$23522 ( \23837 , \23339 , \23428 );
or \U$23523 ( \23838 , \23835 , \23836 , \23837 );
xor \U$23524 ( \23839 , \23834 , \23838 );
xor \U$23525 ( \23840 , \23825 , \23839 );
and \U$23526 ( \23841 , \23578 , \23840 );
and \U$23527 ( \23842 , \23295 , \23840 );
or \U$23528 ( \23843 , \23579 , \23841 , \23842 );
and \U$23529 ( \23844 , \23662 , \23666 );
and \U$23530 ( \23845 , \23666 , \23671 );
and \U$23531 ( \23846 , \23662 , \23671 );
or \U$23532 ( \23847 , \23844 , \23845 , \23846 );
and \U$23533 ( \23848 , \23647 , \23651 );
and \U$23534 ( \23849 , \23651 , \23656 );
and \U$23535 ( \23850 , \23647 , \23656 );
or \U$23536 ( \23851 , \23848 , \23849 , \23850 );
xor \U$23537 ( \23852 , \23847 , \23851 );
and \U$23538 ( \23853 , \23583 , \23597 );
and \U$23539 ( \23854 , \23597 , \23642 );
and \U$23540 ( \23855 , \23583 , \23642 );
or \U$23541 ( \23856 , \23853 , \23854 , \23855 );
xor \U$23542 ( \23857 , \23852 , \23856 );
and \U$23543 ( \23858 , \23815 , \23816 );
and \U$23544 ( \23859 , \23816 , \23821 );
and \U$23545 ( \23860 , \23815 , \23821 );
or \U$23546 ( \23861 , \23858 , \23859 , \23860 );
and \U$23547 ( \23862 , \23780 , \23794 );
and \U$23548 ( \23863 , \23794 , \23809 );
and \U$23549 ( \23864 , \23780 , \23809 );
or \U$23550 ( \23865 , \23862 , \23863 , \23864 );
xor \U$23551 ( \23866 , \23861 , \23865 );
and \U$23552 ( \23867 , \23736 , \23750 );
and \U$23553 ( \23868 , \23750 , \23765 );
and \U$23554 ( \23869 , \23736 , \23765 );
or \U$23555 ( \23870 , \23867 , \23868 , \23869 );
xor \U$23556 ( \23871 , \23866 , \23870 );
and \U$23557 ( \23872 , \23710 , \23714 );
and \U$23558 ( \23873 , \23714 , \23719 );
and \U$23559 ( \23874 , \23710 , \23719 );
or \U$23560 ( \23875 , \23872 , \23873 , \23874 );
and \U$23561 ( \23876 , \23695 , \23699 );
and \U$23562 ( \23877 , \23699 , \23704 );
and \U$23563 ( \23878 , \23695 , \23704 );
or \U$23564 ( \23879 , \23876 , \23877 , \23878 );
xor \U$23565 ( \23880 , \23875 , \23879 );
and \U$23566 ( \23881 , \23681 , \23685 );
and \U$23567 ( \23882 , \23685 , \23690 );
and \U$23568 ( \23883 , \23681 , \23690 );
or \U$23569 ( \23884 , \23881 , \23882 , \23883 );
xor \U$23570 ( \23885 , \23880 , \23884 );
xor \U$23571 ( \23886 , \23871 , \23885 );
and \U$23572 ( \23887 , \23587 , \23591 );
and \U$23573 ( \23888 , \23591 , \23596 );
and \U$23574 ( \23889 , \23587 , \23596 );
or \U$23575 ( \23890 , \23887 , \23888 , \23889 );
and \U$23576 ( \23891 , \23631 , \23635 );
and \U$23577 ( \23892 , \23635 , \23640 );
and \U$23578 ( \23893 , \23631 , \23640 );
or \U$23579 ( \23894 , \23891 , \23892 , \23893 );
xor \U$23580 ( \23895 , \23890 , \23894 );
and \U$23581 ( \23896 , \23616 , \23620 );
and \U$23582 ( \23897 , \23620 , \23625 );
and \U$23583 ( \23898 , \23616 , \23625 );
or \U$23584 ( \23899 , \23896 , \23897 , \23898 );
xor \U$23585 ( \23900 , \23895 , \23899 );
and \U$23586 ( \23901 , \22524 , \22598 );
and \U$23587 ( \23902 , \22535 , \22596 );
nor \U$23588 ( \23903 , \23901 , \23902 );
xnor \U$23589 ( \23904 , \23903 , \22608 );
and \U$23590 ( \23905 , \22545 , \22619 );
and \U$23591 ( \23906 , \22556 , \22617 );
nor \U$23592 ( \23907 , \23905 , \23906 );
xnor \U$23593 ( \23908 , \23907 , \22629 );
xor \U$23594 ( \23909 , \23904 , \23908 );
and \U$23595 ( \23910 , \22567 , \22641 );
and \U$23596 ( \23911 , \22578 , \22639 );
nor \U$23597 ( \23912 , \23910 , \23911 );
xnor \U$23598 ( \23913 , \23912 , \22651 );
xor \U$23599 ( \23914 , \23909 , \23913 );
and \U$23600 ( \23915 , \22457 , \22530 );
and \U$23601 ( \23916 , \22468 , \22528 );
nor \U$23602 ( \23917 , \23915 , \23916 );
xnor \U$23603 ( \23918 , \23917 , \22540 );
and \U$23604 ( \23919 , \22478 , \22551 );
and \U$23605 ( \23920 , \22489 , \22549 );
nor \U$23606 ( \23921 , \23919 , \23920 );
xnor \U$23607 ( \23922 , \23921 , \22561 );
xor \U$23608 ( \23923 , \23918 , \23922 );
and \U$23609 ( \23924 , \22500 , \22573 );
and \U$23610 ( \23925 , \22511 , \22571 );
nor \U$23611 ( \23926 , \23924 , \23925 );
xnor \U$23612 ( \23927 , \23926 , \22583 );
xor \U$23613 ( \23928 , \23923 , \23927 );
xor \U$23614 ( \23929 , \23914 , \23928 );
and \U$23615 ( \23930 , \22386 , \22463 );
and \U$23616 ( \23931 , \22397 , \22461 );
nor \U$23617 ( \23932 , \23930 , \23931 );
xnor \U$23618 ( \23933 , \23932 , \22473 );
and \U$23619 ( \23934 , \22407 , \22484 );
and \U$23620 ( \23935 , \22418 , \22482 );
nor \U$23621 ( \23936 , \23934 , \23935 );
xnor \U$23622 ( \23937 , \23936 , \22494 );
xor \U$23623 ( \23938 , \23933 , \23937 );
and \U$23624 ( \23939 , \22429 , \22506 );
and \U$23625 ( \23940 , \22440 , \22504 );
nor \U$23626 ( \23941 , \23939 , \23940 );
xnor \U$23627 ( \23942 , \23941 , \22516 );
xor \U$23628 ( \23943 , \23938 , \23942 );
xor \U$23629 ( \23944 , \23929 , \23943 );
and \U$23630 ( \23945 , \23770 , \23774 );
and \U$23631 ( \23946 , \23774 , \23779 );
and \U$23632 ( \23947 , \23770 , \23779 );
or \U$23633 ( \23948 , \23945 , \23946 , \23947 );
and \U$23634 ( \23949 , \22665 , \23173 );
and \U$23635 ( \23950 , \22676 , \22999 );
nor \U$23636 ( \23951 , \23949 , \23950 );
xnor \U$23637 ( \23952 , \23951 , \22016 );
and \U$23638 ( \23953 , \22686 , \22021 );
and \U$23639 ( \23954 , \22696 , \22019 );
nor \U$23640 ( \23955 , \23953 , \23954 );
xnor \U$23641 ( \23956 , \23955 , \21595 );
xor \U$23642 ( \23957 , \23952 , \23956 );
nand \U$23643 ( \23958 , \22706 , \21981 );
xnor \U$23644 ( \23959 , \23958 , \21995 );
xor \U$23645 ( \23960 , \23957 , \23959 );
xor \U$23646 ( \23961 , \23948 , \23960 );
and \U$23647 ( \23962 , \22592 , \22671 );
and \U$23648 ( \23963 , \22603 , \22669 );
nor \U$23649 ( \23964 , \23962 , \23963 );
xnor \U$23650 ( \23965 , \23964 , \22681 );
and \U$23651 ( \23966 , \22613 , \22691 );
and \U$23652 ( \23967 , \22624 , \22689 );
nor \U$23653 ( \23968 , \23966 , \23967 );
xnor \U$23654 ( \23969 , \23968 , \22701 );
xor \U$23655 ( \23970 , \23965 , \23969 );
and \U$23656 ( \23971 , \22635 , \22720 );
and \U$23657 ( \23972 , \22646 , \22707 );
nor \U$23658 ( \23973 , \23971 , \23972 );
xnor \U$23659 ( \23974 , \23973 , \22067 );
xor \U$23660 ( \23975 , \23970 , \23974 );
xor \U$23661 ( \23976 , \23961 , \23975 );
xor \U$23662 ( \23977 , \23944 , \23976 );
and \U$23663 ( \23978 , \23726 , \23730 );
and \U$23664 ( \23979 , \23730 , \23735 );
and \U$23665 ( \23980 , \23726 , \23735 );
or \U$23666 ( \23981 , \23978 , \23979 , \23980 );
and \U$23667 ( \23982 , \23799 , \23803 );
and \U$23668 ( \23983 , \23803 , \23808 );
and \U$23669 ( \23984 , \23799 , \23808 );
or \U$23670 ( \23985 , \23982 , \23983 , \23984 );
xor \U$23671 ( \23986 , \23981 , \23985 );
and \U$23672 ( \23987 , \23784 , \23788 );
and \U$23673 ( \23988 , \23788 , \23793 );
and \U$23674 ( \23989 , \23784 , \23793 );
or \U$23675 ( \23990 , \23987 , \23988 , \23989 );
xor \U$23676 ( \23991 , \23986 , \23990 );
xor \U$23677 ( \23992 , \23977 , \23991 );
xor \U$23678 ( \23993 , \23900 , \23992 );
and \U$23679 ( \23994 , \23612 , \23626 );
and \U$23680 ( \23995 , \23626 , \23641 );
and \U$23681 ( \23996 , \23612 , \23641 );
or \U$23682 ( \23997 , \23994 , \23995 , \23996 );
and \U$23683 ( \23998 , \22113 , \22187 );
and \U$23684 ( \23999 , \22124 , \22185 );
nor \U$23685 ( \24000 , \23998 , \23999 );
xnor \U$23686 ( \24001 , \24000 , \22197 );
and \U$23687 ( \24002 , \22134 , \22208 );
and \U$23688 ( \24003 , \22145 , \22206 );
nor \U$23689 ( \24004 , \24002 , \24003 );
xnor \U$23690 ( \24005 , \24004 , \22218 );
xor \U$23691 ( \24006 , \24001 , \24005 );
and \U$23692 ( \24007 , \22156 , \22230 );
and \U$23693 ( \24008 , \22167 , \22228 );
nor \U$23694 ( \24009 , \24007 , \24008 );
xnor \U$23695 ( \24010 , \24009 , \22240 );
xor \U$23696 ( \24011 , \24006 , \24010 );
and \U$23697 ( \24012 , \22858 , \22119 );
and \U$23698 ( \24013 , \22894 , \22117 );
nor \U$23699 ( \24014 , \24012 , \24013 );
xnor \U$23700 ( \24015 , \24014 , \22129 );
and \U$23701 ( \24016 , \22071 , \22140 );
and \U$23702 ( \24017 , \22081 , \22138 );
nor \U$23703 ( \24018 , \24016 , \24017 );
xnor \U$23704 ( \24019 , \24018 , \22150 );
xor \U$23705 ( \24020 , \24015 , \24019 );
and \U$23706 ( \24021 , \22089 , \22162 );
and \U$23707 ( \24022 , \22100 , \22160 );
nor \U$23708 ( \24023 , \24021 , \24022 );
xnor \U$23709 ( \24024 , \24023 , \22172 );
xor \U$23710 ( \24025 , \24020 , \24024 );
xor \U$23711 ( \24026 , \24011 , \24025 );
and \U$23712 ( \24027 , \22030 , \22076 );
and \U$23713 ( \24028 , \22001 , \22073 );
nor \U$23714 ( \24029 , \24027 , \24028 );
xnor \U$23715 ( \24030 , \24029 , \22072 );
xor \U$23716 ( \24031 , \21995 , \24030 );
and \U$23717 ( \24032 , \23230 , \22095 );
and \U$23718 ( \24033 , \23329 , \22093 );
nor \U$23719 ( \24034 , \24032 , \24033 );
xnor \U$23720 ( \24035 , \24034 , \22105 );
xor \U$23721 ( \24036 , \24031 , \24035 );
xor \U$23722 ( \24037 , \24026 , \24036 );
xor \U$23723 ( \24038 , \23997 , \24037 );
and \U$23724 ( \24039 , \22318 , \22392 );
and \U$23725 ( \24040 , \22329 , \22390 );
nor \U$23726 ( \24041 , \24039 , \24040 );
xnor \U$23727 ( \24042 , \24041 , \22402 );
and \U$23728 ( \24043 , \22339 , \22413 );
and \U$23729 ( \24044 , \22350 , \22411 );
nor \U$23730 ( \24045 , \24043 , \24044 );
xnor \U$23731 ( \24046 , \24045 , \22423 );
xor \U$23732 ( \24047 , \24042 , \24046 );
and \U$23733 ( \24048 , \22361 , \22435 );
and \U$23734 ( \24049 , \22372 , \22433 );
nor \U$23735 ( \24050 , \24048 , \24049 );
xnor \U$23736 ( \24051 , \24050 , \22445 );
xor \U$23737 ( \24052 , \24047 , \24051 );
and \U$23738 ( \24053 , \22251 , \22324 );
and \U$23739 ( \24054 , \22262 , \22322 );
nor \U$23740 ( \24055 , \24053 , \24054 );
xnor \U$23741 ( \24056 , \24055 , \22334 );
and \U$23742 ( \24057 , \22272 , \22345 );
and \U$23743 ( \24058 , \22283 , \22343 );
nor \U$23744 ( \24059 , \24057 , \24058 );
xnor \U$23745 ( \24060 , \24059 , \22355 );
xor \U$23746 ( \24061 , \24056 , \24060 );
and \U$23747 ( \24062 , \22294 , \22367 );
and \U$23748 ( \24063 , \22305 , \22365 );
nor \U$23749 ( \24064 , \24062 , \24063 );
xnor \U$23750 ( \24065 , \24064 , \22377 );
xor \U$23751 ( \24066 , \24061 , \24065 );
xor \U$23752 ( \24067 , \24052 , \24066 );
and \U$23753 ( \24068 , \22181 , \22257 );
and \U$23754 ( \24069 , \22192 , \22255 );
nor \U$23755 ( \24070 , \24068 , \24069 );
xnor \U$23756 ( \24071 , \24070 , \22267 );
and \U$23757 ( \24072 , \22202 , \22278 );
and \U$23758 ( \24073 , \22213 , \22276 );
nor \U$23759 ( \24074 , \24072 , \24073 );
xnor \U$23760 ( \24075 , \24074 , \22288 );
xor \U$23761 ( \24076 , \24071 , \24075 );
and \U$23762 ( \24077 , \22224 , \22300 );
and \U$23763 ( \24078 , \22235 , \22298 );
nor \U$23764 ( \24079 , \24077 , \24078 );
xnor \U$23765 ( \24080 , \24079 , \22310 );
xor \U$23766 ( \24081 , \24076 , \24080 );
xor \U$23767 ( \24082 , \24067 , \24081 );
xor \U$23768 ( \24083 , \24038 , \24082 );
xor \U$23769 ( \24084 , \23993 , \24083 );
xor \U$23770 ( \24085 , \23886 , \24084 );
xor \U$23771 ( \24086 , \23857 , \24085 );
and \U$23772 ( \24087 , \23829 , \23833 );
and \U$23773 ( \24088 , \23833 , \23838 );
and \U$23774 ( \24089 , \23829 , \23838 );
or \U$23775 ( \24090 , \24087 , \24088 , \24089 );
and \U$23776 ( \24091 , \23677 , \23721 );
and \U$23777 ( \24092 , \23721 , \23823 );
and \U$23778 ( \24093 , \23677 , \23823 );
or \U$23779 ( \24094 , \24091 , \24092 , \24093 );
xor \U$23780 ( \24095 , \24090 , \24094 );
and \U$23781 ( \24096 , \23643 , \23657 );
and \U$23782 ( \24097 , \23657 , \23672 );
and \U$23783 ( \24098 , \23643 , \23672 );
or \U$23784 ( \24099 , \24096 , \24097 , \24098 );
xor \U$23785 ( \24100 , \24095 , \24099 );
xor \U$23786 ( \24101 , \24086 , \24100 );
and \U$23787 ( \24102 , \23843 , \24101 );
and \U$23788 ( \24103 , \23553 , \23569 );
and \U$23789 ( \24104 , \23569 , \23574 );
and \U$23790 ( \24105 , \23553 , \23574 );
or \U$23791 ( \24106 , \24103 , \24104 , \24105 );
and \U$23792 ( \24107 , \23463 , \23477 );
and \U$23793 ( \24108 , \23477 , \23535 );
and \U$23794 ( \24109 , \23463 , \23535 );
or \U$23795 ( \24110 , \24107 , \24108 , \24109 );
and \U$23796 ( \24111 , \24106 , \24110 );
and \U$23797 ( \24112 , \23429 , \23443 );
and \U$23798 ( \24113 , \23443 , \23458 );
and \U$23799 ( \24114 , \23429 , \23458 );
or \U$23800 ( \24115 , \24112 , \24113 , \24114 );
and \U$23801 ( \24116 , \24110 , \24115 );
and \U$23802 ( \24117 , \24106 , \24115 );
or \U$23803 ( \24118 , \24111 , \24116 , \24117 );
and \U$23804 ( \24119 , \23673 , \23824 );
and \U$23805 ( \24120 , \23824 , \23839 );
and \U$23806 ( \24121 , \23673 , \23839 );
or \U$23807 ( \24122 , \24119 , \24120 , \24121 );
xor \U$23808 ( \24123 , \24118 , \24122 );
and \U$23809 ( \24124 , \23766 , \23810 );
and \U$23810 ( \24125 , \23810 , \23822 );
and \U$23811 ( \24126 , \23766 , \23822 );
or \U$23812 ( \24127 , \24124 , \24125 , \24126 );
and \U$23813 ( \24128 , \23691 , \23705 );
and \U$23814 ( \24129 , \23705 , \23720 );
and \U$23815 ( \24130 , \23691 , \23720 );
or \U$23816 ( \24131 , \24128 , \24129 , \24130 );
xor \U$23817 ( \24132 , \24127 , \24131 );
and \U$23818 ( \24133 , \23602 , \23606 );
and \U$23819 ( \24134 , \23606 , \23611 );
and \U$23820 ( \24135 , \23602 , \23611 );
or \U$23821 ( \24136 , \24133 , \24134 , \24135 );
and \U$23822 ( \24137 , \23755 , \23759 );
and \U$23823 ( \24138 , \23759 , \23764 );
and \U$23824 ( \24139 , \23755 , \23764 );
or \U$23825 ( \24140 , \24137 , \24138 , \24139 );
xor \U$23826 ( \24141 , \24136 , \24140 );
and \U$23827 ( \24142 , \23740 , \23744 );
and \U$23828 ( \24143 , \23744 , \23749 );
and \U$23829 ( \24144 , \23740 , \23749 );
or \U$23830 ( \24145 , \24142 , \24143 , \24144 );
xor \U$23831 ( \24146 , \24141 , \24145 );
xor \U$23832 ( \24147 , \24132 , \24146 );
xor \U$23833 ( \24148 , \24123 , \24147 );
and \U$23834 ( \24149 , \24101 , \24148 );
and \U$23835 ( \24150 , \23843 , \24148 );
or \U$23836 ( \24151 , \24102 , \24149 , \24150 );
and \U$23837 ( \24152 , \24090 , \24094 );
and \U$23838 ( \24153 , \24094 , \24099 );
and \U$23839 ( \24154 , \24090 , \24099 );
or \U$23840 ( \24155 , \24152 , \24153 , \24154 );
and \U$23841 ( \24156 , \23871 , \23885 );
and \U$23842 ( \24157 , \23885 , \24084 );
and \U$23843 ( \24158 , \23871 , \24084 );
or \U$23844 ( \24159 , \24156 , \24157 , \24158 );
xor \U$23845 ( \24160 , \24155 , \24159 );
and \U$23846 ( \24161 , \24011 , \24025 );
and \U$23847 ( \24162 , \24025 , \24036 );
and \U$23848 ( \24163 , \24011 , \24036 );
or \U$23849 ( \24164 , \24161 , \24162 , \24163 );
and \U$23850 ( \24165 , \22081 , \22140 );
and \U$23851 ( \24166 , \22858 , \22138 );
nor \U$23852 ( \24167 , \24165 , \24166 );
xnor \U$23853 ( \24168 , \24167 , \22150 );
and \U$23854 ( \24169 , \22100 , \22162 );
and \U$23855 ( \24170 , \22071 , \22160 );
nor \U$23856 ( \24171 , \24169 , \24170 );
xnor \U$23857 ( \24172 , \24171 , \22172 );
xor \U$23858 ( \24173 , \24168 , \24172 );
and \U$23859 ( \24174 , \22124 , \22187 );
and \U$23860 ( \24175 , \22089 , \22185 );
nor \U$23861 ( \24176 , \24174 , \24175 );
xnor \U$23862 ( \24177 , \24176 , \22197 );
xor \U$23863 ( \24178 , \24173 , \24177 );
and \U$23864 ( \24179 , \22001 , \22076 );
and \U$23865 ( \24180 , \21977 , \22073 );
nor \U$23866 ( \24181 , \24179 , \24180 );
xnor \U$23867 ( \24182 , \24181 , \22072 );
and \U$23868 ( \24183 , \23329 , \22095 );
and \U$23869 ( \24184 , \22030 , \22093 );
nor \U$23870 ( \24185 , \24183 , \24184 );
xnor \U$23871 ( \24186 , \24185 , \22105 );
xor \U$23872 ( \24187 , \24182 , \24186 );
and \U$23873 ( \24188 , \22894 , \22119 );
and \U$23874 ( \24189 , \23230 , \22117 );
nor \U$23875 ( \24190 , \24188 , \24189 );
xnor \U$23876 ( \24191 , \24190 , \22129 );
xor \U$23877 ( \24192 , \24187 , \24191 );
xor \U$23878 ( \24193 , \24178 , \24192 );
xor \U$23879 ( \24194 , \24164 , \24193 );
and \U$23880 ( \24195 , \22283 , \22345 );
and \U$23881 ( \24196 , \22251 , \22343 );
nor \U$23882 ( \24197 , \24195 , \24196 );
xnor \U$23883 ( \24198 , \24197 , \22355 );
and \U$23884 ( \24199 , \22305 , \22367 );
and \U$23885 ( \24200 , \22272 , \22365 );
nor \U$23886 ( \24201 , \24199 , \24200 );
xnor \U$23887 ( \24202 , \24201 , \22377 );
xor \U$23888 ( \24203 , \24198 , \24202 );
and \U$23889 ( \24204 , \22329 , \22392 );
and \U$23890 ( \24205 , \22294 , \22390 );
nor \U$23891 ( \24206 , \24204 , \24205 );
xnor \U$23892 ( \24207 , \24206 , \22402 );
xor \U$23893 ( \24208 , \24203 , \24207 );
and \U$23894 ( \24209 , \22213 , \22278 );
and \U$23895 ( \24210 , \22181 , \22276 );
nor \U$23896 ( \24211 , \24209 , \24210 );
xnor \U$23897 ( \24212 , \24211 , \22288 );
and \U$23898 ( \24213 , \22235 , \22300 );
and \U$23899 ( \24214 , \22202 , \22298 );
nor \U$23900 ( \24215 , \24213 , \24214 );
xnor \U$23901 ( \24216 , \24215 , \22310 );
xor \U$23902 ( \24217 , \24212 , \24216 );
and \U$23903 ( \24218 , \22262 , \22324 );
and \U$23904 ( \24219 , \22224 , \22322 );
nor \U$23905 ( \24220 , \24218 , \24219 );
xnor \U$23906 ( \24221 , \24220 , \22334 );
xor \U$23907 ( \24222 , \24217 , \24221 );
xor \U$23908 ( \24223 , \24208 , \24222 );
and \U$23909 ( \24224 , \22145 , \22208 );
and \U$23910 ( \24225 , \22113 , \22206 );
nor \U$23911 ( \24226 , \24224 , \24225 );
xnor \U$23912 ( \24227 , \24226 , \22218 );
and \U$23913 ( \24228 , \22167 , \22230 );
and \U$23914 ( \24229 , \22134 , \22228 );
nor \U$23915 ( \24230 , \24228 , \24229 );
xnor \U$23916 ( \24231 , \24230 , \22240 );
xor \U$23917 ( \24232 , \24227 , \24231 );
and \U$23918 ( \24233 , \22192 , \22257 );
and \U$23919 ( \24234 , \22156 , \22255 );
nor \U$23920 ( \24235 , \24233 , \24234 );
xnor \U$23921 ( \24236 , \24235 , \22267 );
xor \U$23922 ( \24237 , \24232 , \24236 );
xor \U$23923 ( \24238 , \24223 , \24237 );
xor \U$23924 ( \24239 , \24194 , \24238 );
and \U$23925 ( \24240 , \23948 , \23960 );
and \U$23926 ( \24241 , \23960 , \23975 );
and \U$23927 ( \24242 , \23948 , \23975 );
or \U$23928 ( \24243 , \24240 , \24241 , \24242 );
and \U$23929 ( \24244 , \23914 , \23928 );
and \U$23930 ( \24245 , \23928 , \23943 );
and \U$23931 ( \24246 , \23914 , \23943 );
or \U$23932 ( \24247 , \24244 , \24245 , \24246 );
xor \U$23933 ( \24248 , \24243 , \24247 );
and \U$23934 ( \24249 , \24052 , \24066 );
and \U$23935 ( \24250 , \24066 , \24081 );
and \U$23936 ( \24251 , \24052 , \24081 );
or \U$23937 ( \24252 , \24249 , \24250 , \24251 );
xor \U$23938 ( \24253 , \24248 , \24252 );
xor \U$23939 ( \24254 , \24239 , \24253 );
and \U$23940 ( \24255 , \23890 , \23894 );
and \U$23941 ( \24256 , \23894 , \23899 );
and \U$23942 ( \24257 , \23890 , \23899 );
or \U$23943 ( \24258 , \24255 , \24256 , \24257 );
and \U$23944 ( \24259 , \24136 , \24140 );
and \U$23945 ( \24260 , \24140 , \24145 );
and \U$23946 ( \24261 , \24136 , \24145 );
or \U$23947 ( \24262 , \24259 , \24260 , \24261 );
xor \U$23948 ( \24263 , \24258 , \24262 );
and \U$23949 ( \24264 , \23981 , \23985 );
and \U$23950 ( \24265 , \23985 , \23990 );
and \U$23951 ( \24266 , \23981 , \23990 );
or \U$23952 ( \24267 , \24264 , \24265 , \24266 );
xor \U$23953 ( \24268 , \24263 , \24267 );
xor \U$23954 ( \24269 , \24254 , \24268 );
and \U$23955 ( \24270 , \23944 , \23976 );
and \U$23956 ( \24271 , \23976 , \23991 );
and \U$23957 ( \24272 , \23944 , \23991 );
or \U$23958 ( \24273 , \24270 , \24271 , \24272 );
and \U$23959 ( \24274 , \23933 , \23937 );
and \U$23960 ( \24275 , \23937 , \23942 );
and \U$23961 ( \24276 , \23933 , \23942 );
or \U$23962 ( \24277 , \24274 , \24275 , \24276 );
and \U$23963 ( \24278 , \23918 , \23922 );
and \U$23964 ( \24279 , \23922 , \23927 );
and \U$23965 ( \24280 , \23918 , \23927 );
or \U$23966 ( \24281 , \24278 , \24279 , \24280 );
xor \U$23967 ( \24282 , \24277 , \24281 );
and \U$23968 ( \24283 , \23904 , \23908 );
and \U$23969 ( \24284 , \23908 , \23913 );
and \U$23970 ( \24285 , \23904 , \23913 );
or \U$23971 ( \24286 , \24283 , \24284 , \24285 );
xor \U$23972 ( \24287 , \24282 , \24286 );
and \U$23973 ( \24288 , \24071 , \24075 );
and \U$23974 ( \24289 , \24075 , \24080 );
and \U$23975 ( \24290 , \24071 , \24080 );
or \U$23976 ( \24291 , \24288 , \24289 , \24290 );
and \U$23977 ( \24292 , \24056 , \24060 );
and \U$23978 ( \24293 , \24060 , \24065 );
and \U$23979 ( \24294 , \24056 , \24065 );
or \U$23980 ( \24295 , \24292 , \24293 , \24294 );
xor \U$23981 ( \24296 , \24291 , \24295 );
and \U$23982 ( \24297 , \24042 , \24046 );
and \U$23983 ( \24298 , \24046 , \24051 );
and \U$23984 ( \24299 , \24042 , \24051 );
or \U$23985 ( \24300 , \24297 , \24298 , \24299 );
xor \U$23986 ( \24301 , \24296 , \24300 );
xor \U$23987 ( \24302 , \24287 , \24301 );
and \U$23988 ( \24303 , \21995 , \24030 );
and \U$23989 ( \24304 , \24030 , \24035 );
and \U$23990 ( \24305 , \21995 , \24035 );
or \U$23991 ( \24306 , \24303 , \24304 , \24305 );
and \U$23992 ( \24307 , \24015 , \24019 );
and \U$23993 ( \24308 , \24019 , \24024 );
and \U$23994 ( \24309 , \24015 , \24024 );
or \U$23995 ( \24310 , \24307 , \24308 , \24309 );
xor \U$23996 ( \24311 , \24306 , \24310 );
and \U$23997 ( \24312 , \24001 , \24005 );
and \U$23998 ( \24313 , \24005 , \24010 );
and \U$23999 ( \24314 , \24001 , \24010 );
or \U$24000 ( \24315 , \24312 , \24313 , \24314 );
xor \U$24001 ( \24316 , \24311 , \24315 );
xor \U$24002 ( \24317 , \24302 , \24316 );
xor \U$24003 ( \24318 , \24273 , \24317 );
and \U$24004 ( \24319 , \22489 , \22551 );
and \U$24005 ( \24320 , \22457 , \22549 );
nor \U$24006 ( \24321 , \24319 , \24320 );
xnor \U$24007 ( \24322 , \24321 , \22561 );
and \U$24008 ( \24323 , \22511 , \22573 );
and \U$24009 ( \24324 , \22478 , \22571 );
nor \U$24010 ( \24325 , \24323 , \24324 );
xnor \U$24011 ( \24326 , \24325 , \22583 );
xor \U$24012 ( \24327 , \24322 , \24326 );
and \U$24013 ( \24328 , \22535 , \22598 );
and \U$24014 ( \24329 , \22500 , \22596 );
nor \U$24015 ( \24330 , \24328 , \24329 );
xnor \U$24016 ( \24331 , \24330 , \22608 );
xor \U$24017 ( \24332 , \24327 , \24331 );
and \U$24018 ( \24333 , \22418 , \22484 );
and \U$24019 ( \24334 , \22386 , \22482 );
nor \U$24020 ( \24335 , \24333 , \24334 );
xnor \U$24021 ( \24336 , \24335 , \22494 );
and \U$24022 ( \24337 , \22440 , \22506 );
and \U$24023 ( \24338 , \22407 , \22504 );
nor \U$24024 ( \24339 , \24337 , \24338 );
xnor \U$24025 ( \24340 , \24339 , \22516 );
xor \U$24026 ( \24341 , \24336 , \24340 );
and \U$24027 ( \24342 , \22468 , \22530 );
and \U$24028 ( \24343 , \22429 , \22528 );
nor \U$24029 ( \24344 , \24342 , \24343 );
xnor \U$24030 ( \24345 , \24344 , \22540 );
xor \U$24031 ( \24346 , \24341 , \24345 );
xor \U$24032 ( \24347 , \24332 , \24346 );
and \U$24033 ( \24348 , \22350 , \22413 );
and \U$24034 ( \24349 , \22318 , \22411 );
nor \U$24035 ( \24350 , \24348 , \24349 );
xnor \U$24036 ( \24351 , \24350 , \22423 );
and \U$24037 ( \24352 , \22372 , \22435 );
and \U$24038 ( \24353 , \22339 , \22433 );
nor \U$24039 ( \24354 , \24352 , \24353 );
xnor \U$24040 ( \24355 , \24354 , \22445 );
xor \U$24041 ( \24356 , \24351 , \24355 );
and \U$24042 ( \24357 , \22397 , \22463 );
and \U$24043 ( \24358 , \22361 , \22461 );
nor \U$24044 ( \24359 , \24357 , \24358 );
xnor \U$24045 ( \24360 , \24359 , \22473 );
xor \U$24046 ( \24361 , \24356 , \24360 );
xor \U$24047 ( \24362 , \24347 , \24361 );
and \U$24048 ( \24363 , \22706 , \21983 );
and \U$24049 ( \24364 , \22686 , \21981 );
nor \U$24050 ( \24365 , \24363 , \24364 );
xnor \U$24051 ( \24366 , \24365 , \21995 );
and \U$24052 ( \24367 , \22624 , \22691 );
and \U$24053 ( \24368 , \22592 , \22689 );
nor \U$24054 ( \24369 , \24367 , \24368 );
xnor \U$24055 ( \24370 , \24369 , \22701 );
and \U$24056 ( \24371 , \22646 , \22720 );
and \U$24057 ( \24372 , \22613 , \22707 );
nor \U$24058 ( \24373 , \24371 , \24372 );
xnor \U$24059 ( \24374 , \24373 , \22067 );
xor \U$24060 ( \24375 , \24370 , \24374 );
and \U$24061 ( \24376 , \22676 , \23173 );
and \U$24062 ( \24377 , \22635 , \22999 );
nor \U$24063 ( \24378 , \24376 , \24377 );
xnor \U$24064 ( \24379 , \24378 , \22016 );
xor \U$24065 ( \24380 , \24375 , \24379 );
xor \U$24066 ( \24381 , \24366 , \24380 );
and \U$24067 ( \24382 , \22556 , \22619 );
and \U$24068 ( \24383 , \22524 , \22617 );
nor \U$24069 ( \24384 , \24382 , \24383 );
xnor \U$24070 ( \24385 , \24384 , \22629 );
and \U$24071 ( \24386 , \22578 , \22641 );
and \U$24072 ( \24387 , \22545 , \22639 );
nor \U$24073 ( \24388 , \24386 , \24387 );
xnor \U$24074 ( \24389 , \24388 , \22651 );
xor \U$24075 ( \24390 , \24385 , \24389 );
and \U$24076 ( \24391 , \22603 , \22671 );
and \U$24077 ( \24392 , \22567 , \22669 );
nor \U$24078 ( \24393 , \24391 , \24392 );
xnor \U$24079 ( \24394 , \24393 , \22681 );
xor \U$24080 ( \24395 , \24390 , \24394 );
xor \U$24081 ( \24396 , \24381 , \24395 );
xor \U$24082 ( \24397 , \24362 , \24396 );
and \U$24083 ( \24398 , \23965 , \23969 );
and \U$24084 ( \24399 , \23969 , \23974 );
and \U$24085 ( \24400 , \23965 , \23974 );
or \U$24086 ( \24401 , \24398 , \24399 , \24400 );
and \U$24087 ( \24402 , \23952 , \23956 );
and \U$24088 ( \24403 , \23956 , \23959 );
and \U$24089 ( \24404 , \23952 , \23959 );
or \U$24090 ( \24405 , \24402 , \24403 , \24404 );
xor \U$24091 ( \24406 , \24401 , \24405 );
and \U$24092 ( \24407 , \22696 , \22021 );
and \U$24093 ( \24408 , \22665 , \22019 );
nor \U$24094 ( \24409 , \24407 , \24408 );
xnor \U$24095 ( \24410 , \24409 , \21595 );
xor \U$24096 ( \24411 , \24406 , \24410 );
xor \U$24097 ( \24412 , \24397 , \24411 );
xor \U$24098 ( \24413 , \24318 , \24412 );
xor \U$24099 ( \24414 , \24269 , \24413 );
and \U$24100 ( \24415 , \23875 , \23879 );
and \U$24101 ( \24416 , \23879 , \23884 );
and \U$24102 ( \24417 , \23875 , \23884 );
or \U$24103 ( \24418 , \24415 , \24416 , \24417 );
and \U$24104 ( \24419 , \23861 , \23865 );
and \U$24105 ( \24420 , \23865 , \23870 );
and \U$24106 ( \24421 , \23861 , \23870 );
or \U$24107 ( \24422 , \24419 , \24420 , \24421 );
xor \U$24108 ( \24423 , \24418 , \24422 );
and \U$24109 ( \24424 , \23997 , \24037 );
and \U$24110 ( \24425 , \24037 , \24082 );
and \U$24111 ( \24426 , \23997 , \24082 );
or \U$24112 ( \24427 , \24424 , \24425 , \24426 );
xor \U$24113 ( \24428 , \24423 , \24427 );
xor \U$24114 ( \24429 , \24414 , \24428 );
xor \U$24115 ( \24430 , \24160 , \24429 );
xor \U$24116 ( \24431 , \24151 , \24430 );
and \U$24117 ( \24432 , \24118 , \24122 );
and \U$24118 ( \24433 , \24122 , \24147 );
and \U$24119 ( \24434 , \24118 , \24147 );
or \U$24120 ( \24435 , \24432 , \24433 , \24434 );
and \U$24121 ( \24436 , \23857 , \24085 );
and \U$24122 ( \24437 , \24085 , \24100 );
and \U$24123 ( \24438 , \23857 , \24100 );
or \U$24124 ( \24439 , \24436 , \24437 , \24438 );
xor \U$24125 ( \24440 , \24435 , \24439 );
and \U$24126 ( \24441 , \23847 , \23851 );
and \U$24127 ( \24442 , \23851 , \23856 );
and \U$24128 ( \24443 , \23847 , \23856 );
or \U$24129 ( \24444 , \24441 , \24442 , \24443 );
and \U$24130 ( \24445 , \24127 , \24131 );
and \U$24131 ( \24446 , \24131 , \24146 );
and \U$24132 ( \24447 , \24127 , \24146 );
or \U$24133 ( \24448 , \24445 , \24446 , \24447 );
xor \U$24134 ( \24449 , \24444 , \24448 );
and \U$24135 ( \24450 , \23900 , \23992 );
and \U$24136 ( \24451 , \23992 , \24083 );
and \U$24137 ( \24452 , \23900 , \24083 );
or \U$24138 ( \24453 , \24450 , \24451 , \24452 );
xor \U$24139 ( \24454 , \24449 , \24453 );
xor \U$24140 ( \24455 , \24440 , \24454 );
xor \U$24141 ( \24456 , \24431 , \24455 );
and \U$24142 ( \24457 , \22100 , \22076 );
and \U$24143 ( \24458 , \22071 , \22073 );
nor \U$24144 ( \24459 , \24457 , \24458 );
xnor \U$24145 ( \24460 , \24459 , \22072 );
and \U$24146 ( \24461 , \22124 , \22095 );
and \U$24147 ( \24462 , \22089 , \22093 );
nor \U$24148 ( \24463 , \24461 , \24462 );
xnor \U$24149 ( \24464 , \24463 , \22105 );
and \U$24150 ( \24465 , \24460 , \24464 );
and \U$24151 ( \24466 , \22145 , \22119 );
and \U$24152 ( \24467 , \22113 , \22117 );
nor \U$24153 ( \24468 , \24466 , \24467 );
xnor \U$24154 ( \24469 , \24468 , \22129 );
and \U$24155 ( \24470 , \24464 , \24469 );
and \U$24156 ( \24471 , \24460 , \24469 );
or \U$24157 ( \24472 , \24465 , \24470 , \24471 );
and \U$24158 ( \24473 , \22167 , \22140 );
and \U$24159 ( \24474 , \22134 , \22138 );
nor \U$24160 ( \24475 , \24473 , \24474 );
xnor \U$24161 ( \24476 , \24475 , \22150 );
and \U$24162 ( \24477 , \22192 , \22162 );
and \U$24163 ( \24478 , \22156 , \22160 );
nor \U$24164 ( \24479 , \24477 , \24478 );
xnor \U$24165 ( \24480 , \24479 , \22172 );
and \U$24166 ( \24481 , \24476 , \24480 );
and \U$24167 ( \24482 , \22213 , \22187 );
and \U$24168 ( \24483 , \22181 , \22185 );
nor \U$24169 ( \24484 , \24482 , \24483 );
xnor \U$24170 ( \24485 , \24484 , \22197 );
and \U$24171 ( \24486 , \24480 , \24485 );
and \U$24172 ( \24487 , \24476 , \24485 );
or \U$24173 ( \24488 , \24481 , \24486 , \24487 );
and \U$24174 ( \24489 , \24472 , \24488 );
and \U$24175 ( \24490 , \22235 , \22208 );
and \U$24176 ( \24491 , \22202 , \22206 );
nor \U$24177 ( \24492 , \24490 , \24491 );
xnor \U$24178 ( \24493 , \24492 , \22218 );
and \U$24179 ( \24494 , \22262 , \22230 );
and \U$24180 ( \24495 , \22224 , \22228 );
nor \U$24181 ( \24496 , \24494 , \24495 );
xnor \U$24182 ( \24497 , \24496 , \22240 );
and \U$24183 ( \24498 , \24493 , \24497 );
and \U$24184 ( \24499 , \22283 , \22257 );
and \U$24185 ( \24500 , \22251 , \22255 );
nor \U$24186 ( \24501 , \24499 , \24500 );
xnor \U$24187 ( \24502 , \24501 , \22267 );
and \U$24188 ( \24503 , \24497 , \24502 );
and \U$24189 ( \24504 , \24493 , \24502 );
or \U$24190 ( \24505 , \24498 , \24503 , \24504 );
and \U$24191 ( \24506 , \24488 , \24505 );
and \U$24192 ( \24507 , \24472 , \24505 );
or \U$24193 ( \24508 , \24489 , \24506 , \24507 );
and \U$24194 ( \24509 , \22305 , \22278 );
and \U$24195 ( \24510 , \22272 , \22276 );
nor \U$24196 ( \24511 , \24509 , \24510 );
xnor \U$24197 ( \24512 , \24511 , \22288 );
and \U$24198 ( \24513 , \22329 , \22300 );
and \U$24199 ( \24514 , \22294 , \22298 );
nor \U$24200 ( \24515 , \24513 , \24514 );
xnor \U$24201 ( \24516 , \24515 , \22310 );
and \U$24202 ( \24517 , \24512 , \24516 );
and \U$24203 ( \24518 , \22350 , \22324 );
and \U$24204 ( \24519 , \22318 , \22322 );
nor \U$24205 ( \24520 , \24518 , \24519 );
xnor \U$24206 ( \24521 , \24520 , \22334 );
and \U$24207 ( \24522 , \24516 , \24521 );
and \U$24208 ( \24523 , \24512 , \24521 );
or \U$24209 ( \24524 , \24517 , \24522 , \24523 );
and \U$24210 ( \24525 , \22372 , \22345 );
and \U$24211 ( \24526 , \22339 , \22343 );
nor \U$24212 ( \24527 , \24525 , \24526 );
xnor \U$24213 ( \24528 , \24527 , \22355 );
and \U$24214 ( \24529 , \22397 , \22367 );
and \U$24215 ( \24530 , \22361 , \22365 );
nor \U$24216 ( \24531 , \24529 , \24530 );
xnor \U$24217 ( \24532 , \24531 , \22377 );
and \U$24218 ( \24533 , \24528 , \24532 );
and \U$24219 ( \24534 , \22418 , \22392 );
and \U$24220 ( \24535 , \22386 , \22390 );
nor \U$24221 ( \24536 , \24534 , \24535 );
xnor \U$24222 ( \24537 , \24536 , \22402 );
and \U$24223 ( \24538 , \24532 , \24537 );
and \U$24224 ( \24539 , \24528 , \24537 );
or \U$24225 ( \24540 , \24533 , \24538 , \24539 );
and \U$24226 ( \24541 , \24524 , \24540 );
and \U$24227 ( \24542 , \22440 , \22413 );
and \U$24228 ( \24543 , \22407 , \22411 );
nor \U$24229 ( \24544 , \24542 , \24543 );
xnor \U$24230 ( \24545 , \24544 , \22423 );
and \U$24231 ( \24546 , \22468 , \22435 );
and \U$24232 ( \24547 , \22429 , \22433 );
nor \U$24233 ( \24548 , \24546 , \24547 );
xnor \U$24234 ( \24549 , \24548 , \22445 );
and \U$24235 ( \24550 , \24545 , \24549 );
and \U$24236 ( \24551 , \22489 , \22463 );
and \U$24237 ( \24552 , \22457 , \22461 );
nor \U$24238 ( \24553 , \24551 , \24552 );
xnor \U$24239 ( \24554 , \24553 , \22473 );
and \U$24240 ( \24555 , \24549 , \24554 );
and \U$24241 ( \24556 , \24545 , \24554 );
or \U$24242 ( \24557 , \24550 , \24555 , \24556 );
and \U$24243 ( \24558 , \24540 , \24557 );
and \U$24244 ( \24559 , \24524 , \24557 );
or \U$24245 ( \24560 , \24541 , \24558 , \24559 );
and \U$24246 ( \24561 , \24508 , \24560 );
and \U$24247 ( \24562 , \22511 , \22484 );
and \U$24248 ( \24563 , \22478 , \22482 );
nor \U$24249 ( \24564 , \24562 , \24563 );
xnor \U$24250 ( \24565 , \24564 , \22494 );
and \U$24251 ( \24566 , \22535 , \22506 );
and \U$24252 ( \24567 , \22500 , \22504 );
nor \U$24253 ( \24568 , \24566 , \24567 );
xnor \U$24254 ( \24569 , \24568 , \22516 );
and \U$24255 ( \24570 , \24565 , \24569 );
and \U$24256 ( \24571 , \22556 , \22530 );
and \U$24257 ( \24572 , \22524 , \22528 );
nor \U$24258 ( \24573 , \24571 , \24572 );
xnor \U$24259 ( \24574 , \24573 , \22540 );
and \U$24260 ( \24575 , \24569 , \24574 );
and \U$24261 ( \24576 , \24565 , \24574 );
or \U$24262 ( \24577 , \24570 , \24575 , \24576 );
and \U$24263 ( \24578 , \22578 , \22551 );
and \U$24264 ( \24579 , \22545 , \22549 );
nor \U$24265 ( \24580 , \24578 , \24579 );
xnor \U$24266 ( \24581 , \24580 , \22561 );
and \U$24267 ( \24582 , \22603 , \22573 );
and \U$24268 ( \24583 , \22567 , \22571 );
nor \U$24269 ( \24584 , \24582 , \24583 );
xnor \U$24270 ( \24585 , \24584 , \22583 );
and \U$24271 ( \24586 , \24581 , \24585 );
and \U$24272 ( \24587 , \22624 , \22598 );
and \U$24273 ( \24588 , \22592 , \22596 );
nor \U$24274 ( \24589 , \24587 , \24588 );
xnor \U$24275 ( \24590 , \24589 , \22608 );
and \U$24276 ( \24591 , \24585 , \24590 );
and \U$24277 ( \24592 , \24581 , \24590 );
or \U$24278 ( \24593 , \24586 , \24591 , \24592 );
and \U$24279 ( \24594 , \24577 , \24593 );
and \U$24280 ( \24595 , \22646 , \22619 );
and \U$24281 ( \24596 , \22613 , \22617 );
nor \U$24282 ( \24597 , \24595 , \24596 );
xnor \U$24283 ( \24598 , \24597 , \22629 );
and \U$24284 ( \24599 , \22676 , \22641 );
and \U$24285 ( \24600 , \22635 , \22639 );
nor \U$24286 ( \24601 , \24599 , \24600 );
xnor \U$24287 ( \24602 , \24601 , \22651 );
and \U$24288 ( \24603 , \24598 , \24602 );
and \U$24289 ( \24604 , \22696 , \22671 );
and \U$24290 ( \24605 , \22665 , \22669 );
nor \U$24291 ( \24606 , \24604 , \24605 );
xnor \U$24292 ( \24607 , \24606 , \22681 );
and \U$24293 ( \24608 , \24602 , \24607 );
and \U$24294 ( \24609 , \24598 , \24607 );
or \U$24295 ( \24610 , \24603 , \24608 , \24609 );
and \U$24296 ( \24611 , \24593 , \24610 );
and \U$24297 ( \24612 , \24577 , \24610 );
or \U$24298 ( \24613 , \24594 , \24611 , \24612 );
and \U$24299 ( \24614 , \24560 , \24613 );
and \U$24300 ( \24615 , \24508 , \24613 );
or \U$24301 ( \24616 , \24561 , \24614 , \24615 );
xor \U$24302 ( \24617 , \22682 , \22702 );
xor \U$24303 ( \24618 , \24617 , \22709 );
xor \U$24304 ( \24619 , \22609 , \22630 );
xor \U$24305 ( \24620 , \24619 , \22652 );
and \U$24306 ( \24621 , \24618 , \24620 );
xor \U$24307 ( \24622 , \22541 , \22562 );
xor \U$24308 ( \24623 , \24622 , \22584 );
and \U$24309 ( \24624 , \24620 , \24623 );
and \U$24310 ( \24625 , \24618 , \24623 );
or \U$24311 ( \24626 , \24621 , \24624 , \24625 );
xor \U$24312 ( \24627 , \22474 , \22495 );
xor \U$24313 ( \24628 , \24627 , \22517 );
xor \U$24314 ( \24629 , \22403 , \22424 );
xor \U$24315 ( \24630 , \24629 , \22446 );
and \U$24316 ( \24631 , \24628 , \24630 );
xor \U$24317 ( \24632 , \22335 , \22356 );
xor \U$24318 ( \24633 , \24632 , \22378 );
and \U$24319 ( \24634 , \24630 , \24633 );
and \U$24320 ( \24635 , \24628 , \24633 );
or \U$24321 ( \24636 , \24631 , \24634 , \24635 );
and \U$24322 ( \24637 , \24626 , \24636 );
xor \U$24323 ( \24638 , \22268 , \22289 );
xor \U$24324 ( \24639 , \24638 , \22311 );
xor \U$24325 ( \24640 , \22198 , \22219 );
xor \U$24326 ( \24641 , \24640 , \22241 );
and \U$24327 ( \24642 , \24639 , \24641 );
xor \U$24328 ( \24643 , \22130 , \22151 );
xor \U$24329 ( \24644 , \24643 , \22173 );
and \U$24330 ( \24645 , \24641 , \24644 );
and \U$24331 ( \24646 , \24639 , \24644 );
or \U$24332 ( \24647 , \24642 , \24645 , \24646 );
and \U$24333 ( \24648 , \24636 , \24647 );
and \U$24334 ( \24649 , \24626 , \24647 );
or \U$24335 ( \24650 , \24637 , \24648 , \24649 );
and \U$24336 ( \24651 , \24616 , \24650 );
xor \U$24337 ( \24652 , \22838 , \22852 );
xor \U$24338 ( \24653 , \24652 , \22871 );
xor \U$24339 ( \24654 , \22788 , \22802 );
xor \U$24340 ( \24655 , \24654 , \22817 );
and \U$24341 ( \24656 , \24653 , \24655 );
xor \U$24342 ( \24657 , \22741 , \22755 );
xor \U$24343 ( \24658 , \24657 , \22770 );
and \U$24344 ( \24659 , \24655 , \24658 );
and \U$24345 ( \24660 , \24653 , \24658 );
or \U$24346 ( \24661 , \24656 , \24659 , \24660 );
and \U$24347 ( \24662 , \24650 , \24661 );
and \U$24348 ( \24663 , \24616 , \24661 );
or \U$24349 ( \24664 , \24651 , \24662 , \24663 );
xor \U$24350 ( \24665 , \22712 , \22716 );
xor \U$24351 ( \24666 , \24665 , \22724 );
xor \U$24352 ( \24667 , \22520 , \22587 );
xor \U$24353 ( \24668 , \24667 , \22655 );
and \U$24354 ( \24669 , \24666 , \24668 );
xor \U$24355 ( \24670 , \22314 , \22381 );
xor \U$24356 ( \24671 , \24670 , \22449 );
and \U$24357 ( \24672 , \24668 , \24671 );
and \U$24358 ( \24673 , \24666 , \24671 );
or \U$24359 ( \24674 , \24669 , \24672 , \24673 );
xor \U$24360 ( \24675 , \23048 , \23062 );
xor \U$24361 ( \24676 , \24675 , \23077 );
and \U$24362 ( \24677 , \24674 , \24676 );
xor \U$24363 ( \24678 , \22953 , \22997 );
xor \U$24364 ( \24679 , \24678 , \23031 );
and \U$24365 ( \24680 , \24676 , \24679 );
and \U$24366 ( \24681 , \24674 , \24679 );
or \U$24367 ( \24682 , \24677 , \24680 , \24681 );
and \U$24368 ( \24683 , \24664 , \24682 );
xor \U$24369 ( \24684 , \22874 , \22888 );
xor \U$24370 ( \24685 , \24684 , \22903 );
xor \U$24371 ( \24686 , \22727 , \22773 );
xor \U$24372 ( \24687 , \24686 , \22820 );
and \U$24373 ( \24688 , \24685 , \24687 );
xor \U$24374 ( \24689 , \22247 , \22452 );
xor \U$24375 ( \24690 , \24689 , \22658 );
and \U$24376 ( \24691 , \24687 , \24690 );
and \U$24377 ( \24692 , \24685 , \24690 );
or \U$24378 ( \24693 , \24688 , \24691 , \24692 );
and \U$24379 ( \24694 , \24682 , \24693 );
and \U$24380 ( \24695 , \24664 , \24693 );
or \U$24381 ( \24696 , \24683 , \24694 , \24695 );
xor \U$24382 ( \24697 , \23557 , \23561 );
xor \U$24383 ( \24698 , \24697 , \23566 );
xor \U$24384 ( \24699 , \23541 , \23545 );
xor \U$24385 ( \24700 , \24699 , \23550 );
and \U$24386 ( \24701 , \24698 , \24700 );
xor \U$24387 ( \24702 , \23113 , \23210 );
xor \U$24388 ( \24703 , \24702 , \23289 );
and \U$24389 ( \24704 , \24700 , \24703 );
and \U$24390 ( \24705 , \24698 , \24703 );
or \U$24391 ( \24706 , \24701 , \24704 , \24705 );
and \U$24392 ( \24707 , \24696 , \24706 );
xor \U$24393 ( \24708 , \23459 , \23536 );
xor \U$24394 ( \24709 , \24708 , \23575 );
and \U$24395 ( \24710 , \24706 , \24709 );
and \U$24396 ( \24711 , \24696 , \24709 );
or \U$24397 ( \24712 , \24707 , \24710 , \24711 );
xor \U$24398 ( \24713 , \24106 , \24110 );
xor \U$24399 ( \24714 , \24713 , \24115 );
and \U$24400 ( \24715 , \24712 , \24714 );
xor \U$24401 ( \24716 , \23295 , \23578 );
xor \U$24402 ( \24717 , \24716 , \23840 );
and \U$24403 ( \24718 , \24714 , \24717 );
and \U$24404 ( \24719 , \24712 , \24717 );
or \U$24405 ( \24720 , \24715 , \24718 , \24719 );
xor \U$24406 ( \24721 , \23843 , \24101 );
xor \U$24407 ( \24722 , \24721 , \24148 );
and \U$24408 ( \24723 , \24720 , \24722 );
nor \U$24409 ( \24724 , \24456 , \24723 );
and \U$24410 ( \24725 , \24435 , \24439 );
and \U$24411 ( \24726 , \24439 , \24454 );
and \U$24412 ( \24727 , \24435 , \24454 );
or \U$24413 ( \24728 , \24725 , \24726 , \24727 );
and \U$24414 ( \24729 , \24155 , \24159 );
and \U$24415 ( \24730 , \24159 , \24429 );
and \U$24416 ( \24731 , \24155 , \24429 );
or \U$24417 ( \24732 , \24729 , \24730 , \24731 );
and \U$24418 ( \24733 , \24258 , \24262 );
and \U$24419 ( \24734 , \24262 , \24267 );
and \U$24420 ( \24735 , \24258 , \24267 );
or \U$24421 ( \24736 , \24733 , \24734 , \24735 );
and \U$24422 ( \24737 , \24243 , \24247 );
and \U$24423 ( \24738 , \24247 , \24252 );
and \U$24424 ( \24739 , \24243 , \24252 );
or \U$24425 ( \24740 , \24737 , \24738 , \24739 );
xor \U$24426 ( \24741 , \24736 , \24740 );
and \U$24427 ( \24742 , \24164 , \24193 );
and \U$24428 ( \24743 , \24193 , \24238 );
and \U$24429 ( \24744 , \24164 , \24238 );
or \U$24430 ( \24745 , \24742 , \24743 , \24744 );
xor \U$24431 ( \24746 , \24741 , \24745 );
and \U$24432 ( \24747 , \24401 , \24405 );
and \U$24433 ( \24748 , \24405 , \24410 );
and \U$24434 ( \24749 , \24401 , \24410 );
or \U$24435 ( \24750 , \24747 , \24748 , \24749 );
and \U$24436 ( \24751 , \24366 , \24380 );
and \U$24437 ( \24752 , \24380 , \24395 );
and \U$24438 ( \24753 , \24366 , \24395 );
or \U$24439 ( \24754 , \24751 , \24752 , \24753 );
xor \U$24440 ( \24755 , \24750 , \24754 );
and \U$24441 ( \24756 , \24332 , \24346 );
and \U$24442 ( \24757 , \24346 , \24361 );
and \U$24443 ( \24758 , \24332 , \24361 );
or \U$24444 ( \24759 , \24756 , \24757 , \24758 );
xor \U$24445 ( \24760 , \24755 , \24759 );
and \U$24446 ( \24761 , \24306 , \24310 );
and \U$24447 ( \24762 , \24310 , \24315 );
and \U$24448 ( \24763 , \24306 , \24315 );
or \U$24449 ( \24764 , \24761 , \24762 , \24763 );
and \U$24450 ( \24765 , \24291 , \24295 );
and \U$24451 ( \24766 , \24295 , \24300 );
and \U$24452 ( \24767 , \24291 , \24300 );
or \U$24453 ( \24768 , \24765 , \24766 , \24767 );
xor \U$24454 ( \24769 , \24764 , \24768 );
and \U$24455 ( \24770 , \24277 , \24281 );
and \U$24456 ( \24771 , \24281 , \24286 );
and \U$24457 ( \24772 , \24277 , \24286 );
or \U$24458 ( \24773 , \24770 , \24771 , \24772 );
xor \U$24459 ( \24774 , \24769 , \24773 );
xor \U$24460 ( \24775 , \24760 , \24774 );
and \U$24461 ( \24776 , \24370 , \24374 );
and \U$24462 ( \24777 , \24374 , \24379 );
and \U$24463 ( \24778 , \24370 , \24379 );
or \U$24464 ( \24779 , \24776 , \24777 , \24778 );
nand \U$24465 ( \24780 , \22706 , \21978 );
not \U$24466 ( \24781 , \24780 );
xor \U$24467 ( \24782 , \24779 , \24781 );
and \U$24468 ( \24783 , \22635 , \23173 );
and \U$24469 ( \24784 , \22646 , \22999 );
nor \U$24470 ( \24785 , \24783 , \24784 );
xnor \U$24471 ( \24786 , \24785 , \22016 );
and \U$24472 ( \24787 , \22665 , \22021 );
and \U$24473 ( \24788 , \22676 , \22019 );
nor \U$24474 ( \24789 , \24787 , \24788 );
xnor \U$24475 ( \24790 , \24789 , \21595 );
xor \U$24476 ( \24791 , \24786 , \24790 );
and \U$24477 ( \24792 , \22686 , \21983 );
and \U$24478 ( \24793 , \22696 , \21981 );
nor \U$24479 ( \24794 , \24792 , \24793 );
xnor \U$24480 ( \24795 , \24794 , \21995 );
xor \U$24481 ( \24796 , \24791 , \24795 );
xor \U$24482 ( \24797 , \24782 , \24796 );
and \U$24483 ( \24798 , \24336 , \24340 );
and \U$24484 ( \24799 , \24340 , \24345 );
and \U$24485 ( \24800 , \24336 , \24345 );
or \U$24486 ( \24801 , \24798 , \24799 , \24800 );
and \U$24487 ( \24802 , \24322 , \24326 );
and \U$24488 ( \24803 , \24326 , \24331 );
and \U$24489 ( \24804 , \24322 , \24331 );
or \U$24490 ( \24805 , \24802 , \24803 , \24804 );
xor \U$24491 ( \24806 , \24801 , \24805 );
and \U$24492 ( \24807 , \24385 , \24389 );
and \U$24493 ( \24808 , \24389 , \24394 );
and \U$24494 ( \24809 , \24385 , \24394 );
or \U$24495 ( \24810 , \24807 , \24808 , \24809 );
xor \U$24496 ( \24811 , \24806 , \24810 );
xor \U$24497 ( \24812 , \24797 , \24811 );
and \U$24498 ( \24813 , \24212 , \24216 );
and \U$24499 ( \24814 , \24216 , \24221 );
and \U$24500 ( \24815 , \24212 , \24221 );
or \U$24501 ( \24816 , \24813 , \24814 , \24815 );
and \U$24502 ( \24817 , \24198 , \24202 );
and \U$24503 ( \24818 , \24202 , \24207 );
and \U$24504 ( \24819 , \24198 , \24207 );
or \U$24505 ( \24820 , \24817 , \24818 , \24819 );
xor \U$24506 ( \24821 , \24816 , \24820 );
and \U$24507 ( \24822 , \24351 , \24355 );
and \U$24508 ( \24823 , \24355 , \24360 );
and \U$24509 ( \24824 , \24351 , \24360 );
or \U$24510 ( \24825 , \24822 , \24823 , \24824 );
xor \U$24511 ( \24826 , \24821 , \24825 );
xor \U$24512 ( \24827 , \24812 , \24826 );
and \U$24513 ( \24828 , \22156 , \22257 );
and \U$24514 ( \24829 , \22167 , \22255 );
nor \U$24515 ( \24830 , \24828 , \24829 );
xnor \U$24516 ( \24831 , \24830 , \22267 );
and \U$24517 ( \24832 , \22181 , \22278 );
and \U$24518 ( \24833 , \22192 , \22276 );
nor \U$24519 ( \24834 , \24832 , \24833 );
xnor \U$24520 ( \24835 , \24834 , \22288 );
xor \U$24521 ( \24836 , \24831 , \24835 );
and \U$24522 ( \24837 , \22202 , \22300 );
and \U$24523 ( \24838 , \22213 , \22298 );
nor \U$24524 ( \24839 , \24837 , \24838 );
xnor \U$24525 ( \24840 , \24839 , \22310 );
xor \U$24526 ( \24841 , \24836 , \24840 );
and \U$24527 ( \24842 , \22089 , \22187 );
and \U$24528 ( \24843 , \22100 , \22185 );
nor \U$24529 ( \24844 , \24842 , \24843 );
xnor \U$24530 ( \24845 , \24844 , \22197 );
and \U$24531 ( \24846 , \22113 , \22208 );
and \U$24532 ( \24847 , \22124 , \22206 );
nor \U$24533 ( \24848 , \24846 , \24847 );
xnor \U$24534 ( \24849 , \24848 , \22218 );
xor \U$24535 ( \24850 , \24845 , \24849 );
and \U$24536 ( \24851 , \22134 , \22230 );
and \U$24537 ( \24852 , \22145 , \22228 );
nor \U$24538 ( \24853 , \24851 , \24852 );
xnor \U$24539 ( \24854 , \24853 , \22240 );
xor \U$24540 ( \24855 , \24850 , \24854 );
xor \U$24541 ( \24856 , \24841 , \24855 );
and \U$24542 ( \24857 , \23230 , \22119 );
and \U$24543 ( \24858 , \23329 , \22117 );
nor \U$24544 ( \24859 , \24857 , \24858 );
xnor \U$24545 ( \24860 , \24859 , \22129 );
and \U$24546 ( \24861 , \22858 , \22140 );
and \U$24547 ( \24862 , \22894 , \22138 );
nor \U$24548 ( \24863 , \24861 , \24862 );
xnor \U$24549 ( \24864 , \24863 , \22150 );
xor \U$24550 ( \24865 , \24860 , \24864 );
and \U$24551 ( \24866 , \22071 , \22162 );
and \U$24552 ( \24867 , \22081 , \22160 );
nor \U$24553 ( \24868 , \24866 , \24867 );
xnor \U$24554 ( \24869 , \24868 , \22172 );
xor \U$24555 ( \24870 , \24865 , \24869 );
xor \U$24556 ( \24871 , \24856 , \24870 );
and \U$24557 ( \24872 , \22361 , \22463 );
and \U$24558 ( \24873 , \22372 , \22461 );
nor \U$24559 ( \24874 , \24872 , \24873 );
xnor \U$24560 ( \24875 , \24874 , \22473 );
and \U$24561 ( \24876 , \22386 , \22484 );
and \U$24562 ( \24877 , \22397 , \22482 );
nor \U$24563 ( \24878 , \24876 , \24877 );
xnor \U$24564 ( \24879 , \24878 , \22494 );
xor \U$24565 ( \24880 , \24875 , \24879 );
and \U$24566 ( \24881 , \22407 , \22506 );
and \U$24567 ( \24882 , \22418 , \22504 );
nor \U$24568 ( \24883 , \24881 , \24882 );
xnor \U$24569 ( \24884 , \24883 , \22516 );
xor \U$24570 ( \24885 , \24880 , \24884 );
and \U$24571 ( \24886 , \22294 , \22392 );
and \U$24572 ( \24887 , \22305 , \22390 );
nor \U$24573 ( \24888 , \24886 , \24887 );
xnor \U$24574 ( \24889 , \24888 , \22402 );
and \U$24575 ( \24890 , \22318 , \22413 );
and \U$24576 ( \24891 , \22329 , \22411 );
nor \U$24577 ( \24892 , \24890 , \24891 );
xnor \U$24578 ( \24893 , \24892 , \22423 );
xor \U$24579 ( \24894 , \24889 , \24893 );
and \U$24580 ( \24895 , \22339 , \22435 );
and \U$24581 ( \24896 , \22350 , \22433 );
nor \U$24582 ( \24897 , \24895 , \24896 );
xnor \U$24583 ( \24898 , \24897 , \22445 );
xor \U$24584 ( \24899 , \24894 , \24898 );
xor \U$24585 ( \24900 , \24885 , \24899 );
and \U$24586 ( \24901 , \22224 , \22324 );
and \U$24587 ( \24902 , \22235 , \22322 );
nor \U$24588 ( \24903 , \24901 , \24902 );
xnor \U$24589 ( \24904 , \24903 , \22334 );
and \U$24590 ( \24905 , \22251 , \22345 );
and \U$24591 ( \24906 , \22262 , \22343 );
nor \U$24592 ( \24907 , \24905 , \24906 );
xnor \U$24593 ( \24908 , \24907 , \22355 );
xor \U$24594 ( \24909 , \24904 , \24908 );
and \U$24595 ( \24910 , \22272 , \22367 );
and \U$24596 ( \24911 , \22283 , \22365 );
nor \U$24597 ( \24912 , \24910 , \24911 );
xnor \U$24598 ( \24913 , \24912 , \22377 );
xor \U$24599 ( \24914 , \24909 , \24913 );
xor \U$24600 ( \24915 , \24900 , \24914 );
xor \U$24601 ( \24916 , \24871 , \24915 );
and \U$24602 ( \24917 , \22567 , \22671 );
and \U$24603 ( \24918 , \22578 , \22669 );
nor \U$24604 ( \24919 , \24917 , \24918 );
xnor \U$24605 ( \24920 , \24919 , \22681 );
and \U$24606 ( \24921 , \22592 , \22691 );
and \U$24607 ( \24922 , \22603 , \22689 );
nor \U$24608 ( \24923 , \24921 , \24922 );
xnor \U$24609 ( \24924 , \24923 , \22701 );
xor \U$24610 ( \24925 , \24920 , \24924 );
and \U$24611 ( \24926 , \22613 , \22720 );
and \U$24612 ( \24927 , \22624 , \22707 );
nor \U$24613 ( \24928 , \24926 , \24927 );
xnor \U$24614 ( \24929 , \24928 , \22067 );
xor \U$24615 ( \24930 , \24925 , \24929 );
and \U$24616 ( \24931 , \22500 , \22598 );
and \U$24617 ( \24932 , \22511 , \22596 );
nor \U$24618 ( \24933 , \24931 , \24932 );
xnor \U$24619 ( \24934 , \24933 , \22608 );
and \U$24620 ( \24935 , \22524 , \22619 );
and \U$24621 ( \24936 , \22535 , \22617 );
nor \U$24622 ( \24937 , \24935 , \24936 );
xnor \U$24623 ( \24938 , \24937 , \22629 );
xor \U$24624 ( \24939 , \24934 , \24938 );
and \U$24625 ( \24940 , \22545 , \22641 );
and \U$24626 ( \24941 , \22556 , \22639 );
nor \U$24627 ( \24942 , \24940 , \24941 );
xnor \U$24628 ( \24943 , \24942 , \22651 );
xor \U$24629 ( \24944 , \24939 , \24943 );
xor \U$24630 ( \24945 , \24930 , \24944 );
and \U$24631 ( \24946 , \22429 , \22530 );
and \U$24632 ( \24947 , \22440 , \22528 );
nor \U$24633 ( \24948 , \24946 , \24947 );
xnor \U$24634 ( \24949 , \24948 , \22540 );
and \U$24635 ( \24950 , \22457 , \22551 );
and \U$24636 ( \24951 , \22468 , \22549 );
nor \U$24637 ( \24952 , \24950 , \24951 );
xnor \U$24638 ( \24953 , \24952 , \22561 );
xor \U$24639 ( \24954 , \24949 , \24953 );
and \U$24640 ( \24955 , \22478 , \22573 );
and \U$24641 ( \24956 , \22489 , \22571 );
nor \U$24642 ( \24957 , \24955 , \24956 );
xnor \U$24643 ( \24958 , \24957 , \22583 );
xor \U$24644 ( \24959 , \24954 , \24958 );
xor \U$24645 ( \24960 , \24945 , \24959 );
xor \U$24646 ( \24961 , \24916 , \24960 );
xor \U$24647 ( \24962 , \24827 , \24961 );
and \U$24648 ( \24963 , \24208 , \24222 );
and \U$24649 ( \24964 , \24222 , \24237 );
and \U$24650 ( \24965 , \24208 , \24237 );
or \U$24651 ( \24966 , \24963 , \24964 , \24965 );
and \U$24652 ( \24967 , \24178 , \24192 );
xor \U$24653 ( \24968 , \24966 , \24967 );
and \U$24654 ( \24969 , \21977 , \22076 );
and \U$24655 ( \24970 , \21990 , \22073 );
nor \U$24656 ( \24971 , \24969 , \24970 );
xnor \U$24657 ( \24972 , \24971 , \22072 );
and \U$24658 ( \24973 , \22030 , \22095 );
and \U$24659 ( \24974 , \22001 , \22093 );
nor \U$24660 ( \24975 , \24973 , \24974 );
xnor \U$24661 ( \24976 , \24975 , \22105 );
xor \U$24662 ( \24977 , \24972 , \24976 );
xor \U$24663 ( \24978 , \24968 , \24977 );
xor \U$24664 ( \24979 , \24962 , \24978 );
xor \U$24665 ( \24980 , \24775 , \24979 );
xor \U$24666 ( \24981 , \24746 , \24980 );
and \U$24667 ( \24982 , \24418 , \24422 );
and \U$24668 ( \24983 , \24422 , \24427 );
and \U$24669 ( \24984 , \24418 , \24427 );
or \U$24670 ( \24985 , \24982 , \24983 , \24984 );
and \U$24671 ( \24986 , \24273 , \24317 );
and \U$24672 ( \24987 , \24317 , \24412 );
and \U$24673 ( \24988 , \24273 , \24412 );
or \U$24674 ( \24989 , \24986 , \24987 , \24988 );
xor \U$24675 ( \24990 , \24985 , \24989 );
and \U$24676 ( \24991 , \24239 , \24253 );
and \U$24677 ( \24992 , \24253 , \24268 );
and \U$24678 ( \24993 , \24239 , \24268 );
or \U$24679 ( \24994 , \24991 , \24992 , \24993 );
xor \U$24680 ( \24995 , \24990 , \24994 );
xor \U$24681 ( \24996 , \24981 , \24995 );
xor \U$24682 ( \24997 , \24732 , \24996 );
and \U$24683 ( \24998 , \24444 , \24448 );
and \U$24684 ( \24999 , \24448 , \24453 );
and \U$24685 ( \25000 , \24444 , \24453 );
or \U$24686 ( \25001 , \24998 , \24999 , \25000 );
and \U$24687 ( \25002 , \24269 , \24413 );
and \U$24688 ( \25003 , \24413 , \24428 );
and \U$24689 ( \25004 , \24269 , \24428 );
or \U$24690 ( \25005 , \25002 , \25003 , \25004 );
xor \U$24691 ( \25006 , \25001 , \25005 );
and \U$24692 ( \25007 , \24362 , \24396 );
and \U$24693 ( \25008 , \24396 , \24411 );
and \U$24694 ( \25009 , \24362 , \24411 );
or \U$24695 ( \25010 , \25007 , \25008 , \25009 );
and \U$24696 ( \25011 , \24287 , \24301 );
and \U$24697 ( \25012 , \24301 , \24316 );
and \U$24698 ( \25013 , \24287 , \24316 );
or \U$24699 ( \25014 , \25011 , \25012 , \25013 );
xor \U$24700 ( \25015 , \25010 , \25014 );
and \U$24701 ( \25016 , \24182 , \24186 );
and \U$24702 ( \25017 , \24186 , \24191 );
and \U$24703 ( \25018 , \24182 , \24191 );
or \U$24704 ( \25019 , \25016 , \25017 , \25018 );
and \U$24705 ( \25020 , \24168 , \24172 );
and \U$24706 ( \25021 , \24172 , \24177 );
and \U$24707 ( \25022 , \24168 , \24177 );
or \U$24708 ( \25023 , \25020 , \25021 , \25022 );
xor \U$24709 ( \25024 , \25019 , \25023 );
and \U$24710 ( \25025 , \24227 , \24231 );
and \U$24711 ( \25026 , \24231 , \24236 );
and \U$24712 ( \25027 , \24227 , \24236 );
or \U$24713 ( \25028 , \25025 , \25026 , \25027 );
xor \U$24714 ( \25029 , \25024 , \25028 );
xor \U$24715 ( \25030 , \25015 , \25029 );
xor \U$24716 ( \25031 , \25006 , \25030 );
xor \U$24717 ( \25032 , \24997 , \25031 );
xor \U$24718 ( \25033 , \24728 , \25032 );
and \U$24719 ( \25034 , \24151 , \24430 );
and \U$24720 ( \25035 , \24430 , \24455 );
and \U$24721 ( \25036 , \24151 , \24455 );
or \U$24722 ( \25037 , \25034 , \25035 , \25036 );
nor \U$24723 ( \25038 , \25033 , \25037 );
nor \U$24724 ( \25039 , \24724 , \25038 );
and \U$24725 ( \25040 , \24732 , \24996 );
and \U$24726 ( \25041 , \24996 , \25031 );
and \U$24727 ( \25042 , \24732 , \25031 );
or \U$24728 ( \25043 , \25040 , \25041 , \25042 );
and \U$24729 ( \25044 , \24736 , \24740 );
and \U$24730 ( \25045 , \24740 , \24745 );
and \U$24731 ( \25046 , \24736 , \24745 );
or \U$24732 ( \25047 , \25044 , \25045 , \25046 );
and \U$24733 ( \25048 , \25010 , \25014 );
and \U$24734 ( \25049 , \25014 , \25029 );
and \U$24735 ( \25050 , \25010 , \25029 );
or \U$24736 ( \25051 , \25048 , \25049 , \25050 );
xor \U$24737 ( \25052 , \25047 , \25051 );
and \U$24738 ( \25053 , \24827 , \24961 );
and \U$24739 ( \25054 , \24961 , \24978 );
and \U$24740 ( \25055 , \24827 , \24978 );
or \U$24741 ( \25056 , \25053 , \25054 , \25055 );
xor \U$24742 ( \25057 , \25052 , \25056 );
and \U$24743 ( \25058 , \24985 , \24989 );
and \U$24744 ( \25059 , \24989 , \24994 );
and \U$24745 ( \25060 , \24985 , \24994 );
or \U$24746 ( \25061 , \25058 , \25059 , \25060 );
and \U$24747 ( \25062 , \24760 , \24774 );
and \U$24748 ( \25063 , \24774 , \24979 );
and \U$24749 ( \25064 , \24760 , \24979 );
or \U$24750 ( \25065 , \25062 , \25063 , \25064 );
xor \U$24751 ( \25066 , \25061 , \25065 );
and \U$24752 ( \25067 , \24764 , \24768 );
and \U$24753 ( \25068 , \24768 , \24773 );
and \U$24754 ( \25069 , \24764 , \24773 );
or \U$24755 ( \25070 , \25067 , \25068 , \25069 );
and \U$24756 ( \25071 , \24750 , \24754 );
and \U$24757 ( \25072 , \24754 , \24759 );
and \U$24758 ( \25073 , \24750 , \24759 );
or \U$24759 ( \25074 , \25071 , \25072 , \25073 );
xor \U$24760 ( \25075 , \25070 , \25074 );
and \U$24761 ( \25076 , \24966 , \24967 );
and \U$24762 ( \25077 , \24967 , \24977 );
and \U$24763 ( \25078 , \24966 , \24977 );
or \U$24764 ( \25079 , \25076 , \25077 , \25078 );
xor \U$24765 ( \25080 , \25075 , \25079 );
xor \U$24766 ( \25081 , \25066 , \25080 );
xor \U$24767 ( \25082 , \25057 , \25081 );
xor \U$24768 ( \25083 , \25043 , \25082 );
and \U$24769 ( \25084 , \25001 , \25005 );
and \U$24770 ( \25085 , \25005 , \25030 );
and \U$24771 ( \25086 , \25001 , \25030 );
or \U$24772 ( \25087 , \25084 , \25085 , \25086 );
and \U$24773 ( \25088 , \24746 , \24980 );
and \U$24774 ( \25089 , \24980 , \24995 );
and \U$24775 ( \25090 , \24746 , \24995 );
or \U$24776 ( \25091 , \25088 , \25089 , \25090 );
xor \U$24777 ( \25092 , \25087 , \25091 );
and \U$24778 ( \25093 , \25019 , \25023 );
and \U$24779 ( \25094 , \25023 , \25028 );
and \U$24780 ( \25095 , \25019 , \25028 );
or \U$24781 ( \25096 , \25093 , \25094 , \25095 );
and \U$24782 ( \25097 , \24816 , \24820 );
and \U$24783 ( \25098 , \24820 , \24825 );
and \U$24784 ( \25099 , \24816 , \24825 );
or \U$24785 ( \25100 , \25097 , \25098 , \25099 );
xor \U$24786 ( \25101 , \25096 , \25100 );
and \U$24787 ( \25102 , \24801 , \24805 );
and \U$24788 ( \25103 , \24805 , \24810 );
and \U$24789 ( \25104 , \24801 , \24810 );
or \U$24790 ( \25105 , \25102 , \25103 , \25104 );
xor \U$24791 ( \25106 , \25101 , \25105 );
and \U$24792 ( \25107 , \22397 , \22484 );
and \U$24793 ( \25108 , \22361 , \22482 );
nor \U$24794 ( \25109 , \25107 , \25108 );
xnor \U$24795 ( \25110 , \25109 , \22494 );
and \U$24796 ( \25111 , \22418 , \22506 );
and \U$24797 ( \25112 , \22386 , \22504 );
nor \U$24798 ( \25113 , \25111 , \25112 );
xnor \U$24799 ( \25114 , \25113 , \22516 );
xor \U$24800 ( \25115 , \25110 , \25114 );
and \U$24801 ( \25116 , \22440 , \22530 );
and \U$24802 ( \25117 , \22407 , \22528 );
nor \U$24803 ( \25118 , \25116 , \25117 );
xnor \U$24804 ( \25119 , \25118 , \22540 );
xor \U$24805 ( \25120 , \25115 , \25119 );
and \U$24806 ( \25121 , \22329 , \22413 );
and \U$24807 ( \25122 , \22294 , \22411 );
nor \U$24808 ( \25123 , \25121 , \25122 );
xnor \U$24809 ( \25124 , \25123 , \22423 );
and \U$24810 ( \25125 , \22350 , \22435 );
and \U$24811 ( \25126 , \22318 , \22433 );
nor \U$24812 ( \25127 , \25125 , \25126 );
xnor \U$24813 ( \25128 , \25127 , \22445 );
xor \U$24814 ( \25129 , \25124 , \25128 );
and \U$24815 ( \25130 , \22372 , \22463 );
and \U$24816 ( \25131 , \22339 , \22461 );
nor \U$24817 ( \25132 , \25130 , \25131 );
xnor \U$24818 ( \25133 , \25132 , \22473 );
xor \U$24819 ( \25134 , \25129 , \25133 );
xor \U$24820 ( \25135 , \25120 , \25134 );
and \U$24821 ( \25136 , \22262 , \22345 );
and \U$24822 ( \25137 , \22224 , \22343 );
nor \U$24823 ( \25138 , \25136 , \25137 );
xnor \U$24824 ( \25139 , \25138 , \22355 );
and \U$24825 ( \25140 , \22283 , \22367 );
and \U$24826 ( \25141 , \22251 , \22365 );
nor \U$24827 ( \25142 , \25140 , \25141 );
xnor \U$24828 ( \25143 , \25142 , \22377 );
xor \U$24829 ( \25144 , \25139 , \25143 );
and \U$24830 ( \25145 , \22305 , \22392 );
and \U$24831 ( \25146 , \22272 , \22390 );
nor \U$24832 ( \25147 , \25145 , \25146 );
xnor \U$24833 ( \25148 , \25147 , \22402 );
xor \U$24834 ( \25149 , \25144 , \25148 );
xor \U$24835 ( \25150 , \25135 , \25149 );
and \U$24836 ( \25151 , \22603 , \22691 );
and \U$24837 ( \25152 , \22567 , \22689 );
nor \U$24838 ( \25153 , \25151 , \25152 );
xnor \U$24839 ( \25154 , \25153 , \22701 );
and \U$24840 ( \25155 , \22624 , \22720 );
and \U$24841 ( \25156 , \22592 , \22707 );
nor \U$24842 ( \25157 , \25155 , \25156 );
xnor \U$24843 ( \25158 , \25157 , \22067 );
xor \U$24844 ( \25159 , \25154 , \25158 );
and \U$24845 ( \25160 , \22646 , \23173 );
and \U$24846 ( \25161 , \22613 , \22999 );
nor \U$24847 ( \25162 , \25160 , \25161 );
xnor \U$24848 ( \25163 , \25162 , \22016 );
xor \U$24849 ( \25164 , \25159 , \25163 );
and \U$24850 ( \25165 , \22535 , \22619 );
and \U$24851 ( \25166 , \22500 , \22617 );
nor \U$24852 ( \25167 , \25165 , \25166 );
xnor \U$24853 ( \25168 , \25167 , \22629 );
and \U$24854 ( \25169 , \22556 , \22641 );
and \U$24855 ( \25170 , \22524 , \22639 );
nor \U$24856 ( \25171 , \25169 , \25170 );
xnor \U$24857 ( \25172 , \25171 , \22651 );
xor \U$24858 ( \25173 , \25168 , \25172 );
and \U$24859 ( \25174 , \22578 , \22671 );
and \U$24860 ( \25175 , \22545 , \22669 );
nor \U$24861 ( \25176 , \25174 , \25175 );
xnor \U$24862 ( \25177 , \25176 , \22681 );
xor \U$24863 ( \25178 , \25173 , \25177 );
xor \U$24864 ( \25179 , \25164 , \25178 );
and \U$24865 ( \25180 , \22468 , \22551 );
and \U$24866 ( \25181 , \22429 , \22549 );
nor \U$24867 ( \25182 , \25180 , \25181 );
xnor \U$24868 ( \25183 , \25182 , \22561 );
and \U$24869 ( \25184 , \22489 , \22573 );
and \U$24870 ( \25185 , \22457 , \22571 );
nor \U$24871 ( \25186 , \25184 , \25185 );
xnor \U$24872 ( \25187 , \25186 , \22583 );
xor \U$24873 ( \25188 , \25183 , \25187 );
and \U$24874 ( \25189 , \22511 , \22598 );
and \U$24875 ( \25190 , \22478 , \22596 );
nor \U$24876 ( \25191 , \25189 , \25190 );
xnor \U$24877 ( \25192 , \25191 , \22608 );
xor \U$24878 ( \25193 , \25188 , \25192 );
xor \U$24879 ( \25194 , \25179 , \25193 );
xor \U$24880 ( \25195 , \25150 , \25194 );
and \U$24881 ( \25196 , \24920 , \24924 );
and \U$24882 ( \25197 , \24924 , \24929 );
and \U$24883 ( \25198 , \24920 , \24929 );
or \U$24884 ( \25199 , \25196 , \25197 , \25198 );
and \U$24885 ( \25200 , \24786 , \24790 );
and \U$24886 ( \25201 , \24790 , \24795 );
and \U$24887 ( \25202 , \24786 , \24795 );
or \U$24888 ( \25203 , \25200 , \25201 , \25202 );
xor \U$24889 ( \25204 , \25199 , \25203 );
and \U$24890 ( \25205 , \22676 , \22021 );
and \U$24891 ( \25206 , \22635 , \22019 );
nor \U$24892 ( \25207 , \25205 , \25206 );
xnor \U$24893 ( \25208 , \25207 , \21595 );
and \U$24894 ( \25209 , \22696 , \21983 );
and \U$24895 ( \25210 , \22665 , \21981 );
nor \U$24896 ( \25211 , \25209 , \25210 );
xnor \U$24897 ( \25212 , \25211 , \21995 );
xor \U$24898 ( \25213 , \25208 , \25212 );
and \U$24899 ( \25214 , \22686 , \21978 );
xor \U$24900 ( \25215 , \25213 , \25214 );
xor \U$24901 ( \25216 , \25204 , \25215 );
xor \U$24902 ( \25217 , \25195 , \25216 );
and \U$24903 ( \25218 , \24841 , \24855 );
and \U$24904 ( \25219 , \24855 , \24870 );
and \U$24905 ( \25220 , \24841 , \24870 );
or \U$24906 ( \25221 , \25218 , \25219 , \25220 );
and \U$24907 ( \25222 , \21990 , \22076 );
not \U$24908 ( \25223 , \25222 );
xnor \U$24909 ( \25224 , \25223 , \22072 );
and \U$24910 ( \25225 , \22001 , \22095 );
and \U$24911 ( \25226 , \21977 , \22093 );
nor \U$24912 ( \25227 , \25225 , \25226 );
xnor \U$24913 ( \25228 , \25227 , \22105 );
xor \U$24914 ( \25229 , \25224 , \25228 );
and \U$24915 ( \25230 , \23329 , \22119 );
and \U$24916 ( \25231 , \22030 , \22117 );
nor \U$24917 ( \25232 , \25230 , \25231 );
xnor \U$24918 ( \25233 , \25232 , \22129 );
xor \U$24919 ( \25234 , \25229 , \25233 );
xor \U$24920 ( \25235 , \25221 , \25234 );
and \U$24921 ( \25236 , \22192 , \22278 );
and \U$24922 ( \25237 , \22156 , \22276 );
nor \U$24923 ( \25238 , \25236 , \25237 );
xnor \U$24924 ( \25239 , \25238 , \22288 );
and \U$24925 ( \25240 , \22213 , \22300 );
and \U$24926 ( \25241 , \22181 , \22298 );
nor \U$24927 ( \25242 , \25240 , \25241 );
xnor \U$24928 ( \25243 , \25242 , \22310 );
xor \U$24929 ( \25244 , \25239 , \25243 );
and \U$24930 ( \25245 , \22235 , \22324 );
and \U$24931 ( \25246 , \22202 , \22322 );
nor \U$24932 ( \25247 , \25245 , \25246 );
xnor \U$24933 ( \25248 , \25247 , \22334 );
xor \U$24934 ( \25249 , \25244 , \25248 );
and \U$24935 ( \25250 , \22124 , \22208 );
and \U$24936 ( \25251 , \22089 , \22206 );
nor \U$24937 ( \25252 , \25250 , \25251 );
xnor \U$24938 ( \25253 , \25252 , \22218 );
and \U$24939 ( \25254 , \22145 , \22230 );
and \U$24940 ( \25255 , \22113 , \22228 );
nor \U$24941 ( \25256 , \25254 , \25255 );
xnor \U$24942 ( \25257 , \25256 , \22240 );
xor \U$24943 ( \25258 , \25253 , \25257 );
and \U$24944 ( \25259 , \22167 , \22257 );
and \U$24945 ( \25260 , \22134 , \22255 );
nor \U$24946 ( \25261 , \25259 , \25260 );
xnor \U$24947 ( \25262 , \25261 , \22267 );
xor \U$24948 ( \25263 , \25258 , \25262 );
xor \U$24949 ( \25264 , \25249 , \25263 );
and \U$24950 ( \25265 , \22894 , \22140 );
and \U$24951 ( \25266 , \23230 , \22138 );
nor \U$24952 ( \25267 , \25265 , \25266 );
xnor \U$24953 ( \25268 , \25267 , \22150 );
and \U$24954 ( \25269 , \22081 , \22162 );
and \U$24955 ( \25270 , \22858 , \22160 );
nor \U$24956 ( \25271 , \25269 , \25270 );
xnor \U$24957 ( \25272 , \25271 , \22172 );
xor \U$24958 ( \25273 , \25268 , \25272 );
and \U$24959 ( \25274 , \22100 , \22187 );
and \U$24960 ( \25275 , \22071 , \22185 );
nor \U$24961 ( \25276 , \25274 , \25275 );
xnor \U$24962 ( \25277 , \25276 , \22197 );
xor \U$24963 ( \25278 , \25273 , \25277 );
xor \U$24964 ( \25279 , \25264 , \25278 );
xor \U$24965 ( \25280 , \25235 , \25279 );
xor \U$24966 ( \25281 , \25217 , \25280 );
and \U$24967 ( \25282 , \24779 , \24781 );
and \U$24968 ( \25283 , \24781 , \24796 );
and \U$24969 ( \25284 , \24779 , \24796 );
or \U$24970 ( \25285 , \25282 , \25283 , \25284 );
and \U$24971 ( \25286 , \24930 , \24944 );
and \U$24972 ( \25287 , \24944 , \24959 );
and \U$24973 ( \25288 , \24930 , \24959 );
or \U$24974 ( \25289 , \25286 , \25287 , \25288 );
xor \U$24975 ( \25290 , \25285 , \25289 );
and \U$24976 ( \25291 , \24885 , \24899 );
and \U$24977 ( \25292 , \24899 , \24914 );
and \U$24978 ( \25293 , \24885 , \24914 );
or \U$24979 ( \25294 , \25291 , \25292 , \25293 );
xor \U$24980 ( \25295 , \25290 , \25294 );
xor \U$24981 ( \25296 , \25281 , \25295 );
xor \U$24982 ( \25297 , \25106 , \25296 );
and \U$24983 ( \25298 , \24871 , \24915 );
and \U$24984 ( \25299 , \24915 , \24960 );
and \U$24985 ( \25300 , \24871 , \24960 );
or \U$24986 ( \25301 , \25298 , \25299 , \25300 );
and \U$24987 ( \25302 , \24797 , \24811 );
and \U$24988 ( \25303 , \24811 , \24826 );
and \U$24989 ( \25304 , \24797 , \24826 );
or \U$24990 ( \25305 , \25302 , \25303 , \25304 );
xor \U$24991 ( \25306 , \25301 , \25305 );
and \U$24992 ( \25307 , \24875 , \24879 );
and \U$24993 ( \25308 , \24879 , \24884 );
and \U$24994 ( \25309 , \24875 , \24884 );
or \U$24995 ( \25310 , \25307 , \25308 , \25309 );
and \U$24996 ( \25311 , \24949 , \24953 );
and \U$24997 ( \25312 , \24953 , \24958 );
and \U$24998 ( \25313 , \24949 , \24958 );
or \U$24999 ( \25314 , \25311 , \25312 , \25313 );
xor \U$25000 ( \25315 , \25310 , \25314 );
and \U$25001 ( \25316 , \24934 , \24938 );
and \U$25002 ( \25317 , \24938 , \24943 );
and \U$25003 ( \25318 , \24934 , \24943 );
or \U$25004 ( \25319 , \25316 , \25317 , \25318 );
xor \U$25005 ( \25320 , \25315 , \25319 );
and \U$25006 ( \25321 , \24831 , \24835 );
and \U$25007 ( \25322 , \24835 , \24840 );
and \U$25008 ( \25323 , \24831 , \24840 );
or \U$25009 ( \25324 , \25321 , \25322 , \25323 );
and \U$25010 ( \25325 , \24904 , \24908 );
and \U$25011 ( \25326 , \24908 , \24913 );
and \U$25012 ( \25327 , \24904 , \24913 );
or \U$25013 ( \25328 , \25325 , \25326 , \25327 );
xor \U$25014 ( \25329 , \25324 , \25328 );
and \U$25015 ( \25330 , \24889 , \24893 );
and \U$25016 ( \25331 , \24893 , \24898 );
and \U$25017 ( \25332 , \24889 , \24898 );
or \U$25018 ( \25333 , \25330 , \25331 , \25332 );
xor \U$25019 ( \25334 , \25329 , \25333 );
xor \U$25020 ( \25335 , \25320 , \25334 );
and \U$25021 ( \25336 , \24972 , \24976 );
and \U$25022 ( \25337 , \24860 , \24864 );
and \U$25023 ( \25338 , \24864 , \24869 );
and \U$25024 ( \25339 , \24860 , \24869 );
or \U$25025 ( \25340 , \25337 , \25338 , \25339 );
xor \U$25026 ( \25341 , \25336 , \25340 );
and \U$25027 ( \25342 , \24845 , \24849 );
and \U$25028 ( \25343 , \24849 , \24854 );
and \U$25029 ( \25344 , \24845 , \24854 );
or \U$25030 ( \25345 , \25342 , \25343 , \25344 );
xor \U$25031 ( \25346 , \25341 , \25345 );
xor \U$25032 ( \25347 , \25335 , \25346 );
xor \U$25033 ( \25348 , \25306 , \25347 );
xor \U$25034 ( \25349 , \25297 , \25348 );
xor \U$25035 ( \25350 , \25092 , \25349 );
xor \U$25036 ( \25351 , \25083 , \25350 );
and \U$25037 ( \25352 , \24728 , \25032 );
nor \U$25038 ( \25353 , \25351 , \25352 );
and \U$25039 ( \25354 , \25087 , \25091 );
and \U$25040 ( \25355 , \25091 , \25349 );
and \U$25041 ( \25356 , \25087 , \25349 );
or \U$25042 ( \25357 , \25354 , \25355 , \25356 );
and \U$25043 ( \25358 , \25057 , \25081 );
xor \U$25044 ( \25359 , \25357 , \25358 );
and \U$25045 ( \25360 , \25061 , \25065 );
and \U$25046 ( \25361 , \25065 , \25080 );
and \U$25047 ( \25362 , \25061 , \25080 );
or \U$25048 ( \25363 , \25360 , \25361 , \25362 );
and \U$25049 ( \25364 , \25336 , \25340 );
and \U$25050 ( \25365 , \25340 , \25345 );
and \U$25051 ( \25366 , \25336 , \25345 );
or \U$25052 ( \25367 , \25364 , \25365 , \25366 );
and \U$25053 ( \25368 , \25324 , \25328 );
and \U$25054 ( \25369 , \25328 , \25333 );
and \U$25055 ( \25370 , \25324 , \25333 );
or \U$25056 ( \25371 , \25368 , \25369 , \25370 );
xor \U$25057 ( \25372 , \25367 , \25371 );
and \U$25058 ( \25373 , \25310 , \25314 );
and \U$25059 ( \25374 , \25314 , \25319 );
and \U$25060 ( \25375 , \25310 , \25319 );
or \U$25061 ( \25376 , \25373 , \25374 , \25375 );
xor \U$25062 ( \25377 , \25372 , \25376 );
and \U$25063 ( \25378 , \22429 , \22551 );
and \U$25064 ( \25379 , \22440 , \22549 );
nor \U$25065 ( \25380 , \25378 , \25379 );
xnor \U$25066 ( \25381 , \25380 , \22561 );
and \U$25067 ( \25382 , \22457 , \22573 );
and \U$25068 ( \25383 , \22468 , \22571 );
nor \U$25069 ( \25384 , \25382 , \25383 );
xnor \U$25070 ( \25385 , \25384 , \22583 );
xor \U$25071 ( \25386 , \25381 , \25385 );
and \U$25072 ( \25387 , \22478 , \22598 );
and \U$25073 ( \25388 , \22489 , \22596 );
nor \U$25074 ( \25389 , \25387 , \25388 );
xnor \U$25075 ( \25390 , \25389 , \22608 );
xor \U$25076 ( \25391 , \25386 , \25390 );
and \U$25077 ( \25392 , \22361 , \22484 );
and \U$25078 ( \25393 , \22372 , \22482 );
nor \U$25079 ( \25394 , \25392 , \25393 );
xnor \U$25080 ( \25395 , \25394 , \22494 );
and \U$25081 ( \25396 , \22386 , \22506 );
and \U$25082 ( \25397 , \22397 , \22504 );
nor \U$25083 ( \25398 , \25396 , \25397 );
xnor \U$25084 ( \25399 , \25398 , \22516 );
xor \U$25085 ( \25400 , \25395 , \25399 );
and \U$25086 ( \25401 , \22407 , \22530 );
and \U$25087 ( \25402 , \22418 , \22528 );
nor \U$25088 ( \25403 , \25401 , \25402 );
xnor \U$25089 ( \25404 , \25403 , \22540 );
xor \U$25090 ( \25405 , \25400 , \25404 );
xor \U$25091 ( \25406 , \25391 , \25405 );
and \U$25092 ( \25407 , \22294 , \22413 );
and \U$25093 ( \25408 , \22305 , \22411 );
nor \U$25094 ( \25409 , \25407 , \25408 );
xnor \U$25095 ( \25410 , \25409 , \22423 );
and \U$25096 ( \25411 , \22318 , \22435 );
and \U$25097 ( \25412 , \22329 , \22433 );
nor \U$25098 ( \25413 , \25411 , \25412 );
xnor \U$25099 ( \25414 , \25413 , \22445 );
xor \U$25100 ( \25415 , \25410 , \25414 );
and \U$25101 ( \25416 , \22339 , \22463 );
and \U$25102 ( \25417 , \22350 , \22461 );
nor \U$25103 ( \25418 , \25416 , \25417 );
xnor \U$25104 ( \25419 , \25418 , \22473 );
xor \U$25105 ( \25420 , \25415 , \25419 );
xor \U$25106 ( \25421 , \25406 , \25420 );
and \U$25107 ( \25422 , \22635 , \22021 );
and \U$25108 ( \25423 , \22646 , \22019 );
nor \U$25109 ( \25424 , \25422 , \25423 );
xnor \U$25110 ( \25425 , \25424 , \21595 );
and \U$25111 ( \25426 , \22665 , \21983 );
and \U$25112 ( \25427 , \22676 , \21981 );
nor \U$25113 ( \25428 , \25426 , \25427 );
xnor \U$25114 ( \25429 , \25428 , \21995 );
xor \U$25115 ( \25430 , \25425 , \25429 );
and \U$25116 ( \25431 , \22696 , \21978 );
xor \U$25117 ( \25432 , \25430 , \25431 );
and \U$25118 ( \25433 , \22567 , \22691 );
and \U$25119 ( \25434 , \22578 , \22689 );
nor \U$25120 ( \25435 , \25433 , \25434 );
xnor \U$25121 ( \25436 , \25435 , \22701 );
and \U$25122 ( \25437 , \22592 , \22720 );
and \U$25123 ( \25438 , \22603 , \22707 );
nor \U$25124 ( \25439 , \25437 , \25438 );
xnor \U$25125 ( \25440 , \25439 , \22067 );
xor \U$25126 ( \25441 , \25436 , \25440 );
and \U$25127 ( \25442 , \22613 , \23173 );
and \U$25128 ( \25443 , \22624 , \22999 );
nor \U$25129 ( \25444 , \25442 , \25443 );
xnor \U$25130 ( \25445 , \25444 , \22016 );
xor \U$25131 ( \25446 , \25441 , \25445 );
xor \U$25132 ( \25447 , \25432 , \25446 );
and \U$25133 ( \25448 , \22500 , \22619 );
and \U$25134 ( \25449 , \22511 , \22617 );
nor \U$25135 ( \25450 , \25448 , \25449 );
xnor \U$25136 ( \25451 , \25450 , \22629 );
and \U$25137 ( \25452 , \22524 , \22641 );
and \U$25138 ( \25453 , \22535 , \22639 );
nor \U$25139 ( \25454 , \25452 , \25453 );
xnor \U$25140 ( \25455 , \25454 , \22651 );
xor \U$25141 ( \25456 , \25451 , \25455 );
and \U$25142 ( \25457 , \22545 , \22671 );
and \U$25143 ( \25458 , \22556 , \22669 );
nor \U$25144 ( \25459 , \25457 , \25458 );
xnor \U$25145 ( \25460 , \25459 , \22681 );
xor \U$25146 ( \25461 , \25456 , \25460 );
xor \U$25147 ( \25462 , \25447 , \25461 );
xor \U$25148 ( \25463 , \25421 , \25462 );
and \U$25149 ( \25464 , \25154 , \25158 );
and \U$25150 ( \25465 , \25158 , \25163 );
and \U$25151 ( \25466 , \25154 , \25163 );
or \U$25152 ( \25467 , \25464 , \25465 , \25466 );
and \U$25153 ( \25468 , \25208 , \25212 );
and \U$25154 ( \25469 , \25212 , \25214 );
and \U$25155 ( \25470 , \25208 , \25214 );
or \U$25156 ( \25471 , \25468 , \25469 , \25470 );
xnor \U$25157 ( \25472 , \25467 , \25471 );
xor \U$25158 ( \25473 , \25463 , \25472 );
and \U$25159 ( \25474 , \25249 , \25263 );
and \U$25160 ( \25475 , \25263 , \25278 );
and \U$25161 ( \25476 , \25249 , \25278 );
or \U$25162 ( \25477 , \25474 , \25475 , \25476 );
and \U$25163 ( \25478 , \23230 , \22140 );
and \U$25164 ( \25479 , \23329 , \22138 );
nor \U$25165 ( \25480 , \25478 , \25479 );
xnor \U$25166 ( \25481 , \25480 , \22150 );
and \U$25167 ( \25482 , \22858 , \22162 );
and \U$25168 ( \25483 , \22894 , \22160 );
nor \U$25169 ( \25484 , \25482 , \25483 );
xnor \U$25170 ( \25485 , \25484 , \22172 );
xor \U$25171 ( \25486 , \25481 , \25485 );
and \U$25172 ( \25487 , \22071 , \22187 );
and \U$25173 ( \25488 , \22081 , \22185 );
nor \U$25174 ( \25489 , \25487 , \25488 );
xnor \U$25175 ( \25490 , \25489 , \22197 );
xor \U$25176 ( \25491 , \25486 , \25490 );
not \U$25177 ( \25492 , \22072 );
and \U$25178 ( \25493 , \21977 , \22095 );
and \U$25179 ( \25494 , \21990 , \22093 );
nor \U$25180 ( \25495 , \25493 , \25494 );
xnor \U$25181 ( \25496 , \25495 , \22105 );
xor \U$25182 ( \25497 , \25492 , \25496 );
and \U$25183 ( \25498 , \22030 , \22119 );
and \U$25184 ( \25499 , \22001 , \22117 );
nor \U$25185 ( \25500 , \25498 , \25499 );
xnor \U$25186 ( \25501 , \25500 , \22129 );
xor \U$25187 ( \25502 , \25497 , \25501 );
xor \U$25188 ( \25503 , \25491 , \25502 );
xor \U$25189 ( \25504 , \25477 , \25503 );
and \U$25190 ( \25505 , \22224 , \22345 );
and \U$25191 ( \25506 , \22235 , \22343 );
nor \U$25192 ( \25507 , \25505 , \25506 );
xnor \U$25193 ( \25508 , \25507 , \22355 );
and \U$25194 ( \25509 , \22251 , \22367 );
and \U$25195 ( \25510 , \22262 , \22365 );
nor \U$25196 ( \25511 , \25509 , \25510 );
xnor \U$25197 ( \25512 , \25511 , \22377 );
xor \U$25198 ( \25513 , \25508 , \25512 );
and \U$25199 ( \25514 , \22272 , \22392 );
and \U$25200 ( \25515 , \22283 , \22390 );
nor \U$25201 ( \25516 , \25514 , \25515 );
xnor \U$25202 ( \25517 , \25516 , \22402 );
xor \U$25203 ( \25518 , \25513 , \25517 );
and \U$25204 ( \25519 , \22156 , \22278 );
and \U$25205 ( \25520 , \22167 , \22276 );
nor \U$25206 ( \25521 , \25519 , \25520 );
xnor \U$25207 ( \25522 , \25521 , \22288 );
and \U$25208 ( \25523 , \22181 , \22300 );
and \U$25209 ( \25524 , \22192 , \22298 );
nor \U$25210 ( \25525 , \25523 , \25524 );
xnor \U$25211 ( \25526 , \25525 , \22310 );
xor \U$25212 ( \25527 , \25522 , \25526 );
and \U$25213 ( \25528 , \22202 , \22324 );
and \U$25214 ( \25529 , \22213 , \22322 );
nor \U$25215 ( \25530 , \25528 , \25529 );
xnor \U$25216 ( \25531 , \25530 , \22334 );
xor \U$25217 ( \25532 , \25527 , \25531 );
xor \U$25218 ( \25533 , \25518 , \25532 );
and \U$25219 ( \25534 , \22089 , \22208 );
and \U$25220 ( \25535 , \22100 , \22206 );
nor \U$25221 ( \25536 , \25534 , \25535 );
xnor \U$25222 ( \25537 , \25536 , \22218 );
and \U$25223 ( \25538 , \22113 , \22230 );
and \U$25224 ( \25539 , \22124 , \22228 );
nor \U$25225 ( \25540 , \25538 , \25539 );
xnor \U$25226 ( \25541 , \25540 , \22240 );
xor \U$25227 ( \25542 , \25537 , \25541 );
and \U$25228 ( \25543 , \22134 , \22257 );
and \U$25229 ( \25544 , \22145 , \22255 );
nor \U$25230 ( \25545 , \25543 , \25544 );
xnor \U$25231 ( \25546 , \25545 , \22267 );
xor \U$25232 ( \25547 , \25542 , \25546 );
xor \U$25233 ( \25548 , \25533 , \25547 );
xor \U$25234 ( \25549 , \25504 , \25548 );
xor \U$25235 ( \25550 , \25473 , \25549 );
and \U$25236 ( \25551 , \25199 , \25203 );
and \U$25237 ( \25552 , \25203 , \25215 );
and \U$25238 ( \25553 , \25199 , \25215 );
or \U$25239 ( \25554 , \25551 , \25552 , \25553 );
and \U$25240 ( \25555 , \25164 , \25178 );
and \U$25241 ( \25556 , \25178 , \25193 );
and \U$25242 ( \25557 , \25164 , \25193 );
or \U$25243 ( \25558 , \25555 , \25556 , \25557 );
xor \U$25244 ( \25559 , \25554 , \25558 );
and \U$25245 ( \25560 , \25120 , \25134 );
and \U$25246 ( \25561 , \25134 , \25149 );
and \U$25247 ( \25562 , \25120 , \25149 );
or \U$25248 ( \25563 , \25560 , \25561 , \25562 );
xor \U$25249 ( \25564 , \25559 , \25563 );
xor \U$25250 ( \25565 , \25550 , \25564 );
xor \U$25251 ( \25566 , \25377 , \25565 );
and \U$25252 ( \25567 , \25150 , \25194 );
and \U$25253 ( \25568 , \25194 , \25216 );
and \U$25254 ( \25569 , \25150 , \25216 );
or \U$25255 ( \25570 , \25567 , \25568 , \25569 );
and \U$25256 ( \25571 , \25320 , \25334 );
and \U$25257 ( \25572 , \25334 , \25346 );
and \U$25258 ( \25573 , \25320 , \25346 );
or \U$25259 ( \25574 , \25571 , \25572 , \25573 );
xor \U$25260 ( \25575 , \25570 , \25574 );
and \U$25261 ( \25576 , \25110 , \25114 );
and \U$25262 ( \25577 , \25114 , \25119 );
and \U$25263 ( \25578 , \25110 , \25119 );
or \U$25264 ( \25579 , \25576 , \25577 , \25578 );
and \U$25265 ( \25580 , \25183 , \25187 );
and \U$25266 ( \25581 , \25187 , \25192 );
and \U$25267 ( \25582 , \25183 , \25192 );
or \U$25268 ( \25583 , \25580 , \25581 , \25582 );
xor \U$25269 ( \25584 , \25579 , \25583 );
and \U$25270 ( \25585 , \25168 , \25172 );
and \U$25271 ( \25586 , \25172 , \25177 );
and \U$25272 ( \25587 , \25168 , \25177 );
or \U$25273 ( \25588 , \25585 , \25586 , \25587 );
xor \U$25274 ( \25589 , \25584 , \25588 );
and \U$25275 ( \25590 , \25239 , \25243 );
and \U$25276 ( \25591 , \25243 , \25248 );
and \U$25277 ( \25592 , \25239 , \25248 );
or \U$25278 ( \25593 , \25590 , \25591 , \25592 );
and \U$25279 ( \25594 , \25139 , \25143 );
and \U$25280 ( \25595 , \25143 , \25148 );
and \U$25281 ( \25596 , \25139 , \25148 );
or \U$25282 ( \25597 , \25594 , \25595 , \25596 );
xor \U$25283 ( \25598 , \25593 , \25597 );
and \U$25284 ( \25599 , \25124 , \25128 );
and \U$25285 ( \25600 , \25128 , \25133 );
and \U$25286 ( \25601 , \25124 , \25133 );
or \U$25287 ( \25602 , \25599 , \25600 , \25601 );
xor \U$25288 ( \25603 , \25598 , \25602 );
xor \U$25289 ( \25604 , \25589 , \25603 );
and \U$25290 ( \25605 , \25224 , \25228 );
and \U$25291 ( \25606 , \25228 , \25233 );
and \U$25292 ( \25607 , \25224 , \25233 );
or \U$25293 ( \25608 , \25605 , \25606 , \25607 );
and \U$25294 ( \25609 , \25268 , \25272 );
and \U$25295 ( \25610 , \25272 , \25277 );
and \U$25296 ( \25611 , \25268 , \25277 );
or \U$25297 ( \25612 , \25609 , \25610 , \25611 );
xor \U$25298 ( \25613 , \25608 , \25612 );
and \U$25299 ( \25614 , \25253 , \25257 );
and \U$25300 ( \25615 , \25257 , \25262 );
and \U$25301 ( \25616 , \25253 , \25262 );
or \U$25302 ( \25617 , \25614 , \25615 , \25616 );
xor \U$25303 ( \25618 , \25613 , \25617 );
xor \U$25304 ( \25619 , \25604 , \25618 );
xor \U$25305 ( \25620 , \25575 , \25619 );
xor \U$25306 ( \25621 , \25566 , \25620 );
and \U$25307 ( \25622 , \25070 , \25074 );
and \U$25308 ( \25623 , \25074 , \25079 );
and \U$25309 ( \25624 , \25070 , \25079 );
or \U$25310 ( \25625 , \25622 , \25623 , \25624 );
and \U$25311 ( \25626 , \25301 , \25305 );
and \U$25312 ( \25627 , \25305 , \25347 );
and \U$25313 ( \25628 , \25301 , \25347 );
or \U$25314 ( \25629 , \25626 , \25627 , \25628 );
xor \U$25315 ( \25630 , \25625 , \25629 );
and \U$25316 ( \25631 , \25217 , \25280 );
and \U$25317 ( \25632 , \25280 , \25295 );
and \U$25318 ( \25633 , \25217 , \25295 );
or \U$25319 ( \25634 , \25631 , \25632 , \25633 );
xor \U$25320 ( \25635 , \25630 , \25634 );
xor \U$25321 ( \25636 , \25621 , \25635 );
xor \U$25322 ( \25637 , \25363 , \25636 );
and \U$25323 ( \25638 , \25047 , \25051 );
and \U$25324 ( \25639 , \25051 , \25056 );
and \U$25325 ( \25640 , \25047 , \25056 );
or \U$25326 ( \25641 , \25638 , \25639 , \25640 );
and \U$25327 ( \25642 , \25106 , \25296 );
and \U$25328 ( \25643 , \25296 , \25348 );
and \U$25329 ( \25644 , \25106 , \25348 );
or \U$25330 ( \25645 , \25642 , \25643 , \25644 );
xor \U$25331 ( \25646 , \25641 , \25645 );
and \U$25332 ( \25647 , \25096 , \25100 );
and \U$25333 ( \25648 , \25100 , \25105 );
and \U$25334 ( \25649 , \25096 , \25105 );
or \U$25335 ( \25650 , \25647 , \25648 , \25649 );
and \U$25336 ( \25651 , \25285 , \25289 );
and \U$25337 ( \25652 , \25289 , \25294 );
and \U$25338 ( \25653 , \25285 , \25294 );
or \U$25339 ( \25654 , \25651 , \25652 , \25653 );
xor \U$25340 ( \25655 , \25650 , \25654 );
and \U$25341 ( \25656 , \25221 , \25234 );
and \U$25342 ( \25657 , \25234 , \25279 );
and \U$25343 ( \25658 , \25221 , \25279 );
or \U$25344 ( \25659 , \25656 , \25657 , \25658 );
xor \U$25345 ( \25660 , \25655 , \25659 );
xor \U$25346 ( \25661 , \25646 , \25660 );
xor \U$25347 ( \25662 , \25637 , \25661 );
xor \U$25348 ( \25663 , \25359 , \25662 );
and \U$25349 ( \25664 , \25043 , \25082 );
and \U$25350 ( \25665 , \25082 , \25350 );
and \U$25351 ( \25666 , \25043 , \25350 );
or \U$25352 ( \25667 , \25664 , \25665 , \25666 );
nor \U$25353 ( \25668 , \25663 , \25667 );
nor \U$25354 ( \25669 , \25353 , \25668 );
nand \U$25355 ( \25670 , \25039 , \25669 );
and \U$25356 ( \25671 , \25363 , \25636 );
and \U$25357 ( \25672 , \25636 , \25661 );
and \U$25358 ( \25673 , \25363 , \25661 );
or \U$25359 ( \25674 , \25671 , \25672 , \25673 );
and \U$25360 ( \25675 , \25625 , \25629 );
and \U$25361 ( \25676 , \25629 , \25634 );
and \U$25362 ( \25677 , \25625 , \25634 );
or \U$25363 ( \25678 , \25675 , \25676 , \25677 );
and \U$25364 ( \25679 , \25377 , \25565 );
and \U$25365 ( \25680 , \25565 , \25620 );
and \U$25366 ( \25681 , \25377 , \25620 );
or \U$25367 ( \25682 , \25679 , \25680 , \25681 );
xor \U$25368 ( \25683 , \25678 , \25682 );
and \U$25369 ( \25684 , \25421 , \25462 );
and \U$25370 ( \25685 , \25462 , \25472 );
and \U$25371 ( \25686 , \25421 , \25472 );
or \U$25372 ( \25687 , \25684 , \25685 , \25686 );
and \U$25373 ( \25688 , \25589 , \25603 );
and \U$25374 ( \25689 , \25603 , \25618 );
and \U$25375 ( \25690 , \25589 , \25618 );
or \U$25376 ( \25691 , \25688 , \25689 , \25690 );
xor \U$25377 ( \25692 , \25687 , \25691 );
and \U$25378 ( \25693 , \25492 , \25496 );
and \U$25379 ( \25694 , \25496 , \25501 );
and \U$25380 ( \25695 , \25492 , \25501 );
or \U$25381 ( \25696 , \25693 , \25694 , \25695 );
and \U$25382 ( \25697 , \25481 , \25485 );
and \U$25383 ( \25698 , \25485 , \25490 );
and \U$25384 ( \25699 , \25481 , \25490 );
or \U$25385 ( \25700 , \25697 , \25698 , \25699 );
xor \U$25386 ( \25701 , \25696 , \25700 );
and \U$25387 ( \25702 , \25537 , \25541 );
and \U$25388 ( \25703 , \25541 , \25546 );
and \U$25389 ( \25704 , \25537 , \25546 );
or \U$25390 ( \25705 , \25702 , \25703 , \25704 );
xor \U$25391 ( \25706 , \25701 , \25705 );
xor \U$25392 ( \25707 , \25692 , \25706 );
xor \U$25393 ( \25708 , \25683 , \25707 );
xor \U$25394 ( \25709 , \25674 , \25708 );
and \U$25395 ( \25710 , \25641 , \25645 );
and \U$25396 ( \25711 , \25645 , \25660 );
and \U$25397 ( \25712 , \25641 , \25660 );
or \U$25398 ( \25713 , \25710 , \25711 , \25712 );
and \U$25399 ( \25714 , \25621 , \25635 );
xor \U$25400 ( \25715 , \25713 , \25714 );
and \U$25401 ( \25716 , \25367 , \25371 );
and \U$25402 ( \25717 , \25371 , \25376 );
and \U$25403 ( \25718 , \25367 , \25376 );
or \U$25404 ( \25719 , \25716 , \25717 , \25718 );
and \U$25405 ( \25720 , \25554 , \25558 );
and \U$25406 ( \25721 , \25558 , \25563 );
and \U$25407 ( \25722 , \25554 , \25563 );
or \U$25408 ( \25723 , \25720 , \25721 , \25722 );
xor \U$25409 ( \25724 , \25719 , \25723 );
and \U$25410 ( \25725 , \25477 , \25503 );
and \U$25411 ( \25726 , \25503 , \25548 );
and \U$25412 ( \25727 , \25477 , \25548 );
or \U$25413 ( \25728 , \25725 , \25726 , \25727 );
xor \U$25414 ( \25729 , \25724 , \25728 );
or \U$25415 ( \25730 , \25467 , \25471 );
and \U$25416 ( \25731 , \25432 , \25446 );
and \U$25417 ( \25732 , \25446 , \25461 );
and \U$25418 ( \25733 , \25432 , \25461 );
or \U$25419 ( \25734 , \25731 , \25732 , \25733 );
xor \U$25420 ( \25735 , \25730 , \25734 );
and \U$25421 ( \25736 , \25391 , \25405 );
and \U$25422 ( \25737 , \25405 , \25420 );
and \U$25423 ( \25738 , \25391 , \25420 );
or \U$25424 ( \25739 , \25736 , \25737 , \25738 );
xor \U$25425 ( \25740 , \25735 , \25739 );
and \U$25426 ( \25741 , \25608 , \25612 );
and \U$25427 ( \25742 , \25612 , \25617 );
and \U$25428 ( \25743 , \25608 , \25617 );
or \U$25429 ( \25744 , \25741 , \25742 , \25743 );
and \U$25430 ( \25745 , \25593 , \25597 );
and \U$25431 ( \25746 , \25597 , \25602 );
and \U$25432 ( \25747 , \25593 , \25602 );
or \U$25433 ( \25748 , \25745 , \25746 , \25747 );
xor \U$25434 ( \25749 , \25744 , \25748 );
and \U$25435 ( \25750 , \25579 , \25583 );
and \U$25436 ( \25751 , \25583 , \25588 );
and \U$25437 ( \25752 , \25579 , \25588 );
or \U$25438 ( \25753 , \25750 , \25751 , \25752 );
xor \U$25439 ( \25754 , \25749 , \25753 );
xor \U$25440 ( \25755 , \25740 , \25754 );
and \U$25441 ( \25756 , \25436 , \25440 );
and \U$25442 ( \25757 , \25440 , \25445 );
and \U$25443 ( \25758 , \25436 , \25445 );
or \U$25444 ( \25759 , \25756 , \25757 , \25758 );
and \U$25445 ( \25760 , \25425 , \25429 );
and \U$25446 ( \25761 , \25429 , \25431 );
and \U$25447 ( \25762 , \25425 , \25431 );
or \U$25448 ( \25763 , \25760 , \25761 , \25762 );
xor \U$25449 ( \25764 , \25759 , \25763 );
and \U$25450 ( \25765 , \22676 , \21983 );
and \U$25451 ( \25766 , \22635 , \21981 );
nor \U$25452 ( \25767 , \25765 , \25766 );
xnor \U$25453 ( \25768 , \25767 , \21995 );
and \U$25454 ( \25769 , \22665 , \21978 );
xnor \U$25455 ( \25770 , \25768 , \25769 );
xor \U$25456 ( \25771 , \25764 , \25770 );
and \U$25457 ( \25772 , \25395 , \25399 );
and \U$25458 ( \25773 , \25399 , \25404 );
and \U$25459 ( \25774 , \25395 , \25404 );
or \U$25460 ( \25775 , \25772 , \25773 , \25774 );
and \U$25461 ( \25776 , \25381 , \25385 );
and \U$25462 ( \25777 , \25385 , \25390 );
and \U$25463 ( \25778 , \25381 , \25390 );
or \U$25464 ( \25779 , \25776 , \25777 , \25778 );
xor \U$25465 ( \25780 , \25775 , \25779 );
and \U$25466 ( \25781 , \25451 , \25455 );
and \U$25467 ( \25782 , \25455 , \25460 );
and \U$25468 ( \25783 , \25451 , \25460 );
or \U$25469 ( \25784 , \25781 , \25782 , \25783 );
xor \U$25470 ( \25785 , \25780 , \25784 );
xor \U$25471 ( \25786 , \25771 , \25785 );
and \U$25472 ( \25787 , \25522 , \25526 );
and \U$25473 ( \25788 , \25526 , \25531 );
and \U$25474 ( \25789 , \25522 , \25531 );
or \U$25475 ( \25790 , \25787 , \25788 , \25789 );
and \U$25476 ( \25791 , \25508 , \25512 );
and \U$25477 ( \25792 , \25512 , \25517 );
and \U$25478 ( \25793 , \25508 , \25517 );
or \U$25479 ( \25794 , \25791 , \25792 , \25793 );
xor \U$25480 ( \25795 , \25790 , \25794 );
and \U$25481 ( \25796 , \25410 , \25414 );
and \U$25482 ( \25797 , \25414 , \25419 );
and \U$25483 ( \25798 , \25410 , \25419 );
or \U$25484 ( \25799 , \25796 , \25797 , \25798 );
xor \U$25485 ( \25800 , \25795 , \25799 );
xor \U$25486 ( \25801 , \25786 , \25800 );
and \U$25487 ( \25802 , \22192 , \22300 );
and \U$25488 ( \25803 , \22156 , \22298 );
nor \U$25489 ( \25804 , \25802 , \25803 );
xnor \U$25490 ( \25805 , \25804 , \22310 );
and \U$25491 ( \25806 , \22213 , \22324 );
and \U$25492 ( \25807 , \22181 , \22322 );
nor \U$25493 ( \25808 , \25806 , \25807 );
xnor \U$25494 ( \25809 , \25808 , \22334 );
xor \U$25495 ( \25810 , \25805 , \25809 );
and \U$25496 ( \25811 , \22235 , \22345 );
and \U$25497 ( \25812 , \22202 , \22343 );
nor \U$25498 ( \25813 , \25811 , \25812 );
xnor \U$25499 ( \25814 , \25813 , \22355 );
xor \U$25500 ( \25815 , \25810 , \25814 );
and \U$25501 ( \25816 , \22124 , \22230 );
and \U$25502 ( \25817 , \22089 , \22228 );
nor \U$25503 ( \25818 , \25816 , \25817 );
xnor \U$25504 ( \25819 , \25818 , \22240 );
and \U$25505 ( \25820 , \22145 , \22257 );
and \U$25506 ( \25821 , \22113 , \22255 );
nor \U$25507 ( \25822 , \25820 , \25821 );
xnor \U$25508 ( \25823 , \25822 , \22267 );
xor \U$25509 ( \25824 , \25819 , \25823 );
and \U$25510 ( \25825 , \22167 , \22278 );
and \U$25511 ( \25826 , \22134 , \22276 );
nor \U$25512 ( \25827 , \25825 , \25826 );
xnor \U$25513 ( \25828 , \25827 , \22288 );
xor \U$25514 ( \25829 , \25824 , \25828 );
xor \U$25515 ( \25830 , \25815 , \25829 );
and \U$25516 ( \25831 , \22894 , \22162 );
and \U$25517 ( \25832 , \23230 , \22160 );
nor \U$25518 ( \25833 , \25831 , \25832 );
xnor \U$25519 ( \25834 , \25833 , \22172 );
and \U$25520 ( \25835 , \22081 , \22187 );
and \U$25521 ( \25836 , \22858 , \22185 );
nor \U$25522 ( \25837 , \25835 , \25836 );
xnor \U$25523 ( \25838 , \25837 , \22197 );
xor \U$25524 ( \25839 , \25834 , \25838 );
and \U$25525 ( \25840 , \22100 , \22208 );
and \U$25526 ( \25841 , \22071 , \22206 );
nor \U$25527 ( \25842 , \25840 , \25841 );
xnor \U$25528 ( \25843 , \25842 , \22218 );
xor \U$25529 ( \25844 , \25839 , \25843 );
xor \U$25530 ( \25845 , \25830 , \25844 );
and \U$25531 ( \25846 , \22397 , \22506 );
and \U$25532 ( \25847 , \22361 , \22504 );
nor \U$25533 ( \25848 , \25846 , \25847 );
xnor \U$25534 ( \25849 , \25848 , \22516 );
and \U$25535 ( \25850 , \22418 , \22530 );
and \U$25536 ( \25851 , \22386 , \22528 );
nor \U$25537 ( \25852 , \25850 , \25851 );
xnor \U$25538 ( \25853 , \25852 , \22540 );
xor \U$25539 ( \25854 , \25849 , \25853 );
and \U$25540 ( \25855 , \22440 , \22551 );
and \U$25541 ( \25856 , \22407 , \22549 );
nor \U$25542 ( \25857 , \25855 , \25856 );
xnor \U$25543 ( \25858 , \25857 , \22561 );
xor \U$25544 ( \25859 , \25854 , \25858 );
and \U$25545 ( \25860 , \22329 , \22435 );
and \U$25546 ( \25861 , \22294 , \22433 );
nor \U$25547 ( \25862 , \25860 , \25861 );
xnor \U$25548 ( \25863 , \25862 , \22445 );
and \U$25549 ( \25864 , \22350 , \22463 );
and \U$25550 ( \25865 , \22318 , \22461 );
nor \U$25551 ( \25866 , \25864 , \25865 );
xnor \U$25552 ( \25867 , \25866 , \22473 );
xor \U$25553 ( \25868 , \25863 , \25867 );
and \U$25554 ( \25869 , \22372 , \22484 );
and \U$25555 ( \25870 , \22339 , \22482 );
nor \U$25556 ( \25871 , \25869 , \25870 );
xnor \U$25557 ( \25872 , \25871 , \22494 );
xor \U$25558 ( \25873 , \25868 , \25872 );
xor \U$25559 ( \25874 , \25859 , \25873 );
and \U$25560 ( \25875 , \22262 , \22367 );
and \U$25561 ( \25876 , \22224 , \22365 );
nor \U$25562 ( \25877 , \25875 , \25876 );
xnor \U$25563 ( \25878 , \25877 , \22377 );
and \U$25564 ( \25879 , \22283 , \22392 );
and \U$25565 ( \25880 , \22251 , \22390 );
nor \U$25566 ( \25881 , \25879 , \25880 );
xnor \U$25567 ( \25882 , \25881 , \22402 );
xor \U$25568 ( \25883 , \25878 , \25882 );
and \U$25569 ( \25884 , \22305 , \22413 );
and \U$25570 ( \25885 , \22272 , \22411 );
nor \U$25571 ( \25886 , \25884 , \25885 );
xnor \U$25572 ( \25887 , \25886 , \22423 );
xor \U$25573 ( \25888 , \25883 , \25887 );
xor \U$25574 ( \25889 , \25874 , \25888 );
xor \U$25575 ( \25890 , \25845 , \25889 );
and \U$25576 ( \25891 , \22603 , \22720 );
and \U$25577 ( \25892 , \22567 , \22707 );
nor \U$25578 ( \25893 , \25891 , \25892 );
xnor \U$25579 ( \25894 , \25893 , \22067 );
and \U$25580 ( \25895 , \22624 , \23173 );
and \U$25581 ( \25896 , \22592 , \22999 );
nor \U$25582 ( \25897 , \25895 , \25896 );
xnor \U$25583 ( \25898 , \25897 , \22016 );
xor \U$25584 ( \25899 , \25894 , \25898 );
and \U$25585 ( \25900 , \22646 , \22021 );
and \U$25586 ( \25901 , \22613 , \22019 );
nor \U$25587 ( \25902 , \25900 , \25901 );
xnor \U$25588 ( \25903 , \25902 , \21595 );
xor \U$25589 ( \25904 , \25899 , \25903 );
and \U$25590 ( \25905 , \22535 , \22641 );
and \U$25591 ( \25906 , \22500 , \22639 );
nor \U$25592 ( \25907 , \25905 , \25906 );
xnor \U$25593 ( \25908 , \25907 , \22651 );
and \U$25594 ( \25909 , \22556 , \22671 );
and \U$25595 ( \25910 , \22524 , \22669 );
nor \U$25596 ( \25911 , \25909 , \25910 );
xnor \U$25597 ( \25912 , \25911 , \22681 );
xor \U$25598 ( \25913 , \25908 , \25912 );
and \U$25599 ( \25914 , \22578 , \22691 );
and \U$25600 ( \25915 , \22545 , \22689 );
nor \U$25601 ( \25916 , \25914 , \25915 );
xnor \U$25602 ( \25917 , \25916 , \22701 );
xor \U$25603 ( \25918 , \25913 , \25917 );
xor \U$25604 ( \25919 , \25904 , \25918 );
and \U$25605 ( \25920 , \22468 , \22573 );
and \U$25606 ( \25921 , \22429 , \22571 );
nor \U$25607 ( \25922 , \25920 , \25921 );
xnor \U$25608 ( \25923 , \25922 , \22583 );
and \U$25609 ( \25924 , \22489 , \22598 );
and \U$25610 ( \25925 , \22457 , \22596 );
nor \U$25611 ( \25926 , \25924 , \25925 );
xnor \U$25612 ( \25927 , \25926 , \22608 );
xor \U$25613 ( \25928 , \25923 , \25927 );
and \U$25614 ( \25929 , \22511 , \22619 );
and \U$25615 ( \25930 , \22478 , \22617 );
nor \U$25616 ( \25931 , \25929 , \25930 );
xnor \U$25617 ( \25932 , \25931 , \22629 );
xor \U$25618 ( \25933 , \25928 , \25932 );
xor \U$25619 ( \25934 , \25919 , \25933 );
xor \U$25620 ( \25935 , \25890 , \25934 );
xor \U$25621 ( \25936 , \25801 , \25935 );
and \U$25622 ( \25937 , \25518 , \25532 );
and \U$25623 ( \25938 , \25532 , \25547 );
and \U$25624 ( \25939 , \25518 , \25547 );
or \U$25625 ( \25940 , \25937 , \25938 , \25939 );
and \U$25626 ( \25941 , \25491 , \25502 );
xor \U$25627 ( \25942 , \25940 , \25941 );
and \U$25628 ( \25943 , \21990 , \22095 );
not \U$25629 ( \25944 , \25943 );
xnor \U$25630 ( \25945 , \25944 , \22105 );
and \U$25631 ( \25946 , \22001 , \22119 );
and \U$25632 ( \25947 , \21977 , \22117 );
nor \U$25633 ( \25948 , \25946 , \25947 );
xnor \U$25634 ( \25949 , \25948 , \22129 );
xor \U$25635 ( \25950 , \25945 , \25949 );
and \U$25636 ( \25951 , \23329 , \22140 );
and \U$25637 ( \25952 , \22030 , \22138 );
nor \U$25638 ( \25953 , \25951 , \25952 );
xnor \U$25639 ( \25954 , \25953 , \22150 );
xor \U$25640 ( \25955 , \25950 , \25954 );
xor \U$25641 ( \25956 , \25942 , \25955 );
xor \U$25642 ( \25957 , \25936 , \25956 );
xor \U$25643 ( \25958 , \25755 , \25957 );
xor \U$25644 ( \25959 , \25729 , \25958 );
and \U$25645 ( \25960 , \25650 , \25654 );
and \U$25646 ( \25961 , \25654 , \25659 );
and \U$25647 ( \25962 , \25650 , \25659 );
or \U$25648 ( \25963 , \25960 , \25961 , \25962 );
and \U$25649 ( \25964 , \25570 , \25574 );
and \U$25650 ( \25965 , \25574 , \25619 );
and \U$25651 ( \25966 , \25570 , \25619 );
or \U$25652 ( \25967 , \25964 , \25965 , \25966 );
xor \U$25653 ( \25968 , \25963 , \25967 );
and \U$25654 ( \25969 , \25473 , \25549 );
and \U$25655 ( \25970 , \25549 , \25564 );
and \U$25656 ( \25971 , \25473 , \25564 );
or \U$25657 ( \25972 , \25969 , \25970 , \25971 );
xor \U$25658 ( \25973 , \25968 , \25972 );
xor \U$25659 ( \25974 , \25959 , \25973 );
xor \U$25660 ( \25975 , \25715 , \25974 );
xor \U$25661 ( \25976 , \25709 , \25975 );
and \U$25662 ( \25977 , \25357 , \25358 );
and \U$25663 ( \25978 , \25358 , \25662 );
and \U$25664 ( \25979 , \25357 , \25662 );
or \U$25665 ( \25980 , \25977 , \25978 , \25979 );
nor \U$25666 ( \25981 , \25976 , \25980 );
and \U$25667 ( \25982 , \25713 , \25714 );
and \U$25668 ( \25983 , \25714 , \25974 );
and \U$25669 ( \25984 , \25713 , \25974 );
or \U$25670 ( \25985 , \25982 , \25983 , \25984 );
and \U$25671 ( \25986 , \25719 , \25723 );
and \U$25672 ( \25987 , \25723 , \25728 );
and \U$25673 ( \25988 , \25719 , \25728 );
or \U$25674 ( \25989 , \25986 , \25987 , \25988 );
and \U$25675 ( \25990 , \25687 , \25691 );
and \U$25676 ( \25991 , \25691 , \25706 );
and \U$25677 ( \25992 , \25687 , \25706 );
or \U$25678 ( \25993 , \25990 , \25991 , \25992 );
xor \U$25679 ( \25994 , \25989 , \25993 );
and \U$25680 ( \25995 , \25801 , \25935 );
and \U$25681 ( \25996 , \25935 , \25956 );
and \U$25682 ( \25997 , \25801 , \25956 );
or \U$25683 ( \25998 , \25995 , \25996 , \25997 );
xor \U$25684 ( \25999 , \25994 , \25998 );
and \U$25685 ( \26000 , \25963 , \25967 );
and \U$25686 ( \26001 , \25967 , \25972 );
and \U$25687 ( \26002 , \25963 , \25972 );
or \U$25688 ( \26003 , \26000 , \26001 , \26002 );
and \U$25689 ( \26004 , \25740 , \25754 );
and \U$25690 ( \26005 , \25754 , \25957 );
and \U$25691 ( \26006 , \25740 , \25957 );
or \U$25692 ( \26007 , \26004 , \26005 , \26006 );
xor \U$25693 ( \26008 , \26003 , \26007 );
and \U$25694 ( \26009 , \25744 , \25748 );
and \U$25695 ( \26010 , \25748 , \25753 );
and \U$25696 ( \26011 , \25744 , \25753 );
or \U$25697 ( \26012 , \26009 , \26010 , \26011 );
and \U$25698 ( \26013 , \25730 , \25734 );
and \U$25699 ( \26014 , \25734 , \25739 );
and \U$25700 ( \26015 , \25730 , \25739 );
or \U$25701 ( \26016 , \26013 , \26014 , \26015 );
xor \U$25702 ( \26017 , \26012 , \26016 );
and \U$25703 ( \26018 , \25940 , \25941 );
and \U$25704 ( \26019 , \25941 , \25955 );
and \U$25705 ( \26020 , \25940 , \25955 );
or \U$25706 ( \26021 , \26018 , \26019 , \26020 );
xor \U$25707 ( \26022 , \26017 , \26021 );
xor \U$25708 ( \26023 , \26008 , \26022 );
xor \U$25709 ( \26024 , \25999 , \26023 );
xor \U$25710 ( \26025 , \25985 , \26024 );
and \U$25711 ( \26026 , \25678 , \25682 );
and \U$25712 ( \26027 , \25682 , \25707 );
and \U$25713 ( \26028 , \25678 , \25707 );
or \U$25714 ( \26029 , \26026 , \26027 , \26028 );
and \U$25715 ( \26030 , \25729 , \25958 );
and \U$25716 ( \26031 , \25958 , \25973 );
and \U$25717 ( \26032 , \25729 , \25973 );
or \U$25718 ( \26033 , \26030 , \26031 , \26032 );
xor \U$25719 ( \26034 , \26029 , \26033 );
and \U$25720 ( \26035 , \25696 , \25700 );
and \U$25721 ( \26036 , \25700 , \25705 );
and \U$25722 ( \26037 , \25696 , \25705 );
or \U$25723 ( \26038 , \26035 , \26036 , \26037 );
and \U$25724 ( \26039 , \25790 , \25794 );
and \U$25725 ( \26040 , \25794 , \25799 );
and \U$25726 ( \26041 , \25790 , \25799 );
or \U$25727 ( \26042 , \26039 , \26040 , \26041 );
xor \U$25728 ( \26043 , \26038 , \26042 );
and \U$25729 ( \26044 , \25775 , \25779 );
and \U$25730 ( \26045 , \25779 , \25784 );
and \U$25731 ( \26046 , \25775 , \25784 );
or \U$25732 ( \26047 , \26044 , \26045 , \26046 );
xor \U$25733 ( \26048 , \26043 , \26047 );
and \U$25734 ( \26049 , \22429 , \22573 );
and \U$25735 ( \26050 , \22440 , \22571 );
nor \U$25736 ( \26051 , \26049 , \26050 );
xnor \U$25737 ( \26052 , \26051 , \22583 );
and \U$25738 ( \26053 , \22457 , \22598 );
and \U$25739 ( \26054 , \22468 , \22596 );
nor \U$25740 ( \26055 , \26053 , \26054 );
xnor \U$25741 ( \26056 , \26055 , \22608 );
xor \U$25742 ( \26057 , \26052 , \26056 );
and \U$25743 ( \26058 , \22478 , \22619 );
and \U$25744 ( \26059 , \22489 , \22617 );
nor \U$25745 ( \26060 , \26058 , \26059 );
xnor \U$25746 ( \26061 , \26060 , \22629 );
xor \U$25747 ( \26062 , \26057 , \26061 );
and \U$25748 ( \26063 , \22361 , \22506 );
and \U$25749 ( \26064 , \22372 , \22504 );
nor \U$25750 ( \26065 , \26063 , \26064 );
xnor \U$25751 ( \26066 , \26065 , \22516 );
and \U$25752 ( \26067 , \22386 , \22530 );
and \U$25753 ( \26068 , \22397 , \22528 );
nor \U$25754 ( \26069 , \26067 , \26068 );
xnor \U$25755 ( \26070 , \26069 , \22540 );
xor \U$25756 ( \26071 , \26066 , \26070 );
and \U$25757 ( \26072 , \22407 , \22551 );
and \U$25758 ( \26073 , \22418 , \22549 );
nor \U$25759 ( \26074 , \26072 , \26073 );
xnor \U$25760 ( \26075 , \26074 , \22561 );
xor \U$25761 ( \26076 , \26071 , \26075 );
xor \U$25762 ( \26077 , \26062 , \26076 );
and \U$25763 ( \26078 , \22294 , \22435 );
and \U$25764 ( \26079 , \22305 , \22433 );
nor \U$25765 ( \26080 , \26078 , \26079 );
xnor \U$25766 ( \26081 , \26080 , \22445 );
and \U$25767 ( \26082 , \22318 , \22463 );
and \U$25768 ( \26083 , \22329 , \22461 );
nor \U$25769 ( \26084 , \26082 , \26083 );
xnor \U$25770 ( \26085 , \26084 , \22473 );
xor \U$25771 ( \26086 , \26081 , \26085 );
and \U$25772 ( \26087 , \22339 , \22484 );
and \U$25773 ( \26088 , \22350 , \22482 );
nor \U$25774 ( \26089 , \26087 , \26088 );
xnor \U$25775 ( \26090 , \26089 , \22494 );
xor \U$25776 ( \26091 , \26086 , \26090 );
xor \U$25777 ( \26092 , \26077 , \26091 );
and \U$25778 ( \26093 , \22676 , \21978 );
and \U$25779 ( \26094 , \22567 , \22720 );
and \U$25780 ( \26095 , \22578 , \22707 );
nor \U$25781 ( \26096 , \26094 , \26095 );
xnor \U$25782 ( \26097 , \26096 , \22067 );
and \U$25783 ( \26098 , \22592 , \23173 );
and \U$25784 ( \26099 , \22603 , \22999 );
nor \U$25785 ( \26100 , \26098 , \26099 );
xnor \U$25786 ( \26101 , \26100 , \22016 );
xor \U$25787 ( \26102 , \26097 , \26101 );
and \U$25788 ( \26103 , \22613 , \22021 );
and \U$25789 ( \26104 , \22624 , \22019 );
nor \U$25790 ( \26105 , \26103 , \26104 );
xnor \U$25791 ( \26106 , \26105 , \21595 );
xor \U$25792 ( \26107 , \26102 , \26106 );
xor \U$25793 ( \26108 , \26093 , \26107 );
and \U$25794 ( \26109 , \22500 , \22641 );
and \U$25795 ( \26110 , \22511 , \22639 );
nor \U$25796 ( \26111 , \26109 , \26110 );
xnor \U$25797 ( \26112 , \26111 , \22651 );
and \U$25798 ( \26113 , \22524 , \22671 );
and \U$25799 ( \26114 , \22535 , \22669 );
nor \U$25800 ( \26115 , \26113 , \26114 );
xnor \U$25801 ( \26116 , \26115 , \22681 );
xor \U$25802 ( \26117 , \26112 , \26116 );
and \U$25803 ( \26118 , \22545 , \22691 );
and \U$25804 ( \26119 , \22556 , \22689 );
nor \U$25805 ( \26120 , \26118 , \26119 );
xnor \U$25806 ( \26121 , \26120 , \22701 );
xor \U$25807 ( \26122 , \26117 , \26121 );
xor \U$25808 ( \26123 , \26108 , \26122 );
xor \U$25809 ( \26124 , \26092 , \26123 );
and \U$25810 ( \26125 , \25894 , \25898 );
and \U$25811 ( \26126 , \25898 , \25903 );
and \U$25812 ( \26127 , \25894 , \25903 );
or \U$25813 ( \26128 , \26125 , \26126 , \26127 );
or \U$25814 ( \26129 , \25768 , \25769 );
xor \U$25815 ( \26130 , \26128 , \26129 );
and \U$25816 ( \26131 , \22635 , \21983 );
and \U$25817 ( \26132 , \22646 , \21981 );
nor \U$25818 ( \26133 , \26131 , \26132 );
xnor \U$25819 ( \26134 , \26133 , \21995 );
xor \U$25820 ( \26135 , \26130 , \26134 );
xor \U$25821 ( \26136 , \26124 , \26135 );
and \U$25822 ( \26137 , \25815 , \25829 );
and \U$25823 ( \26138 , \25829 , \25844 );
and \U$25824 ( \26139 , \25815 , \25844 );
or \U$25825 ( \26140 , \26137 , \26138 , \26139 );
and \U$25826 ( \26141 , \23230 , \22162 );
and \U$25827 ( \26142 , \23329 , \22160 );
nor \U$25828 ( \26143 , \26141 , \26142 );
xnor \U$25829 ( \26144 , \26143 , \22172 );
and \U$25830 ( \26145 , \22858 , \22187 );
and \U$25831 ( \26146 , \22894 , \22185 );
nor \U$25832 ( \26147 , \26145 , \26146 );
xnor \U$25833 ( \26148 , \26147 , \22197 );
xor \U$25834 ( \26149 , \26144 , \26148 );
and \U$25835 ( \26150 , \22071 , \22208 );
and \U$25836 ( \26151 , \22081 , \22206 );
nor \U$25837 ( \26152 , \26150 , \26151 );
xnor \U$25838 ( \26153 , \26152 , \22218 );
xor \U$25839 ( \26154 , \26149 , \26153 );
not \U$25840 ( \26155 , \22105 );
and \U$25841 ( \26156 , \21977 , \22119 );
and \U$25842 ( \26157 , \21990 , \22117 );
nor \U$25843 ( \26158 , \26156 , \26157 );
xnor \U$25844 ( \26159 , \26158 , \22129 );
xor \U$25845 ( \26160 , \26155 , \26159 );
and \U$25846 ( \26161 , \22030 , \22140 );
and \U$25847 ( \26162 , \22001 , \22138 );
nor \U$25848 ( \26163 , \26161 , \26162 );
xnor \U$25849 ( \26164 , \26163 , \22150 );
xor \U$25850 ( \26165 , \26160 , \26164 );
xor \U$25851 ( \26166 , \26154 , \26165 );
xor \U$25852 ( \26167 , \26140 , \26166 );
and \U$25853 ( \26168 , \22224 , \22367 );
and \U$25854 ( \26169 , \22235 , \22365 );
nor \U$25855 ( \26170 , \26168 , \26169 );
xnor \U$25856 ( \26171 , \26170 , \22377 );
and \U$25857 ( \26172 , \22251 , \22392 );
and \U$25858 ( \26173 , \22262 , \22390 );
nor \U$25859 ( \26174 , \26172 , \26173 );
xnor \U$25860 ( \26175 , \26174 , \22402 );
xor \U$25861 ( \26176 , \26171 , \26175 );
and \U$25862 ( \26177 , \22272 , \22413 );
and \U$25863 ( \26178 , \22283 , \22411 );
nor \U$25864 ( \26179 , \26177 , \26178 );
xnor \U$25865 ( \26180 , \26179 , \22423 );
xor \U$25866 ( \26181 , \26176 , \26180 );
and \U$25867 ( \26182 , \22156 , \22300 );
and \U$25868 ( \26183 , \22167 , \22298 );
nor \U$25869 ( \26184 , \26182 , \26183 );
xnor \U$25870 ( \26185 , \26184 , \22310 );
and \U$25871 ( \26186 , \22181 , \22324 );
and \U$25872 ( \26187 , \22192 , \22322 );
nor \U$25873 ( \26188 , \26186 , \26187 );
xnor \U$25874 ( \26189 , \26188 , \22334 );
xor \U$25875 ( \26190 , \26185 , \26189 );
and \U$25876 ( \26191 , \22202 , \22345 );
and \U$25877 ( \26192 , \22213 , \22343 );
nor \U$25878 ( \26193 , \26191 , \26192 );
xnor \U$25879 ( \26194 , \26193 , \22355 );
xor \U$25880 ( \26195 , \26190 , \26194 );
xor \U$25881 ( \26196 , \26181 , \26195 );
and \U$25882 ( \26197 , \22089 , \22230 );
and \U$25883 ( \26198 , \22100 , \22228 );
nor \U$25884 ( \26199 , \26197 , \26198 );
xnor \U$25885 ( \26200 , \26199 , \22240 );
and \U$25886 ( \26201 , \22113 , \22257 );
and \U$25887 ( \26202 , \22124 , \22255 );
nor \U$25888 ( \26203 , \26201 , \26202 );
xnor \U$25889 ( \26204 , \26203 , \22267 );
xor \U$25890 ( \26205 , \26200 , \26204 );
and \U$25891 ( \26206 , \22134 , \22278 );
and \U$25892 ( \26207 , \22145 , \22276 );
nor \U$25893 ( \26208 , \26206 , \26207 );
xnor \U$25894 ( \26209 , \26208 , \22288 );
xor \U$25895 ( \26210 , \26205 , \26209 );
xor \U$25896 ( \26211 , \26196 , \26210 );
xor \U$25897 ( \26212 , \26167 , \26211 );
xor \U$25898 ( \26213 , \26136 , \26212 );
and \U$25899 ( \26214 , \25759 , \25763 );
and \U$25900 ( \26215 , \25763 , \25770 );
and \U$25901 ( \26216 , \25759 , \25770 );
or \U$25902 ( \26217 , \26214 , \26215 , \26216 );
and \U$25903 ( \26218 , \25904 , \25918 );
and \U$25904 ( \26219 , \25918 , \25933 );
and \U$25905 ( \26220 , \25904 , \25933 );
or \U$25906 ( \26221 , \26218 , \26219 , \26220 );
xor \U$25907 ( \26222 , \26217 , \26221 );
and \U$25908 ( \26223 , \25859 , \25873 );
and \U$25909 ( \26224 , \25873 , \25888 );
and \U$25910 ( \26225 , \25859 , \25888 );
or \U$25911 ( \26226 , \26223 , \26224 , \26225 );
xor \U$25912 ( \26227 , \26222 , \26226 );
xor \U$25913 ( \26228 , \26213 , \26227 );
xor \U$25914 ( \26229 , \26048 , \26228 );
and \U$25915 ( \26230 , \25845 , \25889 );
and \U$25916 ( \26231 , \25889 , \25934 );
and \U$25917 ( \26232 , \25845 , \25934 );
or \U$25918 ( \26233 , \26230 , \26231 , \26232 );
and \U$25919 ( \26234 , \25771 , \25785 );
and \U$25920 ( \26235 , \25785 , \25800 );
and \U$25921 ( \26236 , \25771 , \25800 );
or \U$25922 ( \26237 , \26234 , \26235 , \26236 );
xor \U$25923 ( \26238 , \26233 , \26237 );
and \U$25924 ( \26239 , \25849 , \25853 );
and \U$25925 ( \26240 , \25853 , \25858 );
and \U$25926 ( \26241 , \25849 , \25858 );
or \U$25927 ( \26242 , \26239 , \26240 , \26241 );
and \U$25928 ( \26243 , \25923 , \25927 );
and \U$25929 ( \26244 , \25927 , \25932 );
and \U$25930 ( \26245 , \25923 , \25932 );
or \U$25931 ( \26246 , \26243 , \26244 , \26245 );
xor \U$25932 ( \26247 , \26242 , \26246 );
and \U$25933 ( \26248 , \25908 , \25912 );
and \U$25934 ( \26249 , \25912 , \25917 );
and \U$25935 ( \26250 , \25908 , \25917 );
or \U$25936 ( \26251 , \26248 , \26249 , \26250 );
xor \U$25937 ( \26252 , \26247 , \26251 );
and \U$25938 ( \26253 , \25805 , \25809 );
and \U$25939 ( \26254 , \25809 , \25814 );
and \U$25940 ( \26255 , \25805 , \25814 );
or \U$25941 ( \26256 , \26253 , \26254 , \26255 );
and \U$25942 ( \26257 , \25878 , \25882 );
and \U$25943 ( \26258 , \25882 , \25887 );
and \U$25944 ( \26259 , \25878 , \25887 );
or \U$25945 ( \26260 , \26257 , \26258 , \26259 );
xor \U$25946 ( \26261 , \26256 , \26260 );
and \U$25947 ( \26262 , \25863 , \25867 );
and \U$25948 ( \26263 , \25867 , \25872 );
and \U$25949 ( \26264 , \25863 , \25872 );
or \U$25950 ( \26265 , \26262 , \26263 , \26264 );
xor \U$25951 ( \26266 , \26261 , \26265 );
xor \U$25952 ( \26267 , \26252 , \26266 );
and \U$25953 ( \26268 , \25945 , \25949 );
and \U$25954 ( \26269 , \25949 , \25954 );
and \U$25955 ( \26270 , \25945 , \25954 );
or \U$25956 ( \26271 , \26268 , \26269 , \26270 );
and \U$25957 ( \26272 , \25834 , \25838 );
and \U$25958 ( \26273 , \25838 , \25843 );
and \U$25959 ( \26274 , \25834 , \25843 );
or \U$25960 ( \26275 , \26272 , \26273 , \26274 );
xor \U$25961 ( \26276 , \26271 , \26275 );
and \U$25962 ( \26277 , \25819 , \25823 );
and \U$25963 ( \26278 , \25823 , \25828 );
and \U$25964 ( \26279 , \25819 , \25828 );
or \U$25965 ( \26280 , \26277 , \26278 , \26279 );
xor \U$25966 ( \26281 , \26276 , \26280 );
xor \U$25967 ( \26282 , \26267 , \26281 );
xor \U$25968 ( \26283 , \26238 , \26282 );
xor \U$25969 ( \26284 , \26229 , \26283 );
xor \U$25970 ( \26285 , \26034 , \26284 );
xor \U$25971 ( \26286 , \26025 , \26285 );
and \U$25972 ( \26287 , \25674 , \25708 );
and \U$25973 ( \26288 , \25708 , \25975 );
and \U$25974 ( \26289 , \25674 , \25975 );
or \U$25975 ( \26290 , \26287 , \26288 , \26289 );
nor \U$25976 ( \26291 , \26286 , \26290 );
nor \U$25977 ( \26292 , \25981 , \26291 );
and \U$25978 ( \26293 , \26029 , \26033 );
and \U$25979 ( \26294 , \26033 , \26284 );
and \U$25980 ( \26295 , \26029 , \26284 );
or \U$25981 ( \26296 , \26293 , \26294 , \26295 );
and \U$25982 ( \26297 , \25999 , \26023 );
xor \U$25983 ( \26298 , \26296 , \26297 );
and \U$25984 ( \26299 , \26003 , \26007 );
and \U$25985 ( \26300 , \26007 , \26022 );
and \U$25986 ( \26301 , \26003 , \26022 );
or \U$25987 ( \26302 , \26299 , \26300 , \26301 );
and \U$25988 ( \26303 , \26271 , \26275 );
and \U$25989 ( \26304 , \26275 , \26280 );
and \U$25990 ( \26305 , \26271 , \26280 );
or \U$25991 ( \26306 , \26303 , \26304 , \26305 );
and \U$25992 ( \26307 , \26256 , \26260 );
and \U$25993 ( \26308 , \26260 , \26265 );
and \U$25994 ( \26309 , \26256 , \26265 );
or \U$25995 ( \26310 , \26307 , \26308 , \26309 );
xor \U$25996 ( \26311 , \26306 , \26310 );
and \U$25997 ( \26312 , \26242 , \26246 );
and \U$25998 ( \26313 , \26246 , \26251 );
and \U$25999 ( \26314 , \26242 , \26251 );
or \U$26000 ( \26315 , \26312 , \26313 , \26314 );
xor \U$26001 ( \26316 , \26311 , \26315 );
and \U$26002 ( \26317 , \22329 , \22463 );
and \U$26003 ( \26318 , \22294 , \22461 );
nor \U$26004 ( \26319 , \26317 , \26318 );
xnor \U$26005 ( \26320 , \26319 , \22473 );
and \U$26006 ( \26321 , \22350 , \22484 );
and \U$26007 ( \26322 , \22318 , \22482 );
nor \U$26008 ( \26323 , \26321 , \26322 );
xnor \U$26009 ( \26324 , \26323 , \22494 );
xor \U$26010 ( \26325 , \26320 , \26324 );
and \U$26011 ( \26326 , \22372 , \22506 );
and \U$26012 ( \26327 , \22339 , \22504 );
nor \U$26013 ( \26328 , \26326 , \26327 );
xnor \U$26014 ( \26329 , \26328 , \22516 );
xor \U$26015 ( \26330 , \26325 , \26329 );
and \U$26016 ( \26331 , \22262 , \22392 );
and \U$26017 ( \26332 , \22224 , \22390 );
nor \U$26018 ( \26333 , \26331 , \26332 );
xnor \U$26019 ( \26334 , \26333 , \22402 );
and \U$26020 ( \26335 , \22283 , \22413 );
and \U$26021 ( \26336 , \22251 , \22411 );
nor \U$26022 ( \26337 , \26335 , \26336 );
xnor \U$26023 ( \26338 , \26337 , \22423 );
xor \U$26024 ( \26339 , \26334 , \26338 );
and \U$26025 ( \26340 , \22305 , \22435 );
and \U$26026 ( \26341 , \22272 , \22433 );
nor \U$26027 ( \26342 , \26340 , \26341 );
xnor \U$26028 ( \26343 , \26342 , \22445 );
xor \U$26029 ( \26344 , \26339 , \26343 );
xor \U$26030 ( \26345 , \26330 , \26344 );
and \U$26031 ( \26346 , \22192 , \22324 );
and \U$26032 ( \26347 , \22156 , \22322 );
nor \U$26033 ( \26348 , \26346 , \26347 );
xnor \U$26034 ( \26349 , \26348 , \22334 );
and \U$26035 ( \26350 , \22213 , \22345 );
and \U$26036 ( \26351 , \22181 , \22343 );
nor \U$26037 ( \26352 , \26350 , \26351 );
xnor \U$26038 ( \26353 , \26352 , \22355 );
xor \U$26039 ( \26354 , \26349 , \26353 );
and \U$26040 ( \26355 , \22235 , \22367 );
and \U$26041 ( \26356 , \22202 , \22365 );
nor \U$26042 ( \26357 , \26355 , \26356 );
xnor \U$26043 ( \26358 , \26357 , \22377 );
xor \U$26044 ( \26359 , \26354 , \26358 );
xor \U$26045 ( \26360 , \26345 , \26359 );
and \U$26046 ( \26361 , \22535 , \22671 );
and \U$26047 ( \26362 , \22500 , \22669 );
nor \U$26048 ( \26363 , \26361 , \26362 );
xnor \U$26049 ( \26364 , \26363 , \22681 );
and \U$26050 ( \26365 , \22556 , \22691 );
and \U$26051 ( \26366 , \22524 , \22689 );
nor \U$26052 ( \26367 , \26365 , \26366 );
xnor \U$26053 ( \26368 , \26367 , \22701 );
xor \U$26054 ( \26369 , \26364 , \26368 );
and \U$26055 ( \26370 , \22578 , \22720 );
and \U$26056 ( \26371 , \22545 , \22707 );
nor \U$26057 ( \26372 , \26370 , \26371 );
xnor \U$26058 ( \26373 , \26372 , \22067 );
xor \U$26059 ( \26374 , \26369 , \26373 );
and \U$26060 ( \26375 , \22468 , \22598 );
and \U$26061 ( \26376 , \22429 , \22596 );
nor \U$26062 ( \26377 , \26375 , \26376 );
xnor \U$26063 ( \26378 , \26377 , \22608 );
and \U$26064 ( \26379 , \22489 , \22619 );
and \U$26065 ( \26380 , \22457 , \22617 );
nor \U$26066 ( \26381 , \26379 , \26380 );
xnor \U$26067 ( \26382 , \26381 , \22629 );
xor \U$26068 ( \26383 , \26378 , \26382 );
and \U$26069 ( \26384 , \22511 , \22641 );
and \U$26070 ( \26385 , \22478 , \22639 );
nor \U$26071 ( \26386 , \26384 , \26385 );
xnor \U$26072 ( \26387 , \26386 , \22651 );
xor \U$26073 ( \26388 , \26383 , \26387 );
xor \U$26074 ( \26389 , \26374 , \26388 );
and \U$26075 ( \26390 , \22397 , \22530 );
and \U$26076 ( \26391 , \22361 , \22528 );
nor \U$26077 ( \26392 , \26390 , \26391 );
xnor \U$26078 ( \26393 , \26392 , \22540 );
and \U$26079 ( \26394 , \22418 , \22551 );
and \U$26080 ( \26395 , \22386 , \22549 );
nor \U$26081 ( \26396 , \26394 , \26395 );
xnor \U$26082 ( \26397 , \26396 , \22561 );
xor \U$26083 ( \26398 , \26393 , \26397 );
and \U$26084 ( \26399 , \22440 , \22573 );
and \U$26085 ( \26400 , \22407 , \22571 );
nor \U$26086 ( \26401 , \26399 , \26400 );
xnor \U$26087 ( \26402 , \26401 , \22583 );
xor \U$26088 ( \26403 , \26398 , \26402 );
xor \U$26089 ( \26404 , \26389 , \26403 );
xor \U$26090 ( \26405 , \26360 , \26404 );
and \U$26091 ( \26406 , \26097 , \26101 );
and \U$26092 ( \26407 , \26101 , \26106 );
and \U$26093 ( \26408 , \26097 , \26106 );
or \U$26094 ( \26409 , \26406 , \26407 , \26408 );
and \U$26095 ( \26410 , \22635 , \21978 );
not \U$26096 ( \26411 , \26410 );
xor \U$26097 ( \26412 , \26409 , \26411 );
and \U$26098 ( \26413 , \22603 , \23173 );
and \U$26099 ( \26414 , \22567 , \22999 );
nor \U$26100 ( \26415 , \26413 , \26414 );
xnor \U$26101 ( \26416 , \26415 , \22016 );
and \U$26102 ( \26417 , \22624 , \22021 );
and \U$26103 ( \26418 , \22592 , \22019 );
nor \U$26104 ( \26419 , \26417 , \26418 );
xnor \U$26105 ( \26420 , \26419 , \21595 );
xor \U$26106 ( \26421 , \26416 , \26420 );
and \U$26107 ( \26422 , \22646 , \21983 );
and \U$26108 ( \26423 , \22613 , \21981 );
nor \U$26109 ( \26424 , \26422 , \26423 );
xnor \U$26110 ( \26425 , \26424 , \21995 );
xor \U$26111 ( \26426 , \26421 , \26425 );
xor \U$26112 ( \26427 , \26412 , \26426 );
xor \U$26113 ( \26428 , \26405 , \26427 );
and \U$26114 ( \26429 , \26181 , \26195 );
and \U$26115 ( \26430 , \26195 , \26210 );
and \U$26116 ( \26431 , \26181 , \26210 );
or \U$26117 ( \26432 , \26429 , \26430 , \26431 );
and \U$26118 ( \26433 , \26154 , \26165 );
xor \U$26119 ( \26434 , \26432 , \26433 );
and \U$26120 ( \26435 , \22124 , \22257 );
and \U$26121 ( \26436 , \22089 , \22255 );
nor \U$26122 ( \26437 , \26435 , \26436 );
xnor \U$26123 ( \26438 , \26437 , \22267 );
and \U$26124 ( \26439 , \22145 , \22278 );
and \U$26125 ( \26440 , \22113 , \22276 );
nor \U$26126 ( \26441 , \26439 , \26440 );
xnor \U$26127 ( \26442 , \26441 , \22288 );
xor \U$26128 ( \26443 , \26438 , \26442 );
and \U$26129 ( \26444 , \22167 , \22300 );
and \U$26130 ( \26445 , \22134 , \22298 );
nor \U$26131 ( \26446 , \26444 , \26445 );
xnor \U$26132 ( \26447 , \26446 , \22310 );
xor \U$26133 ( \26448 , \26443 , \26447 );
and \U$26134 ( \26449 , \22894 , \22187 );
and \U$26135 ( \26450 , \23230 , \22185 );
nor \U$26136 ( \26451 , \26449 , \26450 );
xnor \U$26137 ( \26452 , \26451 , \22197 );
and \U$26138 ( \26453 , \22081 , \22208 );
and \U$26139 ( \26454 , \22858 , \22206 );
nor \U$26140 ( \26455 , \26453 , \26454 );
xnor \U$26141 ( \26456 , \26455 , \22218 );
xor \U$26142 ( \26457 , \26452 , \26456 );
and \U$26143 ( \26458 , \22100 , \22230 );
and \U$26144 ( \26459 , \22071 , \22228 );
nor \U$26145 ( \26460 , \26458 , \26459 );
xnor \U$26146 ( \26461 , \26460 , \22240 );
xor \U$26147 ( \26462 , \26457 , \26461 );
xor \U$26148 ( \26463 , \26448 , \26462 );
and \U$26149 ( \26464 , \21990 , \22119 );
not \U$26150 ( \26465 , \26464 );
xnor \U$26151 ( \26466 , \26465 , \22129 );
and \U$26152 ( \26467 , \22001 , \22140 );
and \U$26153 ( \26468 , \21977 , \22138 );
nor \U$26154 ( \26469 , \26467 , \26468 );
xnor \U$26155 ( \26470 , \26469 , \22150 );
xor \U$26156 ( \26471 , \26466 , \26470 );
and \U$26157 ( \26472 , \23329 , \22162 );
and \U$26158 ( \26473 , \22030 , \22160 );
nor \U$26159 ( \26474 , \26472 , \26473 );
xnor \U$26160 ( \26475 , \26474 , \22172 );
xor \U$26161 ( \26476 , \26471 , \26475 );
xor \U$26162 ( \26477 , \26463 , \26476 );
xor \U$26163 ( \26478 , \26434 , \26477 );
xor \U$26164 ( \26479 , \26428 , \26478 );
and \U$26165 ( \26480 , \26128 , \26129 );
and \U$26166 ( \26481 , \26129 , \26134 );
and \U$26167 ( \26482 , \26128 , \26134 );
or \U$26168 ( \26483 , \26480 , \26481 , \26482 );
and \U$26169 ( \26484 , \26093 , \26107 );
and \U$26170 ( \26485 , \26107 , \26122 );
and \U$26171 ( \26486 , \26093 , \26122 );
or \U$26172 ( \26487 , \26484 , \26485 , \26486 );
xor \U$26173 ( \26488 , \26483 , \26487 );
and \U$26174 ( \26489 , \26062 , \26076 );
and \U$26175 ( \26490 , \26076 , \26091 );
and \U$26176 ( \26491 , \26062 , \26091 );
or \U$26177 ( \26492 , \26489 , \26490 , \26491 );
xor \U$26178 ( \26493 , \26488 , \26492 );
xor \U$26179 ( \26494 , \26479 , \26493 );
xor \U$26180 ( \26495 , \26316 , \26494 );
and \U$26181 ( \26496 , \26092 , \26123 );
and \U$26182 ( \26497 , \26123 , \26135 );
and \U$26183 ( \26498 , \26092 , \26135 );
or \U$26184 ( \26499 , \26496 , \26497 , \26498 );
and \U$26185 ( \26500 , \26252 , \26266 );
and \U$26186 ( \26501 , \26266 , \26281 );
and \U$26187 ( \26502 , \26252 , \26281 );
or \U$26188 ( \26503 , \26500 , \26501 , \26502 );
xor \U$26189 ( \26504 , \26499 , \26503 );
and \U$26190 ( \26505 , \26066 , \26070 );
and \U$26191 ( \26506 , \26070 , \26075 );
and \U$26192 ( \26507 , \26066 , \26075 );
or \U$26193 ( \26508 , \26505 , \26506 , \26507 );
and \U$26194 ( \26509 , \26052 , \26056 );
and \U$26195 ( \26510 , \26056 , \26061 );
and \U$26196 ( \26511 , \26052 , \26061 );
or \U$26197 ( \26512 , \26509 , \26510 , \26511 );
xor \U$26198 ( \26513 , \26508 , \26512 );
and \U$26199 ( \26514 , \26112 , \26116 );
and \U$26200 ( \26515 , \26116 , \26121 );
and \U$26201 ( \26516 , \26112 , \26121 );
or \U$26202 ( \26517 , \26514 , \26515 , \26516 );
xor \U$26203 ( \26518 , \26513 , \26517 );
and \U$26204 ( \26519 , \26185 , \26189 );
and \U$26205 ( \26520 , \26189 , \26194 );
and \U$26206 ( \26521 , \26185 , \26194 );
or \U$26207 ( \26522 , \26519 , \26520 , \26521 );
and \U$26208 ( \26523 , \26171 , \26175 );
and \U$26209 ( \26524 , \26175 , \26180 );
and \U$26210 ( \26525 , \26171 , \26180 );
or \U$26211 ( \26526 , \26523 , \26524 , \26525 );
xor \U$26212 ( \26527 , \26522 , \26526 );
and \U$26213 ( \26528 , \26081 , \26085 );
and \U$26214 ( \26529 , \26085 , \26090 );
and \U$26215 ( \26530 , \26081 , \26090 );
or \U$26216 ( \26531 , \26528 , \26529 , \26530 );
xor \U$26217 ( \26532 , \26527 , \26531 );
xor \U$26218 ( \26533 , \26518 , \26532 );
and \U$26219 ( \26534 , \26155 , \26159 );
and \U$26220 ( \26535 , \26159 , \26164 );
and \U$26221 ( \26536 , \26155 , \26164 );
or \U$26222 ( \26537 , \26534 , \26535 , \26536 );
and \U$26223 ( \26538 , \26144 , \26148 );
and \U$26224 ( \26539 , \26148 , \26153 );
and \U$26225 ( \26540 , \26144 , \26153 );
or \U$26226 ( \26541 , \26538 , \26539 , \26540 );
xor \U$26227 ( \26542 , \26537 , \26541 );
and \U$26228 ( \26543 , \26200 , \26204 );
and \U$26229 ( \26544 , \26204 , \26209 );
and \U$26230 ( \26545 , \26200 , \26209 );
or \U$26231 ( \26546 , \26543 , \26544 , \26545 );
xor \U$26232 ( \26547 , \26542 , \26546 );
xor \U$26233 ( \26548 , \26533 , \26547 );
xor \U$26234 ( \26549 , \26504 , \26548 );
xor \U$26235 ( \26550 , \26495 , \26549 );
and \U$26236 ( \26551 , \26012 , \26016 );
and \U$26237 ( \26552 , \26016 , \26021 );
and \U$26238 ( \26553 , \26012 , \26021 );
or \U$26239 ( \26554 , \26551 , \26552 , \26553 );
and \U$26240 ( \26555 , \26233 , \26237 );
and \U$26241 ( \26556 , \26237 , \26282 );
and \U$26242 ( \26557 , \26233 , \26282 );
or \U$26243 ( \26558 , \26555 , \26556 , \26557 );
xor \U$26244 ( \26559 , \26554 , \26558 );
and \U$26245 ( \26560 , \26136 , \26212 );
and \U$26246 ( \26561 , \26212 , \26227 );
and \U$26247 ( \26562 , \26136 , \26227 );
or \U$26248 ( \26563 , \26560 , \26561 , \26562 );
xor \U$26249 ( \26564 , \26559 , \26563 );
xor \U$26250 ( \26565 , \26550 , \26564 );
xor \U$26251 ( \26566 , \26302 , \26565 );
and \U$26252 ( \26567 , \25989 , \25993 );
and \U$26253 ( \26568 , \25993 , \25998 );
and \U$26254 ( \26569 , \25989 , \25998 );
or \U$26255 ( \26570 , \26567 , \26568 , \26569 );
and \U$26256 ( \26571 , \26048 , \26228 );
and \U$26257 ( \26572 , \26228 , \26283 );
and \U$26258 ( \26573 , \26048 , \26283 );
or \U$26259 ( \26574 , \26571 , \26572 , \26573 );
xor \U$26260 ( \26575 , \26570 , \26574 );
and \U$26261 ( \26576 , \26038 , \26042 );
and \U$26262 ( \26577 , \26042 , \26047 );
and \U$26263 ( \26578 , \26038 , \26047 );
or \U$26264 ( \26579 , \26576 , \26577 , \26578 );
and \U$26265 ( \26580 , \26217 , \26221 );
and \U$26266 ( \26581 , \26221 , \26226 );
and \U$26267 ( \26582 , \26217 , \26226 );
or \U$26268 ( \26583 , \26580 , \26581 , \26582 );
xor \U$26269 ( \26584 , \26579 , \26583 );
and \U$26270 ( \26585 , \26140 , \26166 );
and \U$26271 ( \26586 , \26166 , \26211 );
and \U$26272 ( \26587 , \26140 , \26211 );
or \U$26273 ( \26588 , \26585 , \26586 , \26587 );
xor \U$26274 ( \26589 , \26584 , \26588 );
xor \U$26275 ( \26590 , \26575 , \26589 );
xor \U$26276 ( \26591 , \26566 , \26590 );
xor \U$26277 ( \26592 , \26298 , \26591 );
and \U$26278 ( \26593 , \25985 , \26024 );
and \U$26279 ( \26594 , \26024 , \26285 );
and \U$26280 ( \26595 , \25985 , \26285 );
or \U$26281 ( \26596 , \26593 , \26594 , \26595 );
nor \U$26282 ( \26597 , \26592 , \26596 );
and \U$26283 ( \26598 , \26302 , \26565 );
and \U$26284 ( \26599 , \26565 , \26590 );
and \U$26285 ( \26600 , \26302 , \26590 );
or \U$26286 ( \26601 , \26598 , \26599 , \26600 );
and \U$26287 ( \26602 , \26579 , \26583 );
and \U$26288 ( \26603 , \26583 , \26588 );
and \U$26289 ( \26604 , \26579 , \26588 );
or \U$26290 ( \26605 , \26602 , \26603 , \26604 );
and \U$26291 ( \26606 , \26499 , \26503 );
and \U$26292 ( \26607 , \26503 , \26548 );
and \U$26293 ( \26608 , \26499 , \26548 );
or \U$26294 ( \26609 , \26606 , \26607 , \26608 );
xor \U$26295 ( \26610 , \26605 , \26609 );
and \U$26296 ( \26611 , \26428 , \26478 );
and \U$26297 ( \26612 , \26478 , \26493 );
and \U$26298 ( \26613 , \26428 , \26493 );
or \U$26299 ( \26614 , \26611 , \26612 , \26613 );
xor \U$26300 ( \26615 , \26610 , \26614 );
and \U$26301 ( \26616 , \26554 , \26558 );
and \U$26302 ( \26617 , \26558 , \26563 );
and \U$26303 ( \26618 , \26554 , \26563 );
or \U$26304 ( \26619 , \26616 , \26617 , \26618 );
and \U$26305 ( \26620 , \26316 , \26494 );
and \U$26306 ( \26621 , \26494 , \26549 );
and \U$26307 ( \26622 , \26316 , \26549 );
or \U$26308 ( \26623 , \26620 , \26621 , \26622 );
xor \U$26309 ( \26624 , \26619 , \26623 );
and \U$26310 ( \26625 , \26306 , \26310 );
and \U$26311 ( \26626 , \26310 , \26315 );
and \U$26312 ( \26627 , \26306 , \26315 );
or \U$26313 ( \26628 , \26625 , \26626 , \26627 );
and \U$26314 ( \26629 , \26483 , \26487 );
and \U$26315 ( \26630 , \26487 , \26492 );
and \U$26316 ( \26631 , \26483 , \26492 );
or \U$26317 ( \26632 , \26629 , \26630 , \26631 );
xor \U$26318 ( \26633 , \26628 , \26632 );
and \U$26319 ( \26634 , \26432 , \26433 );
and \U$26320 ( \26635 , \26433 , \26477 );
and \U$26321 ( \26636 , \26432 , \26477 );
or \U$26322 ( \26637 , \26634 , \26635 , \26636 );
xor \U$26323 ( \26638 , \26633 , \26637 );
xor \U$26324 ( \26639 , \26624 , \26638 );
xor \U$26325 ( \26640 , \26615 , \26639 );
xor \U$26326 ( \26641 , \26601 , \26640 );
and \U$26327 ( \26642 , \26570 , \26574 );
and \U$26328 ( \26643 , \26574 , \26589 );
and \U$26329 ( \26644 , \26570 , \26589 );
or \U$26330 ( \26645 , \26642 , \26643 , \26644 );
and \U$26331 ( \26646 , \26550 , \26564 );
xor \U$26332 ( \26647 , \26645 , \26646 );
and \U$26333 ( \26648 , \26537 , \26541 );
and \U$26334 ( \26649 , \26541 , \26546 );
and \U$26335 ( \26650 , \26537 , \26546 );
or \U$26336 ( \26651 , \26648 , \26649 , \26650 );
and \U$26337 ( \26652 , \26522 , \26526 );
and \U$26338 ( \26653 , \26526 , \26531 );
and \U$26339 ( \26654 , \26522 , \26531 );
or \U$26340 ( \26655 , \26652 , \26653 , \26654 );
xor \U$26341 ( \26656 , \26651 , \26655 );
and \U$26342 ( \26657 , \26508 , \26512 );
and \U$26343 ( \26658 , \26512 , \26517 );
and \U$26344 ( \26659 , \26508 , \26517 );
or \U$26345 ( \26660 , \26657 , \26658 , \26659 );
xor \U$26346 ( \26661 , \26656 , \26660 );
and \U$26347 ( \26662 , \22361 , \22530 );
and \U$26348 ( \26663 , \22372 , \22528 );
nor \U$26349 ( \26664 , \26662 , \26663 );
xnor \U$26350 ( \26665 , \26664 , \22540 );
and \U$26351 ( \26666 , \22386 , \22551 );
and \U$26352 ( \26667 , \22397 , \22549 );
nor \U$26353 ( \26668 , \26666 , \26667 );
xnor \U$26354 ( \26669 , \26668 , \22561 );
xor \U$26355 ( \26670 , \26665 , \26669 );
and \U$26356 ( \26671 , \22407 , \22573 );
and \U$26357 ( \26672 , \22418 , \22571 );
nor \U$26358 ( \26673 , \26671 , \26672 );
xnor \U$26359 ( \26674 , \26673 , \22583 );
xor \U$26360 ( \26675 , \26670 , \26674 );
and \U$26361 ( \26676 , \22294 , \22463 );
and \U$26362 ( \26677 , \22305 , \22461 );
nor \U$26363 ( \26678 , \26676 , \26677 );
xnor \U$26364 ( \26679 , \26678 , \22473 );
and \U$26365 ( \26680 , \22318 , \22484 );
and \U$26366 ( \26681 , \22329 , \22482 );
nor \U$26367 ( \26682 , \26680 , \26681 );
xnor \U$26368 ( \26683 , \26682 , \22494 );
xor \U$26369 ( \26684 , \26679 , \26683 );
and \U$26370 ( \26685 , \22339 , \22506 );
and \U$26371 ( \26686 , \22350 , \22504 );
nor \U$26372 ( \26687 , \26685 , \26686 );
xnor \U$26373 ( \26688 , \26687 , \22516 );
xor \U$26374 ( \26689 , \26684 , \26688 );
xor \U$26375 ( \26690 , \26675 , \26689 );
and \U$26376 ( \26691 , \22224 , \22392 );
and \U$26377 ( \26692 , \22235 , \22390 );
nor \U$26378 ( \26693 , \26691 , \26692 );
xnor \U$26379 ( \26694 , \26693 , \22402 );
and \U$26380 ( \26695 , \22251 , \22413 );
and \U$26381 ( \26696 , \22262 , \22411 );
nor \U$26382 ( \26697 , \26695 , \26696 );
xnor \U$26383 ( \26698 , \26697 , \22423 );
xor \U$26384 ( \26699 , \26694 , \26698 );
and \U$26385 ( \26700 , \22272 , \22435 );
and \U$26386 ( \26701 , \22283 , \22433 );
nor \U$26387 ( \26702 , \26700 , \26701 );
xnor \U$26388 ( \26703 , \26702 , \22445 );
xor \U$26389 ( \26704 , \26699 , \26703 );
xor \U$26390 ( \26705 , \26690 , \26704 );
and \U$26391 ( \26706 , \22567 , \23173 );
and \U$26392 ( \26707 , \22578 , \22999 );
nor \U$26393 ( \26708 , \26706 , \26707 );
xnor \U$26394 ( \26709 , \26708 , \22016 );
and \U$26395 ( \26710 , \22592 , \22021 );
and \U$26396 ( \26711 , \22603 , \22019 );
nor \U$26397 ( \26712 , \26710 , \26711 );
xnor \U$26398 ( \26713 , \26712 , \21595 );
xor \U$26399 ( \26714 , \26709 , \26713 );
and \U$26400 ( \26715 , \22613 , \21983 );
and \U$26401 ( \26716 , \22624 , \21981 );
nor \U$26402 ( \26717 , \26715 , \26716 );
xnor \U$26403 ( \26718 , \26717 , \21995 );
xor \U$26404 ( \26719 , \26714 , \26718 );
and \U$26405 ( \26720 , \22500 , \22671 );
and \U$26406 ( \26721 , \22511 , \22669 );
nor \U$26407 ( \26722 , \26720 , \26721 );
xnor \U$26408 ( \26723 , \26722 , \22681 );
and \U$26409 ( \26724 , \22524 , \22691 );
and \U$26410 ( \26725 , \22535 , \22689 );
nor \U$26411 ( \26726 , \26724 , \26725 );
xnor \U$26412 ( \26727 , \26726 , \22701 );
xor \U$26413 ( \26728 , \26723 , \26727 );
and \U$26414 ( \26729 , \22545 , \22720 );
and \U$26415 ( \26730 , \22556 , \22707 );
nor \U$26416 ( \26731 , \26729 , \26730 );
xnor \U$26417 ( \26732 , \26731 , \22067 );
xor \U$26418 ( \26733 , \26728 , \26732 );
xor \U$26419 ( \26734 , \26719 , \26733 );
and \U$26420 ( \26735 , \22429 , \22598 );
and \U$26421 ( \26736 , \22440 , \22596 );
nor \U$26422 ( \26737 , \26735 , \26736 );
xnor \U$26423 ( \26738 , \26737 , \22608 );
and \U$26424 ( \26739 , \22457 , \22619 );
and \U$26425 ( \26740 , \22468 , \22617 );
nor \U$26426 ( \26741 , \26739 , \26740 );
xnor \U$26427 ( \26742 , \26741 , \22629 );
xor \U$26428 ( \26743 , \26738 , \26742 );
and \U$26429 ( \26744 , \22478 , \22641 );
and \U$26430 ( \26745 , \22489 , \22639 );
nor \U$26431 ( \26746 , \26744 , \26745 );
xnor \U$26432 ( \26747 , \26746 , \22651 );
xor \U$26433 ( \26748 , \26743 , \26747 );
xor \U$26434 ( \26749 , \26734 , \26748 );
xor \U$26435 ( \26750 , \26705 , \26749 );
and \U$26436 ( \26751 , \26416 , \26420 );
and \U$26437 ( \26752 , \26420 , \26425 );
and \U$26438 ( \26753 , \26416 , \26425 );
or \U$26439 ( \26754 , \26751 , \26752 , \26753 );
xor \U$26440 ( \26755 , \26754 , \26410 );
and \U$26441 ( \26756 , \22646 , \21978 );
xor \U$26442 ( \26757 , \26755 , \26756 );
xor \U$26443 ( \26758 , \26750 , \26757 );
and \U$26444 ( \26759 , \26448 , \26462 );
and \U$26445 ( \26760 , \26462 , \26476 );
and \U$26446 ( \26761 , \26448 , \26476 );
or \U$26447 ( \26762 , \26759 , \26760 , \26761 );
not \U$26448 ( \26763 , \22129 );
and \U$26449 ( \26764 , \21977 , \22140 );
and \U$26450 ( \26765 , \21990 , \22138 );
nor \U$26451 ( \26766 , \26764 , \26765 );
xnor \U$26452 ( \26767 , \26766 , \22150 );
xor \U$26453 ( \26768 , \26763 , \26767 );
and \U$26454 ( \26769 , \22030 , \22162 );
and \U$26455 ( \26770 , \22001 , \22160 );
nor \U$26456 ( \26771 , \26769 , \26770 );
xnor \U$26457 ( \26772 , \26771 , \22172 );
xor \U$26458 ( \26773 , \26768 , \26772 );
xor \U$26459 ( \26774 , \26762 , \26773 );
and \U$26460 ( \26775 , \22156 , \22324 );
and \U$26461 ( \26776 , \22167 , \22322 );
nor \U$26462 ( \26777 , \26775 , \26776 );
xnor \U$26463 ( \26778 , \26777 , \22334 );
and \U$26464 ( \26779 , \22181 , \22345 );
and \U$26465 ( \26780 , \22192 , \22343 );
nor \U$26466 ( \26781 , \26779 , \26780 );
xnor \U$26467 ( \26782 , \26781 , \22355 );
xor \U$26468 ( \26783 , \26778 , \26782 );
and \U$26469 ( \26784 , \22202 , \22367 );
and \U$26470 ( \26785 , \22213 , \22365 );
nor \U$26471 ( \26786 , \26784 , \26785 );
xnor \U$26472 ( \26787 , \26786 , \22377 );
xor \U$26473 ( \26788 , \26783 , \26787 );
and \U$26474 ( \26789 , \22089 , \22257 );
and \U$26475 ( \26790 , \22100 , \22255 );
nor \U$26476 ( \26791 , \26789 , \26790 );
xnor \U$26477 ( \26792 , \26791 , \22267 );
and \U$26478 ( \26793 , \22113 , \22278 );
and \U$26479 ( \26794 , \22124 , \22276 );
nor \U$26480 ( \26795 , \26793 , \26794 );
xnor \U$26481 ( \26796 , \26795 , \22288 );
xor \U$26482 ( \26797 , \26792 , \26796 );
and \U$26483 ( \26798 , \22134 , \22300 );
and \U$26484 ( \26799 , \22145 , \22298 );
nor \U$26485 ( \26800 , \26798 , \26799 );
xnor \U$26486 ( \26801 , \26800 , \22310 );
xor \U$26487 ( \26802 , \26797 , \26801 );
xor \U$26488 ( \26803 , \26788 , \26802 );
and \U$26489 ( \26804 , \23230 , \22187 );
and \U$26490 ( \26805 , \23329 , \22185 );
nor \U$26491 ( \26806 , \26804 , \26805 );
xnor \U$26492 ( \26807 , \26806 , \22197 );
and \U$26493 ( \26808 , \22858 , \22208 );
and \U$26494 ( \26809 , \22894 , \22206 );
nor \U$26495 ( \26810 , \26808 , \26809 );
xnor \U$26496 ( \26811 , \26810 , \22218 );
xor \U$26497 ( \26812 , \26807 , \26811 );
and \U$26498 ( \26813 , \22071 , \22230 );
and \U$26499 ( \26814 , \22081 , \22228 );
nor \U$26500 ( \26815 , \26813 , \26814 );
xnor \U$26501 ( \26816 , \26815 , \22240 );
xor \U$26502 ( \26817 , \26812 , \26816 );
xor \U$26503 ( \26818 , \26803 , \26817 );
xor \U$26504 ( \26819 , \26774 , \26818 );
xor \U$26505 ( \26820 , \26758 , \26819 );
and \U$26506 ( \26821 , \26409 , \26411 );
and \U$26507 ( \26822 , \26411 , \26426 );
and \U$26508 ( \26823 , \26409 , \26426 );
or \U$26509 ( \26824 , \26821 , \26822 , \26823 );
and \U$26510 ( \26825 , \26374 , \26388 );
and \U$26511 ( \26826 , \26388 , \26403 );
and \U$26512 ( \26827 , \26374 , \26403 );
or \U$26513 ( \26828 , \26825 , \26826 , \26827 );
xor \U$26514 ( \26829 , \26824 , \26828 );
and \U$26515 ( \26830 , \26330 , \26344 );
and \U$26516 ( \26831 , \26344 , \26359 );
and \U$26517 ( \26832 , \26330 , \26359 );
or \U$26518 ( \26833 , \26830 , \26831 , \26832 );
xor \U$26519 ( \26834 , \26829 , \26833 );
xor \U$26520 ( \26835 , \26820 , \26834 );
xor \U$26521 ( \26836 , \26661 , \26835 );
and \U$26522 ( \26837 , \26360 , \26404 );
and \U$26523 ( \26838 , \26404 , \26427 );
and \U$26524 ( \26839 , \26360 , \26427 );
or \U$26525 ( \26840 , \26837 , \26838 , \26839 );
and \U$26526 ( \26841 , \26518 , \26532 );
and \U$26527 ( \26842 , \26532 , \26547 );
and \U$26528 ( \26843 , \26518 , \26547 );
or \U$26529 ( \26844 , \26841 , \26842 , \26843 );
xor \U$26530 ( \26845 , \26840 , \26844 );
and \U$26531 ( \26846 , \26393 , \26397 );
and \U$26532 ( \26847 , \26397 , \26402 );
and \U$26533 ( \26848 , \26393 , \26402 );
or \U$26534 ( \26849 , \26846 , \26847 , \26848 );
and \U$26535 ( \26850 , \26378 , \26382 );
and \U$26536 ( \26851 , \26382 , \26387 );
and \U$26537 ( \26852 , \26378 , \26387 );
or \U$26538 ( \26853 , \26850 , \26851 , \26852 );
xor \U$26539 ( \26854 , \26849 , \26853 );
and \U$26540 ( \26855 , \26364 , \26368 );
and \U$26541 ( \26856 , \26368 , \26373 );
and \U$26542 ( \26857 , \26364 , \26373 );
or \U$26543 ( \26858 , \26855 , \26856 , \26857 );
xor \U$26544 ( \26859 , \26854 , \26858 );
and \U$26545 ( \26860 , \26349 , \26353 );
and \U$26546 ( \26861 , \26353 , \26358 );
and \U$26547 ( \26862 , \26349 , \26358 );
or \U$26548 ( \26863 , \26860 , \26861 , \26862 );
and \U$26549 ( \26864 , \26334 , \26338 );
and \U$26550 ( \26865 , \26338 , \26343 );
and \U$26551 ( \26866 , \26334 , \26343 );
or \U$26552 ( \26867 , \26864 , \26865 , \26866 );
xor \U$26553 ( \26868 , \26863 , \26867 );
and \U$26554 ( \26869 , \26320 , \26324 );
and \U$26555 ( \26870 , \26324 , \26329 );
and \U$26556 ( \26871 , \26320 , \26329 );
or \U$26557 ( \26872 , \26869 , \26870 , \26871 );
xor \U$26558 ( \26873 , \26868 , \26872 );
xor \U$26559 ( \26874 , \26859 , \26873 );
and \U$26560 ( \26875 , \26466 , \26470 );
and \U$26561 ( \26876 , \26470 , \26475 );
and \U$26562 ( \26877 , \26466 , \26475 );
or \U$26563 ( \26878 , \26875 , \26876 , \26877 );
and \U$26564 ( \26879 , \26452 , \26456 );
and \U$26565 ( \26880 , \26456 , \26461 );
and \U$26566 ( \26881 , \26452 , \26461 );
or \U$26567 ( \26882 , \26879 , \26880 , \26881 );
xor \U$26568 ( \26883 , \26878 , \26882 );
and \U$26569 ( \26884 , \26438 , \26442 );
and \U$26570 ( \26885 , \26442 , \26447 );
and \U$26571 ( \26886 , \26438 , \26447 );
or \U$26572 ( \26887 , \26884 , \26885 , \26886 );
xor \U$26573 ( \26888 , \26883 , \26887 );
xor \U$26574 ( \26889 , \26874 , \26888 );
xor \U$26575 ( \26890 , \26845 , \26889 );
xor \U$26576 ( \26891 , \26836 , \26890 );
xor \U$26577 ( \26892 , \26647 , \26891 );
xor \U$26578 ( \26893 , \26641 , \26892 );
and \U$26579 ( \26894 , \26296 , \26297 );
and \U$26580 ( \26895 , \26297 , \26591 );
and \U$26581 ( \26896 , \26296 , \26591 );
or \U$26582 ( \26897 , \26894 , \26895 , \26896 );
nor \U$26583 ( \26898 , \26893 , \26897 );
nor \U$26584 ( \26899 , \26597 , \26898 );
nand \U$26585 ( \26900 , \26292 , \26899 );
nor \U$26586 ( \26901 , \25670 , \26900 );
and \U$26587 ( \26902 , \26645 , \26646 );
and \U$26588 ( \26903 , \26646 , \26891 );
and \U$26589 ( \26904 , \26645 , \26891 );
or \U$26590 ( \26905 , \26902 , \26903 , \26904 );
and \U$26591 ( \26906 , \26615 , \26639 );
xor \U$26592 ( \26907 , \26905 , \26906 );
and \U$26593 ( \26908 , \26619 , \26623 );
and \U$26594 ( \26909 , \26623 , \26638 );
and \U$26595 ( \26910 , \26619 , \26638 );
or \U$26596 ( \26911 , \26908 , \26909 , \26910 );
and \U$26597 ( \26912 , \26651 , \26655 );
and \U$26598 ( \26913 , \26655 , \26660 );
and \U$26599 ( \26914 , \26651 , \26660 );
or \U$26600 ( \26915 , \26912 , \26913 , \26914 );
and \U$26601 ( \26916 , \26824 , \26828 );
and \U$26602 ( \26917 , \26828 , \26833 );
and \U$26603 ( \26918 , \26824 , \26833 );
or \U$26604 ( \26919 , \26916 , \26917 , \26918 );
xor \U$26605 ( \26920 , \26915 , \26919 );
and \U$26606 ( \26921 , \26762 , \26773 );
and \U$26607 ( \26922 , \26773 , \26818 );
and \U$26608 ( \26923 , \26762 , \26818 );
or \U$26609 ( \26924 , \26921 , \26922 , \26923 );
xor \U$26610 ( \26925 , \26920 , \26924 );
and \U$26611 ( \26926 , \26754 , \26410 );
and \U$26612 ( \26927 , \26410 , \26756 );
and \U$26613 ( \26928 , \26754 , \26756 );
or \U$26614 ( \26929 , \26926 , \26927 , \26928 );
and \U$26615 ( \26930 , \26719 , \26733 );
and \U$26616 ( \26931 , \26733 , \26748 );
and \U$26617 ( \26932 , \26719 , \26748 );
or \U$26618 ( \26933 , \26930 , \26931 , \26932 );
xor \U$26619 ( \26934 , \26929 , \26933 );
and \U$26620 ( \26935 , \26675 , \26689 );
and \U$26621 ( \26936 , \26689 , \26704 );
and \U$26622 ( \26937 , \26675 , \26704 );
or \U$26623 ( \26938 , \26935 , \26936 , \26937 );
xor \U$26624 ( \26939 , \26934 , \26938 );
and \U$26625 ( \26940 , \26878 , \26882 );
and \U$26626 ( \26941 , \26882 , \26887 );
and \U$26627 ( \26942 , \26878 , \26887 );
or \U$26628 ( \26943 , \26940 , \26941 , \26942 );
and \U$26629 ( \26944 , \26863 , \26867 );
and \U$26630 ( \26945 , \26867 , \26872 );
and \U$26631 ( \26946 , \26863 , \26872 );
or \U$26632 ( \26947 , \26944 , \26945 , \26946 );
xor \U$26633 ( \26948 , \26943 , \26947 );
and \U$26634 ( \26949 , \26849 , \26853 );
and \U$26635 ( \26950 , \26853 , \26858 );
and \U$26636 ( \26951 , \26849 , \26858 );
or \U$26637 ( \26952 , \26949 , \26950 , \26951 );
xor \U$26638 ( \26953 , \26948 , \26952 );
xor \U$26639 ( \26954 , \26939 , \26953 );
and \U$26640 ( \26955 , \26763 , \26767 );
and \U$26641 ( \26956 , \26767 , \26772 );
and \U$26642 ( \26957 , \26763 , \26772 );
or \U$26643 ( \26958 , \26955 , \26956 , \26957 );
and \U$26644 ( \26959 , \26807 , \26811 );
and \U$26645 ( \26960 , \26811 , \26816 );
and \U$26646 ( \26961 , \26807 , \26816 );
or \U$26647 ( \26962 , \26959 , \26960 , \26961 );
xor \U$26648 ( \26963 , \26958 , \26962 );
and \U$26649 ( \26964 , \26792 , \26796 );
and \U$26650 ( \26965 , \26796 , \26801 );
and \U$26651 ( \26966 , \26792 , \26801 );
or \U$26652 ( \26967 , \26964 , \26965 , \26966 );
xor \U$26653 ( \26968 , \26963 , \26967 );
and \U$26654 ( \26969 , \22535 , \22691 );
and \U$26655 ( \26970 , \22500 , \22689 );
nor \U$26656 ( \26971 , \26969 , \26970 );
xnor \U$26657 ( \26972 , \26971 , \22701 );
and \U$26658 ( \26973 , \22556 , \22720 );
and \U$26659 ( \26974 , \22524 , \22707 );
nor \U$26660 ( \26975 , \26973 , \26974 );
xnor \U$26661 ( \26976 , \26975 , \22067 );
xor \U$26662 ( \26977 , \26972 , \26976 );
and \U$26663 ( \26978 , \22578 , \23173 );
and \U$26664 ( \26979 , \22545 , \22999 );
nor \U$26665 ( \26980 , \26978 , \26979 );
xnor \U$26666 ( \26981 , \26980 , \22016 );
xor \U$26667 ( \26982 , \26977 , \26981 );
and \U$26668 ( \26983 , \22468 , \22619 );
and \U$26669 ( \26984 , \22429 , \22617 );
nor \U$26670 ( \26985 , \26983 , \26984 );
xnor \U$26671 ( \26986 , \26985 , \22629 );
and \U$26672 ( \26987 , \22489 , \22641 );
and \U$26673 ( \26988 , \22457 , \22639 );
nor \U$26674 ( \26989 , \26987 , \26988 );
xnor \U$26675 ( \26990 , \26989 , \22651 );
xor \U$26676 ( \26991 , \26986 , \26990 );
and \U$26677 ( \26992 , \22511 , \22671 );
and \U$26678 ( \26993 , \22478 , \22669 );
nor \U$26679 ( \26994 , \26992 , \26993 );
xnor \U$26680 ( \26995 , \26994 , \22681 );
xor \U$26681 ( \26996 , \26991 , \26995 );
xor \U$26682 ( \26997 , \26982 , \26996 );
and \U$26683 ( \26998 , \22397 , \22551 );
and \U$26684 ( \26999 , \22361 , \22549 );
nor \U$26685 ( \27000 , \26998 , \26999 );
xnor \U$26686 ( \27001 , \27000 , \22561 );
and \U$26687 ( \27002 , \22418 , \22573 );
and \U$26688 ( \27003 , \22386 , \22571 );
nor \U$26689 ( \27004 , \27002 , \27003 );
xnor \U$26690 ( \27005 , \27004 , \22583 );
xor \U$26691 ( \27006 , \27001 , \27005 );
and \U$26692 ( \27007 , \22440 , \22598 );
and \U$26693 ( \27008 , \22407 , \22596 );
nor \U$26694 ( \27009 , \27007 , \27008 );
xnor \U$26695 ( \27010 , \27009 , \22608 );
xor \U$26696 ( \27011 , \27006 , \27010 );
xor \U$26697 ( \27012 , \26997 , \27011 );
and \U$26698 ( \27013 , \26709 , \26713 );
and \U$26699 ( \27014 , \26713 , \26718 );
and \U$26700 ( \27015 , \26709 , \26718 );
or \U$26701 ( \27016 , \27013 , \27014 , \27015 );
and \U$26702 ( \27017 , \22603 , \22021 );
and \U$26703 ( \27018 , \22567 , \22019 );
nor \U$26704 ( \27019 , \27017 , \27018 );
xnor \U$26705 ( \27020 , \27019 , \21595 );
and \U$26706 ( \27021 , \22624 , \21983 );
and \U$26707 ( \27022 , \22592 , \21981 );
nor \U$26708 ( \27023 , \27021 , \27022 );
xnor \U$26709 ( \27024 , \27023 , \21995 );
xor \U$26710 ( \27025 , \27020 , \27024 );
and \U$26711 ( \27026 , \22613 , \21978 );
xor \U$26712 ( \27027 , \27025 , \27026 );
xnor \U$26713 ( \27028 , \27016 , \27027 );
xor \U$26714 ( \27029 , \27012 , \27028 );
and \U$26715 ( \27030 , \26665 , \26669 );
and \U$26716 ( \27031 , \26669 , \26674 );
and \U$26717 ( \27032 , \26665 , \26674 );
or \U$26718 ( \27033 , \27030 , \27031 , \27032 );
and \U$26719 ( \27034 , \26738 , \26742 );
and \U$26720 ( \27035 , \26742 , \26747 );
and \U$26721 ( \27036 , \26738 , \26747 );
or \U$26722 ( \27037 , \27034 , \27035 , \27036 );
xor \U$26723 ( \27038 , \27033 , \27037 );
and \U$26724 ( \27039 , \26723 , \26727 );
and \U$26725 ( \27040 , \26727 , \26732 );
and \U$26726 ( \27041 , \26723 , \26732 );
or \U$26727 ( \27042 , \27039 , \27040 , \27041 );
xor \U$26728 ( \27043 , \27038 , \27042 );
xor \U$26729 ( \27044 , \27029 , \27043 );
xor \U$26730 ( \27045 , \26968 , \27044 );
and \U$26731 ( \27046 , \26788 , \26802 );
and \U$26732 ( \27047 , \26802 , \26817 );
and \U$26733 ( \27048 , \26788 , \26817 );
or \U$26734 ( \27049 , \27046 , \27047 , \27048 );
and \U$26735 ( \27050 , \22124 , \22278 );
and \U$26736 ( \27051 , \22089 , \22276 );
nor \U$26737 ( \27052 , \27050 , \27051 );
xnor \U$26738 ( \27053 , \27052 , \22288 );
and \U$26739 ( \27054 , \22145 , \22300 );
and \U$26740 ( \27055 , \22113 , \22298 );
nor \U$26741 ( \27056 , \27054 , \27055 );
xnor \U$26742 ( \27057 , \27056 , \22310 );
xor \U$26743 ( \27058 , \27053 , \27057 );
and \U$26744 ( \27059 , \22167 , \22324 );
and \U$26745 ( \27060 , \22134 , \22322 );
nor \U$26746 ( \27061 , \27059 , \27060 );
xnor \U$26747 ( \27062 , \27061 , \22334 );
xor \U$26748 ( \27063 , \27058 , \27062 );
and \U$26749 ( \27064 , \22894 , \22208 );
and \U$26750 ( \27065 , \23230 , \22206 );
nor \U$26751 ( \27066 , \27064 , \27065 );
xnor \U$26752 ( \27067 , \27066 , \22218 );
and \U$26753 ( \27068 , \22081 , \22230 );
and \U$26754 ( \27069 , \22858 , \22228 );
nor \U$26755 ( \27070 , \27068 , \27069 );
xnor \U$26756 ( \27071 , \27070 , \22240 );
xor \U$26757 ( \27072 , \27067 , \27071 );
and \U$26758 ( \27073 , \22100 , \22257 );
and \U$26759 ( \27074 , \22071 , \22255 );
nor \U$26760 ( \27075 , \27073 , \27074 );
xnor \U$26761 ( \27076 , \27075 , \22267 );
xor \U$26762 ( \27077 , \27072 , \27076 );
xor \U$26763 ( \27078 , \27063 , \27077 );
and \U$26764 ( \27079 , \21990 , \22140 );
not \U$26765 ( \27080 , \27079 );
xnor \U$26766 ( \27081 , \27080 , \22150 );
and \U$26767 ( \27082 , \22001 , \22162 );
and \U$26768 ( \27083 , \21977 , \22160 );
nor \U$26769 ( \27084 , \27082 , \27083 );
xnor \U$26770 ( \27085 , \27084 , \22172 );
xor \U$26771 ( \27086 , \27081 , \27085 );
and \U$26772 ( \27087 , \23329 , \22187 );
and \U$26773 ( \27088 , \22030 , \22185 );
nor \U$26774 ( \27089 , \27087 , \27088 );
xnor \U$26775 ( \27090 , \27089 , \22197 );
xor \U$26776 ( \27091 , \27086 , \27090 );
xor \U$26777 ( \27092 , \27078 , \27091 );
xor \U$26778 ( \27093 , \27049 , \27092 );
and \U$26779 ( \27094 , \22329 , \22484 );
and \U$26780 ( \27095 , \22294 , \22482 );
nor \U$26781 ( \27096 , \27094 , \27095 );
xnor \U$26782 ( \27097 , \27096 , \22494 );
and \U$26783 ( \27098 , \22350 , \22506 );
and \U$26784 ( \27099 , \22318 , \22504 );
nor \U$26785 ( \27100 , \27098 , \27099 );
xnor \U$26786 ( \27101 , \27100 , \22516 );
xor \U$26787 ( \27102 , \27097 , \27101 );
and \U$26788 ( \27103 , \22372 , \22530 );
and \U$26789 ( \27104 , \22339 , \22528 );
nor \U$26790 ( \27105 , \27103 , \27104 );
xnor \U$26791 ( \27106 , \27105 , \22540 );
xor \U$26792 ( \27107 , \27102 , \27106 );
and \U$26793 ( \27108 , \22262 , \22413 );
and \U$26794 ( \27109 , \22224 , \22411 );
nor \U$26795 ( \27110 , \27108 , \27109 );
xnor \U$26796 ( \27111 , \27110 , \22423 );
and \U$26797 ( \27112 , \22283 , \22435 );
and \U$26798 ( \27113 , \22251 , \22433 );
nor \U$26799 ( \27114 , \27112 , \27113 );
xnor \U$26800 ( \27115 , \27114 , \22445 );
xor \U$26801 ( \27116 , \27111 , \27115 );
and \U$26802 ( \27117 , \22305 , \22463 );
and \U$26803 ( \27118 , \22272 , \22461 );
nor \U$26804 ( \27119 , \27117 , \27118 );
xnor \U$26805 ( \27120 , \27119 , \22473 );
xor \U$26806 ( \27121 , \27116 , \27120 );
xor \U$26807 ( \27122 , \27107 , \27121 );
and \U$26808 ( \27123 , \22192 , \22345 );
and \U$26809 ( \27124 , \22156 , \22343 );
nor \U$26810 ( \27125 , \27123 , \27124 );
xnor \U$26811 ( \27126 , \27125 , \22355 );
and \U$26812 ( \27127 , \22213 , \22367 );
and \U$26813 ( \27128 , \22181 , \22365 );
nor \U$26814 ( \27129 , \27127 , \27128 );
xnor \U$26815 ( \27130 , \27129 , \22377 );
xor \U$26816 ( \27131 , \27126 , \27130 );
and \U$26817 ( \27132 , \22235 , \22392 );
and \U$26818 ( \27133 , \22202 , \22390 );
nor \U$26819 ( \27134 , \27132 , \27133 );
xnor \U$26820 ( \27135 , \27134 , \22402 );
xor \U$26821 ( \27136 , \27131 , \27135 );
xor \U$26822 ( \27137 , \27122 , \27136 );
xor \U$26823 ( \27138 , \27093 , \27137 );
xor \U$26824 ( \27139 , \27045 , \27138 );
xor \U$26825 ( \27140 , \26954 , \27139 );
xor \U$26826 ( \27141 , \26925 , \27140 );
and \U$26827 ( \27142 , \26628 , \26632 );
and \U$26828 ( \27143 , \26632 , \26637 );
and \U$26829 ( \27144 , \26628 , \26637 );
or \U$26830 ( \27145 , \27142 , \27143 , \27144 );
and \U$26831 ( \27146 , \26840 , \26844 );
and \U$26832 ( \27147 , \26844 , \26889 );
and \U$26833 ( \27148 , \26840 , \26889 );
or \U$26834 ( \27149 , \27146 , \27147 , \27148 );
xor \U$26835 ( \27150 , \27145 , \27149 );
and \U$26836 ( \27151 , \26758 , \26819 );
and \U$26837 ( \27152 , \26819 , \26834 );
and \U$26838 ( \27153 , \26758 , \26834 );
or \U$26839 ( \27154 , \27151 , \27152 , \27153 );
xor \U$26840 ( \27155 , \27150 , \27154 );
xor \U$26841 ( \27156 , \27141 , \27155 );
xor \U$26842 ( \27157 , \26911 , \27156 );
and \U$26843 ( \27158 , \26605 , \26609 );
and \U$26844 ( \27159 , \26609 , \26614 );
and \U$26845 ( \27160 , \26605 , \26614 );
or \U$26846 ( \27161 , \27158 , \27159 , \27160 );
and \U$26847 ( \27162 , \26661 , \26835 );
and \U$26848 ( \27163 , \26835 , \26890 );
and \U$26849 ( \27164 , \26661 , \26890 );
or \U$26850 ( \27165 , \27162 , \27163 , \27164 );
xor \U$26851 ( \27166 , \27161 , \27165 );
and \U$26852 ( \27167 , \26705 , \26749 );
and \U$26853 ( \27168 , \26749 , \26757 );
and \U$26854 ( \27169 , \26705 , \26757 );
or \U$26855 ( \27170 , \27167 , \27168 , \27169 );
and \U$26856 ( \27171 , \26859 , \26873 );
and \U$26857 ( \27172 , \26873 , \26888 );
and \U$26858 ( \27173 , \26859 , \26888 );
or \U$26859 ( \27174 , \27171 , \27172 , \27173 );
xor \U$26860 ( \27175 , \27170 , \27174 );
and \U$26861 ( \27176 , \26778 , \26782 );
and \U$26862 ( \27177 , \26782 , \26787 );
and \U$26863 ( \27178 , \26778 , \26787 );
or \U$26864 ( \27179 , \27176 , \27177 , \27178 );
and \U$26865 ( \27180 , \26694 , \26698 );
and \U$26866 ( \27181 , \26698 , \26703 );
and \U$26867 ( \27182 , \26694 , \26703 );
or \U$26868 ( \27183 , \27180 , \27181 , \27182 );
xor \U$26869 ( \27184 , \27179 , \27183 );
and \U$26870 ( \27185 , \26679 , \26683 );
and \U$26871 ( \27186 , \26683 , \26688 );
and \U$26872 ( \27187 , \26679 , \26688 );
or \U$26873 ( \27188 , \27185 , \27186 , \27187 );
xor \U$26874 ( \27189 , \27184 , \27188 );
xor \U$26875 ( \27190 , \27175 , \27189 );
xor \U$26876 ( \27191 , \27166 , \27190 );
xor \U$26877 ( \27192 , \27157 , \27191 );
xor \U$26878 ( \27193 , \26907 , \27192 );
and \U$26879 ( \27194 , \26601 , \26640 );
and \U$26880 ( \27195 , \26640 , \26892 );
and \U$26881 ( \27196 , \26601 , \26892 );
or \U$26882 ( \27197 , \27194 , \27195 , \27196 );
nor \U$26883 ( \27198 , \27193 , \27197 );
and \U$26884 ( \27199 , \26911 , \27156 );
and \U$26885 ( \27200 , \27156 , \27191 );
and \U$26886 ( \27201 , \26911 , \27191 );
or \U$26887 ( \27202 , \27199 , \27200 , \27201 );
and \U$26888 ( \27203 , \27145 , \27149 );
and \U$26889 ( \27204 , \27149 , \27154 );
and \U$26890 ( \27205 , \27145 , \27154 );
or \U$26891 ( \27206 , \27203 , \27204 , \27205 );
and \U$26892 ( \27207 , \26939 , \26953 );
and \U$26893 ( \27208 , \26953 , \27139 );
and \U$26894 ( \27209 , \26939 , \27139 );
or \U$26895 ( \27210 , \27207 , \27208 , \27209 );
xor \U$26896 ( \27211 , \27206 , \27210 );
and \U$26897 ( \27212 , \27063 , \27077 );
and \U$26898 ( \27213 , \27077 , \27091 );
and \U$26899 ( \27214 , \27063 , \27091 );
or \U$26900 ( \27215 , \27212 , \27213 , \27214 );
and \U$26901 ( \27216 , \23230 , \22208 );
and \U$26902 ( \27217 , \23329 , \22206 );
nor \U$26903 ( \27218 , \27216 , \27217 );
xnor \U$26904 ( \27219 , \27218 , \22218 );
and \U$26905 ( \27220 , \22858 , \22230 );
and \U$26906 ( \27221 , \22894 , \22228 );
nor \U$26907 ( \27222 , \27220 , \27221 );
xnor \U$26908 ( \27223 , \27222 , \22240 );
xor \U$26909 ( \27224 , \27219 , \27223 );
and \U$26910 ( \27225 , \22071 , \22257 );
and \U$26911 ( \27226 , \22081 , \22255 );
nor \U$26912 ( \27227 , \27225 , \27226 );
xnor \U$26913 ( \27228 , \27227 , \22267 );
xor \U$26914 ( \27229 , \27224 , \27228 );
xor \U$26915 ( \27230 , \27215 , \27229 );
not \U$26916 ( \27231 , \22150 );
and \U$26917 ( \27232 , \21977 , \22162 );
and \U$26918 ( \27233 , \21990 , \22160 );
nor \U$26919 ( \27234 , \27232 , \27233 );
xnor \U$26920 ( \27235 , \27234 , \22172 );
xor \U$26921 ( \27236 , \27231 , \27235 );
and \U$26922 ( \27237 , \22030 , \22187 );
and \U$26923 ( \27238 , \22001 , \22185 );
nor \U$26924 ( \27239 , \27237 , \27238 );
xnor \U$26925 ( \27240 , \27239 , \22197 );
xor \U$26926 ( \27241 , \27236 , \27240 );
xor \U$26927 ( \27242 , \27230 , \27241 );
or \U$26928 ( \27243 , \27016 , \27027 );
and \U$26929 ( \27244 , \26982 , \26996 );
and \U$26930 ( \27245 , \26996 , \27011 );
and \U$26931 ( \27246 , \26982 , \27011 );
or \U$26932 ( \27247 , \27244 , \27245 , \27246 );
xor \U$26933 ( \27248 , \27243 , \27247 );
and \U$26934 ( \27249 , \27107 , \27121 );
and \U$26935 ( \27250 , \27121 , \27136 );
and \U$26936 ( \27251 , \27107 , \27136 );
or \U$26937 ( \27252 , \27249 , \27250 , \27251 );
xor \U$26938 ( \27253 , \27248 , \27252 );
xor \U$26939 ( \27254 , \27242 , \27253 );
and \U$26940 ( \27255 , \26958 , \26962 );
and \U$26941 ( \27256 , \26962 , \26967 );
and \U$26942 ( \27257 , \26958 , \26967 );
or \U$26943 ( \27258 , \27255 , \27256 , \27257 );
and \U$26944 ( \27259 , \27179 , \27183 );
and \U$26945 ( \27260 , \27183 , \27188 );
and \U$26946 ( \27261 , \27179 , \27188 );
or \U$26947 ( \27262 , \27259 , \27260 , \27261 );
xor \U$26948 ( \27263 , \27258 , \27262 );
and \U$26949 ( \27264 , \27033 , \27037 );
and \U$26950 ( \27265 , \27037 , \27042 );
and \U$26951 ( \27266 , \27033 , \27042 );
or \U$26952 ( \27267 , \27264 , \27265 , \27266 );
xor \U$26953 ( \27268 , \27263 , \27267 );
xor \U$26954 ( \27269 , \27254 , \27268 );
and \U$26955 ( \27270 , \27012 , \27028 );
and \U$26956 ( \27271 , \27028 , \27043 );
and \U$26957 ( \27272 , \27012 , \27043 );
or \U$26958 ( \27273 , \27270 , \27271 , \27272 );
and \U$26959 ( \27274 , \27001 , \27005 );
and \U$26960 ( \27275 , \27005 , \27010 );
and \U$26961 ( \27276 , \27001 , \27010 );
or \U$26962 ( \27277 , \27274 , \27275 , \27276 );
and \U$26963 ( \27278 , \26986 , \26990 );
and \U$26964 ( \27279 , \26990 , \26995 );
and \U$26965 ( \27280 , \26986 , \26995 );
or \U$26966 ( \27281 , \27278 , \27279 , \27280 );
xor \U$26967 ( \27282 , \27277 , \27281 );
and \U$26968 ( \27283 , \26972 , \26976 );
and \U$26969 ( \27284 , \26976 , \26981 );
and \U$26970 ( \27285 , \26972 , \26981 );
or \U$26971 ( \27286 , \27283 , \27284 , \27285 );
xor \U$26972 ( \27287 , \27282 , \27286 );
and \U$26973 ( \27288 , \27126 , \27130 );
and \U$26974 ( \27289 , \27130 , \27135 );
and \U$26975 ( \27290 , \27126 , \27135 );
or \U$26976 ( \27291 , \27288 , \27289 , \27290 );
and \U$26977 ( \27292 , \27111 , \27115 );
and \U$26978 ( \27293 , \27115 , \27120 );
and \U$26979 ( \27294 , \27111 , \27120 );
or \U$26980 ( \27295 , \27292 , \27293 , \27294 );
xor \U$26981 ( \27296 , \27291 , \27295 );
and \U$26982 ( \27297 , \27097 , \27101 );
and \U$26983 ( \27298 , \27101 , \27106 );
and \U$26984 ( \27299 , \27097 , \27106 );
or \U$26985 ( \27300 , \27297 , \27298 , \27299 );
xor \U$26986 ( \27301 , \27296 , \27300 );
xor \U$26987 ( \27302 , \27287 , \27301 );
and \U$26988 ( \27303 , \27081 , \27085 );
and \U$26989 ( \27304 , \27085 , \27090 );
and \U$26990 ( \27305 , \27081 , \27090 );
or \U$26991 ( \27306 , \27303 , \27304 , \27305 );
and \U$26992 ( \27307 , \27067 , \27071 );
and \U$26993 ( \27308 , \27071 , \27076 );
and \U$26994 ( \27309 , \27067 , \27076 );
or \U$26995 ( \27310 , \27307 , \27308 , \27309 );
xor \U$26996 ( \27311 , \27306 , \27310 );
and \U$26997 ( \27312 , \27053 , \27057 );
and \U$26998 ( \27313 , \27057 , \27062 );
and \U$26999 ( \27314 , \27053 , \27062 );
or \U$27000 ( \27315 , \27312 , \27313 , \27314 );
xor \U$27001 ( \27316 , \27311 , \27315 );
xor \U$27002 ( \27317 , \27302 , \27316 );
xor \U$27003 ( \27318 , \27273 , \27317 );
and \U$27004 ( \27319 , \22224 , \22413 );
and \U$27005 ( \27320 , \22235 , \22411 );
nor \U$27006 ( \27321 , \27319 , \27320 );
xnor \U$27007 ( \27322 , \27321 , \22423 );
and \U$27008 ( \27323 , \22251 , \22435 );
and \U$27009 ( \27324 , \22262 , \22433 );
nor \U$27010 ( \27325 , \27323 , \27324 );
xnor \U$27011 ( \27326 , \27325 , \22445 );
xor \U$27012 ( \27327 , \27322 , \27326 );
and \U$27013 ( \27328 , \22272 , \22463 );
and \U$27014 ( \27329 , \22283 , \22461 );
nor \U$27015 ( \27330 , \27328 , \27329 );
xnor \U$27016 ( \27331 , \27330 , \22473 );
xor \U$27017 ( \27332 , \27327 , \27331 );
and \U$27018 ( \27333 , \22156 , \22345 );
and \U$27019 ( \27334 , \22167 , \22343 );
nor \U$27020 ( \27335 , \27333 , \27334 );
xnor \U$27021 ( \27336 , \27335 , \22355 );
and \U$27022 ( \27337 , \22181 , \22367 );
and \U$27023 ( \27338 , \22192 , \22365 );
nor \U$27024 ( \27339 , \27337 , \27338 );
xnor \U$27025 ( \27340 , \27339 , \22377 );
xor \U$27026 ( \27341 , \27336 , \27340 );
and \U$27027 ( \27342 , \22202 , \22392 );
and \U$27028 ( \27343 , \22213 , \22390 );
nor \U$27029 ( \27344 , \27342 , \27343 );
xnor \U$27030 ( \27345 , \27344 , \22402 );
xor \U$27031 ( \27346 , \27341 , \27345 );
xor \U$27032 ( \27347 , \27332 , \27346 );
and \U$27033 ( \27348 , \22089 , \22278 );
and \U$27034 ( \27349 , \22100 , \22276 );
nor \U$27035 ( \27350 , \27348 , \27349 );
xnor \U$27036 ( \27351 , \27350 , \22288 );
and \U$27037 ( \27352 , \22113 , \22300 );
and \U$27038 ( \27353 , \22124 , \22298 );
nor \U$27039 ( \27354 , \27352 , \27353 );
xnor \U$27040 ( \27355 , \27354 , \22310 );
xor \U$27041 ( \27356 , \27351 , \27355 );
and \U$27042 ( \27357 , \22134 , \22324 );
and \U$27043 ( \27358 , \22145 , \22322 );
nor \U$27044 ( \27359 , \27357 , \27358 );
xnor \U$27045 ( \27360 , \27359 , \22334 );
xor \U$27046 ( \27361 , \27356 , \27360 );
xor \U$27047 ( \27362 , \27347 , \27361 );
and \U$27048 ( \27363 , \22429 , \22619 );
and \U$27049 ( \27364 , \22440 , \22617 );
nor \U$27050 ( \27365 , \27363 , \27364 );
xnor \U$27051 ( \27366 , \27365 , \22629 );
and \U$27052 ( \27367 , \22457 , \22641 );
and \U$27053 ( \27368 , \22468 , \22639 );
nor \U$27054 ( \27369 , \27367 , \27368 );
xnor \U$27055 ( \27370 , \27369 , \22651 );
xor \U$27056 ( \27371 , \27366 , \27370 );
and \U$27057 ( \27372 , \22478 , \22671 );
and \U$27058 ( \27373 , \22489 , \22669 );
nor \U$27059 ( \27374 , \27372 , \27373 );
xnor \U$27060 ( \27375 , \27374 , \22681 );
xor \U$27061 ( \27376 , \27371 , \27375 );
and \U$27062 ( \27377 , \22361 , \22551 );
and \U$27063 ( \27378 , \22372 , \22549 );
nor \U$27064 ( \27379 , \27377 , \27378 );
xnor \U$27065 ( \27380 , \27379 , \22561 );
and \U$27066 ( \27381 , \22386 , \22573 );
and \U$27067 ( \27382 , \22397 , \22571 );
nor \U$27068 ( \27383 , \27381 , \27382 );
xnor \U$27069 ( \27384 , \27383 , \22583 );
xor \U$27070 ( \27385 , \27380 , \27384 );
and \U$27071 ( \27386 , \22407 , \22598 );
and \U$27072 ( \27387 , \22418 , \22596 );
nor \U$27073 ( \27388 , \27386 , \27387 );
xnor \U$27074 ( \27389 , \27388 , \22608 );
xor \U$27075 ( \27390 , \27385 , \27389 );
xor \U$27076 ( \27391 , \27376 , \27390 );
and \U$27077 ( \27392 , \22294 , \22484 );
and \U$27078 ( \27393 , \22305 , \22482 );
nor \U$27079 ( \27394 , \27392 , \27393 );
xnor \U$27080 ( \27395 , \27394 , \22494 );
and \U$27081 ( \27396 , \22318 , \22506 );
and \U$27082 ( \27397 , \22329 , \22504 );
nor \U$27083 ( \27398 , \27396 , \27397 );
xnor \U$27084 ( \27399 , \27398 , \22516 );
xor \U$27085 ( \27400 , \27395 , \27399 );
and \U$27086 ( \27401 , \22339 , \22530 );
and \U$27087 ( \27402 , \22350 , \22528 );
nor \U$27088 ( \27403 , \27401 , \27402 );
xnor \U$27089 ( \27404 , \27403 , \22540 );
xor \U$27090 ( \27405 , \27400 , \27404 );
xor \U$27091 ( \27406 , \27391 , \27405 );
xor \U$27092 ( \27407 , \27362 , \27406 );
and \U$27093 ( \27408 , \27020 , \27024 );
and \U$27094 ( \27409 , \27024 , \27026 );
and \U$27095 ( \27410 , \27020 , \27026 );
or \U$27096 ( \27411 , \27408 , \27409 , \27410 );
and \U$27097 ( \27412 , \22567 , \22021 );
and \U$27098 ( \27413 , \22578 , \22019 );
nor \U$27099 ( \27414 , \27412 , \27413 );
xnor \U$27100 ( \27415 , \27414 , \21595 );
and \U$27101 ( \27416 , \22592 , \21983 );
and \U$27102 ( \27417 , \22603 , \21981 );
nor \U$27103 ( \27418 , \27416 , \27417 );
xnor \U$27104 ( \27419 , \27418 , \21995 );
xor \U$27105 ( \27420 , \27415 , \27419 );
and \U$27106 ( \27421 , \22624 , \21978 );
xor \U$27107 ( \27422 , \27420 , \27421 );
xor \U$27108 ( \27423 , \27411 , \27422 );
and \U$27109 ( \27424 , \22500 , \22691 );
and \U$27110 ( \27425 , \22511 , \22689 );
nor \U$27111 ( \27426 , \27424 , \27425 );
xnor \U$27112 ( \27427 , \27426 , \22701 );
and \U$27113 ( \27428 , \22524 , \22720 );
and \U$27114 ( \27429 , \22535 , \22707 );
nor \U$27115 ( \27430 , \27428 , \27429 );
xnor \U$27116 ( \27431 , \27430 , \22067 );
xor \U$27117 ( \27432 , \27427 , \27431 );
and \U$27118 ( \27433 , \22545 , \23173 );
and \U$27119 ( \27434 , \22556 , \22999 );
nor \U$27120 ( \27435 , \27433 , \27434 );
xnor \U$27121 ( \27436 , \27435 , \22016 );
xor \U$27122 ( \27437 , \27432 , \27436 );
xor \U$27123 ( \27438 , \27423 , \27437 );
xor \U$27124 ( \27439 , \27407 , \27438 );
xor \U$27125 ( \27440 , \27318 , \27439 );
xor \U$27126 ( \27441 , \27269 , \27440 );
and \U$27127 ( \27442 , \26943 , \26947 );
and \U$27128 ( \27443 , \26947 , \26952 );
and \U$27129 ( \27444 , \26943 , \26952 );
or \U$27130 ( \27445 , \27442 , \27443 , \27444 );
and \U$27131 ( \27446 , \26929 , \26933 );
and \U$27132 ( \27447 , \26933 , \26938 );
and \U$27133 ( \27448 , \26929 , \26938 );
or \U$27134 ( \27449 , \27446 , \27447 , \27448 );
xor \U$27135 ( \27450 , \27445 , \27449 );
and \U$27136 ( \27451 , \27049 , \27092 );
and \U$27137 ( \27452 , \27092 , \27137 );
and \U$27138 ( \27453 , \27049 , \27137 );
or \U$27139 ( \27454 , \27451 , \27452 , \27453 );
xor \U$27140 ( \27455 , \27450 , \27454 );
xor \U$27141 ( \27456 , \27441 , \27455 );
xor \U$27142 ( \27457 , \27211 , \27456 );
xor \U$27143 ( \27458 , \27202 , \27457 );
and \U$27144 ( \27459 , \27161 , \27165 );
and \U$27145 ( \27460 , \27165 , \27190 );
and \U$27146 ( \27461 , \27161 , \27190 );
or \U$27147 ( \27462 , \27459 , \27460 , \27461 );
and \U$27148 ( \27463 , \26925 , \27140 );
and \U$27149 ( \27464 , \27140 , \27155 );
and \U$27150 ( \27465 , \26925 , \27155 );
or \U$27151 ( \27466 , \27463 , \27464 , \27465 );
xor \U$27152 ( \27467 , \27462 , \27466 );
and \U$27153 ( \27468 , \26915 , \26919 );
and \U$27154 ( \27469 , \26919 , \26924 );
and \U$27155 ( \27470 , \26915 , \26924 );
or \U$27156 ( \27471 , \27468 , \27469 , \27470 );
and \U$27157 ( \27472 , \27170 , \27174 );
and \U$27158 ( \27473 , \27174 , \27189 );
and \U$27159 ( \27474 , \27170 , \27189 );
or \U$27160 ( \27475 , \27472 , \27473 , \27474 );
xor \U$27161 ( \27476 , \27471 , \27475 );
and \U$27162 ( \27477 , \26968 , \27044 );
and \U$27163 ( \27478 , \27044 , \27138 );
and \U$27164 ( \27479 , \26968 , \27138 );
or \U$27165 ( \27480 , \27477 , \27478 , \27479 );
xor \U$27166 ( \27481 , \27476 , \27480 );
xor \U$27167 ( \27482 , \27467 , \27481 );
xor \U$27168 ( \27483 , \27458 , \27482 );
and \U$27169 ( \27484 , \26905 , \26906 );
and \U$27170 ( \27485 , \26906 , \27192 );
and \U$27171 ( \27486 , \26905 , \27192 );
or \U$27172 ( \27487 , \27484 , \27485 , \27486 );
nor \U$27173 ( \27488 , \27483 , \27487 );
nor \U$27174 ( \27489 , \27198 , \27488 );
and \U$27175 ( \27490 , \27462 , \27466 );
and \U$27176 ( \27491 , \27466 , \27481 );
and \U$27177 ( \27492 , \27462 , \27481 );
or \U$27178 ( \27493 , \27490 , \27491 , \27492 );
and \U$27179 ( \27494 , \27206 , \27210 );
and \U$27180 ( \27495 , \27210 , \27456 );
and \U$27181 ( \27496 , \27206 , \27456 );
or \U$27182 ( \27497 , \27494 , \27495 , \27496 );
and \U$27183 ( \27498 , \27258 , \27262 );
and \U$27184 ( \27499 , \27262 , \27267 );
and \U$27185 ( \27500 , \27258 , \27267 );
or \U$27186 ( \27501 , \27498 , \27499 , \27500 );
and \U$27187 ( \27502 , \27243 , \27247 );
and \U$27188 ( \27503 , \27247 , \27252 );
and \U$27189 ( \27504 , \27243 , \27252 );
or \U$27190 ( \27505 , \27502 , \27503 , \27504 );
xor \U$27191 ( \27506 , \27501 , \27505 );
and \U$27192 ( \27507 , \27215 , \27229 );
and \U$27193 ( \27508 , \27229 , \27241 );
and \U$27194 ( \27509 , \27215 , \27241 );
or \U$27195 ( \27510 , \27507 , \27508 , \27509 );
xor \U$27196 ( \27511 , \27506 , \27510 );
and \U$27197 ( \27512 , \27411 , \27422 );
and \U$27198 ( \27513 , \27422 , \27437 );
and \U$27199 ( \27514 , \27411 , \27437 );
or \U$27200 ( \27515 , \27512 , \27513 , \27514 );
and \U$27201 ( \27516 , \27376 , \27390 );
and \U$27202 ( \27517 , \27390 , \27405 );
and \U$27203 ( \27518 , \27376 , \27405 );
or \U$27204 ( \27519 , \27516 , \27517 , \27518 );
xor \U$27205 ( \27520 , \27515 , \27519 );
and \U$27206 ( \27521 , \27332 , \27346 );
and \U$27207 ( \27522 , \27346 , \27361 );
and \U$27208 ( \27523 , \27332 , \27361 );
or \U$27209 ( \27524 , \27521 , \27522 , \27523 );
xor \U$27210 ( \27525 , \27520 , \27524 );
and \U$27211 ( \27526 , \27306 , \27310 );
and \U$27212 ( \27527 , \27310 , \27315 );
and \U$27213 ( \27528 , \27306 , \27315 );
or \U$27214 ( \27529 , \27526 , \27527 , \27528 );
and \U$27215 ( \27530 , \27291 , \27295 );
and \U$27216 ( \27531 , \27295 , \27300 );
and \U$27217 ( \27532 , \27291 , \27300 );
or \U$27218 ( \27533 , \27530 , \27531 , \27532 );
xor \U$27219 ( \27534 , \27529 , \27533 );
and \U$27220 ( \27535 , \27277 , \27281 );
and \U$27221 ( \27536 , \27281 , \27286 );
and \U$27222 ( \27537 , \27277 , \27286 );
or \U$27223 ( \27538 , \27535 , \27536 , \27537 );
xor \U$27224 ( \27539 , \27534 , \27538 );
xor \U$27225 ( \27540 , \27525 , \27539 );
and \U$27226 ( \27541 , \27231 , \27235 );
and \U$27227 ( \27542 , \27235 , \27240 );
and \U$27228 ( \27543 , \27231 , \27240 );
or \U$27229 ( \27544 , \27541 , \27542 , \27543 );
and \U$27230 ( \27545 , \27219 , \27223 );
and \U$27231 ( \27546 , \27223 , \27228 );
and \U$27232 ( \27547 , \27219 , \27228 );
or \U$27233 ( \27548 , \27545 , \27546 , \27547 );
xor \U$27234 ( \27549 , \27544 , \27548 );
and \U$27235 ( \27550 , \27351 , \27355 );
and \U$27236 ( \27551 , \27355 , \27360 );
and \U$27237 ( \27552 , \27351 , \27360 );
or \U$27238 ( \27553 , \27550 , \27551 , \27552 );
xor \U$27239 ( \27554 , \27549 , \27553 );
and \U$27240 ( \27555 , \22468 , \22641 );
and \U$27241 ( \27556 , \22429 , \22639 );
nor \U$27242 ( \27557 , \27555 , \27556 );
xnor \U$27243 ( \27558 , \27557 , \22651 );
and \U$27244 ( \27559 , \22489 , \22671 );
and \U$27245 ( \27560 , \22457 , \22669 );
nor \U$27246 ( \27561 , \27559 , \27560 );
xnor \U$27247 ( \27562 , \27561 , \22681 );
xor \U$27248 ( \27563 , \27558 , \27562 );
and \U$27249 ( \27564 , \22511 , \22691 );
and \U$27250 ( \27565 , \22478 , \22689 );
nor \U$27251 ( \27566 , \27564 , \27565 );
xnor \U$27252 ( \27567 , \27566 , \22701 );
xor \U$27253 ( \27568 , \27563 , \27567 );
and \U$27254 ( \27569 , \22397 , \22573 );
and \U$27255 ( \27570 , \22361 , \22571 );
nor \U$27256 ( \27571 , \27569 , \27570 );
xnor \U$27257 ( \27572 , \27571 , \22583 );
and \U$27258 ( \27573 , \22418 , \22598 );
and \U$27259 ( \27574 , \22386 , \22596 );
nor \U$27260 ( \27575 , \27573 , \27574 );
xnor \U$27261 ( \27576 , \27575 , \22608 );
xor \U$27262 ( \27577 , \27572 , \27576 );
and \U$27263 ( \27578 , \22440 , \22619 );
and \U$27264 ( \27579 , \22407 , \22617 );
nor \U$27265 ( \27580 , \27578 , \27579 );
xnor \U$27266 ( \27581 , \27580 , \22629 );
xor \U$27267 ( \27582 , \27577 , \27581 );
xor \U$27268 ( \27583 , \27568 , \27582 );
and \U$27269 ( \27584 , \22329 , \22506 );
and \U$27270 ( \27585 , \22294 , \22504 );
nor \U$27271 ( \27586 , \27584 , \27585 );
xnor \U$27272 ( \27587 , \27586 , \22516 );
and \U$27273 ( \27588 , \22350 , \22530 );
and \U$27274 ( \27589 , \22318 , \22528 );
nor \U$27275 ( \27590 , \27588 , \27589 );
xnor \U$27276 ( \27591 , \27590 , \22540 );
xor \U$27277 ( \27592 , \27587 , \27591 );
and \U$27278 ( \27593 , \22372 , \22551 );
and \U$27279 ( \27594 , \22339 , \22549 );
nor \U$27280 ( \27595 , \27593 , \27594 );
xnor \U$27281 ( \27596 , \27595 , \22561 );
xor \U$27282 ( \27597 , \27592 , \27596 );
xor \U$27283 ( \27598 , \27583 , \27597 );
and \U$27284 ( \27599 , \27415 , \27419 );
and \U$27285 ( \27600 , \27419 , \27421 );
and \U$27286 ( \27601 , \27415 , \27421 );
or \U$27287 ( \27602 , \27599 , \27600 , \27601 );
and \U$27288 ( \27603 , \22603 , \21983 );
and \U$27289 ( \27604 , \22567 , \21981 );
nor \U$27290 ( \27605 , \27603 , \27604 );
xnor \U$27291 ( \27606 , \27605 , \21995 );
and \U$27292 ( \27607 , \22592 , \21978 );
xnor \U$27293 ( \27608 , \27606 , \27607 );
xor \U$27294 ( \27609 , \27602 , \27608 );
and \U$27295 ( \27610 , \22535 , \22720 );
and \U$27296 ( \27611 , \22500 , \22707 );
nor \U$27297 ( \27612 , \27610 , \27611 );
xnor \U$27298 ( \27613 , \27612 , \22067 );
and \U$27299 ( \27614 , \22556 , \23173 );
and \U$27300 ( \27615 , \22524 , \22999 );
nor \U$27301 ( \27616 , \27614 , \27615 );
xnor \U$27302 ( \27617 , \27616 , \22016 );
xor \U$27303 ( \27618 , \27613 , \27617 );
and \U$27304 ( \27619 , \22578 , \22021 );
and \U$27305 ( \27620 , \22545 , \22019 );
nor \U$27306 ( \27621 , \27619 , \27620 );
xnor \U$27307 ( \27622 , \27621 , \21595 );
xor \U$27308 ( \27623 , \27618 , \27622 );
xor \U$27309 ( \27624 , \27609 , \27623 );
xor \U$27310 ( \27625 , \27598 , \27624 );
and \U$27311 ( \27626 , \27380 , \27384 );
and \U$27312 ( \27627 , \27384 , \27389 );
and \U$27313 ( \27628 , \27380 , \27389 );
or \U$27314 ( \27629 , \27626 , \27627 , \27628 );
and \U$27315 ( \27630 , \27366 , \27370 );
and \U$27316 ( \27631 , \27370 , \27375 );
and \U$27317 ( \27632 , \27366 , \27375 );
or \U$27318 ( \27633 , \27630 , \27631 , \27632 );
xor \U$27319 ( \27634 , \27629 , \27633 );
and \U$27320 ( \27635 , \27427 , \27431 );
and \U$27321 ( \27636 , \27431 , \27436 );
and \U$27322 ( \27637 , \27427 , \27436 );
or \U$27323 ( \27638 , \27635 , \27636 , \27637 );
xor \U$27324 ( \27639 , \27634 , \27638 );
xor \U$27325 ( \27640 , \27625 , \27639 );
xor \U$27326 ( \27641 , \27554 , \27640 );
and \U$27327 ( \27642 , \22894 , \22230 );
and \U$27328 ( \27643 , \23230 , \22228 );
nor \U$27329 ( \27644 , \27642 , \27643 );
xnor \U$27330 ( \27645 , \27644 , \22240 );
and \U$27331 ( \27646 , \22081 , \22257 );
and \U$27332 ( \27647 , \22858 , \22255 );
nor \U$27333 ( \27648 , \27646 , \27647 );
xnor \U$27334 ( \27649 , \27648 , \22267 );
xor \U$27335 ( \27650 , \27645 , \27649 );
and \U$27336 ( \27651 , \22100 , \22278 );
and \U$27337 ( \27652 , \22071 , \22276 );
nor \U$27338 ( \27653 , \27651 , \27652 );
xnor \U$27339 ( \27654 , \27653 , \22288 );
xor \U$27340 ( \27655 , \27650 , \27654 );
and \U$27341 ( \27656 , \21990 , \22162 );
not \U$27342 ( \27657 , \27656 );
xnor \U$27343 ( \27658 , \27657 , \22172 );
and \U$27344 ( \27659 , \22001 , \22187 );
and \U$27345 ( \27660 , \21977 , \22185 );
nor \U$27346 ( \27661 , \27659 , \27660 );
xnor \U$27347 ( \27662 , \27661 , \22197 );
xor \U$27348 ( \27663 , \27658 , \27662 );
and \U$27349 ( \27664 , \23329 , \22208 );
and \U$27350 ( \27665 , \22030 , \22206 );
nor \U$27351 ( \27666 , \27664 , \27665 );
xnor \U$27352 ( \27667 , \27666 , \22218 );
xor \U$27353 ( \27668 , \27663 , \27667 );
xor \U$27354 ( \27669 , \27655 , \27668 );
and \U$27355 ( \27670 , \22262 , \22435 );
and \U$27356 ( \27671 , \22224 , \22433 );
nor \U$27357 ( \27672 , \27670 , \27671 );
xnor \U$27358 ( \27673 , \27672 , \22445 );
and \U$27359 ( \27674 , \22283 , \22463 );
and \U$27360 ( \27675 , \22251 , \22461 );
nor \U$27361 ( \27676 , \27674 , \27675 );
xnor \U$27362 ( \27677 , \27676 , \22473 );
xor \U$27363 ( \27678 , \27673 , \27677 );
and \U$27364 ( \27679 , \22305 , \22484 );
and \U$27365 ( \27680 , \22272 , \22482 );
nor \U$27366 ( \27681 , \27679 , \27680 );
xnor \U$27367 ( \27682 , \27681 , \22494 );
xor \U$27368 ( \27683 , \27678 , \27682 );
and \U$27369 ( \27684 , \22192 , \22367 );
and \U$27370 ( \27685 , \22156 , \22365 );
nor \U$27371 ( \27686 , \27684 , \27685 );
xnor \U$27372 ( \27687 , \27686 , \22377 );
and \U$27373 ( \27688 , \22213 , \22392 );
and \U$27374 ( \27689 , \22181 , \22390 );
nor \U$27375 ( \27690 , \27688 , \27689 );
xnor \U$27376 ( \27691 , \27690 , \22402 );
xor \U$27377 ( \27692 , \27687 , \27691 );
and \U$27378 ( \27693 , \22235 , \22413 );
and \U$27379 ( \27694 , \22202 , \22411 );
nor \U$27380 ( \27695 , \27693 , \27694 );
xnor \U$27381 ( \27696 , \27695 , \22423 );
xor \U$27382 ( \27697 , \27692 , \27696 );
xor \U$27383 ( \27698 , \27683 , \27697 );
and \U$27384 ( \27699 , \22124 , \22300 );
and \U$27385 ( \27700 , \22089 , \22298 );
nor \U$27386 ( \27701 , \27699 , \27700 );
xnor \U$27387 ( \27702 , \27701 , \22310 );
and \U$27388 ( \27703 , \22145 , \22324 );
and \U$27389 ( \27704 , \22113 , \22322 );
nor \U$27390 ( \27705 , \27703 , \27704 );
xnor \U$27391 ( \27706 , \27705 , \22334 );
xor \U$27392 ( \27707 , \27702 , \27706 );
and \U$27393 ( \27708 , \22167 , \22345 );
and \U$27394 ( \27709 , \22134 , \22343 );
nor \U$27395 ( \27710 , \27708 , \27709 );
xnor \U$27396 ( \27711 , \27710 , \22355 );
xor \U$27397 ( \27712 , \27707 , \27711 );
xor \U$27398 ( \27713 , \27698 , \27712 );
xor \U$27399 ( \27714 , \27669 , \27713 );
xor \U$27400 ( \27715 , \27641 , \27714 );
xor \U$27401 ( \27716 , \27540 , \27715 );
xor \U$27402 ( \27717 , \27511 , \27716 );
and \U$27403 ( \27718 , \27445 , \27449 );
and \U$27404 ( \27719 , \27449 , \27454 );
and \U$27405 ( \27720 , \27445 , \27454 );
or \U$27406 ( \27721 , \27718 , \27719 , \27720 );
and \U$27407 ( \27722 , \27273 , \27317 );
and \U$27408 ( \27723 , \27317 , \27439 );
and \U$27409 ( \27724 , \27273 , \27439 );
or \U$27410 ( \27725 , \27722 , \27723 , \27724 );
xor \U$27411 ( \27726 , \27721 , \27725 );
and \U$27412 ( \27727 , \27242 , \27253 );
and \U$27413 ( \27728 , \27253 , \27268 );
and \U$27414 ( \27729 , \27242 , \27268 );
or \U$27415 ( \27730 , \27727 , \27728 , \27729 );
xor \U$27416 ( \27731 , \27726 , \27730 );
xor \U$27417 ( \27732 , \27717 , \27731 );
xor \U$27418 ( \27733 , \27497 , \27732 );
and \U$27419 ( \27734 , \27471 , \27475 );
and \U$27420 ( \27735 , \27475 , \27480 );
and \U$27421 ( \27736 , \27471 , \27480 );
or \U$27422 ( \27737 , \27734 , \27735 , \27736 );
and \U$27423 ( \27738 , \27269 , \27440 );
and \U$27424 ( \27739 , \27440 , \27455 );
and \U$27425 ( \27740 , \27269 , \27455 );
or \U$27426 ( \27741 , \27738 , \27739 , \27740 );
xor \U$27427 ( \27742 , \27737 , \27741 );
and \U$27428 ( \27743 , \27362 , \27406 );
and \U$27429 ( \27744 , \27406 , \27438 );
and \U$27430 ( \27745 , \27362 , \27438 );
or \U$27431 ( \27746 , \27743 , \27744 , \27745 );
and \U$27432 ( \27747 , \27287 , \27301 );
and \U$27433 ( \27748 , \27301 , \27316 );
and \U$27434 ( \27749 , \27287 , \27316 );
or \U$27435 ( \27750 , \27747 , \27748 , \27749 );
xor \U$27436 ( \27751 , \27746 , \27750 );
and \U$27437 ( \27752 , \27336 , \27340 );
and \U$27438 ( \27753 , \27340 , \27345 );
and \U$27439 ( \27754 , \27336 , \27345 );
or \U$27440 ( \27755 , \27752 , \27753 , \27754 );
and \U$27441 ( \27756 , \27322 , \27326 );
and \U$27442 ( \27757 , \27326 , \27331 );
and \U$27443 ( \27758 , \27322 , \27331 );
or \U$27444 ( \27759 , \27756 , \27757 , \27758 );
xor \U$27445 ( \27760 , \27755 , \27759 );
and \U$27446 ( \27761 , \27395 , \27399 );
and \U$27447 ( \27762 , \27399 , \27404 );
and \U$27448 ( \27763 , \27395 , \27404 );
or \U$27449 ( \27764 , \27761 , \27762 , \27763 );
xor \U$27450 ( \27765 , \27760 , \27764 );
xor \U$27451 ( \27766 , \27751 , \27765 );
xor \U$27452 ( \27767 , \27742 , \27766 );
xor \U$27453 ( \27768 , \27733 , \27767 );
xor \U$27454 ( \27769 , \27493 , \27768 );
and \U$27455 ( \27770 , \27202 , \27457 );
and \U$27456 ( \27771 , \27457 , \27482 );
and \U$27457 ( \27772 , \27202 , \27482 );
or \U$27458 ( \27773 , \27770 , \27771 , \27772 );
nor \U$27459 ( \27774 , \27769 , \27773 );
and \U$27460 ( \27775 , \27497 , \27732 );
and \U$27461 ( \27776 , \27732 , \27767 );
and \U$27462 ( \27777 , \27497 , \27767 );
or \U$27463 ( \27778 , \27775 , \27776 , \27777 );
and \U$27464 ( \27779 , \27721 , \27725 );
and \U$27465 ( \27780 , \27725 , \27730 );
and \U$27466 ( \27781 , \27721 , \27730 );
or \U$27467 ( \27782 , \27779 , \27780 , \27781 );
and \U$27468 ( \27783 , \27525 , \27539 );
and \U$27469 ( \27784 , \27539 , \27715 );
and \U$27470 ( \27785 , \27525 , \27715 );
or \U$27471 ( \27786 , \27783 , \27784 , \27785 );
xor \U$27472 ( \27787 , \27782 , \27786 );
and \U$27473 ( \27788 , \22089 , \22300 );
and \U$27474 ( \27789 , \22100 , \22298 );
nor \U$27475 ( \27790 , \27788 , \27789 );
xnor \U$27476 ( \27791 , \27790 , \22310 );
and \U$27477 ( \27792 , \22113 , \22324 );
and \U$27478 ( \27793 , \22124 , \22322 );
nor \U$27479 ( \27794 , \27792 , \27793 );
xnor \U$27480 ( \27795 , \27794 , \22334 );
xor \U$27481 ( \27796 , \27791 , \27795 );
and \U$27482 ( \27797 , \22134 , \22345 );
and \U$27483 ( \27798 , \22145 , \22343 );
nor \U$27484 ( \27799 , \27797 , \27798 );
xnor \U$27485 ( \27800 , \27799 , \22355 );
xor \U$27486 ( \27801 , \27796 , \27800 );
and \U$27487 ( \27802 , \23230 , \22230 );
and \U$27488 ( \27803 , \23329 , \22228 );
nor \U$27489 ( \27804 , \27802 , \27803 );
xnor \U$27490 ( \27805 , \27804 , \22240 );
and \U$27491 ( \27806 , \22858 , \22257 );
and \U$27492 ( \27807 , \22894 , \22255 );
nor \U$27493 ( \27808 , \27806 , \27807 );
xnor \U$27494 ( \27809 , \27808 , \22267 );
xor \U$27495 ( \27810 , \27805 , \27809 );
and \U$27496 ( \27811 , \22071 , \22278 );
and \U$27497 ( \27812 , \22081 , \22276 );
nor \U$27498 ( \27813 , \27811 , \27812 );
xnor \U$27499 ( \27814 , \27813 , \22288 );
xor \U$27500 ( \27815 , \27810 , \27814 );
xor \U$27501 ( \27816 , \27801 , \27815 );
not \U$27502 ( \27817 , \22172 );
and \U$27503 ( \27818 , \21977 , \22187 );
and \U$27504 ( \27819 , \21990 , \22185 );
nor \U$27505 ( \27820 , \27818 , \27819 );
xnor \U$27506 ( \27821 , \27820 , \22197 );
xor \U$27507 ( \27822 , \27817 , \27821 );
and \U$27508 ( \27823 , \22030 , \22208 );
and \U$27509 ( \27824 , \22001 , \22206 );
nor \U$27510 ( \27825 , \27823 , \27824 );
xnor \U$27511 ( \27826 , \27825 , \22218 );
xor \U$27512 ( \27827 , \27822 , \27826 );
xor \U$27513 ( \27828 , \27816 , \27827 );
and \U$27514 ( \27829 , \22294 , \22506 );
and \U$27515 ( \27830 , \22305 , \22504 );
nor \U$27516 ( \27831 , \27829 , \27830 );
xnor \U$27517 ( \27832 , \27831 , \22516 );
and \U$27518 ( \27833 , \22318 , \22530 );
and \U$27519 ( \27834 , \22329 , \22528 );
nor \U$27520 ( \27835 , \27833 , \27834 );
xnor \U$27521 ( \27836 , \27835 , \22540 );
xor \U$27522 ( \27837 , \27832 , \27836 );
and \U$27523 ( \27838 , \22339 , \22551 );
and \U$27524 ( \27839 , \22350 , \22549 );
nor \U$27525 ( \27840 , \27838 , \27839 );
xnor \U$27526 ( \27841 , \27840 , \22561 );
xor \U$27527 ( \27842 , \27837 , \27841 );
and \U$27528 ( \27843 , \22224 , \22435 );
and \U$27529 ( \27844 , \22235 , \22433 );
nor \U$27530 ( \27845 , \27843 , \27844 );
xnor \U$27531 ( \27846 , \27845 , \22445 );
and \U$27532 ( \27847 , \22251 , \22463 );
and \U$27533 ( \27848 , \22262 , \22461 );
nor \U$27534 ( \27849 , \27847 , \27848 );
xnor \U$27535 ( \27850 , \27849 , \22473 );
xor \U$27536 ( \27851 , \27846 , \27850 );
and \U$27537 ( \27852 , \22272 , \22484 );
and \U$27538 ( \27853 , \22283 , \22482 );
nor \U$27539 ( \27854 , \27852 , \27853 );
xnor \U$27540 ( \27855 , \27854 , \22494 );
xor \U$27541 ( \27856 , \27851 , \27855 );
xor \U$27542 ( \27857 , \27842 , \27856 );
and \U$27543 ( \27858 , \22156 , \22367 );
and \U$27544 ( \27859 , \22167 , \22365 );
nor \U$27545 ( \27860 , \27858 , \27859 );
xnor \U$27546 ( \27861 , \27860 , \22377 );
and \U$27547 ( \27862 , \22181 , \22392 );
and \U$27548 ( \27863 , \22192 , \22390 );
nor \U$27549 ( \27864 , \27862 , \27863 );
xnor \U$27550 ( \27865 , \27864 , \22402 );
xor \U$27551 ( \27866 , \27861 , \27865 );
and \U$27552 ( \27867 , \22202 , \22413 );
and \U$27553 ( \27868 , \22213 , \22411 );
nor \U$27554 ( \27869 , \27867 , \27868 );
xnor \U$27555 ( \27870 , \27869 , \22423 );
xor \U$27556 ( \27871 , \27866 , \27870 );
xor \U$27557 ( \27872 , \27857 , \27871 );
xor \U$27558 ( \27873 , \27828 , \27872 );
and \U$27559 ( \27874 , \22500 , \22720 );
and \U$27560 ( \27875 , \22511 , \22707 );
nor \U$27561 ( \27876 , \27874 , \27875 );
xnor \U$27562 ( \27877 , \27876 , \22067 );
and \U$27563 ( \27878 , \22524 , \23173 );
and \U$27564 ( \27879 , \22535 , \22999 );
nor \U$27565 ( \27880 , \27878 , \27879 );
xnor \U$27566 ( \27881 , \27880 , \22016 );
xor \U$27567 ( \27882 , \27877 , \27881 );
and \U$27568 ( \27883 , \22545 , \22021 );
and \U$27569 ( \27884 , \22556 , \22019 );
nor \U$27570 ( \27885 , \27883 , \27884 );
xnor \U$27571 ( \27886 , \27885 , \21595 );
xor \U$27572 ( \27887 , \27882 , \27886 );
and \U$27573 ( \27888 , \22429 , \22641 );
and \U$27574 ( \27889 , \22440 , \22639 );
nor \U$27575 ( \27890 , \27888 , \27889 );
xnor \U$27576 ( \27891 , \27890 , \22651 );
and \U$27577 ( \27892 , \22457 , \22671 );
and \U$27578 ( \27893 , \22468 , \22669 );
nor \U$27579 ( \27894 , \27892 , \27893 );
xnor \U$27580 ( \27895 , \27894 , \22681 );
xor \U$27581 ( \27896 , \27891 , \27895 );
and \U$27582 ( \27897 , \22478 , \22691 );
and \U$27583 ( \27898 , \22489 , \22689 );
nor \U$27584 ( \27899 , \27897 , \27898 );
xnor \U$27585 ( \27900 , \27899 , \22701 );
xor \U$27586 ( \27901 , \27896 , \27900 );
xor \U$27587 ( \27902 , \27887 , \27901 );
and \U$27588 ( \27903 , \22361 , \22573 );
and \U$27589 ( \27904 , \22372 , \22571 );
nor \U$27590 ( \27905 , \27903 , \27904 );
xnor \U$27591 ( \27906 , \27905 , \22583 );
and \U$27592 ( \27907 , \22386 , \22598 );
and \U$27593 ( \27908 , \22397 , \22596 );
nor \U$27594 ( \27909 , \27907 , \27908 );
xnor \U$27595 ( \27910 , \27909 , \22608 );
xor \U$27596 ( \27911 , \27906 , \27910 );
and \U$27597 ( \27912 , \22407 , \22619 );
and \U$27598 ( \27913 , \22418 , \22617 );
nor \U$27599 ( \27914 , \27912 , \27913 );
xnor \U$27600 ( \27915 , \27914 , \22629 );
xor \U$27601 ( \27916 , \27911 , \27915 );
xor \U$27602 ( \27917 , \27902 , \27916 );
xor \U$27603 ( \27918 , \27873 , \27917 );
and \U$27604 ( \27919 , \27602 , \27608 );
and \U$27605 ( \27920 , \27608 , \27623 );
and \U$27606 ( \27921 , \27602 , \27623 );
or \U$27607 ( \27922 , \27919 , \27920 , \27921 );
and \U$27608 ( \27923 , \27568 , \27582 );
and \U$27609 ( \27924 , \27582 , \27597 );
and \U$27610 ( \27925 , \27568 , \27597 );
or \U$27611 ( \27926 , \27923 , \27924 , \27925 );
xor \U$27612 ( \27927 , \27922 , \27926 );
and \U$27613 ( \27928 , \27683 , \27697 );
and \U$27614 ( \27929 , \27697 , \27712 );
and \U$27615 ( \27930 , \27683 , \27712 );
or \U$27616 ( \27931 , \27928 , \27929 , \27930 );
xor \U$27617 ( \27932 , \27927 , \27931 );
xor \U$27618 ( \27933 , \27918 , \27932 );
and \U$27619 ( \27934 , \27544 , \27548 );
and \U$27620 ( \27935 , \27548 , \27553 );
and \U$27621 ( \27936 , \27544 , \27553 );
or \U$27622 ( \27937 , \27934 , \27935 , \27936 );
and \U$27623 ( \27938 , \27755 , \27759 );
and \U$27624 ( \27939 , \27759 , \27764 );
and \U$27625 ( \27940 , \27755 , \27764 );
or \U$27626 ( \27941 , \27938 , \27939 , \27940 );
xor \U$27627 ( \27942 , \27937 , \27941 );
and \U$27628 ( \27943 , \27629 , \27633 );
and \U$27629 ( \27944 , \27633 , \27638 );
and \U$27630 ( \27945 , \27629 , \27638 );
or \U$27631 ( \27946 , \27943 , \27944 , \27945 );
xor \U$27632 ( \27947 , \27942 , \27946 );
xor \U$27633 ( \27948 , \27933 , \27947 );
and \U$27634 ( \27949 , \27598 , \27624 );
and \U$27635 ( \27950 , \27624 , \27639 );
and \U$27636 ( \27951 , \27598 , \27639 );
or \U$27637 ( \27952 , \27949 , \27950 , \27951 );
and \U$27638 ( \27953 , \27658 , \27662 );
and \U$27639 ( \27954 , \27662 , \27667 );
and \U$27640 ( \27955 , \27658 , \27667 );
or \U$27641 ( \27956 , \27953 , \27954 , \27955 );
and \U$27642 ( \27957 , \27645 , \27649 );
and \U$27643 ( \27958 , \27649 , \27654 );
and \U$27644 ( \27959 , \27645 , \27654 );
or \U$27645 ( \27960 , \27957 , \27958 , \27959 );
xor \U$27646 ( \27961 , \27956 , \27960 );
and \U$27647 ( \27962 , \27702 , \27706 );
and \U$27648 ( \27963 , \27706 , \27711 );
and \U$27649 ( \27964 , \27702 , \27711 );
or \U$27650 ( \27965 , \27962 , \27963 , \27964 );
xor \U$27651 ( \27966 , \27961 , \27965 );
xor \U$27652 ( \27967 , \27952 , \27966 );
or \U$27653 ( \27968 , \27606 , \27607 );
and \U$27654 ( \27969 , \22567 , \21983 );
and \U$27655 ( \27970 , \22578 , \21981 );
nor \U$27656 ( \27971 , \27969 , \27970 );
xnor \U$27657 ( \27972 , \27971 , \21995 );
xor \U$27658 ( \27973 , \27968 , \27972 );
and \U$27659 ( \27974 , \22603 , \21978 );
xor \U$27660 ( \27975 , \27973 , \27974 );
and \U$27661 ( \27976 , \27572 , \27576 );
and \U$27662 ( \27977 , \27576 , \27581 );
and \U$27663 ( \27978 , \27572 , \27581 );
or \U$27664 ( \27979 , \27976 , \27977 , \27978 );
and \U$27665 ( \27980 , \27558 , \27562 );
and \U$27666 ( \27981 , \27562 , \27567 );
and \U$27667 ( \27982 , \27558 , \27567 );
or \U$27668 ( \27983 , \27980 , \27981 , \27982 );
xor \U$27669 ( \27984 , \27979 , \27983 );
and \U$27670 ( \27985 , \27613 , \27617 );
and \U$27671 ( \27986 , \27617 , \27622 );
and \U$27672 ( \27987 , \27613 , \27622 );
or \U$27673 ( \27988 , \27985 , \27986 , \27987 );
xor \U$27674 ( \27989 , \27984 , \27988 );
xor \U$27675 ( \27990 , \27975 , \27989 );
and \U$27676 ( \27991 , \27687 , \27691 );
and \U$27677 ( \27992 , \27691 , \27696 );
and \U$27678 ( \27993 , \27687 , \27696 );
or \U$27679 ( \27994 , \27991 , \27992 , \27993 );
and \U$27680 ( \27995 , \27673 , \27677 );
and \U$27681 ( \27996 , \27677 , \27682 );
and \U$27682 ( \27997 , \27673 , \27682 );
or \U$27683 ( \27998 , \27995 , \27996 , \27997 );
xor \U$27684 ( \27999 , \27994 , \27998 );
and \U$27685 ( \28000 , \27587 , \27591 );
and \U$27686 ( \28001 , \27591 , \27596 );
and \U$27687 ( \28002 , \27587 , \27596 );
or \U$27688 ( \28003 , \28000 , \28001 , \28002 );
xor \U$27689 ( \28004 , \27999 , \28003 );
xor \U$27690 ( \28005 , \27990 , \28004 );
xor \U$27691 ( \28006 , \27967 , \28005 );
xor \U$27692 ( \28007 , \27948 , \28006 );
and \U$27693 ( \28008 , \27529 , \27533 );
and \U$27694 ( \28009 , \27533 , \27538 );
and \U$27695 ( \28010 , \27529 , \27538 );
or \U$27696 ( \28011 , \28008 , \28009 , \28010 );
and \U$27697 ( \28012 , \27515 , \27519 );
and \U$27698 ( \28013 , \27519 , \27524 );
and \U$27699 ( \28014 , \27515 , \27524 );
or \U$27700 ( \28015 , \28012 , \28013 , \28014 );
xor \U$27701 ( \28016 , \28011 , \28015 );
and \U$27702 ( \28017 , \27655 , \27668 );
and \U$27703 ( \28018 , \27668 , \27713 );
and \U$27704 ( \28019 , \27655 , \27713 );
or \U$27705 ( \28020 , \28017 , \28018 , \28019 );
xor \U$27706 ( \28021 , \28016 , \28020 );
xor \U$27707 ( \28022 , \28007 , \28021 );
xor \U$27708 ( \28023 , \27787 , \28022 );
xor \U$27709 ( \28024 , \27778 , \28023 );
and \U$27710 ( \28025 , \27737 , \27741 );
and \U$27711 ( \28026 , \27741 , \27766 );
and \U$27712 ( \28027 , \27737 , \27766 );
or \U$27713 ( \28028 , \28025 , \28026 , \28027 );
and \U$27714 ( \28029 , \27511 , \27716 );
and \U$27715 ( \28030 , \27716 , \27731 );
and \U$27716 ( \28031 , \27511 , \27731 );
or \U$27717 ( \28032 , \28029 , \28030 , \28031 );
xor \U$27718 ( \28033 , \28028 , \28032 );
and \U$27719 ( \28034 , \27501 , \27505 );
and \U$27720 ( \28035 , \27505 , \27510 );
and \U$27721 ( \28036 , \27501 , \27510 );
or \U$27722 ( \28037 , \28034 , \28035 , \28036 );
and \U$27723 ( \28038 , \27746 , \27750 );
and \U$27724 ( \28039 , \27750 , \27765 );
and \U$27725 ( \28040 , \27746 , \27765 );
or \U$27726 ( \28041 , \28038 , \28039 , \28040 );
xor \U$27727 ( \28042 , \28037 , \28041 );
and \U$27728 ( \28043 , \27554 , \27640 );
and \U$27729 ( \28044 , \27640 , \27714 );
and \U$27730 ( \28045 , \27554 , \27714 );
or \U$27731 ( \28046 , \28043 , \28044 , \28045 );
xor \U$27732 ( \28047 , \28042 , \28046 );
xor \U$27733 ( \28048 , \28033 , \28047 );
xor \U$27734 ( \28049 , \28024 , \28048 );
and \U$27735 ( \28050 , \27493 , \27768 );
nor \U$27736 ( \28051 , \28049 , \28050 );
nor \U$27737 ( \28052 , \27774 , \28051 );
nand \U$27738 ( \28053 , \27489 , \28052 );
and \U$27739 ( \28054 , \28028 , \28032 );
and \U$27740 ( \28055 , \28032 , \28047 );
and \U$27741 ( \28056 , \28028 , \28047 );
or \U$27742 ( \28057 , \28054 , \28055 , \28056 );
and \U$27743 ( \28058 , \27782 , \27786 );
and \U$27744 ( \28059 , \27786 , \28022 );
and \U$27745 ( \28060 , \27782 , \28022 );
or \U$27746 ( \28061 , \28058 , \28059 , \28060 );
and \U$27747 ( \28062 , \28011 , \28015 );
and \U$27748 ( \28063 , \28015 , \28020 );
and \U$27749 ( \28064 , \28011 , \28020 );
or \U$27750 ( \28065 , \28062 , \28063 , \28064 );
and \U$27751 ( \28066 , \27952 , \27966 );
and \U$27752 ( \28067 , \27966 , \28005 );
and \U$27753 ( \28068 , \27952 , \28005 );
or \U$27754 ( \28069 , \28066 , \28067 , \28068 );
xor \U$27755 ( \28070 , \28065 , \28069 );
and \U$27756 ( \28071 , \27918 , \27932 );
and \U$27757 ( \28072 , \27932 , \27947 );
and \U$27758 ( \28073 , \27918 , \27947 );
or \U$27759 ( \28074 , \28071 , \28072 , \28073 );
xor \U$27760 ( \28075 , \28070 , \28074 );
xor \U$27761 ( \28076 , \28061 , \28075 );
and \U$27762 ( \28077 , \28037 , \28041 );
and \U$27763 ( \28078 , \28041 , \28046 );
and \U$27764 ( \28079 , \28037 , \28046 );
or \U$27765 ( \28080 , \28077 , \28078 , \28079 );
and \U$27766 ( \28081 , \27948 , \28006 );
and \U$27767 ( \28082 , \28006 , \28021 );
and \U$27768 ( \28083 , \27948 , \28021 );
or \U$27769 ( \28084 , \28081 , \28082 , \28083 );
xor \U$27770 ( \28085 , \28080 , \28084 );
and \U$27771 ( \28086 , \27801 , \27815 );
and \U$27772 ( \28087 , \27815 , \27827 );
and \U$27773 ( \28088 , \27801 , \27827 );
or \U$27774 ( \28089 , \28086 , \28087 , \28088 );
and \U$27775 ( \28090 , \22894 , \22257 );
and \U$27776 ( \28091 , \23230 , \22255 );
nor \U$27777 ( \28092 , \28090 , \28091 );
xnor \U$27778 ( \28093 , \28092 , \22267 );
and \U$27779 ( \28094 , \22081 , \22278 );
and \U$27780 ( \28095 , \22858 , \22276 );
nor \U$27781 ( \28096 , \28094 , \28095 );
xnor \U$27782 ( \28097 , \28096 , \22288 );
xor \U$27783 ( \28098 , \28093 , \28097 );
and \U$27784 ( \28099 , \22100 , \22300 );
and \U$27785 ( \28100 , \22071 , \22298 );
nor \U$27786 ( \28101 , \28099 , \28100 );
xnor \U$27787 ( \28102 , \28101 , \22310 );
xor \U$27788 ( \28103 , \28098 , \28102 );
xor \U$27789 ( \28104 , \28089 , \28103 );
and \U$27790 ( \28105 , \21990 , \22187 );
not \U$27791 ( \28106 , \28105 );
xnor \U$27792 ( \28107 , \28106 , \22197 );
and \U$27793 ( \28108 , \22001 , \22208 );
and \U$27794 ( \28109 , \21977 , \22206 );
nor \U$27795 ( \28110 , \28108 , \28109 );
xnor \U$27796 ( \28111 , \28110 , \22218 );
xor \U$27797 ( \28112 , \28107 , \28111 );
and \U$27798 ( \28113 , \23329 , \22230 );
and \U$27799 ( \28114 , \22030 , \22228 );
nor \U$27800 ( \28115 , \28113 , \28114 );
xnor \U$27801 ( \28116 , \28115 , \22240 );
xor \U$27802 ( \28117 , \28112 , \28116 );
xor \U$27803 ( \28118 , \28104 , \28117 );
and \U$27804 ( \28119 , \27968 , \27972 );
and \U$27805 ( \28120 , \27972 , \27974 );
and \U$27806 ( \28121 , \27968 , \27974 );
or \U$27807 ( \28122 , \28119 , \28120 , \28121 );
and \U$27808 ( \28123 , \27887 , \27901 );
and \U$27809 ( \28124 , \27901 , \27916 );
and \U$27810 ( \28125 , \27887 , \27916 );
or \U$27811 ( \28126 , \28123 , \28124 , \28125 );
xor \U$27812 ( \28127 , \28122 , \28126 );
and \U$27813 ( \28128 , \27842 , \27856 );
and \U$27814 ( \28129 , \27856 , \27871 );
and \U$27815 ( \28130 , \27842 , \27871 );
or \U$27816 ( \28131 , \28128 , \28129 , \28130 );
xor \U$27817 ( \28132 , \28127 , \28131 );
xor \U$27818 ( \28133 , \28118 , \28132 );
and \U$27819 ( \28134 , \27956 , \27960 );
and \U$27820 ( \28135 , \27960 , \27965 );
and \U$27821 ( \28136 , \27956 , \27965 );
or \U$27822 ( \28137 , \28134 , \28135 , \28136 );
and \U$27823 ( \28138 , \27994 , \27998 );
and \U$27824 ( \28139 , \27998 , \28003 );
and \U$27825 ( \28140 , \27994 , \28003 );
or \U$27826 ( \28141 , \28138 , \28139 , \28140 );
xor \U$27827 ( \28142 , \28137 , \28141 );
and \U$27828 ( \28143 , \27979 , \27983 );
and \U$27829 ( \28144 , \27983 , \27988 );
and \U$27830 ( \28145 , \27979 , \27988 );
or \U$27831 ( \28146 , \28143 , \28144 , \28145 );
xor \U$27832 ( \28147 , \28142 , \28146 );
xor \U$27833 ( \28148 , \28133 , \28147 );
and \U$27834 ( \28149 , \27975 , \27989 );
and \U$27835 ( \28150 , \27989 , \28004 );
and \U$27836 ( \28151 , \27975 , \28004 );
or \U$27837 ( \28152 , \28149 , \28150 , \28151 );
and \U$27838 ( \28153 , \27906 , \27910 );
and \U$27839 ( \28154 , \27910 , \27915 );
and \U$27840 ( \28155 , \27906 , \27915 );
or \U$27841 ( \28156 , \28153 , \28154 , \28155 );
and \U$27842 ( \28157 , \27891 , \27895 );
and \U$27843 ( \28158 , \27895 , \27900 );
and \U$27844 ( \28159 , \27891 , \27900 );
or \U$27845 ( \28160 , \28157 , \28158 , \28159 );
xor \U$27846 ( \28161 , \28156 , \28160 );
and \U$27847 ( \28162 , \27877 , \27881 );
and \U$27848 ( \28163 , \27881 , \27886 );
and \U$27849 ( \28164 , \27877 , \27886 );
or \U$27850 ( \28165 , \28162 , \28163 , \28164 );
xor \U$27851 ( \28166 , \28161 , \28165 );
and \U$27852 ( \28167 , \27861 , \27865 );
and \U$27853 ( \28168 , \27865 , \27870 );
and \U$27854 ( \28169 , \27861 , \27870 );
or \U$27855 ( \28170 , \28167 , \28168 , \28169 );
and \U$27856 ( \28171 , \27846 , \27850 );
and \U$27857 ( \28172 , \27850 , \27855 );
and \U$27858 ( \28173 , \27846 , \27855 );
or \U$27859 ( \28174 , \28171 , \28172 , \28173 );
xor \U$27860 ( \28175 , \28170 , \28174 );
and \U$27861 ( \28176 , \27832 , \27836 );
and \U$27862 ( \28177 , \27836 , \27841 );
and \U$27863 ( \28178 , \27832 , \27841 );
or \U$27864 ( \28179 , \28176 , \28177 , \28178 );
xor \U$27865 ( \28180 , \28175 , \28179 );
xor \U$27866 ( \28181 , \28166 , \28180 );
and \U$27867 ( \28182 , \27817 , \27821 );
and \U$27868 ( \28183 , \27821 , \27826 );
and \U$27869 ( \28184 , \27817 , \27826 );
or \U$27870 ( \28185 , \28182 , \28183 , \28184 );
and \U$27871 ( \28186 , \27805 , \27809 );
and \U$27872 ( \28187 , \27809 , \27814 );
and \U$27873 ( \28188 , \27805 , \27814 );
or \U$27874 ( \28189 , \28186 , \28187 , \28188 );
xor \U$27875 ( \28190 , \28185 , \28189 );
and \U$27876 ( \28191 , \27791 , \27795 );
and \U$27877 ( \28192 , \27795 , \27800 );
and \U$27878 ( \28193 , \27791 , \27800 );
or \U$27879 ( \28194 , \28191 , \28192 , \28193 );
xor \U$27880 ( \28195 , \28190 , \28194 );
xor \U$27881 ( \28196 , \28181 , \28195 );
xor \U$27882 ( \28197 , \28152 , \28196 );
and \U$27883 ( \28198 , \22262 , \22463 );
and \U$27884 ( \28199 , \22224 , \22461 );
nor \U$27885 ( \28200 , \28198 , \28199 );
xnor \U$27886 ( \28201 , \28200 , \22473 );
and \U$27887 ( \28202 , \22283 , \22484 );
and \U$27888 ( \28203 , \22251 , \22482 );
nor \U$27889 ( \28204 , \28202 , \28203 );
xnor \U$27890 ( \28205 , \28204 , \22494 );
xor \U$27891 ( \28206 , \28201 , \28205 );
and \U$27892 ( \28207 , \22305 , \22506 );
and \U$27893 ( \28208 , \22272 , \22504 );
nor \U$27894 ( \28209 , \28207 , \28208 );
xnor \U$27895 ( \28210 , \28209 , \22516 );
xor \U$27896 ( \28211 , \28206 , \28210 );
and \U$27897 ( \28212 , \22192 , \22392 );
and \U$27898 ( \28213 , \22156 , \22390 );
nor \U$27899 ( \28214 , \28212 , \28213 );
xnor \U$27900 ( \28215 , \28214 , \22402 );
and \U$27901 ( \28216 , \22213 , \22413 );
and \U$27902 ( \28217 , \22181 , \22411 );
nor \U$27903 ( \28218 , \28216 , \28217 );
xnor \U$27904 ( \28219 , \28218 , \22423 );
xor \U$27905 ( \28220 , \28215 , \28219 );
and \U$27906 ( \28221 , \22235 , \22435 );
and \U$27907 ( \28222 , \22202 , \22433 );
nor \U$27908 ( \28223 , \28221 , \28222 );
xnor \U$27909 ( \28224 , \28223 , \22445 );
xor \U$27910 ( \28225 , \28220 , \28224 );
xor \U$27911 ( \28226 , \28211 , \28225 );
and \U$27912 ( \28227 , \22124 , \22324 );
and \U$27913 ( \28228 , \22089 , \22322 );
nor \U$27914 ( \28229 , \28227 , \28228 );
xnor \U$27915 ( \28230 , \28229 , \22334 );
and \U$27916 ( \28231 , \22145 , \22345 );
and \U$27917 ( \28232 , \22113 , \22343 );
nor \U$27918 ( \28233 , \28231 , \28232 );
xnor \U$27919 ( \28234 , \28233 , \22355 );
xor \U$27920 ( \28235 , \28230 , \28234 );
and \U$27921 ( \28236 , \22167 , \22367 );
and \U$27922 ( \28237 , \22134 , \22365 );
nor \U$27923 ( \28238 , \28236 , \28237 );
xnor \U$27924 ( \28239 , \28238 , \22377 );
xor \U$27925 ( \28240 , \28235 , \28239 );
xor \U$27926 ( \28241 , \28226 , \28240 );
and \U$27927 ( \28242 , \22468 , \22671 );
and \U$27928 ( \28243 , \22429 , \22669 );
nor \U$27929 ( \28244 , \28242 , \28243 );
xnor \U$27930 ( \28245 , \28244 , \22681 );
and \U$27931 ( \28246 , \22489 , \22691 );
and \U$27932 ( \28247 , \22457 , \22689 );
nor \U$27933 ( \28248 , \28246 , \28247 );
xnor \U$27934 ( \28249 , \28248 , \22701 );
xor \U$27935 ( \28250 , \28245 , \28249 );
and \U$27936 ( \28251 , \22511 , \22720 );
and \U$27937 ( \28252 , \22478 , \22707 );
nor \U$27938 ( \28253 , \28251 , \28252 );
xnor \U$27939 ( \28254 , \28253 , \22067 );
xor \U$27940 ( \28255 , \28250 , \28254 );
and \U$27941 ( \28256 , \22397 , \22598 );
and \U$27942 ( \28257 , \22361 , \22596 );
nor \U$27943 ( \28258 , \28256 , \28257 );
xnor \U$27944 ( \28259 , \28258 , \22608 );
and \U$27945 ( \28260 , \22418 , \22619 );
and \U$27946 ( \28261 , \22386 , \22617 );
nor \U$27947 ( \28262 , \28260 , \28261 );
xnor \U$27948 ( \28263 , \28262 , \22629 );
xor \U$27949 ( \28264 , \28259 , \28263 );
and \U$27950 ( \28265 , \22440 , \22641 );
and \U$27951 ( \28266 , \22407 , \22639 );
nor \U$27952 ( \28267 , \28265 , \28266 );
xnor \U$27953 ( \28268 , \28267 , \22651 );
xor \U$27954 ( \28269 , \28264 , \28268 );
xor \U$27955 ( \28270 , \28255 , \28269 );
and \U$27956 ( \28271 , \22329 , \22530 );
and \U$27957 ( \28272 , \22294 , \22528 );
nor \U$27958 ( \28273 , \28271 , \28272 );
xnor \U$27959 ( \28274 , \28273 , \22540 );
and \U$27960 ( \28275 , \22350 , \22551 );
and \U$27961 ( \28276 , \22318 , \22549 );
nor \U$27962 ( \28277 , \28275 , \28276 );
xnor \U$27963 ( \28278 , \28277 , \22561 );
xor \U$27964 ( \28279 , \28274 , \28278 );
and \U$27965 ( \28280 , \22372 , \22573 );
and \U$27966 ( \28281 , \22339 , \22571 );
nor \U$27967 ( \28282 , \28280 , \28281 );
xnor \U$27968 ( \28283 , \28282 , \22583 );
xor \U$27969 ( \28284 , \28279 , \28283 );
xor \U$27970 ( \28285 , \28270 , \28284 );
xor \U$27971 ( \28286 , \28241 , \28285 );
and \U$27972 ( \28287 , \22567 , \21978 );
and \U$27973 ( \28288 , \22535 , \23173 );
and \U$27974 ( \28289 , \22500 , \22999 );
nor \U$27975 ( \28290 , \28288 , \28289 );
xnor \U$27976 ( \28291 , \28290 , \22016 );
and \U$27977 ( \28292 , \22556 , \22021 );
and \U$27978 ( \28293 , \22524 , \22019 );
nor \U$27979 ( \28294 , \28292 , \28293 );
xnor \U$27980 ( \28295 , \28294 , \21595 );
xor \U$27981 ( \28296 , \28291 , \28295 );
and \U$27982 ( \28297 , \22578 , \21983 );
and \U$27983 ( \28298 , \22545 , \21981 );
nor \U$27984 ( \28299 , \28297 , \28298 );
xnor \U$27985 ( \28300 , \28299 , \21995 );
xor \U$27986 ( \28301 , \28296 , \28300 );
xnor \U$27987 ( \28302 , \28287 , \28301 );
xor \U$27988 ( \28303 , \28286 , \28302 );
xor \U$27989 ( \28304 , \28197 , \28303 );
xor \U$27990 ( \28305 , \28148 , \28304 );
and \U$27991 ( \28306 , \27937 , \27941 );
and \U$27992 ( \28307 , \27941 , \27946 );
and \U$27993 ( \28308 , \27937 , \27946 );
or \U$27994 ( \28309 , \28306 , \28307 , \28308 );
and \U$27995 ( \28310 , \27922 , \27926 );
and \U$27996 ( \28311 , \27926 , \27931 );
and \U$27997 ( \28312 , \27922 , \27931 );
or \U$27998 ( \28313 , \28310 , \28311 , \28312 );
xor \U$27999 ( \28314 , \28309 , \28313 );
and \U$28000 ( \28315 , \27828 , \27872 );
and \U$28001 ( \28316 , \27872 , \27917 );
and \U$28002 ( \28317 , \27828 , \27917 );
or \U$28003 ( \28318 , \28315 , \28316 , \28317 );
xor \U$28004 ( \28319 , \28314 , \28318 );
xor \U$28005 ( \28320 , \28305 , \28319 );
xor \U$28006 ( \28321 , \28085 , \28320 );
xor \U$28007 ( \28322 , \28076 , \28321 );
xor \U$28008 ( \28323 , \28057 , \28322 );
and \U$28009 ( \28324 , \27778 , \28023 );
and \U$28010 ( \28325 , \28023 , \28048 );
and \U$28011 ( \28326 , \27778 , \28048 );
or \U$28012 ( \28327 , \28324 , \28325 , \28326 );
nor \U$28013 ( \28328 , \28323 , \28327 );
and \U$28014 ( \28329 , \28061 , \28075 );
and \U$28015 ( \28330 , \28075 , \28321 );
and \U$28016 ( \28331 , \28061 , \28321 );
or \U$28017 ( \28332 , \28329 , \28330 , \28331 );
and \U$28018 ( \28333 , \28080 , \28084 );
and \U$28019 ( \28334 , \28084 , \28320 );
and \U$28020 ( \28335 , \28080 , \28320 );
or \U$28021 ( \28336 , \28333 , \28334 , \28335 );
and \U$28022 ( \28337 , \28185 , \28189 );
and \U$28023 ( \28338 , \28189 , \28194 );
and \U$28024 ( \28339 , \28185 , \28194 );
or \U$28025 ( \28340 , \28337 , \28338 , \28339 );
and \U$28026 ( \28341 , \28170 , \28174 );
and \U$28027 ( \28342 , \28174 , \28179 );
and \U$28028 ( \28343 , \28170 , \28179 );
or \U$28029 ( \28344 , \28341 , \28342 , \28343 );
xor \U$28030 ( \28345 , \28340 , \28344 );
and \U$28031 ( \28346 , \28156 , \28160 );
and \U$28032 ( \28347 , \28160 , \28165 );
and \U$28033 ( \28348 , \28156 , \28165 );
or \U$28034 ( \28349 , \28346 , \28347 , \28348 );
xor \U$28035 ( \28350 , \28345 , \28349 );
and \U$28036 ( \28351 , \22578 , \21978 );
and \U$28037 ( \28352 , \22500 , \23173 );
and \U$28038 ( \28353 , \22511 , \22999 );
nor \U$28039 ( \28354 , \28352 , \28353 );
xnor \U$28040 ( \28355 , \28354 , \22016 );
and \U$28041 ( \28356 , \22524 , \22021 );
and \U$28042 ( \28357 , \22535 , \22019 );
nor \U$28043 ( \28358 , \28356 , \28357 );
xnor \U$28044 ( \28359 , \28358 , \21595 );
xor \U$28045 ( \28360 , \28355 , \28359 );
and \U$28046 ( \28361 , \22545 , \21983 );
and \U$28047 ( \28362 , \22556 , \21981 );
nor \U$28048 ( \28363 , \28361 , \28362 );
xnor \U$28049 ( \28364 , \28363 , \21995 );
xor \U$28050 ( \28365 , \28360 , \28364 );
xor \U$28051 ( \28366 , \28351 , \28365 );
and \U$28052 ( \28367 , \22429 , \22671 );
and \U$28053 ( \28368 , \22440 , \22669 );
nor \U$28054 ( \28369 , \28367 , \28368 );
xnor \U$28055 ( \28370 , \28369 , \22681 );
and \U$28056 ( \28371 , \22457 , \22691 );
and \U$28057 ( \28372 , \22468 , \22689 );
nor \U$28058 ( \28373 , \28371 , \28372 );
xnor \U$28059 ( \28374 , \28373 , \22701 );
xor \U$28060 ( \28375 , \28370 , \28374 );
and \U$28061 ( \28376 , \22478 , \22720 );
and \U$28062 ( \28377 , \22489 , \22707 );
nor \U$28063 ( \28378 , \28376 , \28377 );
xnor \U$28064 ( \28379 , \28378 , \22067 );
xor \U$28065 ( \28380 , \28375 , \28379 );
xor \U$28066 ( \28381 , \28366 , \28380 );
and \U$28067 ( \28382 , \28259 , \28263 );
and \U$28068 ( \28383 , \28263 , \28268 );
and \U$28069 ( \28384 , \28259 , \28268 );
or \U$28070 ( \28385 , \28382 , \28383 , \28384 );
and \U$28071 ( \28386 , \28245 , \28249 );
and \U$28072 ( \28387 , \28249 , \28254 );
and \U$28073 ( \28388 , \28245 , \28254 );
or \U$28074 ( \28389 , \28386 , \28387 , \28388 );
xor \U$28075 ( \28390 , \28385 , \28389 );
and \U$28076 ( \28391 , \28291 , \28295 );
and \U$28077 ( \28392 , \28295 , \28300 );
and \U$28078 ( \28393 , \28291 , \28300 );
or \U$28079 ( \28394 , \28391 , \28392 , \28393 );
xor \U$28080 ( \28395 , \28390 , \28394 );
xor \U$28081 ( \28396 , \28381 , \28395 );
and \U$28082 ( \28397 , \28215 , \28219 );
and \U$28083 ( \28398 , \28219 , \28224 );
and \U$28084 ( \28399 , \28215 , \28224 );
or \U$28085 ( \28400 , \28397 , \28398 , \28399 );
and \U$28086 ( \28401 , \28201 , \28205 );
and \U$28087 ( \28402 , \28205 , \28210 );
and \U$28088 ( \28403 , \28201 , \28210 );
or \U$28089 ( \28404 , \28401 , \28402 , \28403 );
xor \U$28090 ( \28405 , \28400 , \28404 );
and \U$28091 ( \28406 , \28274 , \28278 );
and \U$28092 ( \28407 , \28278 , \28283 );
and \U$28093 ( \28408 , \28274 , \28283 );
or \U$28094 ( \28409 , \28406 , \28407 , \28408 );
xor \U$28095 ( \28410 , \28405 , \28409 );
xor \U$28096 ( \28411 , \28396 , \28410 );
not \U$28097 ( \28412 , \22197 );
and \U$28098 ( \28413 , \21977 , \22208 );
and \U$28099 ( \28414 , \21990 , \22206 );
nor \U$28100 ( \28415 , \28413 , \28414 );
xnor \U$28101 ( \28416 , \28415 , \22218 );
xor \U$28102 ( \28417 , \28412 , \28416 );
and \U$28103 ( \28418 , \22030 , \22230 );
and \U$28104 ( \28419 , \22001 , \22228 );
nor \U$28105 ( \28420 , \28418 , \28419 );
xnor \U$28106 ( \28421 , \28420 , \22240 );
xor \U$28107 ( \28422 , \28417 , \28421 );
and \U$28108 ( \28423 , \22156 , \22392 );
and \U$28109 ( \28424 , \22167 , \22390 );
nor \U$28110 ( \28425 , \28423 , \28424 );
xnor \U$28111 ( \28426 , \28425 , \22402 );
and \U$28112 ( \28427 , \22181 , \22413 );
and \U$28113 ( \28428 , \22192 , \22411 );
nor \U$28114 ( \28429 , \28427 , \28428 );
xnor \U$28115 ( \28430 , \28429 , \22423 );
xor \U$28116 ( \28431 , \28426 , \28430 );
and \U$28117 ( \28432 , \22202 , \22435 );
and \U$28118 ( \28433 , \22213 , \22433 );
nor \U$28119 ( \28434 , \28432 , \28433 );
xnor \U$28120 ( \28435 , \28434 , \22445 );
xor \U$28121 ( \28436 , \28431 , \28435 );
and \U$28122 ( \28437 , \22089 , \22324 );
and \U$28123 ( \28438 , \22100 , \22322 );
nor \U$28124 ( \28439 , \28437 , \28438 );
xnor \U$28125 ( \28440 , \28439 , \22334 );
and \U$28126 ( \28441 , \22113 , \22345 );
and \U$28127 ( \28442 , \22124 , \22343 );
nor \U$28128 ( \28443 , \28441 , \28442 );
xnor \U$28129 ( \28444 , \28443 , \22355 );
xor \U$28130 ( \28445 , \28440 , \28444 );
and \U$28131 ( \28446 , \22134 , \22367 );
and \U$28132 ( \28447 , \22145 , \22365 );
nor \U$28133 ( \28448 , \28446 , \28447 );
xnor \U$28134 ( \28449 , \28448 , \22377 );
xor \U$28135 ( \28450 , \28445 , \28449 );
xor \U$28136 ( \28451 , \28436 , \28450 );
and \U$28137 ( \28452 , \23230 , \22257 );
and \U$28138 ( \28453 , \23329 , \22255 );
nor \U$28139 ( \28454 , \28452 , \28453 );
xnor \U$28140 ( \28455 , \28454 , \22267 );
and \U$28141 ( \28456 , \22858 , \22278 );
and \U$28142 ( \28457 , \22894 , \22276 );
nor \U$28143 ( \28458 , \28456 , \28457 );
xnor \U$28144 ( \28459 , \28458 , \22288 );
xor \U$28145 ( \28460 , \28455 , \28459 );
and \U$28146 ( \28461 , \22071 , \22300 );
and \U$28147 ( \28462 , \22081 , \22298 );
nor \U$28148 ( \28463 , \28461 , \28462 );
xnor \U$28149 ( \28464 , \28463 , \22310 );
xor \U$28150 ( \28465 , \28460 , \28464 );
xor \U$28151 ( \28466 , \28451 , \28465 );
xor \U$28152 ( \28467 , \28422 , \28466 );
and \U$28153 ( \28468 , \22361 , \22598 );
and \U$28154 ( \28469 , \22372 , \22596 );
nor \U$28155 ( \28470 , \28468 , \28469 );
xnor \U$28156 ( \28471 , \28470 , \22608 );
and \U$28157 ( \28472 , \22386 , \22619 );
and \U$28158 ( \28473 , \22397 , \22617 );
nor \U$28159 ( \28474 , \28472 , \28473 );
xnor \U$28160 ( \28475 , \28474 , \22629 );
xor \U$28161 ( \28476 , \28471 , \28475 );
and \U$28162 ( \28477 , \22407 , \22641 );
and \U$28163 ( \28478 , \22418 , \22639 );
nor \U$28164 ( \28479 , \28477 , \28478 );
xnor \U$28165 ( \28480 , \28479 , \22651 );
xor \U$28166 ( \28481 , \28476 , \28480 );
and \U$28167 ( \28482 , \22294 , \22530 );
and \U$28168 ( \28483 , \22305 , \22528 );
nor \U$28169 ( \28484 , \28482 , \28483 );
xnor \U$28170 ( \28485 , \28484 , \22540 );
and \U$28171 ( \28486 , \22318 , \22551 );
and \U$28172 ( \28487 , \22329 , \22549 );
nor \U$28173 ( \28488 , \28486 , \28487 );
xnor \U$28174 ( \28489 , \28488 , \22561 );
xor \U$28175 ( \28490 , \28485 , \28489 );
and \U$28176 ( \28491 , \22339 , \22573 );
and \U$28177 ( \28492 , \22350 , \22571 );
nor \U$28178 ( \28493 , \28491 , \28492 );
xnor \U$28179 ( \28494 , \28493 , \22583 );
xor \U$28180 ( \28495 , \28490 , \28494 );
xor \U$28181 ( \28496 , \28481 , \28495 );
and \U$28182 ( \28497 , \22224 , \22463 );
and \U$28183 ( \28498 , \22235 , \22461 );
nor \U$28184 ( \28499 , \28497 , \28498 );
xnor \U$28185 ( \28500 , \28499 , \22473 );
and \U$28186 ( \28501 , \22251 , \22484 );
and \U$28187 ( \28502 , \22262 , \22482 );
nor \U$28188 ( \28503 , \28501 , \28502 );
xnor \U$28189 ( \28504 , \28503 , \22494 );
xor \U$28190 ( \28505 , \28500 , \28504 );
and \U$28191 ( \28506 , \22272 , \22506 );
and \U$28192 ( \28507 , \22283 , \22504 );
nor \U$28193 ( \28508 , \28506 , \28507 );
xnor \U$28194 ( \28509 , \28508 , \22516 );
xor \U$28195 ( \28510 , \28505 , \28509 );
xor \U$28196 ( \28511 , \28496 , \28510 );
xor \U$28197 ( \28512 , \28467 , \28511 );
xor \U$28198 ( \28513 , \28411 , \28512 );
or \U$28199 ( \28514 , \28287 , \28301 );
and \U$28200 ( \28515 , \28255 , \28269 );
and \U$28201 ( \28516 , \28269 , \28284 );
and \U$28202 ( \28517 , \28255 , \28284 );
or \U$28203 ( \28518 , \28515 , \28516 , \28517 );
xor \U$28204 ( \28519 , \28514 , \28518 );
and \U$28205 ( \28520 , \28211 , \28225 );
and \U$28206 ( \28521 , \28225 , \28240 );
and \U$28207 ( \28522 , \28211 , \28240 );
or \U$28208 ( \28523 , \28520 , \28521 , \28522 );
xor \U$28209 ( \28524 , \28519 , \28523 );
xor \U$28210 ( \28525 , \28513 , \28524 );
xor \U$28211 ( \28526 , \28350 , \28525 );
and \U$28212 ( \28527 , \28241 , \28285 );
and \U$28213 ( \28528 , \28285 , \28302 );
and \U$28214 ( \28529 , \28241 , \28302 );
or \U$28215 ( \28530 , \28527 , \28528 , \28529 );
and \U$28216 ( \28531 , \28166 , \28180 );
and \U$28217 ( \28532 , \28180 , \28195 );
and \U$28218 ( \28533 , \28166 , \28195 );
or \U$28219 ( \28534 , \28531 , \28532 , \28533 );
xor \U$28220 ( \28535 , \28530 , \28534 );
and \U$28221 ( \28536 , \28107 , \28111 );
and \U$28222 ( \28537 , \28111 , \28116 );
and \U$28223 ( \28538 , \28107 , \28116 );
or \U$28224 ( \28539 , \28536 , \28537 , \28538 );
and \U$28225 ( \28540 , \28093 , \28097 );
and \U$28226 ( \28541 , \28097 , \28102 );
and \U$28227 ( \28542 , \28093 , \28102 );
or \U$28228 ( \28543 , \28540 , \28541 , \28542 );
xor \U$28229 ( \28544 , \28539 , \28543 );
and \U$28230 ( \28545 , \28230 , \28234 );
and \U$28231 ( \28546 , \28234 , \28239 );
and \U$28232 ( \28547 , \28230 , \28239 );
or \U$28233 ( \28548 , \28545 , \28546 , \28547 );
xor \U$28234 ( \28549 , \28544 , \28548 );
xor \U$28235 ( \28550 , \28535 , \28549 );
xor \U$28236 ( \28551 , \28526 , \28550 );
and \U$28237 ( \28552 , \28309 , \28313 );
and \U$28238 ( \28553 , \28313 , \28318 );
and \U$28239 ( \28554 , \28309 , \28318 );
or \U$28240 ( \28555 , \28552 , \28553 , \28554 );
and \U$28241 ( \28556 , \28152 , \28196 );
and \U$28242 ( \28557 , \28196 , \28303 );
and \U$28243 ( \28558 , \28152 , \28303 );
or \U$28244 ( \28559 , \28556 , \28557 , \28558 );
xor \U$28245 ( \28560 , \28555 , \28559 );
and \U$28246 ( \28561 , \28118 , \28132 );
and \U$28247 ( \28562 , \28132 , \28147 );
and \U$28248 ( \28563 , \28118 , \28147 );
or \U$28249 ( \28564 , \28561 , \28562 , \28563 );
xor \U$28250 ( \28565 , \28560 , \28564 );
xor \U$28251 ( \28566 , \28551 , \28565 );
xor \U$28252 ( \28567 , \28336 , \28566 );
and \U$28253 ( \28568 , \28065 , \28069 );
and \U$28254 ( \28569 , \28069 , \28074 );
and \U$28255 ( \28570 , \28065 , \28074 );
or \U$28256 ( \28571 , \28568 , \28569 , \28570 );
and \U$28257 ( \28572 , \28148 , \28304 );
and \U$28258 ( \28573 , \28304 , \28319 );
and \U$28259 ( \28574 , \28148 , \28319 );
or \U$28260 ( \28575 , \28572 , \28573 , \28574 );
xor \U$28261 ( \28576 , \28571 , \28575 );
and \U$28262 ( \28577 , \28137 , \28141 );
and \U$28263 ( \28578 , \28141 , \28146 );
and \U$28264 ( \28579 , \28137 , \28146 );
or \U$28265 ( \28580 , \28577 , \28578 , \28579 );
and \U$28266 ( \28581 , \28122 , \28126 );
and \U$28267 ( \28582 , \28126 , \28131 );
and \U$28268 ( \28583 , \28122 , \28131 );
or \U$28269 ( \28584 , \28581 , \28582 , \28583 );
xor \U$28270 ( \28585 , \28580 , \28584 );
and \U$28271 ( \28586 , \28089 , \28103 );
and \U$28272 ( \28587 , \28103 , \28117 );
and \U$28273 ( \28588 , \28089 , \28117 );
or \U$28274 ( \28589 , \28586 , \28587 , \28588 );
xor \U$28275 ( \28590 , \28585 , \28589 );
xor \U$28276 ( \28591 , \28576 , \28590 );
xor \U$28277 ( \28592 , \28567 , \28591 );
xor \U$28278 ( \28593 , \28332 , \28592 );
and \U$28279 ( \28594 , \28057 , \28322 );
nor \U$28280 ( \28595 , \28593 , \28594 );
nor \U$28281 ( \28596 , \28328 , \28595 );
and \U$28282 ( \28597 , \28336 , \28566 );
and \U$28283 ( \28598 , \28566 , \28591 );
and \U$28284 ( \28599 , \28336 , \28591 );
or \U$28285 ( \28600 , \28597 , \28598 , \28599 );
and \U$28286 ( \28601 , \28555 , \28559 );
and \U$28287 ( \28602 , \28559 , \28564 );
and \U$28288 ( \28603 , \28555 , \28564 );
or \U$28289 ( \28604 , \28601 , \28602 , \28603 );
and \U$28290 ( \28605 , \28350 , \28525 );
and \U$28291 ( \28606 , \28525 , \28550 );
and \U$28292 ( \28607 , \28350 , \28550 );
or \U$28293 ( \28608 , \28605 , \28606 , \28607 );
xor \U$28294 ( \28609 , \28604 , \28608 );
and \U$28295 ( \28610 , \21990 , \22208 );
not \U$28296 ( \28611 , \28610 );
xnor \U$28297 ( \28612 , \28611 , \22218 );
and \U$28298 ( \28613 , \22001 , \22230 );
and \U$28299 ( \28614 , \21977 , \22228 );
nor \U$28300 ( \28615 , \28613 , \28614 );
xnor \U$28301 ( \28616 , \28615 , \22240 );
xor \U$28302 ( \28617 , \28612 , \28616 );
and \U$28303 ( \28618 , \23329 , \22257 );
and \U$28304 ( \28619 , \22030 , \22255 );
nor \U$28305 ( \28620 , \28618 , \28619 );
xnor \U$28306 ( \28621 , \28620 , \22267 );
xor \U$28307 ( \28622 , \28617 , \28621 );
and \U$28308 ( \28623 , \22192 , \22413 );
and \U$28309 ( \28624 , \22156 , \22411 );
nor \U$28310 ( \28625 , \28623 , \28624 );
xnor \U$28311 ( \28626 , \28625 , \22423 );
and \U$28312 ( \28627 , \22213 , \22435 );
and \U$28313 ( \28628 , \22181 , \22433 );
nor \U$28314 ( \28629 , \28627 , \28628 );
xnor \U$28315 ( \28630 , \28629 , \22445 );
xor \U$28316 ( \28631 , \28626 , \28630 );
and \U$28317 ( \28632 , \22235 , \22463 );
and \U$28318 ( \28633 , \22202 , \22461 );
nor \U$28319 ( \28634 , \28632 , \28633 );
xnor \U$28320 ( \28635 , \28634 , \22473 );
xor \U$28321 ( \28636 , \28631 , \28635 );
and \U$28322 ( \28637 , \22124 , \22345 );
and \U$28323 ( \28638 , \22089 , \22343 );
nor \U$28324 ( \28639 , \28637 , \28638 );
xnor \U$28325 ( \28640 , \28639 , \22355 );
and \U$28326 ( \28641 , \22145 , \22367 );
and \U$28327 ( \28642 , \22113 , \22365 );
nor \U$28328 ( \28643 , \28641 , \28642 );
xnor \U$28329 ( \28644 , \28643 , \22377 );
xor \U$28330 ( \28645 , \28640 , \28644 );
and \U$28331 ( \28646 , \22167 , \22392 );
and \U$28332 ( \28647 , \22134 , \22390 );
nor \U$28333 ( \28648 , \28646 , \28647 );
xnor \U$28334 ( \28649 , \28648 , \22402 );
xor \U$28335 ( \28650 , \28645 , \28649 );
xor \U$28336 ( \28651 , \28636 , \28650 );
and \U$28337 ( \28652 , \22894 , \22278 );
and \U$28338 ( \28653 , \23230 , \22276 );
nor \U$28339 ( \28654 , \28652 , \28653 );
xnor \U$28340 ( \28655 , \28654 , \22288 );
and \U$28341 ( \28656 , \22081 , \22300 );
and \U$28342 ( \28657 , \22858 , \22298 );
nor \U$28343 ( \28658 , \28656 , \28657 );
xnor \U$28344 ( \28659 , \28658 , \22310 );
xor \U$28345 ( \28660 , \28655 , \28659 );
and \U$28346 ( \28661 , \22100 , \22324 );
and \U$28347 ( \28662 , \22071 , \22322 );
nor \U$28348 ( \28663 , \28661 , \28662 );
xnor \U$28349 ( \28664 , \28663 , \22334 );
xor \U$28350 ( \28665 , \28660 , \28664 );
xor \U$28351 ( \28666 , \28651 , \28665 );
xor \U$28352 ( \28667 , \28622 , \28666 );
and \U$28353 ( \28668 , \22397 , \22619 );
and \U$28354 ( \28669 , \22361 , \22617 );
nor \U$28355 ( \28670 , \28668 , \28669 );
xnor \U$28356 ( \28671 , \28670 , \22629 );
and \U$28357 ( \28672 , \22418 , \22641 );
and \U$28358 ( \28673 , \22386 , \22639 );
nor \U$28359 ( \28674 , \28672 , \28673 );
xnor \U$28360 ( \28675 , \28674 , \22651 );
xor \U$28361 ( \28676 , \28671 , \28675 );
and \U$28362 ( \28677 , \22440 , \22671 );
and \U$28363 ( \28678 , \22407 , \22669 );
nor \U$28364 ( \28679 , \28677 , \28678 );
xnor \U$28365 ( \28680 , \28679 , \22681 );
xor \U$28366 ( \28681 , \28676 , \28680 );
and \U$28367 ( \28682 , \22329 , \22551 );
and \U$28368 ( \28683 , \22294 , \22549 );
nor \U$28369 ( \28684 , \28682 , \28683 );
xnor \U$28370 ( \28685 , \28684 , \22561 );
and \U$28371 ( \28686 , \22350 , \22573 );
and \U$28372 ( \28687 , \22318 , \22571 );
nor \U$28373 ( \28688 , \28686 , \28687 );
xnor \U$28374 ( \28689 , \28688 , \22583 );
xor \U$28375 ( \28690 , \28685 , \28689 );
and \U$28376 ( \28691 , \22372 , \22598 );
and \U$28377 ( \28692 , \22339 , \22596 );
nor \U$28378 ( \28693 , \28691 , \28692 );
xnor \U$28379 ( \28694 , \28693 , \22608 );
xor \U$28380 ( \28695 , \28690 , \28694 );
xor \U$28381 ( \28696 , \28681 , \28695 );
and \U$28382 ( \28697 , \22262 , \22484 );
and \U$28383 ( \28698 , \22224 , \22482 );
nor \U$28384 ( \28699 , \28697 , \28698 );
xnor \U$28385 ( \28700 , \28699 , \22494 );
and \U$28386 ( \28701 , \22283 , \22506 );
and \U$28387 ( \28702 , \22251 , \22504 );
nor \U$28388 ( \28703 , \28701 , \28702 );
xnor \U$28389 ( \28704 , \28703 , \22516 );
xor \U$28390 ( \28705 , \28700 , \28704 );
and \U$28391 ( \28706 , \22305 , \22530 );
and \U$28392 ( \28707 , \22272 , \22528 );
nor \U$28393 ( \28708 , \28706 , \28707 );
xnor \U$28394 ( \28709 , \28708 , \22540 );
xor \U$28395 ( \28710 , \28705 , \28709 );
xor \U$28396 ( \28711 , \28696 , \28710 );
xor \U$28397 ( \28712 , \28667 , \28711 );
and \U$28398 ( \28713 , \28351 , \28365 );
and \U$28399 ( \28714 , \28365 , \28380 );
and \U$28400 ( \28715 , \28351 , \28380 );
or \U$28401 ( \28716 , \28713 , \28714 , \28715 );
and \U$28402 ( \28717 , \28481 , \28495 );
and \U$28403 ( \28718 , \28495 , \28510 );
and \U$28404 ( \28719 , \28481 , \28510 );
or \U$28405 ( \28720 , \28717 , \28718 , \28719 );
xor \U$28406 ( \28721 , \28716 , \28720 );
and \U$28407 ( \28722 , \28436 , \28450 );
and \U$28408 ( \28723 , \28450 , \28465 );
and \U$28409 ( \28724 , \28436 , \28465 );
or \U$28410 ( \28725 , \28722 , \28723 , \28724 );
xor \U$28411 ( \28726 , \28721 , \28725 );
xor \U$28412 ( \28727 , \28712 , \28726 );
and \U$28413 ( \28728 , \28539 , \28543 );
and \U$28414 ( \28729 , \28543 , \28548 );
and \U$28415 ( \28730 , \28539 , \28548 );
or \U$28416 ( \28731 , \28728 , \28729 , \28730 );
and \U$28417 ( \28732 , \28400 , \28404 );
and \U$28418 ( \28733 , \28404 , \28409 );
and \U$28419 ( \28734 , \28400 , \28409 );
or \U$28420 ( \28735 , \28732 , \28733 , \28734 );
xor \U$28421 ( \28736 , \28731 , \28735 );
and \U$28422 ( \28737 , \28385 , \28389 );
and \U$28423 ( \28738 , \28389 , \28394 );
and \U$28424 ( \28739 , \28385 , \28394 );
or \U$28425 ( \28740 , \28737 , \28738 , \28739 );
xor \U$28426 ( \28741 , \28736 , \28740 );
xor \U$28427 ( \28742 , \28727 , \28741 );
and \U$28428 ( \28743 , \28381 , \28395 );
and \U$28429 ( \28744 , \28395 , \28410 );
and \U$28430 ( \28745 , \28381 , \28410 );
or \U$28431 ( \28746 , \28743 , \28744 , \28745 );
and \U$28432 ( \28747 , \28412 , \28416 );
and \U$28433 ( \28748 , \28416 , \28421 );
and \U$28434 ( \28749 , \28412 , \28421 );
or \U$28435 ( \28750 , \28747 , \28748 , \28749 );
and \U$28436 ( \28751 , \28455 , \28459 );
and \U$28437 ( \28752 , \28459 , \28464 );
and \U$28438 ( \28753 , \28455 , \28464 );
or \U$28439 ( \28754 , \28751 , \28752 , \28753 );
xor \U$28440 ( \28755 , \28750 , \28754 );
and \U$28441 ( \28756 , \28440 , \28444 );
and \U$28442 ( \28757 , \28444 , \28449 );
and \U$28443 ( \28758 , \28440 , \28449 );
or \U$28444 ( \28759 , \28756 , \28757 , \28758 );
xor \U$28445 ( \28760 , \28755 , \28759 );
xor \U$28446 ( \28761 , \28746 , \28760 );
and \U$28447 ( \28762 , \22535 , \22021 );
and \U$28448 ( \28763 , \22500 , \22019 );
nor \U$28449 ( \28764 , \28762 , \28763 );
xnor \U$28450 ( \28765 , \28764 , \21595 );
and \U$28451 ( \28766 , \22556 , \21983 );
and \U$28452 ( \28767 , \22524 , \21981 );
nor \U$28453 ( \28768 , \28766 , \28767 );
xnor \U$28454 ( \28769 , \28768 , \21995 );
xor \U$28455 ( \28770 , \28765 , \28769 );
and \U$28456 ( \28771 , \22545 , \21978 );
xor \U$28457 ( \28772 , \28770 , \28771 );
and \U$28458 ( \28773 , \22468 , \22691 );
and \U$28459 ( \28774 , \22429 , \22689 );
nor \U$28460 ( \28775 , \28773 , \28774 );
xnor \U$28461 ( \28776 , \28775 , \22701 );
and \U$28462 ( \28777 , \22489 , \22720 );
and \U$28463 ( \28778 , \22457 , \22707 );
nor \U$28464 ( \28779 , \28777 , \28778 );
xnor \U$28465 ( \28780 , \28779 , \22067 );
xor \U$28466 ( \28781 , \28776 , \28780 );
and \U$28467 ( \28782 , \22511 , \23173 );
and \U$28468 ( \28783 , \22478 , \22999 );
nor \U$28469 ( \28784 , \28782 , \28783 );
xnor \U$28470 ( \28785 , \28784 , \22016 );
xor \U$28471 ( \28786 , \28781 , \28785 );
xnor \U$28472 ( \28787 , \28772 , \28786 );
and \U$28473 ( \28788 , \28471 , \28475 );
and \U$28474 ( \28789 , \28475 , \28480 );
and \U$28475 ( \28790 , \28471 , \28480 );
or \U$28476 ( \28791 , \28788 , \28789 , \28790 );
and \U$28477 ( \28792 , \28370 , \28374 );
and \U$28478 ( \28793 , \28374 , \28379 );
and \U$28479 ( \28794 , \28370 , \28379 );
or \U$28480 ( \28795 , \28792 , \28793 , \28794 );
xor \U$28481 ( \28796 , \28791 , \28795 );
and \U$28482 ( \28797 , \28355 , \28359 );
and \U$28483 ( \28798 , \28359 , \28364 );
and \U$28484 ( \28799 , \28355 , \28364 );
or \U$28485 ( \28800 , \28797 , \28798 , \28799 );
xor \U$28486 ( \28801 , \28796 , \28800 );
xor \U$28487 ( \28802 , \28787 , \28801 );
and \U$28488 ( \28803 , \28426 , \28430 );
and \U$28489 ( \28804 , \28430 , \28435 );
and \U$28490 ( \28805 , \28426 , \28435 );
or \U$28491 ( \28806 , \28803 , \28804 , \28805 );
and \U$28492 ( \28807 , \28500 , \28504 );
and \U$28493 ( \28808 , \28504 , \28509 );
and \U$28494 ( \28809 , \28500 , \28509 );
or \U$28495 ( \28810 , \28807 , \28808 , \28809 );
xor \U$28496 ( \28811 , \28806 , \28810 );
and \U$28497 ( \28812 , \28485 , \28489 );
and \U$28498 ( \28813 , \28489 , \28494 );
and \U$28499 ( \28814 , \28485 , \28494 );
or \U$28500 ( \28815 , \28812 , \28813 , \28814 );
xor \U$28501 ( \28816 , \28811 , \28815 );
xor \U$28502 ( \28817 , \28802 , \28816 );
xor \U$28503 ( \28818 , \28761 , \28817 );
xor \U$28504 ( \28819 , \28742 , \28818 );
and \U$28505 ( \28820 , \28340 , \28344 );
and \U$28506 ( \28821 , \28344 , \28349 );
and \U$28507 ( \28822 , \28340 , \28349 );
or \U$28508 ( \28823 , \28820 , \28821 , \28822 );
and \U$28509 ( \28824 , \28514 , \28518 );
and \U$28510 ( \28825 , \28518 , \28523 );
and \U$28511 ( \28826 , \28514 , \28523 );
or \U$28512 ( \28827 , \28824 , \28825 , \28826 );
xor \U$28513 ( \28828 , \28823 , \28827 );
and \U$28514 ( \28829 , \28422 , \28466 );
and \U$28515 ( \28830 , \28466 , \28511 );
and \U$28516 ( \28831 , \28422 , \28511 );
or \U$28517 ( \28832 , \28829 , \28830 , \28831 );
xor \U$28518 ( \28833 , \28828 , \28832 );
xor \U$28519 ( \28834 , \28819 , \28833 );
xor \U$28520 ( \28835 , \28609 , \28834 );
xor \U$28521 ( \28836 , \28600 , \28835 );
and \U$28522 ( \28837 , \28571 , \28575 );
and \U$28523 ( \28838 , \28575 , \28590 );
and \U$28524 ( \28839 , \28571 , \28590 );
or \U$28525 ( \28840 , \28837 , \28838 , \28839 );
and \U$28526 ( \28841 , \28551 , \28565 );
xor \U$28527 ( \28842 , \28840 , \28841 );
and \U$28528 ( \28843 , \28580 , \28584 );
and \U$28529 ( \28844 , \28584 , \28589 );
and \U$28530 ( \28845 , \28580 , \28589 );
or \U$28531 ( \28846 , \28843 , \28844 , \28845 );
and \U$28532 ( \28847 , \28530 , \28534 );
and \U$28533 ( \28848 , \28534 , \28549 );
and \U$28534 ( \28849 , \28530 , \28549 );
or \U$28535 ( \28850 , \28847 , \28848 , \28849 );
xor \U$28536 ( \28851 , \28846 , \28850 );
and \U$28537 ( \28852 , \28411 , \28512 );
and \U$28538 ( \28853 , \28512 , \28524 );
and \U$28539 ( \28854 , \28411 , \28524 );
or \U$28540 ( \28855 , \28852 , \28853 , \28854 );
xor \U$28541 ( \28856 , \28851 , \28855 );
xor \U$28542 ( \28857 , \28842 , \28856 );
xor \U$28543 ( \28858 , \28836 , \28857 );
and \U$28544 ( \28859 , \28332 , \28592 );
nor \U$28545 ( \28860 , \28858 , \28859 );
and \U$28546 ( \28861 , \28840 , \28841 );
and \U$28547 ( \28862 , \28841 , \28856 );
and \U$28548 ( \28863 , \28840 , \28856 );
or \U$28549 ( \28864 , \28861 , \28862 , \28863 );
and \U$28550 ( \28865 , \28604 , \28608 );
and \U$28551 ( \28866 , \28608 , \28834 );
and \U$28552 ( \28867 , \28604 , \28834 );
or \U$28553 ( \28868 , \28865 , \28866 , \28867 );
and \U$28554 ( \28869 , \28823 , \28827 );
and \U$28555 ( \28870 , \28827 , \28832 );
and \U$28556 ( \28871 , \28823 , \28832 );
or \U$28557 ( \28872 , \28869 , \28870 , \28871 );
and \U$28558 ( \28873 , \28746 , \28760 );
and \U$28559 ( \28874 , \28760 , \28817 );
and \U$28560 ( \28875 , \28746 , \28817 );
or \U$28561 ( \28876 , \28873 , \28874 , \28875 );
xor \U$28562 ( \28877 , \28872 , \28876 );
and \U$28563 ( \28878 , \28712 , \28726 );
and \U$28564 ( \28879 , \28726 , \28741 );
and \U$28565 ( \28880 , \28712 , \28741 );
or \U$28566 ( \28881 , \28878 , \28879 , \28880 );
xor \U$28567 ( \28882 , \28877 , \28881 );
xor \U$28568 ( \28883 , \28868 , \28882 );
and \U$28569 ( \28884 , \28846 , \28850 );
and \U$28570 ( \28885 , \28850 , \28855 );
and \U$28571 ( \28886 , \28846 , \28855 );
or \U$28572 ( \28887 , \28884 , \28885 , \28886 );
and \U$28573 ( \28888 , \28742 , \28818 );
and \U$28574 ( \28889 , \28818 , \28833 );
and \U$28575 ( \28890 , \28742 , \28833 );
or \U$28576 ( \28891 , \28888 , \28889 , \28890 );
xor \U$28577 ( \28892 , \28887 , \28891 );
or \U$28578 ( \28893 , \28772 , \28786 );
and \U$28579 ( \28894 , \28681 , \28695 );
and \U$28580 ( \28895 , \28695 , \28710 );
and \U$28581 ( \28896 , \28681 , \28710 );
or \U$28582 ( \28897 , \28894 , \28895 , \28896 );
xor \U$28583 ( \28898 , \28893 , \28897 );
and \U$28584 ( \28899 , \28636 , \28650 );
and \U$28585 ( \28900 , \28650 , \28665 );
and \U$28586 ( \28901 , \28636 , \28665 );
or \U$28587 ( \28902 , \28899 , \28900 , \28901 );
xor \U$28588 ( \28903 , \28898 , \28902 );
and \U$28589 ( \28904 , \28750 , \28754 );
and \U$28590 ( \28905 , \28754 , \28759 );
and \U$28591 ( \28906 , \28750 , \28759 );
or \U$28592 ( \28907 , \28904 , \28905 , \28906 );
and \U$28593 ( \28908 , \28806 , \28810 );
and \U$28594 ( \28909 , \28810 , \28815 );
and \U$28595 ( \28910 , \28806 , \28815 );
or \U$28596 ( \28911 , \28908 , \28909 , \28910 );
xor \U$28597 ( \28912 , \28907 , \28911 );
and \U$28598 ( \28913 , \28791 , \28795 );
and \U$28599 ( \28914 , \28795 , \28800 );
and \U$28600 ( \28915 , \28791 , \28800 );
or \U$28601 ( \28916 , \28913 , \28914 , \28915 );
xor \U$28602 ( \28917 , \28912 , \28916 );
xor \U$28603 ( \28918 , \28903 , \28917 );
and \U$28604 ( \28919 , \28787 , \28801 );
and \U$28605 ( \28920 , \28801 , \28816 );
and \U$28606 ( \28921 , \28787 , \28816 );
or \U$28607 ( \28922 , \28919 , \28920 , \28921 );
and \U$28608 ( \28923 , \28671 , \28675 );
and \U$28609 ( \28924 , \28675 , \28680 );
and \U$28610 ( \28925 , \28671 , \28680 );
or \U$28611 ( \28926 , \28923 , \28924 , \28925 );
and \U$28612 ( \28927 , \28776 , \28780 );
and \U$28613 ( \28928 , \28780 , \28785 );
and \U$28614 ( \28929 , \28776 , \28785 );
or \U$28615 ( \28930 , \28927 , \28928 , \28929 );
xor \U$28616 ( \28931 , \28926 , \28930 );
and \U$28617 ( \28932 , \28765 , \28769 );
and \U$28618 ( \28933 , \28769 , \28771 );
and \U$28619 ( \28934 , \28765 , \28771 );
or \U$28620 ( \28935 , \28932 , \28933 , \28934 );
xor \U$28621 ( \28936 , \28931 , \28935 );
and \U$28622 ( \28937 , \28626 , \28630 );
and \U$28623 ( \28938 , \28630 , \28635 );
and \U$28624 ( \28939 , \28626 , \28635 );
or \U$28625 ( \28940 , \28937 , \28938 , \28939 );
and \U$28626 ( \28941 , \28700 , \28704 );
and \U$28627 ( \28942 , \28704 , \28709 );
and \U$28628 ( \28943 , \28700 , \28709 );
or \U$28629 ( \28944 , \28941 , \28942 , \28943 );
xor \U$28630 ( \28945 , \28940 , \28944 );
and \U$28631 ( \28946 , \28685 , \28689 );
and \U$28632 ( \28947 , \28689 , \28694 );
and \U$28633 ( \28948 , \28685 , \28694 );
or \U$28634 ( \28949 , \28946 , \28947 , \28948 );
xor \U$28635 ( \28950 , \28945 , \28949 );
xor \U$28636 ( \28951 , \28936 , \28950 );
and \U$28637 ( \28952 , \28612 , \28616 );
and \U$28638 ( \28953 , \28616 , \28621 );
and \U$28639 ( \28954 , \28612 , \28621 );
or \U$28640 ( \28955 , \28952 , \28953 , \28954 );
and \U$28641 ( \28956 , \28655 , \28659 );
and \U$28642 ( \28957 , \28659 , \28664 );
and \U$28643 ( \28958 , \28655 , \28664 );
or \U$28644 ( \28959 , \28956 , \28957 , \28958 );
xor \U$28645 ( \28960 , \28955 , \28959 );
and \U$28646 ( \28961 , \28640 , \28644 );
and \U$28647 ( \28962 , \28644 , \28649 );
and \U$28648 ( \28963 , \28640 , \28649 );
or \U$28649 ( \28964 , \28961 , \28962 , \28963 );
xor \U$28650 ( \28965 , \28960 , \28964 );
xor \U$28651 ( \28966 , \28951 , \28965 );
xor \U$28652 ( \28967 , \28922 , \28966 );
and \U$28653 ( \28968 , \22089 , \22345 );
and \U$28654 ( \28969 , \22100 , \22343 );
nor \U$28655 ( \28970 , \28968 , \28969 );
xnor \U$28656 ( \28971 , \28970 , \22355 );
and \U$28657 ( \28972 , \22113 , \22367 );
and \U$28658 ( \28973 , \22124 , \22365 );
nor \U$28659 ( \28974 , \28972 , \28973 );
xnor \U$28660 ( \28975 , \28974 , \22377 );
xor \U$28661 ( \28976 , \28971 , \28975 );
and \U$28662 ( \28977 , \22134 , \22392 );
and \U$28663 ( \28978 , \22145 , \22390 );
nor \U$28664 ( \28979 , \28977 , \28978 );
xnor \U$28665 ( \28980 , \28979 , \22402 );
xor \U$28666 ( \28981 , \28976 , \28980 );
and \U$28667 ( \28982 , \23230 , \22278 );
and \U$28668 ( \28983 , \23329 , \22276 );
nor \U$28669 ( \28984 , \28982 , \28983 );
xnor \U$28670 ( \28985 , \28984 , \22288 );
and \U$28671 ( \28986 , \22858 , \22300 );
and \U$28672 ( \28987 , \22894 , \22298 );
nor \U$28673 ( \28988 , \28986 , \28987 );
xnor \U$28674 ( \28989 , \28988 , \22310 );
xor \U$28675 ( \28990 , \28985 , \28989 );
and \U$28676 ( \28991 , \22071 , \22324 );
and \U$28677 ( \28992 , \22081 , \22322 );
nor \U$28678 ( \28993 , \28991 , \28992 );
xnor \U$28679 ( \28994 , \28993 , \22334 );
xor \U$28680 ( \28995 , \28990 , \28994 );
xor \U$28681 ( \28996 , \28981 , \28995 );
not \U$28682 ( \28997 , \22218 );
and \U$28683 ( \28998 , \21977 , \22230 );
and \U$28684 ( \28999 , \21990 , \22228 );
nor \U$28685 ( \29000 , \28998 , \28999 );
xnor \U$28686 ( \29001 , \29000 , \22240 );
xor \U$28687 ( \29002 , \28997 , \29001 );
and \U$28688 ( \29003 , \22030 , \22257 );
and \U$28689 ( \29004 , \22001 , \22255 );
nor \U$28690 ( \29005 , \29003 , \29004 );
xnor \U$28691 ( \29006 , \29005 , \22267 );
xor \U$28692 ( \29007 , \29002 , \29006 );
xor \U$28693 ( \29008 , \28996 , \29007 );
and \U$28694 ( \29009 , \22294 , \22551 );
and \U$28695 ( \29010 , \22305 , \22549 );
nor \U$28696 ( \29011 , \29009 , \29010 );
xnor \U$28697 ( \29012 , \29011 , \22561 );
and \U$28698 ( \29013 , \22318 , \22573 );
and \U$28699 ( \29014 , \22329 , \22571 );
nor \U$28700 ( \29015 , \29013 , \29014 );
xnor \U$28701 ( \29016 , \29015 , \22583 );
xor \U$28702 ( \29017 , \29012 , \29016 );
and \U$28703 ( \29018 , \22339 , \22598 );
and \U$28704 ( \29019 , \22350 , \22596 );
nor \U$28705 ( \29020 , \29018 , \29019 );
xnor \U$28706 ( \29021 , \29020 , \22608 );
xor \U$28707 ( \29022 , \29017 , \29021 );
and \U$28708 ( \29023 , \22224 , \22484 );
and \U$28709 ( \29024 , \22235 , \22482 );
nor \U$28710 ( \29025 , \29023 , \29024 );
xnor \U$28711 ( \29026 , \29025 , \22494 );
and \U$28712 ( \29027 , \22251 , \22506 );
and \U$28713 ( \29028 , \22262 , \22504 );
nor \U$28714 ( \29029 , \29027 , \29028 );
xnor \U$28715 ( \29030 , \29029 , \22516 );
xor \U$28716 ( \29031 , \29026 , \29030 );
and \U$28717 ( \29032 , \22272 , \22530 );
and \U$28718 ( \29033 , \22283 , \22528 );
nor \U$28719 ( \29034 , \29032 , \29033 );
xnor \U$28720 ( \29035 , \29034 , \22540 );
xor \U$28721 ( \29036 , \29031 , \29035 );
xor \U$28722 ( \29037 , \29022 , \29036 );
and \U$28723 ( \29038 , \22156 , \22413 );
and \U$28724 ( \29039 , \22167 , \22411 );
nor \U$28725 ( \29040 , \29038 , \29039 );
xnor \U$28726 ( \29041 , \29040 , \22423 );
and \U$28727 ( \29042 , \22181 , \22435 );
and \U$28728 ( \29043 , \22192 , \22433 );
nor \U$28729 ( \29044 , \29042 , \29043 );
xnor \U$28730 ( \29045 , \29044 , \22445 );
xor \U$28731 ( \29046 , \29041 , \29045 );
and \U$28732 ( \29047 , \22202 , \22463 );
and \U$28733 ( \29048 , \22213 , \22461 );
nor \U$28734 ( \29049 , \29047 , \29048 );
xnor \U$28735 ( \29050 , \29049 , \22473 );
xor \U$28736 ( \29051 , \29046 , \29050 );
xor \U$28737 ( \29052 , \29037 , \29051 );
xor \U$28738 ( \29053 , \29008 , \29052 );
and \U$28739 ( \29054 , \22500 , \22021 );
and \U$28740 ( \29055 , \22511 , \22019 );
nor \U$28741 ( \29056 , \29054 , \29055 );
xnor \U$28742 ( \29057 , \29056 , \21595 );
and \U$28743 ( \29058 , \22524 , \21983 );
and \U$28744 ( \29059 , \22535 , \21981 );
nor \U$28745 ( \29060 , \29058 , \29059 );
xnor \U$28746 ( \29061 , \29060 , \21995 );
xor \U$28747 ( \29062 , \29057 , \29061 );
and \U$28748 ( \29063 , \22556 , \21978 );
xor \U$28749 ( \29064 , \29062 , \29063 );
and \U$28750 ( \29065 , \22429 , \22691 );
and \U$28751 ( \29066 , \22440 , \22689 );
nor \U$28752 ( \29067 , \29065 , \29066 );
xnor \U$28753 ( \29068 , \29067 , \22701 );
and \U$28754 ( \29069 , \22457 , \22720 );
and \U$28755 ( \29070 , \22468 , \22707 );
nor \U$28756 ( \29071 , \29069 , \29070 );
xnor \U$28757 ( \29072 , \29071 , \22067 );
xor \U$28758 ( \29073 , \29068 , \29072 );
and \U$28759 ( \29074 , \22478 , \23173 );
and \U$28760 ( \29075 , \22489 , \22999 );
nor \U$28761 ( \29076 , \29074 , \29075 );
xnor \U$28762 ( \29077 , \29076 , \22016 );
xor \U$28763 ( \29078 , \29073 , \29077 );
xor \U$28764 ( \29079 , \29064 , \29078 );
and \U$28765 ( \29080 , \22361 , \22619 );
and \U$28766 ( \29081 , \22372 , \22617 );
nor \U$28767 ( \29082 , \29080 , \29081 );
xnor \U$28768 ( \29083 , \29082 , \22629 );
and \U$28769 ( \29084 , \22386 , \22641 );
and \U$28770 ( \29085 , \22397 , \22639 );
nor \U$28771 ( \29086 , \29084 , \29085 );
xnor \U$28772 ( \29087 , \29086 , \22651 );
xor \U$28773 ( \29088 , \29083 , \29087 );
and \U$28774 ( \29089 , \22407 , \22671 );
and \U$28775 ( \29090 , \22418 , \22669 );
nor \U$28776 ( \29091 , \29089 , \29090 );
xnor \U$28777 ( \29092 , \29091 , \22681 );
xor \U$28778 ( \29093 , \29088 , \29092 );
xor \U$28779 ( \29094 , \29079 , \29093 );
xor \U$28780 ( \29095 , \29053 , \29094 );
xor \U$28781 ( \29096 , \28967 , \29095 );
xor \U$28782 ( \29097 , \28918 , \29096 );
and \U$28783 ( \29098 , \28731 , \28735 );
and \U$28784 ( \29099 , \28735 , \28740 );
and \U$28785 ( \29100 , \28731 , \28740 );
or \U$28786 ( \29101 , \29098 , \29099 , \29100 );
and \U$28787 ( \29102 , \28716 , \28720 );
and \U$28788 ( \29103 , \28720 , \28725 );
and \U$28789 ( \29104 , \28716 , \28725 );
or \U$28790 ( \29105 , \29102 , \29103 , \29104 );
xor \U$28791 ( \29106 , \29101 , \29105 );
and \U$28792 ( \29107 , \28622 , \28666 );
and \U$28793 ( \29108 , \28666 , \28711 );
and \U$28794 ( \29109 , \28622 , \28711 );
or \U$28795 ( \29110 , \29107 , \29108 , \29109 );
xor \U$28796 ( \29111 , \29106 , \29110 );
xor \U$28797 ( \29112 , \29097 , \29111 );
xor \U$28798 ( \29113 , \28892 , \29112 );
xor \U$28799 ( \29114 , \28883 , \29113 );
xor \U$28800 ( \29115 , \28864 , \29114 );
and \U$28801 ( \29116 , \28600 , \28835 );
and \U$28802 ( \29117 , \28835 , \28857 );
and \U$28803 ( \29118 , \28600 , \28857 );
or \U$28804 ( \29119 , \29116 , \29117 , \29118 );
nor \U$28805 ( \29120 , \29115 , \29119 );
nor \U$28806 ( \29121 , \28860 , \29120 );
nand \U$28807 ( \29122 , \28596 , \29121 );
nor \U$28808 ( \29123 , \28053 , \29122 );
nand \U$28809 ( \29124 , \26901 , \29123 );
and \U$28810 ( \29125 , \28868 , \28882 );
and \U$28811 ( \29126 , \28882 , \29113 );
and \U$28812 ( \29127 , \28868 , \29113 );
or \U$28813 ( \29128 , \29125 , \29126 , \29127 );
and \U$28814 ( \29129 , \28887 , \28891 );
and \U$28815 ( \29130 , \28891 , \29112 );
and \U$28816 ( \29131 , \28887 , \29112 );
or \U$28817 ( \29132 , \29129 , \29130 , \29131 );
and \U$28818 ( \29133 , \29101 , \29105 );
and \U$28819 ( \29134 , \29105 , \29110 );
and \U$28820 ( \29135 , \29101 , \29110 );
or \U$28821 ( \29136 , \29133 , \29134 , \29135 );
and \U$28822 ( \29137 , \28922 , \28966 );
and \U$28823 ( \29138 , \28966 , \29095 );
and \U$28824 ( \29139 , \28922 , \29095 );
or \U$28825 ( \29140 , \29137 , \29138 , \29139 );
xor \U$28826 ( \29141 , \29136 , \29140 );
and \U$28827 ( \29142 , \28903 , \28917 );
xor \U$28828 ( \29143 , \29141 , \29142 );
xor \U$28829 ( \29144 , \29132 , \29143 );
and \U$28830 ( \29145 , \28872 , \28876 );
and \U$28831 ( \29146 , \28876 , \28881 );
and \U$28832 ( \29147 , \28872 , \28881 );
or \U$28833 ( \29148 , \29145 , \29146 , \29147 );
and \U$28834 ( \29149 , \28918 , \29096 );
and \U$28835 ( \29150 , \29096 , \29111 );
and \U$28836 ( \29151 , \28918 , \29111 );
or \U$28837 ( \29152 , \29149 , \29150 , \29151 );
xor \U$28838 ( \29153 , \29148 , \29152 );
and \U$28839 ( \29154 , \29064 , \29078 );
and \U$28840 ( \29155 , \29078 , \29093 );
and \U$28841 ( \29156 , \29064 , \29093 );
or \U$28842 ( \29157 , \29154 , \29155 , \29156 );
and \U$28843 ( \29158 , \29022 , \29036 );
and \U$28844 ( \29159 , \29036 , \29051 );
and \U$28845 ( \29160 , \29022 , \29051 );
or \U$28846 ( \29161 , \29158 , \29159 , \29160 );
xor \U$28847 ( \29162 , \29157 , \29161 );
and \U$28848 ( \29163 , \28981 , \28995 );
and \U$28849 ( \29164 , \28995 , \29007 );
and \U$28850 ( \29165 , \28981 , \29007 );
or \U$28851 ( \29166 , \29163 , \29164 , \29165 );
xor \U$28852 ( \29167 , \29162 , \29166 );
and \U$28853 ( \29168 , \28955 , \28959 );
and \U$28854 ( \29169 , \28959 , \28964 );
and \U$28855 ( \29170 , \28955 , \28964 );
or \U$28856 ( \29171 , \29168 , \29169 , \29170 );
and \U$28857 ( \29172 , \28940 , \28944 );
and \U$28858 ( \29173 , \28944 , \28949 );
and \U$28859 ( \29174 , \28940 , \28949 );
or \U$28860 ( \29175 , \29172 , \29173 , \29174 );
xor \U$28861 ( \29176 , \29171 , \29175 );
and \U$28862 ( \29177 , \28926 , \28930 );
and \U$28863 ( \29178 , \28930 , \28935 );
and \U$28864 ( \29179 , \28926 , \28935 );
or \U$28865 ( \29180 , \29177 , \29178 , \29179 );
xor \U$28866 ( \29181 , \29176 , \29180 );
xor \U$28867 ( \29182 , \29167 , \29181 );
and \U$28868 ( \29183 , \28936 , \28950 );
and \U$28869 ( \29184 , \28950 , \28965 );
and \U$28870 ( \29185 , \28936 , \28965 );
or \U$28871 ( \29186 , \29183 , \29184 , \29185 );
and \U$28872 ( \29187 , \29083 , \29087 );
and \U$28873 ( \29188 , \29087 , \29092 );
and \U$28874 ( \29189 , \29083 , \29092 );
or \U$28875 ( \29190 , \29187 , \29188 , \29189 );
and \U$28876 ( \29191 , \29068 , \29072 );
and \U$28877 ( \29192 , \29072 , \29077 );
and \U$28878 ( \29193 , \29068 , \29077 );
or \U$28879 ( \29194 , \29191 , \29192 , \29193 );
xor \U$28880 ( \29195 , \29190 , \29194 );
and \U$28881 ( \29196 , \29057 , \29061 );
and \U$28882 ( \29197 , \29061 , \29063 );
and \U$28883 ( \29198 , \29057 , \29063 );
or \U$28884 ( \29199 , \29196 , \29197 , \29198 );
xor \U$28885 ( \29200 , \29195 , \29199 );
and \U$28886 ( \29201 , \29041 , \29045 );
and \U$28887 ( \29202 , \29045 , \29050 );
and \U$28888 ( \29203 , \29041 , \29050 );
or \U$28889 ( \29204 , \29201 , \29202 , \29203 );
and \U$28890 ( \29205 , \29026 , \29030 );
and \U$28891 ( \29206 , \29030 , \29035 );
and \U$28892 ( \29207 , \29026 , \29035 );
or \U$28893 ( \29208 , \29205 , \29206 , \29207 );
xor \U$28894 ( \29209 , \29204 , \29208 );
and \U$28895 ( \29210 , \29012 , \29016 );
and \U$28896 ( \29211 , \29016 , \29021 );
and \U$28897 ( \29212 , \29012 , \29021 );
or \U$28898 ( \29213 , \29210 , \29211 , \29212 );
xor \U$28899 ( \29214 , \29209 , \29213 );
xor \U$28900 ( \29215 , \29200 , \29214 );
and \U$28901 ( \29216 , \28997 , \29001 );
and \U$28902 ( \29217 , \29001 , \29006 );
and \U$28903 ( \29218 , \28997 , \29006 );
or \U$28904 ( \29219 , \29216 , \29217 , \29218 );
and \U$28905 ( \29220 , \28985 , \28989 );
and \U$28906 ( \29221 , \28989 , \28994 );
and \U$28907 ( \29222 , \28985 , \28994 );
or \U$28908 ( \29223 , \29220 , \29221 , \29222 );
xor \U$28909 ( \29224 , \29219 , \29223 );
and \U$28910 ( \29225 , \28971 , \28975 );
and \U$28911 ( \29226 , \28975 , \28980 );
and \U$28912 ( \29227 , \28971 , \28980 );
or \U$28913 ( \29228 , \29225 , \29226 , \29227 );
xor \U$28914 ( \29229 , \29224 , \29228 );
xor \U$28915 ( \29230 , \29215 , \29229 );
xor \U$28916 ( \29231 , \29186 , \29230 );
and \U$28917 ( \29232 , \22124 , \22367 );
and \U$28918 ( \29233 , \22089 , \22365 );
nor \U$28919 ( \29234 , \29232 , \29233 );
xnor \U$28920 ( \29235 , \29234 , \22377 );
and \U$28921 ( \29236 , \22145 , \22392 );
and \U$28922 ( \29237 , \22113 , \22390 );
nor \U$28923 ( \29238 , \29236 , \29237 );
xnor \U$28924 ( \29239 , \29238 , \22402 );
xor \U$28925 ( \29240 , \29235 , \29239 );
and \U$28926 ( \29241 , \22167 , \22413 );
and \U$28927 ( \29242 , \22134 , \22411 );
nor \U$28928 ( \29243 , \29241 , \29242 );
xnor \U$28929 ( \29244 , \29243 , \22423 );
xor \U$28930 ( \29245 , \29240 , \29244 );
and \U$28931 ( \29246 , \22894 , \22300 );
and \U$28932 ( \29247 , \23230 , \22298 );
nor \U$28933 ( \29248 , \29246 , \29247 );
xnor \U$28934 ( \29249 , \29248 , \22310 );
and \U$28935 ( \29250 , \22081 , \22324 );
and \U$28936 ( \29251 , \22858 , \22322 );
nor \U$28937 ( \29252 , \29250 , \29251 );
xnor \U$28938 ( \29253 , \29252 , \22334 );
xor \U$28939 ( \29254 , \29249 , \29253 );
and \U$28940 ( \29255 , \22100 , \22345 );
and \U$28941 ( \29256 , \22071 , \22343 );
nor \U$28942 ( \29257 , \29255 , \29256 );
xnor \U$28943 ( \29258 , \29257 , \22355 );
xor \U$28944 ( \29259 , \29254 , \29258 );
xor \U$28945 ( \29260 , \29245 , \29259 );
and \U$28946 ( \29261 , \21990 , \22230 );
not \U$28947 ( \29262 , \29261 );
xnor \U$28948 ( \29263 , \29262 , \22240 );
and \U$28949 ( \29264 , \22001 , \22257 );
and \U$28950 ( \29265 , \21977 , \22255 );
nor \U$28951 ( \29266 , \29264 , \29265 );
xnor \U$28952 ( \29267 , \29266 , \22267 );
xor \U$28953 ( \29268 , \29263 , \29267 );
and \U$28954 ( \29269 , \23329 , \22278 );
and \U$28955 ( \29270 , \22030 , \22276 );
nor \U$28956 ( \29271 , \29269 , \29270 );
xnor \U$28957 ( \29272 , \29271 , \22288 );
xor \U$28958 ( \29273 , \29268 , \29272 );
xor \U$28959 ( \29274 , \29260 , \29273 );
and \U$28960 ( \29275 , \22329 , \22573 );
and \U$28961 ( \29276 , \22294 , \22571 );
nor \U$28962 ( \29277 , \29275 , \29276 );
xnor \U$28963 ( \29278 , \29277 , \22583 );
and \U$28964 ( \29279 , \22350 , \22598 );
and \U$28965 ( \29280 , \22318 , \22596 );
nor \U$28966 ( \29281 , \29279 , \29280 );
xnor \U$28967 ( \29282 , \29281 , \22608 );
xor \U$28968 ( \29283 , \29278 , \29282 );
and \U$28969 ( \29284 , \22372 , \22619 );
and \U$28970 ( \29285 , \22339 , \22617 );
nor \U$28971 ( \29286 , \29284 , \29285 );
xnor \U$28972 ( \29287 , \29286 , \22629 );
xor \U$28973 ( \29288 , \29283 , \29287 );
and \U$28974 ( \29289 , \22262 , \22506 );
and \U$28975 ( \29290 , \22224 , \22504 );
nor \U$28976 ( \29291 , \29289 , \29290 );
xnor \U$28977 ( \29292 , \29291 , \22516 );
and \U$28978 ( \29293 , \22283 , \22530 );
and \U$28979 ( \29294 , \22251 , \22528 );
nor \U$28980 ( \29295 , \29293 , \29294 );
xnor \U$28981 ( \29296 , \29295 , \22540 );
xor \U$28982 ( \29297 , \29292 , \29296 );
and \U$28983 ( \29298 , \22305 , \22551 );
and \U$28984 ( \29299 , \22272 , \22549 );
nor \U$28985 ( \29300 , \29298 , \29299 );
xnor \U$28986 ( \29301 , \29300 , \22561 );
xor \U$28987 ( \29302 , \29297 , \29301 );
xor \U$28988 ( \29303 , \29288 , \29302 );
and \U$28989 ( \29304 , \22192 , \22435 );
and \U$28990 ( \29305 , \22156 , \22433 );
nor \U$28991 ( \29306 , \29304 , \29305 );
xnor \U$28992 ( \29307 , \29306 , \22445 );
and \U$28993 ( \29308 , \22213 , \22463 );
and \U$28994 ( \29309 , \22181 , \22461 );
nor \U$28995 ( \29310 , \29308 , \29309 );
xnor \U$28996 ( \29311 , \29310 , \22473 );
xor \U$28997 ( \29312 , \29307 , \29311 );
and \U$28998 ( \29313 , \22235 , \22484 );
and \U$28999 ( \29314 , \22202 , \22482 );
nor \U$29000 ( \29315 , \29313 , \29314 );
xnor \U$29001 ( \29316 , \29315 , \22494 );
xor \U$29002 ( \29317 , \29312 , \29316 );
xor \U$29003 ( \29318 , \29303 , \29317 );
xor \U$29004 ( \29319 , \29274 , \29318 );
and \U$29005 ( \29320 , \22535 , \21983 );
and \U$29006 ( \29321 , \22500 , \21981 );
nor \U$29007 ( \29322 , \29320 , \29321 );
xnor \U$29008 ( \29323 , \29322 , \21995 );
and \U$29009 ( \29324 , \22524 , \21978 );
xnor \U$29010 ( \29325 , \29323 , \29324 );
and \U$29011 ( \29326 , \22468 , \22720 );
and \U$29012 ( \29327 , \22429 , \22707 );
nor \U$29013 ( \29328 , \29326 , \29327 );
xnor \U$29014 ( \29329 , \29328 , \22067 );
and \U$29015 ( \29330 , \22489 , \23173 );
and \U$29016 ( \29331 , \22457 , \22999 );
nor \U$29017 ( \29332 , \29330 , \29331 );
xnor \U$29018 ( \29333 , \29332 , \22016 );
xor \U$29019 ( \29334 , \29329 , \29333 );
and \U$29020 ( \29335 , \22511 , \22021 );
and \U$29021 ( \29336 , \22478 , \22019 );
nor \U$29022 ( \29337 , \29335 , \29336 );
xnor \U$29023 ( \29338 , \29337 , \21595 );
xor \U$29024 ( \29339 , \29334 , \29338 );
xor \U$29025 ( \29340 , \29325 , \29339 );
and \U$29026 ( \29341 , \22397 , \22641 );
and \U$29027 ( \29342 , \22361 , \22639 );
nor \U$29028 ( \29343 , \29341 , \29342 );
xnor \U$29029 ( \29344 , \29343 , \22651 );
and \U$29030 ( \29345 , \22418 , \22671 );
and \U$29031 ( \29346 , \22386 , \22669 );
nor \U$29032 ( \29347 , \29345 , \29346 );
xnor \U$29033 ( \29348 , \29347 , \22681 );
xor \U$29034 ( \29349 , \29344 , \29348 );
and \U$29035 ( \29350 , \22440 , \22691 );
and \U$29036 ( \29351 , \22407 , \22689 );
nor \U$29037 ( \29352 , \29350 , \29351 );
xnor \U$29038 ( \29353 , \29352 , \22701 );
xor \U$29039 ( \29354 , \29349 , \29353 );
xor \U$29040 ( \29355 , \29340 , \29354 );
xor \U$29041 ( \29356 , \29319 , \29355 );
xor \U$29042 ( \29357 , \29231 , \29356 );
xor \U$29043 ( \29358 , \29182 , \29357 );
and \U$29044 ( \29359 , \28907 , \28911 );
and \U$29045 ( \29360 , \28911 , \28916 );
and \U$29046 ( \29361 , \28907 , \28916 );
or \U$29047 ( \29362 , \29359 , \29360 , \29361 );
and \U$29048 ( \29363 , \28893 , \28897 );
and \U$29049 ( \29364 , \28897 , \28902 );
and \U$29050 ( \29365 , \28893 , \28902 );
or \U$29051 ( \29366 , \29363 , \29364 , \29365 );
xor \U$29052 ( \29367 , \29362 , \29366 );
and \U$29053 ( \29368 , \29008 , \29052 );
and \U$29054 ( \29369 , \29052 , \29094 );
and \U$29055 ( \29370 , \29008 , \29094 );
or \U$29056 ( \29371 , \29368 , \29369 , \29370 );
xor \U$29057 ( \29372 , \29367 , \29371 );
xor \U$29058 ( \29373 , \29358 , \29372 );
xor \U$29059 ( \29374 , \29153 , \29373 );
xor \U$29060 ( \29375 , \29144 , \29374 );
xor \U$29061 ( \29376 , \29128 , \29375 );
and \U$29062 ( \29377 , \28864 , \29114 );
nor \U$29063 ( \29378 , \29376 , \29377 );
and \U$29064 ( \29379 , \29132 , \29143 );
and \U$29065 ( \29380 , \29143 , \29374 );
and \U$29066 ( \29381 , \29132 , \29374 );
or \U$29067 ( \29382 , \29379 , \29380 , \29381 );
and \U$29068 ( \29383 , \29148 , \29152 );
and \U$29069 ( \29384 , \29152 , \29373 );
and \U$29070 ( \29385 , \29148 , \29373 );
or \U$29071 ( \29386 , \29383 , \29384 , \29385 );
and \U$29072 ( \29387 , \29362 , \29366 );
and \U$29073 ( \29388 , \29366 , \29371 );
and \U$29074 ( \29389 , \29362 , \29371 );
or \U$29075 ( \29390 , \29387 , \29388 , \29389 );
and \U$29076 ( \29391 , \29186 , \29230 );
and \U$29077 ( \29392 , \29230 , \29356 );
and \U$29078 ( \29393 , \29186 , \29356 );
or \U$29079 ( \29394 , \29391 , \29392 , \29393 );
xor \U$29080 ( \29395 , \29390 , \29394 );
and \U$29081 ( \29396 , \29167 , \29181 );
xor \U$29082 ( \29397 , \29395 , \29396 );
xor \U$29083 ( \29398 , \29386 , \29397 );
and \U$29084 ( \29399 , \29136 , \29140 );
and \U$29085 ( \29400 , \29140 , \29142 );
and \U$29086 ( \29401 , \29136 , \29142 );
or \U$29087 ( \29402 , \29399 , \29400 , \29401 );
and \U$29088 ( \29403 , \29182 , \29357 );
and \U$29089 ( \29404 , \29357 , \29372 );
and \U$29090 ( \29405 , \29182 , \29372 );
or \U$29091 ( \29406 , \29403 , \29404 , \29405 );
xor \U$29092 ( \29407 , \29402 , \29406 );
and \U$29093 ( \29408 , \29325 , \29339 );
and \U$29094 ( \29409 , \29339 , \29354 );
and \U$29095 ( \29410 , \29325 , \29354 );
or \U$29096 ( \29411 , \29408 , \29409 , \29410 );
and \U$29097 ( \29412 , \29288 , \29302 );
and \U$29098 ( \29413 , \29302 , \29317 );
and \U$29099 ( \29414 , \29288 , \29317 );
or \U$29100 ( \29415 , \29412 , \29413 , \29414 );
xor \U$29101 ( \29416 , \29411 , \29415 );
and \U$29102 ( \29417 , \29245 , \29259 );
and \U$29103 ( \29418 , \29259 , \29273 );
and \U$29104 ( \29419 , \29245 , \29273 );
or \U$29105 ( \29420 , \29417 , \29418 , \29419 );
xor \U$29106 ( \29421 , \29416 , \29420 );
and \U$29107 ( \29422 , \29219 , \29223 );
and \U$29108 ( \29423 , \29223 , \29228 );
and \U$29109 ( \29424 , \29219 , \29228 );
or \U$29110 ( \29425 , \29422 , \29423 , \29424 );
and \U$29111 ( \29426 , \29204 , \29208 );
and \U$29112 ( \29427 , \29208 , \29213 );
and \U$29113 ( \29428 , \29204 , \29213 );
or \U$29114 ( \29429 , \29426 , \29427 , \29428 );
xor \U$29115 ( \29430 , \29425 , \29429 );
and \U$29116 ( \29431 , \29190 , \29194 );
and \U$29117 ( \29432 , \29194 , \29199 );
and \U$29118 ( \29433 , \29190 , \29199 );
or \U$29119 ( \29434 , \29431 , \29432 , \29433 );
xor \U$29120 ( \29435 , \29430 , \29434 );
xor \U$29121 ( \29436 , \29421 , \29435 );
and \U$29122 ( \29437 , \29200 , \29214 );
and \U$29123 ( \29438 , \29214 , \29229 );
and \U$29124 ( \29439 , \29200 , \29229 );
or \U$29125 ( \29440 , \29437 , \29438 , \29439 );
and \U$29126 ( \29441 , \29344 , \29348 );
and \U$29127 ( \29442 , \29348 , \29353 );
and \U$29128 ( \29443 , \29344 , \29353 );
or \U$29129 ( \29444 , \29441 , \29442 , \29443 );
and \U$29130 ( \29445 , \29329 , \29333 );
and \U$29131 ( \29446 , \29333 , \29338 );
and \U$29132 ( \29447 , \29329 , \29338 );
or \U$29133 ( \29448 , \29445 , \29446 , \29447 );
xor \U$29134 ( \29449 , \29444 , \29448 );
or \U$29135 ( \29450 , \29323 , \29324 );
xor \U$29136 ( \29451 , \29449 , \29450 );
and \U$29137 ( \29452 , \29307 , \29311 );
and \U$29138 ( \29453 , \29311 , \29316 );
and \U$29139 ( \29454 , \29307 , \29316 );
or \U$29140 ( \29455 , \29452 , \29453 , \29454 );
and \U$29141 ( \29456 , \29292 , \29296 );
and \U$29142 ( \29457 , \29296 , \29301 );
and \U$29143 ( \29458 , \29292 , \29301 );
or \U$29144 ( \29459 , \29456 , \29457 , \29458 );
xor \U$29145 ( \29460 , \29455 , \29459 );
and \U$29146 ( \29461 , \29278 , \29282 );
and \U$29147 ( \29462 , \29282 , \29287 );
and \U$29148 ( \29463 , \29278 , \29287 );
or \U$29149 ( \29464 , \29461 , \29462 , \29463 );
xor \U$29150 ( \29465 , \29460 , \29464 );
xor \U$29151 ( \29466 , \29451 , \29465 );
and \U$29152 ( \29467 , \29263 , \29267 );
and \U$29153 ( \29468 , \29267 , \29272 );
and \U$29154 ( \29469 , \29263 , \29272 );
or \U$29155 ( \29470 , \29467 , \29468 , \29469 );
and \U$29156 ( \29471 , \29249 , \29253 );
and \U$29157 ( \29472 , \29253 , \29258 );
and \U$29158 ( \29473 , \29249 , \29258 );
or \U$29159 ( \29474 , \29471 , \29472 , \29473 );
xor \U$29160 ( \29475 , \29470 , \29474 );
and \U$29161 ( \29476 , \29235 , \29239 );
and \U$29162 ( \29477 , \29239 , \29244 );
and \U$29163 ( \29478 , \29235 , \29244 );
or \U$29164 ( \29479 , \29476 , \29477 , \29478 );
xor \U$29165 ( \29480 , \29475 , \29479 );
xor \U$29166 ( \29481 , \29466 , \29480 );
xor \U$29167 ( \29482 , \29440 , \29481 );
and \U$29168 ( \29483 , \22089 , \22367 );
and \U$29169 ( \29484 , \22100 , \22365 );
nor \U$29170 ( \29485 , \29483 , \29484 );
xnor \U$29171 ( \29486 , \29485 , \22377 );
and \U$29172 ( \29487 , \22113 , \22392 );
and \U$29173 ( \29488 , \22124 , \22390 );
nor \U$29174 ( \29489 , \29487 , \29488 );
xnor \U$29175 ( \29490 , \29489 , \22402 );
xor \U$29176 ( \29491 , \29486 , \29490 );
and \U$29177 ( \29492 , \22134 , \22413 );
and \U$29178 ( \29493 , \22145 , \22411 );
nor \U$29179 ( \29494 , \29492 , \29493 );
xnor \U$29180 ( \29495 , \29494 , \22423 );
xor \U$29181 ( \29496 , \29491 , \29495 );
and \U$29182 ( \29497 , \23230 , \22300 );
and \U$29183 ( \29498 , \23329 , \22298 );
nor \U$29184 ( \29499 , \29497 , \29498 );
xnor \U$29185 ( \29500 , \29499 , \22310 );
and \U$29186 ( \29501 , \22858 , \22324 );
and \U$29187 ( \29502 , \22894 , \22322 );
nor \U$29188 ( \29503 , \29501 , \29502 );
xnor \U$29189 ( \29504 , \29503 , \22334 );
xor \U$29190 ( \29505 , \29500 , \29504 );
and \U$29191 ( \29506 , \22071 , \22345 );
and \U$29192 ( \29507 , \22081 , \22343 );
nor \U$29193 ( \29508 , \29506 , \29507 );
xnor \U$29194 ( \29509 , \29508 , \22355 );
xor \U$29195 ( \29510 , \29505 , \29509 );
xor \U$29196 ( \29511 , \29496 , \29510 );
not \U$29197 ( \29512 , \22240 );
and \U$29198 ( \29513 , \21977 , \22257 );
and \U$29199 ( \29514 , \21990 , \22255 );
nor \U$29200 ( \29515 , \29513 , \29514 );
xnor \U$29201 ( \29516 , \29515 , \22267 );
xor \U$29202 ( \29517 , \29512 , \29516 );
and \U$29203 ( \29518 , \22030 , \22278 );
and \U$29204 ( \29519 , \22001 , \22276 );
nor \U$29205 ( \29520 , \29518 , \29519 );
xnor \U$29206 ( \29521 , \29520 , \22288 );
xor \U$29207 ( \29522 , \29517 , \29521 );
xor \U$29208 ( \29523 , \29511 , \29522 );
and \U$29209 ( \29524 , \22294 , \22573 );
and \U$29210 ( \29525 , \22305 , \22571 );
nor \U$29211 ( \29526 , \29524 , \29525 );
xnor \U$29212 ( \29527 , \29526 , \22583 );
and \U$29213 ( \29528 , \22318 , \22598 );
and \U$29214 ( \29529 , \22329 , \22596 );
nor \U$29215 ( \29530 , \29528 , \29529 );
xnor \U$29216 ( \29531 , \29530 , \22608 );
xor \U$29217 ( \29532 , \29527 , \29531 );
and \U$29218 ( \29533 , \22339 , \22619 );
and \U$29219 ( \29534 , \22350 , \22617 );
nor \U$29220 ( \29535 , \29533 , \29534 );
xnor \U$29221 ( \29536 , \29535 , \22629 );
xor \U$29222 ( \29537 , \29532 , \29536 );
and \U$29223 ( \29538 , \22224 , \22506 );
and \U$29224 ( \29539 , \22235 , \22504 );
nor \U$29225 ( \29540 , \29538 , \29539 );
xnor \U$29226 ( \29541 , \29540 , \22516 );
and \U$29227 ( \29542 , \22251 , \22530 );
and \U$29228 ( \29543 , \22262 , \22528 );
nor \U$29229 ( \29544 , \29542 , \29543 );
xnor \U$29230 ( \29545 , \29544 , \22540 );
xor \U$29231 ( \29546 , \29541 , \29545 );
and \U$29232 ( \29547 , \22272 , \22551 );
and \U$29233 ( \29548 , \22283 , \22549 );
nor \U$29234 ( \29549 , \29547 , \29548 );
xnor \U$29235 ( \29550 , \29549 , \22561 );
xor \U$29236 ( \29551 , \29546 , \29550 );
xor \U$29237 ( \29552 , \29537 , \29551 );
and \U$29238 ( \29553 , \22156 , \22435 );
and \U$29239 ( \29554 , \22167 , \22433 );
nor \U$29240 ( \29555 , \29553 , \29554 );
xnor \U$29241 ( \29556 , \29555 , \22445 );
and \U$29242 ( \29557 , \22181 , \22463 );
and \U$29243 ( \29558 , \22192 , \22461 );
nor \U$29244 ( \29559 , \29557 , \29558 );
xnor \U$29245 ( \29560 , \29559 , \22473 );
xor \U$29246 ( \29561 , \29556 , \29560 );
and \U$29247 ( \29562 , \22202 , \22484 );
and \U$29248 ( \29563 , \22213 , \22482 );
nor \U$29249 ( \29564 , \29562 , \29563 );
xnor \U$29250 ( \29565 , \29564 , \22494 );
xor \U$29251 ( \29566 , \29561 , \29565 );
xor \U$29252 ( \29567 , \29552 , \29566 );
xor \U$29253 ( \29568 , \29523 , \29567 );
and \U$29254 ( \29569 , \22500 , \21983 );
and \U$29255 ( \29570 , \22511 , \21981 );
nor \U$29256 ( \29571 , \29569 , \29570 );
xnor \U$29257 ( \29572 , \29571 , \21995 );
and \U$29258 ( \29573 , \22535 , \21978 );
xor \U$29259 ( \29574 , \29572 , \29573 );
and \U$29260 ( \29575 , \22429 , \22720 );
and \U$29261 ( \29576 , \22440 , \22707 );
nor \U$29262 ( \29577 , \29575 , \29576 );
xnor \U$29263 ( \29578 , \29577 , \22067 );
and \U$29264 ( \29579 , \22457 , \23173 );
and \U$29265 ( \29580 , \22468 , \22999 );
nor \U$29266 ( \29581 , \29579 , \29580 );
xnor \U$29267 ( \29582 , \29581 , \22016 );
xor \U$29268 ( \29583 , \29578 , \29582 );
and \U$29269 ( \29584 , \22478 , \22021 );
and \U$29270 ( \29585 , \22489 , \22019 );
nor \U$29271 ( \29586 , \29584 , \29585 );
xnor \U$29272 ( \29587 , \29586 , \21595 );
xor \U$29273 ( \29588 , \29583 , \29587 );
xor \U$29274 ( \29589 , \29574 , \29588 );
and \U$29275 ( \29590 , \22361 , \22641 );
and \U$29276 ( \29591 , \22372 , \22639 );
nor \U$29277 ( \29592 , \29590 , \29591 );
xnor \U$29278 ( \29593 , \29592 , \22651 );
and \U$29279 ( \29594 , \22386 , \22671 );
and \U$29280 ( \29595 , \22397 , \22669 );
nor \U$29281 ( \29596 , \29594 , \29595 );
xnor \U$29282 ( \29597 , \29596 , \22681 );
xor \U$29283 ( \29598 , \29593 , \29597 );
and \U$29284 ( \29599 , \22407 , \22691 );
and \U$29285 ( \29600 , \22418 , \22689 );
nor \U$29286 ( \29601 , \29599 , \29600 );
xnor \U$29287 ( \29602 , \29601 , \22701 );
xor \U$29288 ( \29603 , \29598 , \29602 );
xor \U$29289 ( \29604 , \29589 , \29603 );
xor \U$29290 ( \29605 , \29568 , \29604 );
xor \U$29291 ( \29606 , \29482 , \29605 );
xor \U$29292 ( \29607 , \29436 , \29606 );
and \U$29293 ( \29608 , \29171 , \29175 );
and \U$29294 ( \29609 , \29175 , \29180 );
and \U$29295 ( \29610 , \29171 , \29180 );
or \U$29296 ( \29611 , \29608 , \29609 , \29610 );
and \U$29297 ( \29612 , \29157 , \29161 );
and \U$29298 ( \29613 , \29161 , \29166 );
and \U$29299 ( \29614 , \29157 , \29166 );
or \U$29300 ( \29615 , \29612 , \29613 , \29614 );
xor \U$29301 ( \29616 , \29611 , \29615 );
and \U$29302 ( \29617 , \29274 , \29318 );
and \U$29303 ( \29618 , \29318 , \29355 );
and \U$29304 ( \29619 , \29274 , \29355 );
or \U$29305 ( \29620 , \29617 , \29618 , \29619 );
xor \U$29306 ( \29621 , \29616 , \29620 );
xor \U$29307 ( \29622 , \29607 , \29621 );
xor \U$29308 ( \29623 , \29407 , \29622 );
xor \U$29309 ( \29624 , \29398 , \29623 );
xor \U$29310 ( \29625 , \29382 , \29624 );
and \U$29311 ( \29626 , \29128 , \29375 );
nor \U$29312 ( \29627 , \29625 , \29626 );
nor \U$29313 ( \29628 , \29378 , \29627 );
and \U$29314 ( \29629 , \29386 , \29397 );
and \U$29315 ( \29630 , \29397 , \29623 );
and \U$29316 ( \29631 , \29386 , \29623 );
or \U$29317 ( \29632 , \29629 , \29630 , \29631 );
and \U$29318 ( \29633 , \29402 , \29406 );
and \U$29319 ( \29634 , \29406 , \29622 );
and \U$29320 ( \29635 , \29402 , \29622 );
or \U$29321 ( \29636 , \29633 , \29634 , \29635 );
and \U$29322 ( \29637 , \29611 , \29615 );
and \U$29323 ( \29638 , \29615 , \29620 );
and \U$29324 ( \29639 , \29611 , \29620 );
or \U$29325 ( \29640 , \29637 , \29638 , \29639 );
and \U$29326 ( \29641 , \29440 , \29481 );
and \U$29327 ( \29642 , \29481 , \29605 );
and \U$29328 ( \29643 , \29440 , \29605 );
or \U$29329 ( \29644 , \29641 , \29642 , \29643 );
xor \U$29330 ( \29645 , \29640 , \29644 );
and \U$29331 ( \29646 , \29421 , \29435 );
xor \U$29332 ( \29647 , \29645 , \29646 );
xor \U$29333 ( \29648 , \29636 , \29647 );
and \U$29334 ( \29649 , \29390 , \29394 );
and \U$29335 ( \29650 , \29394 , \29396 );
and \U$29336 ( \29651 , \29390 , \29396 );
or \U$29337 ( \29652 , \29649 , \29650 , \29651 );
and \U$29338 ( \29653 , \29436 , \29606 );
and \U$29339 ( \29654 , \29606 , \29621 );
and \U$29340 ( \29655 , \29436 , \29621 );
or \U$29341 ( \29656 , \29653 , \29654 , \29655 );
xor \U$29342 ( \29657 , \29652 , \29656 );
and \U$29343 ( \29658 , \29574 , \29588 );
and \U$29344 ( \29659 , \29588 , \29603 );
and \U$29345 ( \29660 , \29574 , \29603 );
or \U$29346 ( \29661 , \29658 , \29659 , \29660 );
and \U$29347 ( \29662 , \29537 , \29551 );
and \U$29348 ( \29663 , \29551 , \29566 );
and \U$29349 ( \29664 , \29537 , \29566 );
or \U$29350 ( \29665 , \29662 , \29663 , \29664 );
xor \U$29351 ( \29666 , \29661 , \29665 );
and \U$29352 ( \29667 , \29496 , \29510 );
and \U$29353 ( \29668 , \29510 , \29522 );
and \U$29354 ( \29669 , \29496 , \29522 );
or \U$29355 ( \29670 , \29667 , \29668 , \29669 );
xor \U$29356 ( \29671 , \29666 , \29670 );
and \U$29357 ( \29672 , \29470 , \29474 );
and \U$29358 ( \29673 , \29474 , \29479 );
and \U$29359 ( \29674 , \29470 , \29479 );
or \U$29360 ( \29675 , \29672 , \29673 , \29674 );
and \U$29361 ( \29676 , \29455 , \29459 );
and \U$29362 ( \29677 , \29459 , \29464 );
and \U$29363 ( \29678 , \29455 , \29464 );
or \U$29364 ( \29679 , \29676 , \29677 , \29678 );
xor \U$29365 ( \29680 , \29675 , \29679 );
and \U$29366 ( \29681 , \29444 , \29448 );
and \U$29367 ( \29682 , \29448 , \29450 );
and \U$29368 ( \29683 , \29444 , \29450 );
or \U$29369 ( \29684 , \29681 , \29682 , \29683 );
xor \U$29370 ( \29685 , \29680 , \29684 );
xor \U$29371 ( \29686 , \29671 , \29685 );
and \U$29372 ( \29687 , \29451 , \29465 );
and \U$29373 ( \29688 , \29465 , \29480 );
and \U$29374 ( \29689 , \29451 , \29480 );
or \U$29375 ( \29690 , \29687 , \29688 , \29689 );
and \U$29376 ( \29691 , \29593 , \29597 );
and \U$29377 ( \29692 , \29597 , \29602 );
and \U$29378 ( \29693 , \29593 , \29602 );
or \U$29379 ( \29694 , \29691 , \29692 , \29693 );
and \U$29380 ( \29695 , \29578 , \29582 );
and \U$29381 ( \29696 , \29582 , \29587 );
and \U$29382 ( \29697 , \29578 , \29587 );
or \U$29383 ( \29698 , \29695 , \29696 , \29697 );
xor \U$29384 ( \29699 , \29694 , \29698 );
and \U$29385 ( \29700 , \29572 , \29573 );
xor \U$29386 ( \29701 , \29699 , \29700 );
and \U$29387 ( \29702 , \29556 , \29560 );
and \U$29388 ( \29703 , \29560 , \29565 );
and \U$29389 ( \29704 , \29556 , \29565 );
or \U$29390 ( \29705 , \29702 , \29703 , \29704 );
and \U$29391 ( \29706 , \29541 , \29545 );
and \U$29392 ( \29707 , \29545 , \29550 );
and \U$29393 ( \29708 , \29541 , \29550 );
or \U$29394 ( \29709 , \29706 , \29707 , \29708 );
xor \U$29395 ( \29710 , \29705 , \29709 );
and \U$29396 ( \29711 , \29527 , \29531 );
and \U$29397 ( \29712 , \29531 , \29536 );
and \U$29398 ( \29713 , \29527 , \29536 );
or \U$29399 ( \29714 , \29711 , \29712 , \29713 );
xor \U$29400 ( \29715 , \29710 , \29714 );
xor \U$29401 ( \29716 , \29701 , \29715 );
and \U$29402 ( \29717 , \29512 , \29516 );
and \U$29403 ( \29718 , \29516 , \29521 );
and \U$29404 ( \29719 , \29512 , \29521 );
or \U$29405 ( \29720 , \29717 , \29718 , \29719 );
and \U$29406 ( \29721 , \29500 , \29504 );
and \U$29407 ( \29722 , \29504 , \29509 );
and \U$29408 ( \29723 , \29500 , \29509 );
or \U$29409 ( \29724 , \29721 , \29722 , \29723 );
xor \U$29410 ( \29725 , \29720 , \29724 );
and \U$29411 ( \29726 , \29486 , \29490 );
and \U$29412 ( \29727 , \29490 , \29495 );
and \U$29413 ( \29728 , \29486 , \29495 );
or \U$29414 ( \29729 , \29726 , \29727 , \29728 );
xor \U$29415 ( \29730 , \29725 , \29729 );
xor \U$29416 ( \29731 , \29716 , \29730 );
xor \U$29417 ( \29732 , \29690 , \29731 );
and \U$29418 ( \29733 , \22124 , \22392 );
and \U$29419 ( \29734 , \22089 , \22390 );
nor \U$29420 ( \29735 , \29733 , \29734 );
xnor \U$29421 ( \29736 , \29735 , \22402 );
and \U$29422 ( \29737 , \22145 , \22413 );
and \U$29423 ( \29738 , \22113 , \22411 );
nor \U$29424 ( \29739 , \29737 , \29738 );
xnor \U$29425 ( \29740 , \29739 , \22423 );
xor \U$29426 ( \29741 , \29736 , \29740 );
and \U$29427 ( \29742 , \22167 , \22435 );
and \U$29428 ( \29743 , \22134 , \22433 );
nor \U$29429 ( \29744 , \29742 , \29743 );
xnor \U$29430 ( \29745 , \29744 , \22445 );
xor \U$29431 ( \29746 , \29741 , \29745 );
and \U$29432 ( \29747 , \22894 , \22324 );
and \U$29433 ( \29748 , \23230 , \22322 );
nor \U$29434 ( \29749 , \29747 , \29748 );
xnor \U$29435 ( \29750 , \29749 , \22334 );
and \U$29436 ( \29751 , \22081 , \22345 );
and \U$29437 ( \29752 , \22858 , \22343 );
nor \U$29438 ( \29753 , \29751 , \29752 );
xnor \U$29439 ( \29754 , \29753 , \22355 );
xor \U$29440 ( \29755 , \29750 , \29754 );
and \U$29441 ( \29756 , \22100 , \22367 );
and \U$29442 ( \29757 , \22071 , \22365 );
nor \U$29443 ( \29758 , \29756 , \29757 );
xnor \U$29444 ( \29759 , \29758 , \22377 );
xor \U$29445 ( \29760 , \29755 , \29759 );
xor \U$29446 ( \29761 , \29746 , \29760 );
and \U$29447 ( \29762 , \21990 , \22257 );
not \U$29448 ( \29763 , \29762 );
xnor \U$29449 ( \29764 , \29763 , \22267 );
and \U$29450 ( \29765 , \22001 , \22278 );
and \U$29451 ( \29766 , \21977 , \22276 );
nor \U$29452 ( \29767 , \29765 , \29766 );
xnor \U$29453 ( \29768 , \29767 , \22288 );
xor \U$29454 ( \29769 , \29764 , \29768 );
and \U$29455 ( \29770 , \23329 , \22300 );
and \U$29456 ( \29771 , \22030 , \22298 );
nor \U$29457 ( \29772 , \29770 , \29771 );
xnor \U$29458 ( \29773 , \29772 , \22310 );
xor \U$29459 ( \29774 , \29769 , \29773 );
xor \U$29460 ( \29775 , \29761 , \29774 );
and \U$29461 ( \29776 , \22329 , \22598 );
and \U$29462 ( \29777 , \22294 , \22596 );
nor \U$29463 ( \29778 , \29776 , \29777 );
xnor \U$29464 ( \29779 , \29778 , \22608 );
and \U$29465 ( \29780 , \22350 , \22619 );
and \U$29466 ( \29781 , \22318 , \22617 );
nor \U$29467 ( \29782 , \29780 , \29781 );
xnor \U$29468 ( \29783 , \29782 , \22629 );
xor \U$29469 ( \29784 , \29779 , \29783 );
and \U$29470 ( \29785 , \22372 , \22641 );
and \U$29471 ( \29786 , \22339 , \22639 );
nor \U$29472 ( \29787 , \29785 , \29786 );
xnor \U$29473 ( \29788 , \29787 , \22651 );
xor \U$29474 ( \29789 , \29784 , \29788 );
and \U$29475 ( \29790 , \22262 , \22530 );
and \U$29476 ( \29791 , \22224 , \22528 );
nor \U$29477 ( \29792 , \29790 , \29791 );
xnor \U$29478 ( \29793 , \29792 , \22540 );
and \U$29479 ( \29794 , \22283 , \22551 );
and \U$29480 ( \29795 , \22251 , \22549 );
nor \U$29481 ( \29796 , \29794 , \29795 );
xnor \U$29482 ( \29797 , \29796 , \22561 );
xor \U$29483 ( \29798 , \29793 , \29797 );
and \U$29484 ( \29799 , \22305 , \22573 );
and \U$29485 ( \29800 , \22272 , \22571 );
nor \U$29486 ( \29801 , \29799 , \29800 );
xnor \U$29487 ( \29802 , \29801 , \22583 );
xor \U$29488 ( \29803 , \29798 , \29802 );
xor \U$29489 ( \29804 , \29789 , \29803 );
and \U$29490 ( \29805 , \22192 , \22463 );
and \U$29491 ( \29806 , \22156 , \22461 );
nor \U$29492 ( \29807 , \29805 , \29806 );
xnor \U$29493 ( \29808 , \29807 , \22473 );
and \U$29494 ( \29809 , \22213 , \22484 );
and \U$29495 ( \29810 , \22181 , \22482 );
nor \U$29496 ( \29811 , \29809 , \29810 );
xnor \U$29497 ( \29812 , \29811 , \22494 );
xor \U$29498 ( \29813 , \29808 , \29812 );
and \U$29499 ( \29814 , \22235 , \22506 );
and \U$29500 ( \29815 , \22202 , \22504 );
nor \U$29501 ( \29816 , \29814 , \29815 );
xnor \U$29502 ( \29817 , \29816 , \22516 );
xor \U$29503 ( \29818 , \29813 , \29817 );
xor \U$29504 ( \29819 , \29804 , \29818 );
xor \U$29505 ( \29820 , \29775 , \29819 );
and \U$29506 ( \29821 , \22500 , \21978 );
not \U$29507 ( \29822 , \29821 );
and \U$29508 ( \29823 , \22468 , \23173 );
and \U$29509 ( \29824 , \22429 , \22999 );
nor \U$29510 ( \29825 , \29823 , \29824 );
xnor \U$29511 ( \29826 , \29825 , \22016 );
and \U$29512 ( \29827 , \22489 , \22021 );
and \U$29513 ( \29828 , \22457 , \22019 );
nor \U$29514 ( \29829 , \29827 , \29828 );
xnor \U$29515 ( \29830 , \29829 , \21595 );
xor \U$29516 ( \29831 , \29826 , \29830 );
and \U$29517 ( \29832 , \22511 , \21983 );
and \U$29518 ( \29833 , \22478 , \21981 );
nor \U$29519 ( \29834 , \29832 , \29833 );
xnor \U$29520 ( \29835 , \29834 , \21995 );
xor \U$29521 ( \29836 , \29831 , \29835 );
xor \U$29522 ( \29837 , \29822 , \29836 );
and \U$29523 ( \29838 , \22397 , \22671 );
and \U$29524 ( \29839 , \22361 , \22669 );
nor \U$29525 ( \29840 , \29838 , \29839 );
xnor \U$29526 ( \29841 , \29840 , \22681 );
and \U$29527 ( \29842 , \22418 , \22691 );
and \U$29528 ( \29843 , \22386 , \22689 );
nor \U$29529 ( \29844 , \29842 , \29843 );
xnor \U$29530 ( \29845 , \29844 , \22701 );
xor \U$29531 ( \29846 , \29841 , \29845 );
and \U$29532 ( \29847 , \22440 , \22720 );
and \U$29533 ( \29848 , \22407 , \22707 );
nor \U$29534 ( \29849 , \29847 , \29848 );
xnor \U$29535 ( \29850 , \29849 , \22067 );
xor \U$29536 ( \29851 , \29846 , \29850 );
xor \U$29537 ( \29852 , \29837 , \29851 );
xor \U$29538 ( \29853 , \29820 , \29852 );
xor \U$29539 ( \29854 , \29732 , \29853 );
xor \U$29540 ( \29855 , \29686 , \29854 );
and \U$29541 ( \29856 , \29425 , \29429 );
and \U$29542 ( \29857 , \29429 , \29434 );
and \U$29543 ( \29858 , \29425 , \29434 );
or \U$29544 ( \29859 , \29856 , \29857 , \29858 );
and \U$29545 ( \29860 , \29411 , \29415 );
and \U$29546 ( \29861 , \29415 , \29420 );
and \U$29547 ( \29862 , \29411 , \29420 );
or \U$29548 ( \29863 , \29860 , \29861 , \29862 );
xor \U$29549 ( \29864 , \29859 , \29863 );
and \U$29550 ( \29865 , \29523 , \29567 );
and \U$29551 ( \29866 , \29567 , \29604 );
and \U$29552 ( \29867 , \29523 , \29604 );
or \U$29553 ( \29868 , \29865 , \29866 , \29867 );
xor \U$29554 ( \29869 , \29864 , \29868 );
xor \U$29555 ( \29870 , \29855 , \29869 );
xor \U$29556 ( \29871 , \29657 , \29870 );
xor \U$29557 ( \29872 , \29648 , \29871 );
xor \U$29558 ( \29873 , \29632 , \29872 );
and \U$29559 ( \29874 , \29382 , \29624 );
nor \U$29560 ( \29875 , \29873 , \29874 );
and \U$29561 ( \29876 , \29636 , \29647 );
and \U$29562 ( \29877 , \29647 , \29871 );
and \U$29563 ( \29878 , \29636 , \29871 );
or \U$29564 ( \29879 , \29876 , \29877 , \29878 );
and \U$29565 ( \29880 , \29652 , \29656 );
and \U$29566 ( \29881 , \29656 , \29870 );
and \U$29567 ( \29882 , \29652 , \29870 );
or \U$29568 ( \29883 , \29880 , \29881 , \29882 );
and \U$29569 ( \29884 , \29859 , \29863 );
and \U$29570 ( \29885 , \29863 , \29868 );
and \U$29571 ( \29886 , \29859 , \29868 );
or \U$29572 ( \29887 , \29884 , \29885 , \29886 );
and \U$29573 ( \29888 , \29690 , \29731 );
and \U$29574 ( \29889 , \29731 , \29853 );
and \U$29575 ( \29890 , \29690 , \29853 );
or \U$29576 ( \29891 , \29888 , \29889 , \29890 );
xor \U$29577 ( \29892 , \29887 , \29891 );
and \U$29578 ( \29893 , \29671 , \29685 );
xor \U$29579 ( \29894 , \29892 , \29893 );
xor \U$29580 ( \29895 , \29883 , \29894 );
and \U$29581 ( \29896 , \29640 , \29644 );
and \U$29582 ( \29897 , \29644 , \29646 );
and \U$29583 ( \29898 , \29640 , \29646 );
or \U$29584 ( \29899 , \29896 , \29897 , \29898 );
and \U$29585 ( \29900 , \29686 , \29854 );
and \U$29586 ( \29901 , \29854 , \29869 );
and \U$29587 ( \29902 , \29686 , \29869 );
or \U$29588 ( \29903 , \29900 , \29901 , \29902 );
xor \U$29589 ( \29904 , \29899 , \29903 );
and \U$29590 ( \29905 , \29822 , \29836 );
and \U$29591 ( \29906 , \29836 , \29851 );
and \U$29592 ( \29907 , \29822 , \29851 );
or \U$29593 ( \29908 , \29905 , \29906 , \29907 );
and \U$29594 ( \29909 , \29789 , \29803 );
and \U$29595 ( \29910 , \29803 , \29818 );
and \U$29596 ( \29911 , \29789 , \29818 );
or \U$29597 ( \29912 , \29909 , \29910 , \29911 );
xor \U$29598 ( \29913 , \29908 , \29912 );
and \U$29599 ( \29914 , \29746 , \29760 );
and \U$29600 ( \29915 , \29760 , \29774 );
and \U$29601 ( \29916 , \29746 , \29774 );
or \U$29602 ( \29917 , \29914 , \29915 , \29916 );
xor \U$29603 ( \29918 , \29913 , \29917 );
and \U$29604 ( \29919 , \29720 , \29724 );
and \U$29605 ( \29920 , \29724 , \29729 );
and \U$29606 ( \29921 , \29720 , \29729 );
or \U$29607 ( \29922 , \29919 , \29920 , \29921 );
and \U$29608 ( \29923 , \29705 , \29709 );
and \U$29609 ( \29924 , \29709 , \29714 );
and \U$29610 ( \29925 , \29705 , \29714 );
or \U$29611 ( \29926 , \29923 , \29924 , \29925 );
xor \U$29612 ( \29927 , \29922 , \29926 );
and \U$29613 ( \29928 , \29694 , \29698 );
and \U$29614 ( \29929 , \29698 , \29700 );
and \U$29615 ( \29930 , \29694 , \29700 );
or \U$29616 ( \29931 , \29928 , \29929 , \29930 );
xor \U$29617 ( \29932 , \29927 , \29931 );
xor \U$29618 ( \29933 , \29918 , \29932 );
and \U$29619 ( \29934 , \29701 , \29715 );
and \U$29620 ( \29935 , \29715 , \29730 );
and \U$29621 ( \29936 , \29701 , \29730 );
or \U$29622 ( \29937 , \29934 , \29935 , \29936 );
and \U$29623 ( \29938 , \29841 , \29845 );
and \U$29624 ( \29939 , \29845 , \29850 );
and \U$29625 ( \29940 , \29841 , \29850 );
or \U$29626 ( \29941 , \29938 , \29939 , \29940 );
and \U$29627 ( \29942 , \29826 , \29830 );
and \U$29628 ( \29943 , \29830 , \29835 );
and \U$29629 ( \29944 , \29826 , \29835 );
or \U$29630 ( \29945 , \29942 , \29943 , \29944 );
xor \U$29631 ( \29946 , \29941 , \29945 );
xor \U$29632 ( \29947 , \29946 , \29821 );
and \U$29633 ( \29948 , \29808 , \29812 );
and \U$29634 ( \29949 , \29812 , \29817 );
and \U$29635 ( \29950 , \29808 , \29817 );
or \U$29636 ( \29951 , \29948 , \29949 , \29950 );
and \U$29637 ( \29952 , \29793 , \29797 );
and \U$29638 ( \29953 , \29797 , \29802 );
and \U$29639 ( \29954 , \29793 , \29802 );
or \U$29640 ( \29955 , \29952 , \29953 , \29954 );
xor \U$29641 ( \29956 , \29951 , \29955 );
and \U$29642 ( \29957 , \29779 , \29783 );
and \U$29643 ( \29958 , \29783 , \29788 );
and \U$29644 ( \29959 , \29779 , \29788 );
or \U$29645 ( \29960 , \29957 , \29958 , \29959 );
xor \U$29646 ( \29961 , \29956 , \29960 );
xor \U$29647 ( \29962 , \29947 , \29961 );
and \U$29648 ( \29963 , \29764 , \29768 );
and \U$29649 ( \29964 , \29768 , \29773 );
and \U$29650 ( \29965 , \29764 , \29773 );
or \U$29651 ( \29966 , \29963 , \29964 , \29965 );
and \U$29652 ( \29967 , \29750 , \29754 );
and \U$29653 ( \29968 , \29754 , \29759 );
and \U$29654 ( \29969 , \29750 , \29759 );
or \U$29655 ( \29970 , \29967 , \29968 , \29969 );
xor \U$29656 ( \29971 , \29966 , \29970 );
and \U$29657 ( \29972 , \29736 , \29740 );
and \U$29658 ( \29973 , \29740 , \29745 );
and \U$29659 ( \29974 , \29736 , \29745 );
or \U$29660 ( \29975 , \29972 , \29973 , \29974 );
xor \U$29661 ( \29976 , \29971 , \29975 );
xor \U$29662 ( \29977 , \29962 , \29976 );
xor \U$29663 ( \29978 , \29937 , \29977 );
and \U$29664 ( \29979 , \22089 , \22392 );
and \U$29665 ( \29980 , \22100 , \22390 );
nor \U$29666 ( \29981 , \29979 , \29980 );
xnor \U$29667 ( \29982 , \29981 , \22402 );
and \U$29668 ( \29983 , \22113 , \22413 );
and \U$29669 ( \29984 , \22124 , \22411 );
nor \U$29670 ( \29985 , \29983 , \29984 );
xnor \U$29671 ( \29986 , \29985 , \22423 );
xor \U$29672 ( \29987 , \29982 , \29986 );
and \U$29673 ( \29988 , \22134 , \22435 );
and \U$29674 ( \29989 , \22145 , \22433 );
nor \U$29675 ( \29990 , \29988 , \29989 );
xnor \U$29676 ( \29991 , \29990 , \22445 );
xor \U$29677 ( \29992 , \29987 , \29991 );
and \U$29678 ( \29993 , \23230 , \22324 );
and \U$29679 ( \29994 , \23329 , \22322 );
nor \U$29680 ( \29995 , \29993 , \29994 );
xnor \U$29681 ( \29996 , \29995 , \22334 );
and \U$29682 ( \29997 , \22858 , \22345 );
and \U$29683 ( \29998 , \22894 , \22343 );
nor \U$29684 ( \29999 , \29997 , \29998 );
xnor \U$29685 ( \30000 , \29999 , \22355 );
xor \U$29686 ( \30001 , \29996 , \30000 );
and \U$29687 ( \30002 , \22071 , \22367 );
and \U$29688 ( \30003 , \22081 , \22365 );
nor \U$29689 ( \30004 , \30002 , \30003 );
xnor \U$29690 ( \30005 , \30004 , \22377 );
xor \U$29691 ( \30006 , \30001 , \30005 );
xor \U$29692 ( \30007 , \29992 , \30006 );
not \U$29693 ( \30008 , \22267 );
and \U$29694 ( \30009 , \21977 , \22278 );
and \U$29695 ( \30010 , \21990 , \22276 );
nor \U$29696 ( \30011 , \30009 , \30010 );
xnor \U$29697 ( \30012 , \30011 , \22288 );
xor \U$29698 ( \30013 , \30008 , \30012 );
and \U$29699 ( \30014 , \22030 , \22300 );
and \U$29700 ( \30015 , \22001 , \22298 );
nor \U$29701 ( \30016 , \30014 , \30015 );
xnor \U$29702 ( \30017 , \30016 , \22310 );
xor \U$29703 ( \30018 , \30013 , \30017 );
xor \U$29704 ( \30019 , \30007 , \30018 );
and \U$29705 ( \30020 , \22294 , \22598 );
and \U$29706 ( \30021 , \22305 , \22596 );
nor \U$29707 ( \30022 , \30020 , \30021 );
xnor \U$29708 ( \30023 , \30022 , \22608 );
and \U$29709 ( \30024 , \22318 , \22619 );
and \U$29710 ( \30025 , \22329 , \22617 );
nor \U$29711 ( \30026 , \30024 , \30025 );
xnor \U$29712 ( \30027 , \30026 , \22629 );
xor \U$29713 ( \30028 , \30023 , \30027 );
and \U$29714 ( \30029 , \22339 , \22641 );
and \U$29715 ( \30030 , \22350 , \22639 );
nor \U$29716 ( \30031 , \30029 , \30030 );
xnor \U$29717 ( \30032 , \30031 , \22651 );
xor \U$29718 ( \30033 , \30028 , \30032 );
and \U$29719 ( \30034 , \22224 , \22530 );
and \U$29720 ( \30035 , \22235 , \22528 );
nor \U$29721 ( \30036 , \30034 , \30035 );
xnor \U$29722 ( \30037 , \30036 , \22540 );
and \U$29723 ( \30038 , \22251 , \22551 );
and \U$29724 ( \30039 , \22262 , \22549 );
nor \U$29725 ( \30040 , \30038 , \30039 );
xnor \U$29726 ( \30041 , \30040 , \22561 );
xor \U$29727 ( \30042 , \30037 , \30041 );
and \U$29728 ( \30043 , \22272 , \22573 );
and \U$29729 ( \30044 , \22283 , \22571 );
nor \U$29730 ( \30045 , \30043 , \30044 );
xnor \U$29731 ( \30046 , \30045 , \22583 );
xor \U$29732 ( \30047 , \30042 , \30046 );
xor \U$29733 ( \30048 , \30033 , \30047 );
and \U$29734 ( \30049 , \22156 , \22463 );
and \U$29735 ( \30050 , \22167 , \22461 );
nor \U$29736 ( \30051 , \30049 , \30050 );
xnor \U$29737 ( \30052 , \30051 , \22473 );
and \U$29738 ( \30053 , \22181 , \22484 );
and \U$29739 ( \30054 , \22192 , \22482 );
nor \U$29740 ( \30055 , \30053 , \30054 );
xnor \U$29741 ( \30056 , \30055 , \22494 );
xor \U$29742 ( \30057 , \30052 , \30056 );
and \U$29743 ( \30058 , \22202 , \22506 );
and \U$29744 ( \30059 , \22213 , \22504 );
nor \U$29745 ( \30060 , \30058 , \30059 );
xnor \U$29746 ( \30061 , \30060 , \22516 );
xor \U$29747 ( \30062 , \30057 , \30061 );
xor \U$29748 ( \30063 , \30048 , \30062 );
xor \U$29749 ( \30064 , \30019 , \30063 );
and \U$29750 ( \30065 , \22511 , \21978 );
and \U$29751 ( \30066 , \22429 , \23173 );
and \U$29752 ( \30067 , \22440 , \22999 );
nor \U$29753 ( \30068 , \30066 , \30067 );
xnor \U$29754 ( \30069 , \30068 , \22016 );
and \U$29755 ( \30070 , \22457 , \22021 );
and \U$29756 ( \30071 , \22468 , \22019 );
nor \U$29757 ( \30072 , \30070 , \30071 );
xnor \U$29758 ( \30073 , \30072 , \21595 );
xor \U$29759 ( \30074 , \30069 , \30073 );
and \U$29760 ( \30075 , \22478 , \21983 );
and \U$29761 ( \30076 , \22489 , \21981 );
nor \U$29762 ( \30077 , \30075 , \30076 );
xnor \U$29763 ( \30078 , \30077 , \21995 );
xor \U$29764 ( \30079 , \30074 , \30078 );
xor \U$29765 ( \30080 , \30065 , \30079 );
and \U$29766 ( \30081 , \22361 , \22671 );
and \U$29767 ( \30082 , \22372 , \22669 );
nor \U$29768 ( \30083 , \30081 , \30082 );
xnor \U$29769 ( \30084 , \30083 , \22681 );
and \U$29770 ( \30085 , \22386 , \22691 );
and \U$29771 ( \30086 , \22397 , \22689 );
nor \U$29772 ( \30087 , \30085 , \30086 );
xnor \U$29773 ( \30088 , \30087 , \22701 );
xor \U$29774 ( \30089 , \30084 , \30088 );
and \U$29775 ( \30090 , \22407 , \22720 );
and \U$29776 ( \30091 , \22418 , \22707 );
nor \U$29777 ( \30092 , \30090 , \30091 );
xnor \U$29778 ( \30093 , \30092 , \22067 );
xor \U$29779 ( \30094 , \30089 , \30093 );
xor \U$29780 ( \30095 , \30080 , \30094 );
xor \U$29781 ( \30096 , \30064 , \30095 );
xor \U$29782 ( \30097 , \29978 , \30096 );
xor \U$29783 ( \30098 , \29933 , \30097 );
and \U$29784 ( \30099 , \29675 , \29679 );
and \U$29785 ( \30100 , \29679 , \29684 );
and \U$29786 ( \30101 , \29675 , \29684 );
or \U$29787 ( \30102 , \30099 , \30100 , \30101 );
and \U$29788 ( \30103 , \29661 , \29665 );
and \U$29789 ( \30104 , \29665 , \29670 );
and \U$29790 ( \30105 , \29661 , \29670 );
or \U$29791 ( \30106 , \30103 , \30104 , \30105 );
xor \U$29792 ( \30107 , \30102 , \30106 );
and \U$29793 ( \30108 , \29775 , \29819 );
and \U$29794 ( \30109 , \29819 , \29852 );
and \U$29795 ( \30110 , \29775 , \29852 );
or \U$29796 ( \30111 , \30108 , \30109 , \30110 );
xor \U$29797 ( \30112 , \30107 , \30111 );
xor \U$29798 ( \30113 , \30098 , \30112 );
xor \U$29799 ( \30114 , \29904 , \30113 );
xor \U$29800 ( \30115 , \29895 , \30114 );
xor \U$29801 ( \30116 , \29879 , \30115 );
and \U$29802 ( \30117 , \29632 , \29872 );
nor \U$29803 ( \30118 , \30116 , \30117 );
nor \U$29804 ( \30119 , \29875 , \30118 );
nand \U$29805 ( \30120 , \29628 , \30119 );
and \U$29806 ( \30121 , \29883 , \29894 );
and \U$29807 ( \30122 , \29894 , \30114 );
and \U$29808 ( \30123 , \29883 , \30114 );
or \U$29809 ( \30124 , \30121 , \30122 , \30123 );
and \U$29810 ( \30125 , \29899 , \29903 );
and \U$29811 ( \30126 , \29903 , \30113 );
and \U$29812 ( \30127 , \29899 , \30113 );
or \U$29813 ( \30128 , \30125 , \30126 , \30127 );
and \U$29814 ( \30129 , \30102 , \30106 );
and \U$29815 ( \30130 , \30106 , \30111 );
and \U$29816 ( \30131 , \30102 , \30111 );
or \U$29817 ( \30132 , \30129 , \30130 , \30131 );
and \U$29818 ( \30133 , \29937 , \29977 );
and \U$29819 ( \30134 , \29977 , \30096 );
and \U$29820 ( \30135 , \29937 , \30096 );
or \U$29821 ( \30136 , \30133 , \30134 , \30135 );
xor \U$29822 ( \30137 , \30132 , \30136 );
and \U$29823 ( \30138 , \29918 , \29932 );
xor \U$29824 ( \30139 , \30137 , \30138 );
xor \U$29825 ( \30140 , \30128 , \30139 );
and \U$29826 ( \30141 , \29887 , \29891 );
and \U$29827 ( \30142 , \29891 , \29893 );
and \U$29828 ( \30143 , \29887 , \29893 );
or \U$29829 ( \30144 , \30141 , \30142 , \30143 );
and \U$29830 ( \30145 , \29933 , \30097 );
and \U$29831 ( \30146 , \30097 , \30112 );
and \U$29832 ( \30147 , \29933 , \30112 );
or \U$29833 ( \30148 , \30145 , \30146 , \30147 );
xor \U$29834 ( \30149 , \30144 , \30148 );
and \U$29835 ( \30150 , \30065 , \30079 );
and \U$29836 ( \30151 , \30079 , \30094 );
and \U$29837 ( \30152 , \30065 , \30094 );
or \U$29838 ( \30153 , \30150 , \30151 , \30152 );
and \U$29839 ( \30154 , \30033 , \30047 );
and \U$29840 ( \30155 , \30047 , \30062 );
and \U$29841 ( \30156 , \30033 , \30062 );
or \U$29842 ( \30157 , \30154 , \30155 , \30156 );
xor \U$29843 ( \30158 , \30153 , \30157 );
and \U$29844 ( \30159 , \29992 , \30006 );
and \U$29845 ( \30160 , \30006 , \30018 );
and \U$29846 ( \30161 , \29992 , \30018 );
or \U$29847 ( \30162 , \30159 , \30160 , \30161 );
xor \U$29848 ( \30163 , \30158 , \30162 );
and \U$29849 ( \30164 , \29966 , \29970 );
and \U$29850 ( \30165 , \29970 , \29975 );
and \U$29851 ( \30166 , \29966 , \29975 );
or \U$29852 ( \30167 , \30164 , \30165 , \30166 );
and \U$29853 ( \30168 , \29951 , \29955 );
and \U$29854 ( \30169 , \29955 , \29960 );
and \U$29855 ( \30170 , \29951 , \29960 );
or \U$29856 ( \30171 , \30168 , \30169 , \30170 );
xor \U$29857 ( \30172 , \30167 , \30171 );
and \U$29858 ( \30173 , \29941 , \29945 );
and \U$29859 ( \30174 , \29945 , \29821 );
and \U$29860 ( \30175 , \29941 , \29821 );
or \U$29861 ( \30176 , \30173 , \30174 , \30175 );
xor \U$29862 ( \30177 , \30172 , \30176 );
xor \U$29863 ( \30178 , \30163 , \30177 );
and \U$29864 ( \30179 , \29947 , \29961 );
and \U$29865 ( \30180 , \29961 , \29976 );
and \U$29866 ( \30181 , \29947 , \29976 );
or \U$29867 ( \30182 , \30179 , \30180 , \30181 );
and \U$29868 ( \30183 , \30084 , \30088 );
and \U$29869 ( \30184 , \30088 , \30093 );
and \U$29870 ( \30185 , \30084 , \30093 );
or \U$29871 ( \30186 , \30183 , \30184 , \30185 );
and \U$29872 ( \30187 , \30069 , \30073 );
and \U$29873 ( \30188 , \30073 , \30078 );
and \U$29874 ( \30189 , \30069 , \30078 );
or \U$29875 ( \30190 , \30187 , \30188 , \30189 );
xnor \U$29876 ( \30191 , \30186 , \30190 );
and \U$29877 ( \30192 , \30052 , \30056 );
and \U$29878 ( \30193 , \30056 , \30061 );
and \U$29879 ( \30194 , \30052 , \30061 );
or \U$29880 ( \30195 , \30192 , \30193 , \30194 );
and \U$29881 ( \30196 , \30037 , \30041 );
and \U$29882 ( \30197 , \30041 , \30046 );
and \U$29883 ( \30198 , \30037 , \30046 );
or \U$29884 ( \30199 , \30196 , \30197 , \30198 );
xor \U$29885 ( \30200 , \30195 , \30199 );
and \U$29886 ( \30201 , \30023 , \30027 );
and \U$29887 ( \30202 , \30027 , \30032 );
and \U$29888 ( \30203 , \30023 , \30032 );
or \U$29889 ( \30204 , \30201 , \30202 , \30203 );
xor \U$29890 ( \30205 , \30200 , \30204 );
xor \U$29891 ( \30206 , \30191 , \30205 );
and \U$29892 ( \30207 , \30008 , \30012 );
and \U$29893 ( \30208 , \30012 , \30017 );
and \U$29894 ( \30209 , \30008 , \30017 );
or \U$29895 ( \30210 , \30207 , \30208 , \30209 );
and \U$29896 ( \30211 , \29996 , \30000 );
and \U$29897 ( \30212 , \30000 , \30005 );
and \U$29898 ( \30213 , \29996 , \30005 );
or \U$29899 ( \30214 , \30211 , \30212 , \30213 );
xor \U$29900 ( \30215 , \30210 , \30214 );
and \U$29901 ( \30216 , \29982 , \29986 );
and \U$29902 ( \30217 , \29986 , \29991 );
and \U$29903 ( \30218 , \29982 , \29991 );
or \U$29904 ( \30219 , \30216 , \30217 , \30218 );
xor \U$29905 ( \30220 , \30215 , \30219 );
xor \U$29906 ( \30221 , \30206 , \30220 );
xor \U$29907 ( \30222 , \30182 , \30221 );
and \U$29908 ( \30223 , \22894 , \22345 );
and \U$29909 ( \30224 , \23230 , \22343 );
nor \U$29910 ( \30225 , \30223 , \30224 );
xnor \U$29911 ( \30226 , \30225 , \22355 );
and \U$29912 ( \30227 , \22081 , \22367 );
and \U$29913 ( \30228 , \22858 , \22365 );
nor \U$29914 ( \30229 , \30227 , \30228 );
xnor \U$29915 ( \30230 , \30229 , \22377 );
xor \U$29916 ( \30231 , \30226 , \30230 );
and \U$29917 ( \30232 , \22100 , \22392 );
and \U$29918 ( \30233 , \22071 , \22390 );
nor \U$29919 ( \30234 , \30232 , \30233 );
xnor \U$29920 ( \30235 , \30234 , \22402 );
xor \U$29921 ( \30236 , \30231 , \30235 );
and \U$29922 ( \30237 , \21990 , \22278 );
not \U$29923 ( \30238 , \30237 );
xnor \U$29924 ( \30239 , \30238 , \22288 );
and \U$29925 ( \30240 , \22001 , \22300 );
and \U$29926 ( \30241 , \21977 , \22298 );
nor \U$29927 ( \30242 , \30240 , \30241 );
xnor \U$29928 ( \30243 , \30242 , \22310 );
xor \U$29929 ( \30244 , \30239 , \30243 );
and \U$29930 ( \30245 , \23329 , \22324 );
and \U$29931 ( \30246 , \22030 , \22322 );
nor \U$29932 ( \30247 , \30245 , \30246 );
xnor \U$29933 ( \30248 , \30247 , \22334 );
xor \U$29934 ( \30249 , \30244 , \30248 );
xor \U$29935 ( \30250 , \30236 , \30249 );
and \U$29936 ( \30251 , \22262 , \22551 );
and \U$29937 ( \30252 , \22224 , \22549 );
nor \U$29938 ( \30253 , \30251 , \30252 );
xnor \U$29939 ( \30254 , \30253 , \22561 );
and \U$29940 ( \30255 , \22283 , \22573 );
and \U$29941 ( \30256 , \22251 , \22571 );
nor \U$29942 ( \30257 , \30255 , \30256 );
xnor \U$29943 ( \30258 , \30257 , \22583 );
xor \U$29944 ( \30259 , \30254 , \30258 );
and \U$29945 ( \30260 , \22305 , \22598 );
and \U$29946 ( \30261 , \22272 , \22596 );
nor \U$29947 ( \30262 , \30260 , \30261 );
xnor \U$29948 ( \30263 , \30262 , \22608 );
xor \U$29949 ( \30264 , \30259 , \30263 );
and \U$29950 ( \30265 , \22192 , \22484 );
and \U$29951 ( \30266 , \22156 , \22482 );
nor \U$29952 ( \30267 , \30265 , \30266 );
xnor \U$29953 ( \30268 , \30267 , \22494 );
and \U$29954 ( \30269 , \22213 , \22506 );
and \U$29955 ( \30270 , \22181 , \22504 );
nor \U$29956 ( \30271 , \30269 , \30270 );
xnor \U$29957 ( \30272 , \30271 , \22516 );
xor \U$29958 ( \30273 , \30268 , \30272 );
and \U$29959 ( \30274 , \22235 , \22530 );
and \U$29960 ( \30275 , \22202 , \22528 );
nor \U$29961 ( \30276 , \30274 , \30275 );
xnor \U$29962 ( \30277 , \30276 , \22540 );
xor \U$29963 ( \30278 , \30273 , \30277 );
xor \U$29964 ( \30279 , \30264 , \30278 );
and \U$29965 ( \30280 , \22124 , \22413 );
and \U$29966 ( \30281 , \22089 , \22411 );
nor \U$29967 ( \30282 , \30280 , \30281 );
xnor \U$29968 ( \30283 , \30282 , \22423 );
and \U$29969 ( \30284 , \22145 , \22435 );
and \U$29970 ( \30285 , \22113 , \22433 );
nor \U$29971 ( \30286 , \30284 , \30285 );
xnor \U$29972 ( \30287 , \30286 , \22445 );
xor \U$29973 ( \30288 , \30283 , \30287 );
and \U$29974 ( \30289 , \22167 , \22463 );
and \U$29975 ( \30290 , \22134 , \22461 );
nor \U$29976 ( \30291 , \30289 , \30290 );
xnor \U$29977 ( \30292 , \30291 , \22473 );
xor \U$29978 ( \30293 , \30288 , \30292 );
xor \U$29979 ( \30294 , \30279 , \30293 );
xor \U$29980 ( \30295 , \30250 , \30294 );
and \U$29981 ( \30296 , \22468 , \22021 );
and \U$29982 ( \30297 , \22429 , \22019 );
nor \U$29983 ( \30298 , \30296 , \30297 );
xnor \U$29984 ( \30299 , \30298 , \21595 );
and \U$29985 ( \30300 , \22489 , \21983 );
and \U$29986 ( \30301 , \22457 , \21981 );
nor \U$29987 ( \30302 , \30300 , \30301 );
xnor \U$29988 ( \30303 , \30302 , \21995 );
xor \U$29989 ( \30304 , \30299 , \30303 );
and \U$29990 ( \30305 , \22478 , \21978 );
xor \U$29991 ( \30306 , \30304 , \30305 );
and \U$29992 ( \30307 , \22397 , \22691 );
and \U$29993 ( \30308 , \22361 , \22689 );
nor \U$29994 ( \30309 , \30307 , \30308 );
xnor \U$29995 ( \30310 , \30309 , \22701 );
and \U$29996 ( \30311 , \22418 , \22720 );
and \U$29997 ( \30312 , \22386 , \22707 );
nor \U$29998 ( \30313 , \30311 , \30312 );
xnor \U$29999 ( \30314 , \30313 , \22067 );
xor \U$30000 ( \30315 , \30310 , \30314 );
and \U$30001 ( \30316 , \22440 , \23173 );
and \U$30002 ( \30317 , \22407 , \22999 );
nor \U$30003 ( \30318 , \30316 , \30317 );
xnor \U$30004 ( \30319 , \30318 , \22016 );
xor \U$30005 ( \30320 , \30315 , \30319 );
xor \U$30006 ( \30321 , \30306 , \30320 );
and \U$30007 ( \30322 , \22329 , \22619 );
and \U$30008 ( \30323 , \22294 , \22617 );
nor \U$30009 ( \30324 , \30322 , \30323 );
xnor \U$30010 ( \30325 , \30324 , \22629 );
and \U$30011 ( \30326 , \22350 , \22641 );
and \U$30012 ( \30327 , \22318 , \22639 );
nor \U$30013 ( \30328 , \30326 , \30327 );
xnor \U$30014 ( \30329 , \30328 , \22651 );
xor \U$30015 ( \30330 , \30325 , \30329 );
and \U$30016 ( \30331 , \22372 , \22671 );
and \U$30017 ( \30332 , \22339 , \22669 );
nor \U$30018 ( \30333 , \30331 , \30332 );
xnor \U$30019 ( \30334 , \30333 , \22681 );
xor \U$30020 ( \30335 , \30330 , \30334 );
xor \U$30021 ( \30336 , \30321 , \30335 );
xor \U$30022 ( \30337 , \30295 , \30336 );
xor \U$30023 ( \30338 , \30222 , \30337 );
xor \U$30024 ( \30339 , \30178 , \30338 );
and \U$30025 ( \30340 , \29922 , \29926 );
and \U$30026 ( \30341 , \29926 , \29931 );
and \U$30027 ( \30342 , \29922 , \29931 );
or \U$30028 ( \30343 , \30340 , \30341 , \30342 );
and \U$30029 ( \30344 , \29908 , \29912 );
and \U$30030 ( \30345 , \29912 , \29917 );
and \U$30031 ( \30346 , \29908 , \29917 );
or \U$30032 ( \30347 , \30344 , \30345 , \30346 );
xor \U$30033 ( \30348 , \30343 , \30347 );
and \U$30034 ( \30349 , \30019 , \30063 );
and \U$30035 ( \30350 , \30063 , \30095 );
and \U$30036 ( \30351 , \30019 , \30095 );
or \U$30037 ( \30352 , \30349 , \30350 , \30351 );
xor \U$30038 ( \30353 , \30348 , \30352 );
xor \U$30039 ( \30354 , \30339 , \30353 );
xor \U$30040 ( \30355 , \30149 , \30354 );
xor \U$30041 ( \30356 , \30140 , \30355 );
xor \U$30042 ( \30357 , \30124 , \30356 );
and \U$30043 ( \30358 , \29879 , \30115 );
nor \U$30044 ( \30359 , \30357 , \30358 );
and \U$30045 ( \30360 , \30128 , \30139 );
and \U$30046 ( \30361 , \30139 , \30355 );
and \U$30047 ( \30362 , \30128 , \30355 );
or \U$30048 ( \30363 , \30360 , \30361 , \30362 );
and \U$30049 ( \30364 , \30144 , \30148 );
and \U$30050 ( \30365 , \30148 , \30354 );
and \U$30051 ( \30366 , \30144 , \30354 );
or \U$30052 ( \30367 , \30364 , \30365 , \30366 );
and \U$30053 ( \30368 , \30343 , \30347 );
and \U$30054 ( \30369 , \30347 , \30352 );
and \U$30055 ( \30370 , \30343 , \30352 );
or \U$30056 ( \30371 , \30368 , \30369 , \30370 );
and \U$30057 ( \30372 , \30182 , \30221 );
and \U$30058 ( \30373 , \30221 , \30337 );
and \U$30059 ( \30374 , \30182 , \30337 );
or \U$30060 ( \30375 , \30372 , \30373 , \30374 );
xor \U$30061 ( \30376 , \30371 , \30375 );
and \U$30062 ( \30377 , \30163 , \30177 );
xor \U$30063 ( \30378 , \30376 , \30377 );
xor \U$30064 ( \30379 , \30367 , \30378 );
and \U$30065 ( \30380 , \30132 , \30136 );
and \U$30066 ( \30381 , \30136 , \30138 );
and \U$30067 ( \30382 , \30132 , \30138 );
or \U$30068 ( \30383 , \30380 , \30381 , \30382 );
and \U$30069 ( \30384 , \30178 , \30338 );
and \U$30070 ( \30385 , \30338 , \30353 );
and \U$30071 ( \30386 , \30178 , \30353 );
or \U$30072 ( \30387 , \30384 , \30385 , \30386 );
xor \U$30073 ( \30388 , \30383 , \30387 );
and \U$30074 ( \30389 , \30306 , \30320 );
and \U$30075 ( \30390 , \30320 , \30335 );
and \U$30076 ( \30391 , \30306 , \30335 );
or \U$30077 ( \30392 , \30389 , \30390 , \30391 );
and \U$30078 ( \30393 , \30264 , \30278 );
and \U$30079 ( \30394 , \30278 , \30293 );
and \U$30080 ( \30395 , \30264 , \30293 );
or \U$30081 ( \30396 , \30393 , \30394 , \30395 );
xor \U$30082 ( \30397 , \30392 , \30396 );
and \U$30083 ( \30398 , \30236 , \30249 );
xor \U$30084 ( \30399 , \30397 , \30398 );
and \U$30085 ( \30400 , \30210 , \30214 );
and \U$30086 ( \30401 , \30214 , \30219 );
and \U$30087 ( \30402 , \30210 , \30219 );
or \U$30088 ( \30403 , \30400 , \30401 , \30402 );
and \U$30089 ( \30404 , \30195 , \30199 );
and \U$30090 ( \30405 , \30199 , \30204 );
and \U$30091 ( \30406 , \30195 , \30204 );
or \U$30092 ( \30407 , \30404 , \30405 , \30406 );
xor \U$30093 ( \30408 , \30403 , \30407 );
or \U$30094 ( \30409 , \30186 , \30190 );
xor \U$30095 ( \30410 , \30408 , \30409 );
xor \U$30096 ( \30411 , \30399 , \30410 );
and \U$30097 ( \30412 , \30191 , \30205 );
and \U$30098 ( \30413 , \30205 , \30220 );
and \U$30099 ( \30414 , \30191 , \30220 );
or \U$30100 ( \30415 , \30412 , \30413 , \30414 );
and \U$30101 ( \30416 , \30310 , \30314 );
and \U$30102 ( \30417 , \30314 , \30319 );
and \U$30103 ( \30418 , \30310 , \30319 );
or \U$30104 ( \30419 , \30416 , \30417 , \30418 );
and \U$30105 ( \30420 , \30299 , \30303 );
and \U$30106 ( \30421 , \30303 , \30305 );
and \U$30107 ( \30422 , \30299 , \30305 );
or \U$30108 ( \30423 , \30420 , \30421 , \30422 );
xor \U$30109 ( \30424 , \30419 , \30423 );
and \U$30110 ( \30425 , \22429 , \22021 );
and \U$30111 ( \30426 , \22440 , \22019 );
nor \U$30112 ( \30427 , \30425 , \30426 );
xnor \U$30113 ( \30428 , \30427 , \21595 );
and \U$30114 ( \30429 , \22457 , \21983 );
and \U$30115 ( \30430 , \22468 , \21981 );
nor \U$30116 ( \30431 , \30429 , \30430 );
xnor \U$30117 ( \30432 , \30431 , \21995 );
xor \U$30118 ( \30433 , \30428 , \30432 );
and \U$30119 ( \30434 , \22489 , \21978 );
xor \U$30120 ( \30435 , \30433 , \30434 );
xor \U$30121 ( \30436 , \30424 , \30435 );
and \U$30122 ( \30437 , \30268 , \30272 );
and \U$30123 ( \30438 , \30272 , \30277 );
and \U$30124 ( \30439 , \30268 , \30277 );
or \U$30125 ( \30440 , \30437 , \30438 , \30439 );
and \U$30126 ( \30441 , \30254 , \30258 );
and \U$30127 ( \30442 , \30258 , \30263 );
and \U$30128 ( \30443 , \30254 , \30263 );
or \U$30129 ( \30444 , \30441 , \30442 , \30443 );
xor \U$30130 ( \30445 , \30440 , \30444 );
and \U$30131 ( \30446 , \30325 , \30329 );
and \U$30132 ( \30447 , \30329 , \30334 );
and \U$30133 ( \30448 , \30325 , \30334 );
or \U$30134 ( \30449 , \30446 , \30447 , \30448 );
xor \U$30135 ( \30450 , \30445 , \30449 );
xor \U$30136 ( \30451 , \30436 , \30450 );
and \U$30137 ( \30452 , \30239 , \30243 );
and \U$30138 ( \30453 , \30243 , \30248 );
and \U$30139 ( \30454 , \30239 , \30248 );
or \U$30140 ( \30455 , \30452 , \30453 , \30454 );
and \U$30141 ( \30456 , \30226 , \30230 );
and \U$30142 ( \30457 , \30230 , \30235 );
and \U$30143 ( \30458 , \30226 , \30235 );
or \U$30144 ( \30459 , \30456 , \30457 , \30458 );
xor \U$30145 ( \30460 , \30455 , \30459 );
and \U$30146 ( \30461 , \30283 , \30287 );
and \U$30147 ( \30462 , \30287 , \30292 );
and \U$30148 ( \30463 , \30283 , \30292 );
or \U$30149 ( \30464 , \30461 , \30462 , \30463 );
xor \U$30150 ( \30465 , \30460 , \30464 );
xor \U$30151 ( \30466 , \30451 , \30465 );
xor \U$30152 ( \30467 , \30415 , \30466 );
not \U$30153 ( \30468 , \22288 );
and \U$30154 ( \30469 , \21977 , \22300 );
and \U$30155 ( \30470 , \21990 , \22298 );
nor \U$30156 ( \30471 , \30469 , \30470 );
xnor \U$30157 ( \30472 , \30471 , \22310 );
xor \U$30158 ( \30473 , \30468 , \30472 );
and \U$30159 ( \30474 , \22030 , \22324 );
and \U$30160 ( \30475 , \22001 , \22322 );
nor \U$30161 ( \30476 , \30474 , \30475 );
xnor \U$30162 ( \30477 , \30476 , \22334 );
xor \U$30163 ( \30478 , \30473 , \30477 );
and \U$30164 ( \30479 , \22156 , \22484 );
and \U$30165 ( \30480 , \22167 , \22482 );
nor \U$30166 ( \30481 , \30479 , \30480 );
xnor \U$30167 ( \30482 , \30481 , \22494 );
and \U$30168 ( \30483 , \22181 , \22506 );
and \U$30169 ( \30484 , \22192 , \22504 );
nor \U$30170 ( \30485 , \30483 , \30484 );
xnor \U$30171 ( \30486 , \30485 , \22516 );
xor \U$30172 ( \30487 , \30482 , \30486 );
and \U$30173 ( \30488 , \22202 , \22530 );
and \U$30174 ( \30489 , \22213 , \22528 );
nor \U$30175 ( \30490 , \30488 , \30489 );
xnor \U$30176 ( \30491 , \30490 , \22540 );
xor \U$30177 ( \30492 , \30487 , \30491 );
and \U$30178 ( \30493 , \22089 , \22413 );
and \U$30179 ( \30494 , \22100 , \22411 );
nor \U$30180 ( \30495 , \30493 , \30494 );
xnor \U$30181 ( \30496 , \30495 , \22423 );
and \U$30182 ( \30497 , \22113 , \22435 );
and \U$30183 ( \30498 , \22124 , \22433 );
nor \U$30184 ( \30499 , \30497 , \30498 );
xnor \U$30185 ( \30500 , \30499 , \22445 );
xor \U$30186 ( \30501 , \30496 , \30500 );
and \U$30187 ( \30502 , \22134 , \22463 );
and \U$30188 ( \30503 , \22145 , \22461 );
nor \U$30189 ( \30504 , \30502 , \30503 );
xnor \U$30190 ( \30505 , \30504 , \22473 );
xor \U$30191 ( \30506 , \30501 , \30505 );
xor \U$30192 ( \30507 , \30492 , \30506 );
and \U$30193 ( \30508 , \23230 , \22345 );
and \U$30194 ( \30509 , \23329 , \22343 );
nor \U$30195 ( \30510 , \30508 , \30509 );
xnor \U$30196 ( \30511 , \30510 , \22355 );
and \U$30197 ( \30512 , \22858 , \22367 );
and \U$30198 ( \30513 , \22894 , \22365 );
nor \U$30199 ( \30514 , \30512 , \30513 );
xnor \U$30200 ( \30515 , \30514 , \22377 );
xor \U$30201 ( \30516 , \30511 , \30515 );
and \U$30202 ( \30517 , \22071 , \22392 );
and \U$30203 ( \30518 , \22081 , \22390 );
nor \U$30204 ( \30519 , \30517 , \30518 );
xnor \U$30205 ( \30520 , \30519 , \22402 );
xor \U$30206 ( \30521 , \30516 , \30520 );
xor \U$30207 ( \30522 , \30507 , \30521 );
xor \U$30208 ( \30523 , \30478 , \30522 );
and \U$30209 ( \30524 , \22361 , \22691 );
and \U$30210 ( \30525 , \22372 , \22689 );
nor \U$30211 ( \30526 , \30524 , \30525 );
xnor \U$30212 ( \30527 , \30526 , \22701 );
and \U$30213 ( \30528 , \22386 , \22720 );
and \U$30214 ( \30529 , \22397 , \22707 );
nor \U$30215 ( \30530 , \30528 , \30529 );
xnor \U$30216 ( \30531 , \30530 , \22067 );
xor \U$30217 ( \30532 , \30527 , \30531 );
and \U$30218 ( \30533 , \22407 , \23173 );
and \U$30219 ( \30534 , \22418 , \22999 );
nor \U$30220 ( \30535 , \30533 , \30534 );
xnor \U$30221 ( \30536 , \30535 , \22016 );
xor \U$30222 ( \30537 , \30532 , \30536 );
and \U$30223 ( \30538 , \22294 , \22619 );
and \U$30224 ( \30539 , \22305 , \22617 );
nor \U$30225 ( \30540 , \30538 , \30539 );
xnor \U$30226 ( \30541 , \30540 , \22629 );
and \U$30227 ( \30542 , \22318 , \22641 );
and \U$30228 ( \30543 , \22329 , \22639 );
nor \U$30229 ( \30544 , \30542 , \30543 );
xnor \U$30230 ( \30545 , \30544 , \22651 );
xor \U$30231 ( \30546 , \30541 , \30545 );
and \U$30232 ( \30547 , \22339 , \22671 );
and \U$30233 ( \30548 , \22350 , \22669 );
nor \U$30234 ( \30549 , \30547 , \30548 );
xnor \U$30235 ( \30550 , \30549 , \22681 );
xor \U$30236 ( \30551 , \30546 , \30550 );
xor \U$30237 ( \30552 , \30537 , \30551 );
and \U$30238 ( \30553 , \22224 , \22551 );
and \U$30239 ( \30554 , \22235 , \22549 );
nor \U$30240 ( \30555 , \30553 , \30554 );
xnor \U$30241 ( \30556 , \30555 , \22561 );
and \U$30242 ( \30557 , \22251 , \22573 );
and \U$30243 ( \30558 , \22262 , \22571 );
nor \U$30244 ( \30559 , \30557 , \30558 );
xnor \U$30245 ( \30560 , \30559 , \22583 );
xor \U$30246 ( \30561 , \30556 , \30560 );
and \U$30247 ( \30562 , \22272 , \22598 );
and \U$30248 ( \30563 , \22283 , \22596 );
nor \U$30249 ( \30564 , \30562 , \30563 );
xnor \U$30250 ( \30565 , \30564 , \22608 );
xor \U$30251 ( \30566 , \30561 , \30565 );
xor \U$30252 ( \30567 , \30552 , \30566 );
xor \U$30253 ( \30568 , \30523 , \30567 );
xor \U$30254 ( \30569 , \30467 , \30568 );
xor \U$30255 ( \30570 , \30411 , \30569 );
and \U$30256 ( \30571 , \30167 , \30171 );
and \U$30257 ( \30572 , \30171 , \30176 );
and \U$30258 ( \30573 , \30167 , \30176 );
or \U$30259 ( \30574 , \30571 , \30572 , \30573 );
and \U$30260 ( \30575 , \30153 , \30157 );
and \U$30261 ( \30576 , \30157 , \30162 );
and \U$30262 ( \30577 , \30153 , \30162 );
or \U$30263 ( \30578 , \30575 , \30576 , \30577 );
xor \U$30264 ( \30579 , \30574 , \30578 );
and \U$30265 ( \30580 , \30250 , \30294 );
and \U$30266 ( \30581 , \30294 , \30336 );
and \U$30267 ( \30582 , \30250 , \30336 );
or \U$30268 ( \30583 , \30580 , \30581 , \30582 );
xor \U$30269 ( \30584 , \30579 , \30583 );
xor \U$30270 ( \30585 , \30570 , \30584 );
xor \U$30271 ( \30586 , \30388 , \30585 );
xor \U$30272 ( \30587 , \30379 , \30586 );
xor \U$30273 ( \30588 , \30363 , \30587 );
and \U$30274 ( \30589 , \30124 , \30356 );
nor \U$30275 ( \30590 , \30588 , \30589 );
nor \U$30276 ( \30591 , \30359 , \30590 );
and \U$30277 ( \30592 , \30367 , \30378 );
and \U$30278 ( \30593 , \30378 , \30586 );
and \U$30279 ( \30594 , \30367 , \30586 );
or \U$30280 ( \30595 , \30592 , \30593 , \30594 );
and \U$30281 ( \30596 , \30383 , \30387 );
and \U$30282 ( \30597 , \30387 , \30585 );
and \U$30283 ( \30598 , \30383 , \30585 );
or \U$30284 ( \30599 , \30596 , \30597 , \30598 );
and \U$30285 ( \30600 , \30574 , \30578 );
and \U$30286 ( \30601 , \30578 , \30583 );
and \U$30287 ( \30602 , \30574 , \30583 );
or \U$30288 ( \30603 , \30600 , \30601 , \30602 );
and \U$30289 ( \30604 , \30415 , \30466 );
and \U$30290 ( \30605 , \30466 , \30568 );
and \U$30291 ( \30606 , \30415 , \30568 );
or \U$30292 ( \30607 , \30604 , \30605 , \30606 );
xor \U$30293 ( \30608 , \30603 , \30607 );
and \U$30294 ( \30609 , \30399 , \30410 );
xor \U$30295 ( \30610 , \30608 , \30609 );
xor \U$30296 ( \30611 , \30599 , \30610 );
and \U$30297 ( \30612 , \30371 , \30375 );
and \U$30298 ( \30613 , \30375 , \30377 );
and \U$30299 ( \30614 , \30371 , \30377 );
or \U$30300 ( \30615 , \30612 , \30613 , \30614 );
and \U$30301 ( \30616 , \30411 , \30569 );
and \U$30302 ( \30617 , \30569 , \30584 );
and \U$30303 ( \30618 , \30411 , \30584 );
or \U$30304 ( \30619 , \30616 , \30617 , \30618 );
xor \U$30305 ( \30620 , \30615 , \30619 );
and \U$30306 ( \30621 , \22192 , \22506 );
and \U$30307 ( \30622 , \22156 , \22504 );
nor \U$30308 ( \30623 , \30621 , \30622 );
xnor \U$30309 ( \30624 , \30623 , \22516 );
and \U$30310 ( \30625 , \22213 , \22530 );
and \U$30311 ( \30626 , \22181 , \22528 );
nor \U$30312 ( \30627 , \30625 , \30626 );
xnor \U$30313 ( \30628 , \30627 , \22540 );
xor \U$30314 ( \30629 , \30624 , \30628 );
and \U$30315 ( \30630 , \22235 , \22551 );
and \U$30316 ( \30631 , \22202 , \22549 );
nor \U$30317 ( \30632 , \30630 , \30631 );
xnor \U$30318 ( \30633 , \30632 , \22561 );
xor \U$30319 ( \30634 , \30629 , \30633 );
and \U$30320 ( \30635 , \22124 , \22435 );
and \U$30321 ( \30636 , \22089 , \22433 );
nor \U$30322 ( \30637 , \30635 , \30636 );
xnor \U$30323 ( \30638 , \30637 , \22445 );
and \U$30324 ( \30639 , \22145 , \22463 );
and \U$30325 ( \30640 , \22113 , \22461 );
nor \U$30326 ( \30641 , \30639 , \30640 );
xnor \U$30327 ( \30642 , \30641 , \22473 );
xor \U$30328 ( \30643 , \30638 , \30642 );
and \U$30329 ( \30644 , \22167 , \22484 );
and \U$30330 ( \30645 , \22134 , \22482 );
nor \U$30331 ( \30646 , \30644 , \30645 );
xnor \U$30332 ( \30647 , \30646 , \22494 );
xor \U$30333 ( \30648 , \30643 , \30647 );
xor \U$30334 ( \30649 , \30634 , \30648 );
and \U$30335 ( \30650 , \22894 , \22367 );
and \U$30336 ( \30651 , \23230 , \22365 );
nor \U$30337 ( \30652 , \30650 , \30651 );
xnor \U$30338 ( \30653 , \30652 , \22377 );
and \U$30339 ( \30654 , \22081 , \22392 );
and \U$30340 ( \30655 , \22858 , \22390 );
nor \U$30341 ( \30656 , \30654 , \30655 );
xnor \U$30342 ( \30657 , \30656 , \22402 );
xor \U$30343 ( \30658 , \30653 , \30657 );
and \U$30344 ( \30659 , \22100 , \22413 );
and \U$30345 ( \30660 , \22071 , \22411 );
nor \U$30346 ( \30661 , \30659 , \30660 );
xnor \U$30347 ( \30662 , \30661 , \22423 );
xor \U$30348 ( \30663 , \30658 , \30662 );
xor \U$30349 ( \30664 , \30649 , \30663 );
and \U$30350 ( \30665 , \22397 , \22720 );
and \U$30351 ( \30666 , \22361 , \22707 );
nor \U$30352 ( \30667 , \30665 , \30666 );
xnor \U$30353 ( \30668 , \30667 , \22067 );
and \U$30354 ( \30669 , \22418 , \23173 );
and \U$30355 ( \30670 , \22386 , \22999 );
nor \U$30356 ( \30671 , \30669 , \30670 );
xnor \U$30357 ( \30672 , \30671 , \22016 );
xor \U$30358 ( \30673 , \30668 , \30672 );
and \U$30359 ( \30674 , \22440 , \22021 );
and \U$30360 ( \30675 , \22407 , \22019 );
nor \U$30361 ( \30676 , \30674 , \30675 );
xnor \U$30362 ( \30677 , \30676 , \21595 );
xor \U$30363 ( \30678 , \30673 , \30677 );
and \U$30364 ( \30679 , \22329 , \22641 );
and \U$30365 ( \30680 , \22294 , \22639 );
nor \U$30366 ( \30681 , \30679 , \30680 );
xnor \U$30367 ( \30682 , \30681 , \22651 );
and \U$30368 ( \30683 , \22350 , \22671 );
and \U$30369 ( \30684 , \22318 , \22669 );
nor \U$30370 ( \30685 , \30683 , \30684 );
xnor \U$30371 ( \30686 , \30685 , \22681 );
xor \U$30372 ( \30687 , \30682 , \30686 );
and \U$30373 ( \30688 , \22372 , \22691 );
and \U$30374 ( \30689 , \22339 , \22689 );
nor \U$30375 ( \30690 , \30688 , \30689 );
xnor \U$30376 ( \30691 , \30690 , \22701 );
xor \U$30377 ( \30692 , \30687 , \30691 );
xor \U$30378 ( \30693 , \30678 , \30692 );
and \U$30379 ( \30694 , \22262 , \22573 );
and \U$30380 ( \30695 , \22224 , \22571 );
nor \U$30381 ( \30696 , \30694 , \30695 );
xnor \U$30382 ( \30697 , \30696 , \22583 );
and \U$30383 ( \30698 , \22283 , \22598 );
and \U$30384 ( \30699 , \22251 , \22596 );
nor \U$30385 ( \30700 , \30698 , \30699 );
xnor \U$30386 ( \30701 , \30700 , \22608 );
xor \U$30387 ( \30702 , \30697 , \30701 );
and \U$30388 ( \30703 , \22305 , \22619 );
and \U$30389 ( \30704 , \22272 , \22617 );
nor \U$30390 ( \30705 , \30703 , \30704 );
xnor \U$30391 ( \30706 , \30705 , \22629 );
xor \U$30392 ( \30707 , \30702 , \30706 );
xor \U$30393 ( \30708 , \30693 , \30707 );
xor \U$30394 ( \30709 , \30664 , \30708 );
and \U$30395 ( \30710 , \30527 , \30531 );
and \U$30396 ( \30711 , \30531 , \30536 );
and \U$30397 ( \30712 , \30527 , \30536 );
or \U$30398 ( \30713 , \30710 , \30711 , \30712 );
and \U$30399 ( \30714 , \30428 , \30432 );
and \U$30400 ( \30715 , \30432 , \30434 );
and \U$30401 ( \30716 , \30428 , \30434 );
or \U$30402 ( \30717 , \30714 , \30715 , \30716 );
xor \U$30403 ( \30718 , \30713 , \30717 );
and \U$30404 ( \30719 , \22468 , \21983 );
and \U$30405 ( \30720 , \22429 , \21981 );
nor \U$30406 ( \30721 , \30719 , \30720 );
xnor \U$30407 ( \30722 , \30721 , \21995 );
and \U$30408 ( \30723 , \22457 , \21978 );
xnor \U$30409 ( \30724 , \30722 , \30723 );
xor \U$30410 ( \30725 , \30718 , \30724 );
xor \U$30411 ( \30726 , \30709 , \30725 );
and \U$30412 ( \30727 , \30537 , \30551 );
and \U$30413 ( \30728 , \30551 , \30566 );
and \U$30414 ( \30729 , \30537 , \30566 );
or \U$30415 ( \30730 , \30727 , \30728 , \30729 );
and \U$30416 ( \30731 , \30492 , \30506 );
and \U$30417 ( \30732 , \30506 , \30521 );
and \U$30418 ( \30733 , \30492 , \30521 );
or \U$30419 ( \30734 , \30731 , \30732 , \30733 );
xor \U$30420 ( \30735 , \30730 , \30734 );
and \U$30421 ( \30736 , \21990 , \22300 );
not \U$30422 ( \30737 , \30736 );
xnor \U$30423 ( \30738 , \30737 , \22310 );
and \U$30424 ( \30739 , \22001 , \22324 );
and \U$30425 ( \30740 , \21977 , \22322 );
nor \U$30426 ( \30741 , \30739 , \30740 );
xnor \U$30427 ( \30742 , \30741 , \22334 );
xor \U$30428 ( \30743 , \30738 , \30742 );
and \U$30429 ( \30744 , \23329 , \22345 );
and \U$30430 ( \30745 , \22030 , \22343 );
nor \U$30431 ( \30746 , \30744 , \30745 );
xnor \U$30432 ( \30747 , \30746 , \22355 );
xor \U$30433 ( \30748 , \30743 , \30747 );
xor \U$30434 ( \30749 , \30735 , \30748 );
xor \U$30435 ( \30750 , \30726 , \30749 );
and \U$30436 ( \30751 , \30455 , \30459 );
and \U$30437 ( \30752 , \30459 , \30464 );
and \U$30438 ( \30753 , \30455 , \30464 );
or \U$30439 ( \30754 , \30751 , \30752 , \30753 );
and \U$30440 ( \30755 , \30440 , \30444 );
and \U$30441 ( \30756 , \30444 , \30449 );
and \U$30442 ( \30757 , \30440 , \30449 );
or \U$30443 ( \30758 , \30755 , \30756 , \30757 );
xor \U$30444 ( \30759 , \30754 , \30758 );
and \U$30445 ( \30760 , \30419 , \30423 );
and \U$30446 ( \30761 , \30423 , \30435 );
and \U$30447 ( \30762 , \30419 , \30435 );
or \U$30448 ( \30763 , \30760 , \30761 , \30762 );
xor \U$30449 ( \30764 , \30759 , \30763 );
xor \U$30450 ( \30765 , \30750 , \30764 );
and \U$30451 ( \30766 , \30436 , \30450 );
and \U$30452 ( \30767 , \30450 , \30465 );
and \U$30453 ( \30768 , \30436 , \30465 );
or \U$30454 ( \30769 , \30766 , \30767 , \30768 );
and \U$30455 ( \30770 , \30482 , \30486 );
and \U$30456 ( \30771 , \30486 , \30491 );
and \U$30457 ( \30772 , \30482 , \30491 );
or \U$30458 ( \30773 , \30770 , \30771 , \30772 );
and \U$30459 ( \30774 , \30556 , \30560 );
and \U$30460 ( \30775 , \30560 , \30565 );
and \U$30461 ( \30776 , \30556 , \30565 );
or \U$30462 ( \30777 , \30774 , \30775 , \30776 );
xor \U$30463 ( \30778 , \30773 , \30777 );
and \U$30464 ( \30779 , \30541 , \30545 );
and \U$30465 ( \30780 , \30545 , \30550 );
and \U$30466 ( \30781 , \30541 , \30550 );
or \U$30467 ( \30782 , \30779 , \30780 , \30781 );
xor \U$30468 ( \30783 , \30778 , \30782 );
xor \U$30469 ( \30784 , \30769 , \30783 );
and \U$30470 ( \30785 , \30468 , \30472 );
and \U$30471 ( \30786 , \30472 , \30477 );
and \U$30472 ( \30787 , \30468 , \30477 );
or \U$30473 ( \30788 , \30785 , \30786 , \30787 );
and \U$30474 ( \30789 , \30511 , \30515 );
and \U$30475 ( \30790 , \30515 , \30520 );
and \U$30476 ( \30791 , \30511 , \30520 );
or \U$30477 ( \30792 , \30789 , \30790 , \30791 );
xor \U$30478 ( \30793 , \30788 , \30792 );
and \U$30479 ( \30794 , \30496 , \30500 );
and \U$30480 ( \30795 , \30500 , \30505 );
and \U$30481 ( \30796 , \30496 , \30505 );
or \U$30482 ( \30797 , \30794 , \30795 , \30796 );
xor \U$30483 ( \30798 , \30793 , \30797 );
xor \U$30484 ( \30799 , \30784 , \30798 );
xor \U$30485 ( \30800 , \30765 , \30799 );
and \U$30486 ( \30801 , \30403 , \30407 );
and \U$30487 ( \30802 , \30407 , \30409 );
and \U$30488 ( \30803 , \30403 , \30409 );
or \U$30489 ( \30804 , \30801 , \30802 , \30803 );
and \U$30490 ( \30805 , \30392 , \30396 );
and \U$30491 ( \30806 , \30396 , \30398 );
and \U$30492 ( \30807 , \30392 , \30398 );
or \U$30493 ( \30808 , \30805 , \30806 , \30807 );
xor \U$30494 ( \30809 , \30804 , \30808 );
and \U$30495 ( \30810 , \30478 , \30522 );
and \U$30496 ( \30811 , \30522 , \30567 );
and \U$30497 ( \30812 , \30478 , \30567 );
or \U$30498 ( \30813 , \30810 , \30811 , \30812 );
xor \U$30499 ( \30814 , \30809 , \30813 );
xor \U$30500 ( \30815 , \30800 , \30814 );
xor \U$30501 ( \30816 , \30620 , \30815 );
xor \U$30502 ( \30817 , \30611 , \30816 );
xor \U$30503 ( \30818 , \30595 , \30817 );
and \U$30504 ( \30819 , \30363 , \30587 );
nor \U$30505 ( \30820 , \30818 , \30819 );
and \U$30506 ( \30821 , \30599 , \30610 );
and \U$30507 ( \30822 , \30610 , \30816 );
and \U$30508 ( \30823 , \30599 , \30816 );
or \U$30509 ( \30824 , \30821 , \30822 , \30823 );
and \U$30510 ( \30825 , \30615 , \30619 );
and \U$30511 ( \30826 , \30619 , \30815 );
and \U$30512 ( \30827 , \30615 , \30815 );
or \U$30513 ( \30828 , \30825 , \30826 , \30827 );
and \U$30514 ( \30829 , \30804 , \30808 );
and \U$30515 ( \30830 , \30808 , \30813 );
and \U$30516 ( \30831 , \30804 , \30813 );
or \U$30517 ( \30832 , \30829 , \30830 , \30831 );
and \U$30518 ( \30833 , \30769 , \30783 );
and \U$30519 ( \30834 , \30783 , \30798 );
and \U$30520 ( \30835 , \30769 , \30798 );
or \U$30521 ( \30836 , \30833 , \30834 , \30835 );
xor \U$30522 ( \30837 , \30832 , \30836 );
and \U$30523 ( \30838 , \30726 , \30749 );
and \U$30524 ( \30839 , \30749 , \30764 );
and \U$30525 ( \30840 , \30726 , \30764 );
or \U$30526 ( \30841 , \30838 , \30839 , \30840 );
xor \U$30527 ( \30842 , \30837 , \30841 );
xor \U$30528 ( \30843 , \30828 , \30842 );
and \U$30529 ( \30844 , \30603 , \30607 );
and \U$30530 ( \30845 , \30607 , \30609 );
and \U$30531 ( \30846 , \30603 , \30609 );
or \U$30532 ( \30847 , \30844 , \30845 , \30846 );
and \U$30533 ( \30848 , \30765 , \30799 );
and \U$30534 ( \30849 , \30799 , \30814 );
and \U$30535 ( \30850 , \30765 , \30814 );
or \U$30536 ( \30851 , \30848 , \30849 , \30850 );
xor \U$30537 ( \30852 , \30847 , \30851 );
and \U$30538 ( \30853 , \30788 , \30792 );
and \U$30539 ( \30854 , \30792 , \30797 );
and \U$30540 ( \30855 , \30788 , \30797 );
or \U$30541 ( \30856 , \30853 , \30854 , \30855 );
and \U$30542 ( \30857 , \30773 , \30777 );
and \U$30543 ( \30858 , \30777 , \30782 );
and \U$30544 ( \30859 , \30773 , \30782 );
or \U$30545 ( \30860 , \30857 , \30858 , \30859 );
xor \U$30546 ( \30861 , \30856 , \30860 );
and \U$30547 ( \30862 , \30713 , \30717 );
and \U$30548 ( \30863 , \30717 , \30724 );
and \U$30549 ( \30864 , \30713 , \30724 );
or \U$30550 ( \30865 , \30862 , \30863 , \30864 );
xor \U$30551 ( \30866 , \30861 , \30865 );
and \U$30552 ( \30867 , \30668 , \30672 );
and \U$30553 ( \30868 , \30672 , \30677 );
and \U$30554 ( \30869 , \30668 , \30677 );
or \U$30555 ( \30870 , \30867 , \30868 , \30869 );
or \U$30556 ( \30871 , \30722 , \30723 );
xor \U$30557 ( \30872 , \30870 , \30871 );
and \U$30558 ( \30873 , \22429 , \21983 );
and \U$30559 ( \30874 , \22440 , \21981 );
nor \U$30560 ( \30875 , \30873 , \30874 );
xnor \U$30561 ( \30876 , \30875 , \21995 );
xor \U$30562 ( \30877 , \30872 , \30876 );
and \U$30563 ( \30878 , \30624 , \30628 );
and \U$30564 ( \30879 , \30628 , \30633 );
and \U$30565 ( \30880 , \30624 , \30633 );
or \U$30566 ( \30881 , \30878 , \30879 , \30880 );
and \U$30567 ( \30882 , \30697 , \30701 );
and \U$30568 ( \30883 , \30701 , \30706 );
and \U$30569 ( \30884 , \30697 , \30706 );
or \U$30570 ( \30885 , \30882 , \30883 , \30884 );
xor \U$30571 ( \30886 , \30881 , \30885 );
and \U$30572 ( \30887 , \30682 , \30686 );
and \U$30573 ( \30888 , \30686 , \30691 );
and \U$30574 ( \30889 , \30682 , \30691 );
or \U$30575 ( \30890 , \30887 , \30888 , \30889 );
xor \U$30576 ( \30891 , \30886 , \30890 );
xor \U$30577 ( \30892 , \30877 , \30891 );
and \U$30578 ( \30893 , \30738 , \30742 );
and \U$30579 ( \30894 , \30742 , \30747 );
and \U$30580 ( \30895 , \30738 , \30747 );
or \U$30581 ( \30896 , \30893 , \30894 , \30895 );
and \U$30582 ( \30897 , \30653 , \30657 );
and \U$30583 ( \30898 , \30657 , \30662 );
and \U$30584 ( \30899 , \30653 , \30662 );
or \U$30585 ( \30900 , \30897 , \30898 , \30899 );
xor \U$30586 ( \30901 , \30896 , \30900 );
and \U$30587 ( \30902 , \30638 , \30642 );
and \U$30588 ( \30903 , \30642 , \30647 );
and \U$30589 ( \30904 , \30638 , \30647 );
or \U$30590 ( \30905 , \30902 , \30903 , \30904 );
xor \U$30591 ( \30906 , \30901 , \30905 );
xor \U$30592 ( \30907 , \30892 , \30906 );
not \U$30593 ( \30908 , \22310 );
and \U$30594 ( \30909 , \21977 , \22324 );
and \U$30595 ( \30910 , \21990 , \22322 );
nor \U$30596 ( \30911 , \30909 , \30910 );
xnor \U$30597 ( \30912 , \30911 , \22334 );
xor \U$30598 ( \30913 , \30908 , \30912 );
and \U$30599 ( \30914 , \22030 , \22345 );
and \U$30600 ( \30915 , \22001 , \22343 );
nor \U$30601 ( \30916 , \30914 , \30915 );
xnor \U$30602 ( \30917 , \30916 , \22355 );
xor \U$30603 ( \30918 , \30913 , \30917 );
and \U$30604 ( \30919 , \22224 , \22573 );
and \U$30605 ( \30920 , \22235 , \22571 );
nor \U$30606 ( \30921 , \30919 , \30920 );
xnor \U$30607 ( \30922 , \30921 , \22583 );
and \U$30608 ( \30923 , \22251 , \22598 );
and \U$30609 ( \30924 , \22262 , \22596 );
nor \U$30610 ( \30925 , \30923 , \30924 );
xnor \U$30611 ( \30926 , \30925 , \22608 );
xor \U$30612 ( \30927 , \30922 , \30926 );
and \U$30613 ( \30928 , \22272 , \22619 );
and \U$30614 ( \30929 , \22283 , \22617 );
nor \U$30615 ( \30930 , \30928 , \30929 );
xnor \U$30616 ( \30931 , \30930 , \22629 );
xor \U$30617 ( \30932 , \30927 , \30931 );
and \U$30618 ( \30933 , \22156 , \22506 );
and \U$30619 ( \30934 , \22167 , \22504 );
nor \U$30620 ( \30935 , \30933 , \30934 );
xnor \U$30621 ( \30936 , \30935 , \22516 );
and \U$30622 ( \30937 , \22181 , \22530 );
and \U$30623 ( \30938 , \22192 , \22528 );
nor \U$30624 ( \30939 , \30937 , \30938 );
xnor \U$30625 ( \30940 , \30939 , \22540 );
xor \U$30626 ( \30941 , \30936 , \30940 );
and \U$30627 ( \30942 , \22202 , \22551 );
and \U$30628 ( \30943 , \22213 , \22549 );
nor \U$30629 ( \30944 , \30942 , \30943 );
xnor \U$30630 ( \30945 , \30944 , \22561 );
xor \U$30631 ( \30946 , \30941 , \30945 );
xor \U$30632 ( \30947 , \30932 , \30946 );
and \U$30633 ( \30948 , \22089 , \22435 );
and \U$30634 ( \30949 , \22100 , \22433 );
nor \U$30635 ( \30950 , \30948 , \30949 );
xnor \U$30636 ( \30951 , \30950 , \22445 );
and \U$30637 ( \30952 , \22113 , \22463 );
and \U$30638 ( \30953 , \22124 , \22461 );
nor \U$30639 ( \30954 , \30952 , \30953 );
xnor \U$30640 ( \30955 , \30954 , \22473 );
xor \U$30641 ( \30956 , \30951 , \30955 );
and \U$30642 ( \30957 , \22134 , \22484 );
and \U$30643 ( \30958 , \22145 , \22482 );
nor \U$30644 ( \30959 , \30957 , \30958 );
xnor \U$30645 ( \30960 , \30959 , \22494 );
xor \U$30646 ( \30961 , \30956 , \30960 );
xor \U$30647 ( \30962 , \30947 , \30961 );
xor \U$30648 ( \30963 , \30918 , \30962 );
and \U$30649 ( \30964 , \22468 , \21978 );
and \U$30650 ( \30965 , \22361 , \22720 );
and \U$30651 ( \30966 , \22372 , \22707 );
nor \U$30652 ( \30967 , \30965 , \30966 );
xnor \U$30653 ( \30968 , \30967 , \22067 );
and \U$30654 ( \30969 , \22386 , \23173 );
and \U$30655 ( \30970 , \22397 , \22999 );
nor \U$30656 ( \30971 , \30969 , \30970 );
xnor \U$30657 ( \30972 , \30971 , \22016 );
xor \U$30658 ( \30973 , \30968 , \30972 );
and \U$30659 ( \30974 , \22407 , \22021 );
and \U$30660 ( \30975 , \22418 , \22019 );
nor \U$30661 ( \30976 , \30974 , \30975 );
xnor \U$30662 ( \30977 , \30976 , \21595 );
xor \U$30663 ( \30978 , \30973 , \30977 );
xor \U$30664 ( \30979 , \30964 , \30978 );
and \U$30665 ( \30980 , \22294 , \22641 );
and \U$30666 ( \30981 , \22305 , \22639 );
nor \U$30667 ( \30982 , \30980 , \30981 );
xnor \U$30668 ( \30983 , \30982 , \22651 );
and \U$30669 ( \30984 , \22318 , \22671 );
and \U$30670 ( \30985 , \22329 , \22669 );
nor \U$30671 ( \30986 , \30984 , \30985 );
xnor \U$30672 ( \30987 , \30986 , \22681 );
xor \U$30673 ( \30988 , \30983 , \30987 );
and \U$30674 ( \30989 , \22339 , \22691 );
and \U$30675 ( \30990 , \22350 , \22689 );
nor \U$30676 ( \30991 , \30989 , \30990 );
xnor \U$30677 ( \30992 , \30991 , \22701 );
xor \U$30678 ( \30993 , \30988 , \30992 );
xor \U$30679 ( \30994 , \30979 , \30993 );
xor \U$30680 ( \30995 , \30963 , \30994 );
xor \U$30681 ( \30996 , \30907 , \30995 );
and \U$30682 ( \30997 , \30678 , \30692 );
and \U$30683 ( \30998 , \30692 , \30707 );
and \U$30684 ( \30999 , \30678 , \30707 );
or \U$30685 ( \31000 , \30997 , \30998 , \30999 );
and \U$30686 ( \31001 , \30634 , \30648 );
and \U$30687 ( \31002 , \30648 , \30663 );
and \U$30688 ( \31003 , \30634 , \30663 );
or \U$30689 ( \31004 , \31001 , \31002 , \31003 );
xor \U$30690 ( \31005 , \31000 , \31004 );
and \U$30691 ( \31006 , \23230 , \22367 );
and \U$30692 ( \31007 , \23329 , \22365 );
nor \U$30693 ( \31008 , \31006 , \31007 );
xnor \U$30694 ( \31009 , \31008 , \22377 );
and \U$30695 ( \31010 , \22858 , \22392 );
and \U$30696 ( \31011 , \22894 , \22390 );
nor \U$30697 ( \31012 , \31010 , \31011 );
xnor \U$30698 ( \31013 , \31012 , \22402 );
xor \U$30699 ( \31014 , \31009 , \31013 );
and \U$30700 ( \31015 , \22071 , \22413 );
and \U$30701 ( \31016 , \22081 , \22411 );
nor \U$30702 ( \31017 , \31015 , \31016 );
xnor \U$30703 ( \31018 , \31017 , \22423 );
xor \U$30704 ( \31019 , \31014 , \31018 );
xor \U$30705 ( \31020 , \31005 , \31019 );
xor \U$30706 ( \31021 , \30996 , \31020 );
xor \U$30707 ( \31022 , \30866 , \31021 );
and \U$30708 ( \31023 , \30754 , \30758 );
and \U$30709 ( \31024 , \30758 , \30763 );
and \U$30710 ( \31025 , \30754 , \30763 );
or \U$30711 ( \31026 , \31023 , \31024 , \31025 );
and \U$30712 ( \31027 , \30730 , \30734 );
and \U$30713 ( \31028 , \30734 , \30748 );
and \U$30714 ( \31029 , \30730 , \30748 );
or \U$30715 ( \31030 , \31027 , \31028 , \31029 );
xor \U$30716 ( \31031 , \31026 , \31030 );
and \U$30717 ( \31032 , \30664 , \30708 );
and \U$30718 ( \31033 , \30708 , \30725 );
and \U$30719 ( \31034 , \30664 , \30725 );
or \U$30720 ( \31035 , \31032 , \31033 , \31034 );
xor \U$30721 ( \31036 , \31031 , \31035 );
xor \U$30722 ( \31037 , \31022 , \31036 );
xor \U$30723 ( \31038 , \30852 , \31037 );
xor \U$30724 ( \31039 , \30843 , \31038 );
xor \U$30725 ( \31040 , \30824 , \31039 );
and \U$30726 ( \31041 , \30595 , \30817 );
nor \U$30727 ( \31042 , \31040 , \31041 );
nor \U$30728 ( \31043 , \30820 , \31042 );
nand \U$30729 ( \31044 , \30591 , \31043 );
nor \U$30730 ( \31045 , \30120 , \31044 );
and \U$30731 ( \31046 , \30828 , \30842 );
and \U$30732 ( \31047 , \30842 , \31038 );
and \U$30733 ( \31048 , \30828 , \31038 );
or \U$30734 ( \31049 , \31046 , \31047 , \31048 );
and \U$30735 ( \31050 , \30847 , \30851 );
and \U$30736 ( \31051 , \30851 , \31037 );
and \U$30737 ( \31052 , \30847 , \31037 );
or \U$30738 ( \31053 , \31050 , \31051 , \31052 );
and \U$30739 ( \31054 , \31026 , \31030 );
and \U$30740 ( \31055 , \31030 , \31035 );
and \U$30741 ( \31056 , \31026 , \31035 );
or \U$30742 ( \31057 , \31054 , \31055 , \31056 );
and \U$30743 ( \31058 , \30907 , \30995 );
and \U$30744 ( \31059 , \30995 , \31020 );
and \U$30745 ( \31060 , \30907 , \31020 );
or \U$30746 ( \31061 , \31058 , \31059 , \31060 );
xor \U$30747 ( \31062 , \31057 , \31061 );
and \U$30748 ( \31063 , \30964 , \30978 );
and \U$30749 ( \31064 , \30978 , \30993 );
and \U$30750 ( \31065 , \30964 , \30993 );
or \U$30751 ( \31066 , \31063 , \31064 , \31065 );
and \U$30752 ( \31067 , \30932 , \30946 );
and \U$30753 ( \31068 , \30946 , \30961 );
and \U$30754 ( \31069 , \30932 , \30961 );
or \U$30755 ( \31070 , \31067 , \31068 , \31069 );
xor \U$30756 ( \31071 , \31066 , \31070 );
and \U$30757 ( \31072 , \22124 , \22463 );
and \U$30758 ( \31073 , \22089 , \22461 );
nor \U$30759 ( \31074 , \31072 , \31073 );
xnor \U$30760 ( \31075 , \31074 , \22473 );
and \U$30761 ( \31076 , \22145 , \22484 );
and \U$30762 ( \31077 , \22113 , \22482 );
nor \U$30763 ( \31078 , \31076 , \31077 );
xnor \U$30764 ( \31079 , \31078 , \22494 );
xor \U$30765 ( \31080 , \31075 , \31079 );
and \U$30766 ( \31081 , \22167 , \22506 );
and \U$30767 ( \31082 , \22134 , \22504 );
nor \U$30768 ( \31083 , \31081 , \31082 );
xnor \U$30769 ( \31084 , \31083 , \22516 );
xor \U$30770 ( \31085 , \31080 , \31084 );
and \U$30771 ( \31086 , \22894 , \22392 );
and \U$30772 ( \31087 , \23230 , \22390 );
nor \U$30773 ( \31088 , \31086 , \31087 );
xnor \U$30774 ( \31089 , \31088 , \22402 );
and \U$30775 ( \31090 , \22081 , \22413 );
and \U$30776 ( \31091 , \22858 , \22411 );
nor \U$30777 ( \31092 , \31090 , \31091 );
xnor \U$30778 ( \31093 , \31092 , \22423 );
xor \U$30779 ( \31094 , \31089 , \31093 );
and \U$30780 ( \31095 , \22100 , \22435 );
and \U$30781 ( \31096 , \22071 , \22433 );
nor \U$30782 ( \31097 , \31095 , \31096 );
xnor \U$30783 ( \31098 , \31097 , \22445 );
xor \U$30784 ( \31099 , \31094 , \31098 );
xor \U$30785 ( \31100 , \31085 , \31099 );
and \U$30786 ( \31101 , \21990 , \22324 );
not \U$30787 ( \31102 , \31101 );
xnor \U$30788 ( \31103 , \31102 , \22334 );
and \U$30789 ( \31104 , \22001 , \22345 );
and \U$30790 ( \31105 , \21977 , \22343 );
nor \U$30791 ( \31106 , \31104 , \31105 );
xnor \U$30792 ( \31107 , \31106 , \22355 );
xor \U$30793 ( \31108 , \31103 , \31107 );
and \U$30794 ( \31109 , \23329 , \22367 );
and \U$30795 ( \31110 , \22030 , \22365 );
nor \U$30796 ( \31111 , \31109 , \31110 );
xnor \U$30797 ( \31112 , \31111 , \22377 );
xor \U$30798 ( \31113 , \31108 , \31112 );
xor \U$30799 ( \31114 , \31100 , \31113 );
xor \U$30800 ( \31115 , \31071 , \31114 );
xor \U$30801 ( \31116 , \31062 , \31115 );
xor \U$30802 ( \31117 , \31053 , \31116 );
and \U$30803 ( \31118 , \30832 , \30836 );
and \U$30804 ( \31119 , \30836 , \30841 );
and \U$30805 ( \31120 , \30832 , \30841 );
or \U$30806 ( \31121 , \31118 , \31119 , \31120 );
and \U$30807 ( \31122 , \30866 , \31021 );
and \U$30808 ( \31123 , \31021 , \31036 );
and \U$30809 ( \31124 , \30866 , \31036 );
or \U$30810 ( \31125 , \31122 , \31123 , \31124 );
xor \U$30811 ( \31126 , \31121 , \31125 );
and \U$30812 ( \31127 , \30896 , \30900 );
and \U$30813 ( \31128 , \30900 , \30905 );
and \U$30814 ( \31129 , \30896 , \30905 );
or \U$30815 ( \31130 , \31127 , \31128 , \31129 );
and \U$30816 ( \31131 , \30881 , \30885 );
and \U$30817 ( \31132 , \30885 , \30890 );
and \U$30818 ( \31133 , \30881 , \30890 );
or \U$30819 ( \31134 , \31131 , \31132 , \31133 );
xor \U$30820 ( \31135 , \31130 , \31134 );
and \U$30821 ( \31136 , \30870 , \30871 );
and \U$30822 ( \31137 , \30871 , \30876 );
and \U$30823 ( \31138 , \30870 , \30876 );
or \U$30824 ( \31139 , \31136 , \31137 , \31138 );
xor \U$30825 ( \31140 , \31135 , \31139 );
and \U$30826 ( \31141 , \30877 , \30891 );
and \U$30827 ( \31142 , \30891 , \30906 );
and \U$30828 ( \31143 , \30877 , \30906 );
or \U$30829 ( \31144 , \31141 , \31142 , \31143 );
and \U$30830 ( \31145 , \30908 , \30912 );
and \U$30831 ( \31146 , \30912 , \30917 );
and \U$30832 ( \31147 , \30908 , \30917 );
or \U$30833 ( \31148 , \31145 , \31146 , \31147 );
and \U$30834 ( \31149 , \31009 , \31013 );
and \U$30835 ( \31150 , \31013 , \31018 );
and \U$30836 ( \31151 , \31009 , \31018 );
or \U$30837 ( \31152 , \31149 , \31150 , \31151 );
xor \U$30838 ( \31153 , \31148 , \31152 );
and \U$30839 ( \31154 , \30951 , \30955 );
and \U$30840 ( \31155 , \30955 , \30960 );
and \U$30841 ( \31156 , \30951 , \30960 );
or \U$30842 ( \31157 , \31154 , \31155 , \31156 );
xor \U$30843 ( \31158 , \31153 , \31157 );
xor \U$30844 ( \31159 , \31144 , \31158 );
and \U$30845 ( \31160 , \22329 , \22671 );
and \U$30846 ( \31161 , \22294 , \22669 );
nor \U$30847 ( \31162 , \31160 , \31161 );
xnor \U$30848 ( \31163 , \31162 , \22681 );
and \U$30849 ( \31164 , \22350 , \22691 );
and \U$30850 ( \31165 , \22318 , \22689 );
nor \U$30851 ( \31166 , \31164 , \31165 );
xnor \U$30852 ( \31167 , \31166 , \22701 );
xor \U$30853 ( \31168 , \31163 , \31167 );
and \U$30854 ( \31169 , \22372 , \22720 );
and \U$30855 ( \31170 , \22339 , \22707 );
nor \U$30856 ( \31171 , \31169 , \31170 );
xnor \U$30857 ( \31172 , \31171 , \22067 );
xor \U$30858 ( \31173 , \31168 , \31172 );
and \U$30859 ( \31174 , \22262 , \22598 );
and \U$30860 ( \31175 , \22224 , \22596 );
nor \U$30861 ( \31176 , \31174 , \31175 );
xnor \U$30862 ( \31177 , \31176 , \22608 );
and \U$30863 ( \31178 , \22283 , \22619 );
and \U$30864 ( \31179 , \22251 , \22617 );
nor \U$30865 ( \31180 , \31178 , \31179 );
xnor \U$30866 ( \31181 , \31180 , \22629 );
xor \U$30867 ( \31182 , \31177 , \31181 );
and \U$30868 ( \31183 , \22305 , \22641 );
and \U$30869 ( \31184 , \22272 , \22639 );
nor \U$30870 ( \31185 , \31183 , \31184 );
xnor \U$30871 ( \31186 , \31185 , \22651 );
xor \U$30872 ( \31187 , \31182 , \31186 );
xor \U$30873 ( \31188 , \31173 , \31187 );
and \U$30874 ( \31189 , \22192 , \22530 );
and \U$30875 ( \31190 , \22156 , \22528 );
nor \U$30876 ( \31191 , \31189 , \31190 );
xnor \U$30877 ( \31192 , \31191 , \22540 );
and \U$30878 ( \31193 , \22213 , \22551 );
and \U$30879 ( \31194 , \22181 , \22549 );
nor \U$30880 ( \31195 , \31193 , \31194 );
xnor \U$30881 ( \31196 , \31195 , \22561 );
xor \U$30882 ( \31197 , \31192 , \31196 );
and \U$30883 ( \31198 , \22235 , \22573 );
and \U$30884 ( \31199 , \22202 , \22571 );
nor \U$30885 ( \31200 , \31198 , \31199 );
xnor \U$30886 ( \31201 , \31200 , \22583 );
xor \U$30887 ( \31202 , \31197 , \31201 );
xor \U$30888 ( \31203 , \31188 , \31202 );
and \U$30889 ( \31204 , \30968 , \30972 );
and \U$30890 ( \31205 , \30972 , \30977 );
and \U$30891 ( \31206 , \30968 , \30977 );
or \U$30892 ( \31207 , \31204 , \31205 , \31206 );
and \U$30893 ( \31208 , \22429 , \21978 );
not \U$30894 ( \31209 , \31208 );
xor \U$30895 ( \31210 , \31207 , \31209 );
and \U$30896 ( \31211 , \22397 , \23173 );
and \U$30897 ( \31212 , \22361 , \22999 );
nor \U$30898 ( \31213 , \31211 , \31212 );
xnor \U$30899 ( \31214 , \31213 , \22016 );
and \U$30900 ( \31215 , \22418 , \22021 );
and \U$30901 ( \31216 , \22386 , \22019 );
nor \U$30902 ( \31217 , \31215 , \31216 );
xnor \U$30903 ( \31218 , \31217 , \21595 );
xor \U$30904 ( \31219 , \31214 , \31218 );
and \U$30905 ( \31220 , \22440 , \21983 );
and \U$30906 ( \31221 , \22407 , \21981 );
nor \U$30907 ( \31222 , \31220 , \31221 );
xnor \U$30908 ( \31223 , \31222 , \21995 );
xor \U$30909 ( \31224 , \31219 , \31223 );
xor \U$30910 ( \31225 , \31210 , \31224 );
xor \U$30911 ( \31226 , \31203 , \31225 );
and \U$30912 ( \31227 , \30936 , \30940 );
and \U$30913 ( \31228 , \30940 , \30945 );
and \U$30914 ( \31229 , \30936 , \30945 );
or \U$30915 ( \31230 , \31227 , \31228 , \31229 );
and \U$30916 ( \31231 , \30922 , \30926 );
and \U$30917 ( \31232 , \30926 , \30931 );
and \U$30918 ( \31233 , \30922 , \30931 );
or \U$30919 ( \31234 , \31231 , \31232 , \31233 );
xor \U$30920 ( \31235 , \31230 , \31234 );
and \U$30921 ( \31236 , \30983 , \30987 );
and \U$30922 ( \31237 , \30987 , \30992 );
and \U$30923 ( \31238 , \30983 , \30992 );
or \U$30924 ( \31239 , \31236 , \31237 , \31238 );
xor \U$30925 ( \31240 , \31235 , \31239 );
xor \U$30926 ( \31241 , \31226 , \31240 );
xor \U$30927 ( \31242 , \31159 , \31241 );
xor \U$30928 ( \31243 , \31140 , \31242 );
and \U$30929 ( \31244 , \30856 , \30860 );
and \U$30930 ( \31245 , \30860 , \30865 );
and \U$30931 ( \31246 , \30856 , \30865 );
or \U$30932 ( \31247 , \31244 , \31245 , \31246 );
and \U$30933 ( \31248 , \31000 , \31004 );
and \U$30934 ( \31249 , \31004 , \31019 );
and \U$30935 ( \31250 , \31000 , \31019 );
or \U$30936 ( \31251 , \31248 , \31249 , \31250 );
xor \U$30937 ( \31252 , \31247 , \31251 );
and \U$30938 ( \31253 , \30918 , \30962 );
and \U$30939 ( \31254 , \30962 , \30994 );
and \U$30940 ( \31255 , \30918 , \30994 );
or \U$30941 ( \31256 , \31253 , \31254 , \31255 );
xor \U$30942 ( \31257 , \31252 , \31256 );
xor \U$30943 ( \31258 , \31243 , \31257 );
xor \U$30944 ( \31259 , \31126 , \31258 );
xor \U$30945 ( \31260 , \31117 , \31259 );
xor \U$30946 ( \31261 , \31049 , \31260 );
and \U$30947 ( \31262 , \30824 , \31039 );
nor \U$30948 ( \31263 , \31261 , \31262 );
and \U$30949 ( \31264 , \31053 , \31116 );
and \U$30950 ( \31265 , \31116 , \31259 );
and \U$30951 ( \31266 , \31053 , \31259 );
or \U$30952 ( \31267 , \31264 , \31265 , \31266 );
and \U$30953 ( \31268 , \31121 , \31125 );
and \U$30954 ( \31269 , \31125 , \31258 );
and \U$30955 ( \31270 , \31121 , \31258 );
or \U$30956 ( \31271 , \31268 , \31269 , \31270 );
and \U$30957 ( \31272 , \31247 , \31251 );
and \U$30958 ( \31273 , \31251 , \31256 );
and \U$30959 ( \31274 , \31247 , \31256 );
or \U$30960 ( \31275 , \31272 , \31273 , \31274 );
and \U$30961 ( \31276 , \31144 , \31158 );
and \U$30962 ( \31277 , \31158 , \31241 );
and \U$30963 ( \31278 , \31144 , \31241 );
or \U$30964 ( \31279 , \31276 , \31277 , \31278 );
xor \U$30965 ( \31280 , \31275 , \31279 );
and \U$30966 ( \31281 , \31173 , \31187 );
and \U$30967 ( \31282 , \31187 , \31202 );
and \U$30968 ( \31283 , \31173 , \31202 );
or \U$30969 ( \31284 , \31281 , \31282 , \31283 );
and \U$30970 ( \31285 , \31085 , \31099 );
and \U$30971 ( \31286 , \31099 , \31113 );
and \U$30972 ( \31287 , \31085 , \31113 );
or \U$30973 ( \31288 , \31285 , \31286 , \31287 );
xor \U$30974 ( \31289 , \31284 , \31288 );
not \U$30975 ( \31290 , \22334 );
and \U$30976 ( \31291 , \21977 , \22345 );
and \U$30977 ( \31292 , \21990 , \22343 );
nor \U$30978 ( \31293 , \31291 , \31292 );
xnor \U$30979 ( \31294 , \31293 , \22355 );
xor \U$30980 ( \31295 , \31290 , \31294 );
and \U$30981 ( \31296 , \22030 , \22367 );
and \U$30982 ( \31297 , \22001 , \22365 );
nor \U$30983 ( \31298 , \31296 , \31297 );
xnor \U$30984 ( \31299 , \31298 , \22377 );
xor \U$30985 ( \31300 , \31295 , \31299 );
xor \U$30986 ( \31301 , \31289 , \31300 );
xor \U$30987 ( \31302 , \31280 , \31301 );
xor \U$30988 ( \31303 , \31271 , \31302 );
and \U$30989 ( \31304 , \31057 , \31061 );
and \U$30990 ( \31305 , \31061 , \31115 );
and \U$30991 ( \31306 , \31057 , \31115 );
or \U$30992 ( \31307 , \31304 , \31305 , \31306 );
and \U$30993 ( \31308 , \31140 , \31242 );
and \U$30994 ( \31309 , \31242 , \31257 );
and \U$30995 ( \31310 , \31140 , \31257 );
or \U$30996 ( \31311 , \31308 , \31309 , \31310 );
xor \U$30997 ( \31312 , \31307 , \31311 );
and \U$30998 ( \31313 , \31148 , \31152 );
and \U$30999 ( \31314 , \31152 , \31157 );
and \U$31000 ( \31315 , \31148 , \31157 );
or \U$31001 ( \31316 , \31313 , \31314 , \31315 );
and \U$31002 ( \31317 , \31230 , \31234 );
and \U$31003 ( \31318 , \31234 , \31239 );
and \U$31004 ( \31319 , \31230 , \31239 );
or \U$31005 ( \31320 , \31317 , \31318 , \31319 );
xor \U$31006 ( \31321 , \31316 , \31320 );
and \U$31007 ( \31322 , \31207 , \31209 );
and \U$31008 ( \31323 , \31209 , \31224 );
and \U$31009 ( \31324 , \31207 , \31224 );
or \U$31010 ( \31325 , \31322 , \31323 , \31324 );
xor \U$31011 ( \31326 , \31321 , \31325 );
and \U$31012 ( \31327 , \31192 , \31196 );
and \U$31013 ( \31328 , \31196 , \31201 );
and \U$31014 ( \31329 , \31192 , \31201 );
or \U$31015 ( \31330 , \31327 , \31328 , \31329 );
and \U$31016 ( \31331 , \31177 , \31181 );
and \U$31017 ( \31332 , \31181 , \31186 );
and \U$31018 ( \31333 , \31177 , \31186 );
or \U$31019 ( \31334 , \31331 , \31332 , \31333 );
xor \U$31020 ( \31335 , \31330 , \31334 );
and \U$31021 ( \31336 , \31163 , \31167 );
and \U$31022 ( \31337 , \31167 , \31172 );
and \U$31023 ( \31338 , \31163 , \31172 );
or \U$31024 ( \31339 , \31336 , \31337 , \31338 );
xor \U$31025 ( \31340 , \31335 , \31339 );
and \U$31026 ( \31341 , \31103 , \31107 );
and \U$31027 ( \31342 , \31107 , \31112 );
and \U$31028 ( \31343 , \31103 , \31112 );
or \U$31029 ( \31344 , \31341 , \31342 , \31343 );
and \U$31030 ( \31345 , \31089 , \31093 );
and \U$31031 ( \31346 , \31093 , \31098 );
and \U$31032 ( \31347 , \31089 , \31098 );
or \U$31033 ( \31348 , \31345 , \31346 , \31347 );
xor \U$31034 ( \31349 , \31344 , \31348 );
and \U$31035 ( \31350 , \31075 , \31079 );
and \U$31036 ( \31351 , \31079 , \31084 );
and \U$31037 ( \31352 , \31075 , \31084 );
or \U$31038 ( \31353 , \31350 , \31351 , \31352 );
xor \U$31039 ( \31354 , \31349 , \31353 );
xor \U$31040 ( \31355 , \31340 , \31354 );
and \U$31041 ( \31356 , \22156 , \22530 );
and \U$31042 ( \31357 , \22167 , \22528 );
nor \U$31043 ( \31358 , \31356 , \31357 );
xnor \U$31044 ( \31359 , \31358 , \22540 );
and \U$31045 ( \31360 , \22181 , \22551 );
and \U$31046 ( \31361 , \22192 , \22549 );
nor \U$31047 ( \31362 , \31360 , \31361 );
xnor \U$31048 ( \31363 , \31362 , \22561 );
xor \U$31049 ( \31364 , \31359 , \31363 );
and \U$31050 ( \31365 , \22202 , \22573 );
and \U$31051 ( \31366 , \22213 , \22571 );
nor \U$31052 ( \31367 , \31365 , \31366 );
xnor \U$31053 ( \31368 , \31367 , \22583 );
xor \U$31054 ( \31369 , \31364 , \31368 );
and \U$31055 ( \31370 , \22089 , \22463 );
and \U$31056 ( \31371 , \22100 , \22461 );
nor \U$31057 ( \31372 , \31370 , \31371 );
xnor \U$31058 ( \31373 , \31372 , \22473 );
and \U$31059 ( \31374 , \22113 , \22484 );
and \U$31060 ( \31375 , \22124 , \22482 );
nor \U$31061 ( \31376 , \31374 , \31375 );
xnor \U$31062 ( \31377 , \31376 , \22494 );
xor \U$31063 ( \31378 , \31373 , \31377 );
and \U$31064 ( \31379 , \22134 , \22506 );
and \U$31065 ( \31380 , \22145 , \22504 );
nor \U$31066 ( \31381 , \31379 , \31380 );
xnor \U$31067 ( \31382 , \31381 , \22516 );
xor \U$31068 ( \31383 , \31378 , \31382 );
xor \U$31069 ( \31384 , \31369 , \31383 );
and \U$31070 ( \31385 , \23230 , \22392 );
and \U$31071 ( \31386 , \23329 , \22390 );
nor \U$31072 ( \31387 , \31385 , \31386 );
xnor \U$31073 ( \31388 , \31387 , \22402 );
and \U$31074 ( \31389 , \22858 , \22413 );
and \U$31075 ( \31390 , \22894 , \22411 );
nor \U$31076 ( \31391 , \31389 , \31390 );
xnor \U$31077 ( \31392 , \31391 , \22423 );
xor \U$31078 ( \31393 , \31388 , \31392 );
and \U$31079 ( \31394 , \22071 , \22435 );
and \U$31080 ( \31395 , \22081 , \22433 );
nor \U$31081 ( \31396 , \31394 , \31395 );
xnor \U$31082 ( \31397 , \31396 , \22445 );
xor \U$31083 ( \31398 , \31393 , \31397 );
xor \U$31084 ( \31399 , \31384 , \31398 );
and \U$31085 ( \31400 , \22361 , \23173 );
and \U$31086 ( \31401 , \22372 , \22999 );
nor \U$31087 ( \31402 , \31400 , \31401 );
xnor \U$31088 ( \31403 , \31402 , \22016 );
and \U$31089 ( \31404 , \22386 , \22021 );
and \U$31090 ( \31405 , \22397 , \22019 );
nor \U$31091 ( \31406 , \31404 , \31405 );
xnor \U$31092 ( \31407 , \31406 , \21595 );
xor \U$31093 ( \31408 , \31403 , \31407 );
and \U$31094 ( \31409 , \22407 , \21983 );
and \U$31095 ( \31410 , \22418 , \21981 );
nor \U$31096 ( \31411 , \31409 , \31410 );
xnor \U$31097 ( \31412 , \31411 , \21995 );
xor \U$31098 ( \31413 , \31408 , \31412 );
and \U$31099 ( \31414 , \22294 , \22671 );
and \U$31100 ( \31415 , \22305 , \22669 );
nor \U$31101 ( \31416 , \31414 , \31415 );
xnor \U$31102 ( \31417 , \31416 , \22681 );
and \U$31103 ( \31418 , \22318 , \22691 );
and \U$31104 ( \31419 , \22329 , \22689 );
nor \U$31105 ( \31420 , \31418 , \31419 );
xnor \U$31106 ( \31421 , \31420 , \22701 );
xor \U$31107 ( \31422 , \31417 , \31421 );
and \U$31108 ( \31423 , \22339 , \22720 );
and \U$31109 ( \31424 , \22350 , \22707 );
nor \U$31110 ( \31425 , \31423 , \31424 );
xnor \U$31111 ( \31426 , \31425 , \22067 );
xor \U$31112 ( \31427 , \31422 , \31426 );
xor \U$31113 ( \31428 , \31413 , \31427 );
and \U$31114 ( \31429 , \22224 , \22598 );
and \U$31115 ( \31430 , \22235 , \22596 );
nor \U$31116 ( \31431 , \31429 , \31430 );
xnor \U$31117 ( \31432 , \31431 , \22608 );
and \U$31118 ( \31433 , \22251 , \22619 );
and \U$31119 ( \31434 , \22262 , \22617 );
nor \U$31120 ( \31435 , \31433 , \31434 );
xnor \U$31121 ( \31436 , \31435 , \22629 );
xor \U$31122 ( \31437 , \31432 , \31436 );
and \U$31123 ( \31438 , \22272 , \22641 );
and \U$31124 ( \31439 , \22283 , \22639 );
nor \U$31125 ( \31440 , \31438 , \31439 );
xnor \U$31126 ( \31441 , \31440 , \22651 );
xor \U$31127 ( \31442 , \31437 , \31441 );
xor \U$31128 ( \31443 , \31428 , \31442 );
xor \U$31129 ( \31444 , \31399 , \31443 );
and \U$31130 ( \31445 , \31214 , \31218 );
and \U$31131 ( \31446 , \31218 , \31223 );
and \U$31132 ( \31447 , \31214 , \31223 );
or \U$31133 ( \31448 , \31445 , \31446 , \31447 );
xor \U$31134 ( \31449 , \31448 , \31208 );
and \U$31135 ( \31450 , \22440 , \21978 );
xor \U$31136 ( \31451 , \31449 , \31450 );
xor \U$31137 ( \31452 , \31444 , \31451 );
xor \U$31138 ( \31453 , \31355 , \31452 );
xor \U$31139 ( \31454 , \31326 , \31453 );
and \U$31140 ( \31455 , \31130 , \31134 );
and \U$31141 ( \31456 , \31134 , \31139 );
and \U$31142 ( \31457 , \31130 , \31139 );
or \U$31143 ( \31458 , \31455 , \31456 , \31457 );
and \U$31144 ( \31459 , \31066 , \31070 );
and \U$31145 ( \31460 , \31070 , \31114 );
and \U$31146 ( \31461 , \31066 , \31114 );
or \U$31147 ( \31462 , \31459 , \31460 , \31461 );
xor \U$31148 ( \31463 , \31458 , \31462 );
and \U$31149 ( \31464 , \31203 , \31225 );
and \U$31150 ( \31465 , \31225 , \31240 );
and \U$31151 ( \31466 , \31203 , \31240 );
or \U$31152 ( \31467 , \31464 , \31465 , \31466 );
xor \U$31153 ( \31468 , \31463 , \31467 );
xor \U$31154 ( \31469 , \31454 , \31468 );
xor \U$31155 ( \31470 , \31312 , \31469 );
xor \U$31156 ( \31471 , \31303 , \31470 );
xor \U$31157 ( \31472 , \31267 , \31471 );
and \U$31158 ( \31473 , \31049 , \31260 );
nor \U$31159 ( \31474 , \31472 , \31473 );
nor \U$31160 ( \31475 , \31263 , \31474 );
and \U$31161 ( \31476 , \31271 , \31302 );
and \U$31162 ( \31477 , \31302 , \31470 );
and \U$31163 ( \31478 , \31271 , \31470 );
or \U$31164 ( \31479 , \31476 , \31477 , \31478 );
and \U$31165 ( \31480 , \31307 , \31311 );
and \U$31166 ( \31481 , \31311 , \31469 );
and \U$31167 ( \31482 , \31307 , \31469 );
or \U$31168 ( \31483 , \31480 , \31481 , \31482 );
and \U$31169 ( \31484 , \31316 , \31320 );
and \U$31170 ( \31485 , \31320 , \31325 );
and \U$31171 ( \31486 , \31316 , \31325 );
or \U$31172 ( \31487 , \31484 , \31485 , \31486 );
and \U$31173 ( \31488 , \31284 , \31288 );
and \U$31174 ( \31489 , \31288 , \31300 );
and \U$31175 ( \31490 , \31284 , \31300 );
or \U$31176 ( \31491 , \31488 , \31489 , \31490 );
xor \U$31177 ( \31492 , \31487 , \31491 );
and \U$31178 ( \31493 , \31399 , \31443 );
and \U$31179 ( \31494 , \31443 , \31451 );
and \U$31180 ( \31495 , \31399 , \31451 );
or \U$31181 ( \31496 , \31493 , \31494 , \31495 );
xor \U$31182 ( \31497 , \31492 , \31496 );
and \U$31183 ( \31498 , \31458 , \31462 );
and \U$31184 ( \31499 , \31462 , \31467 );
and \U$31185 ( \31500 , \31458 , \31467 );
or \U$31186 ( \31501 , \31498 , \31499 , \31500 );
and \U$31187 ( \31502 , \31340 , \31354 );
and \U$31188 ( \31503 , \31354 , \31452 );
and \U$31189 ( \31504 , \31340 , \31452 );
or \U$31190 ( \31505 , \31502 , \31503 , \31504 );
xor \U$31191 ( \31506 , \31501 , \31505 );
and \U$31192 ( \31507 , \31344 , \31348 );
and \U$31193 ( \31508 , \31348 , \31353 );
and \U$31194 ( \31509 , \31344 , \31353 );
or \U$31195 ( \31510 , \31507 , \31508 , \31509 );
and \U$31196 ( \31511 , \31330 , \31334 );
and \U$31197 ( \31512 , \31334 , \31339 );
and \U$31198 ( \31513 , \31330 , \31339 );
or \U$31199 ( \31514 , \31511 , \31512 , \31513 );
xor \U$31200 ( \31515 , \31510 , \31514 );
and \U$31201 ( \31516 , \31448 , \31208 );
and \U$31202 ( \31517 , \31208 , \31450 );
and \U$31203 ( \31518 , \31448 , \31450 );
or \U$31204 ( \31519 , \31516 , \31517 , \31518 );
xor \U$31205 ( \31520 , \31515 , \31519 );
xor \U$31206 ( \31521 , \31506 , \31520 );
xor \U$31207 ( \31522 , \31497 , \31521 );
xor \U$31208 ( \31523 , \31483 , \31522 );
and \U$31209 ( \31524 , \31275 , \31279 );
and \U$31210 ( \31525 , \31279 , \31301 );
and \U$31211 ( \31526 , \31275 , \31301 );
or \U$31212 ( \31527 , \31524 , \31525 , \31526 );
and \U$31213 ( \31528 , \31326 , \31453 );
and \U$31214 ( \31529 , \31453 , \31468 );
and \U$31215 ( \31530 , \31326 , \31468 );
or \U$31216 ( \31531 , \31528 , \31529 , \31530 );
xor \U$31217 ( \31532 , \31527 , \31531 );
and \U$31218 ( \31533 , \31290 , \31294 );
and \U$31219 ( \31534 , \31294 , \31299 );
and \U$31220 ( \31535 , \31290 , \31299 );
or \U$31221 ( \31536 , \31533 , \31534 , \31535 );
and \U$31222 ( \31537 , \31388 , \31392 );
and \U$31223 ( \31538 , \31392 , \31397 );
and \U$31224 ( \31539 , \31388 , \31397 );
or \U$31225 ( \31540 , \31537 , \31538 , \31539 );
xor \U$31226 ( \31541 , \31536 , \31540 );
and \U$31227 ( \31542 , \31373 , \31377 );
and \U$31228 ( \31543 , \31377 , \31382 );
and \U$31229 ( \31544 , \31373 , \31382 );
or \U$31230 ( \31545 , \31542 , \31543 , \31544 );
xor \U$31231 ( \31546 , \31541 , \31545 );
and \U$31232 ( \31547 , \22329 , \22691 );
and \U$31233 ( \31548 , \22294 , \22689 );
nor \U$31234 ( \31549 , \31547 , \31548 );
xnor \U$31235 ( \31550 , \31549 , \22701 );
and \U$31236 ( \31551 , \22350 , \22720 );
and \U$31237 ( \31552 , \22318 , \22707 );
nor \U$31238 ( \31553 , \31551 , \31552 );
xnor \U$31239 ( \31554 , \31553 , \22067 );
xor \U$31240 ( \31555 , \31550 , \31554 );
and \U$31241 ( \31556 , \22372 , \23173 );
and \U$31242 ( \31557 , \22339 , \22999 );
nor \U$31243 ( \31558 , \31556 , \31557 );
xnor \U$31244 ( \31559 , \31558 , \22016 );
xor \U$31245 ( \31560 , \31555 , \31559 );
and \U$31246 ( \31561 , \22262 , \22619 );
and \U$31247 ( \31562 , \22224 , \22617 );
nor \U$31248 ( \31563 , \31561 , \31562 );
xnor \U$31249 ( \31564 , \31563 , \22629 );
and \U$31250 ( \31565 , \22283 , \22641 );
and \U$31251 ( \31566 , \22251 , \22639 );
nor \U$31252 ( \31567 , \31565 , \31566 );
xnor \U$31253 ( \31568 , \31567 , \22651 );
xor \U$31254 ( \31569 , \31564 , \31568 );
and \U$31255 ( \31570 , \22305 , \22671 );
and \U$31256 ( \31571 , \22272 , \22669 );
nor \U$31257 ( \31572 , \31570 , \31571 );
xnor \U$31258 ( \31573 , \31572 , \22681 );
xor \U$31259 ( \31574 , \31569 , \31573 );
xor \U$31260 ( \31575 , \31560 , \31574 );
and \U$31261 ( \31576 , \22192 , \22551 );
and \U$31262 ( \31577 , \22156 , \22549 );
nor \U$31263 ( \31578 , \31576 , \31577 );
xnor \U$31264 ( \31579 , \31578 , \22561 );
and \U$31265 ( \31580 , \22213 , \22573 );
and \U$31266 ( \31581 , \22181 , \22571 );
nor \U$31267 ( \31582 , \31580 , \31581 );
xnor \U$31268 ( \31583 , \31582 , \22583 );
xor \U$31269 ( \31584 , \31579 , \31583 );
and \U$31270 ( \31585 , \22235 , \22598 );
and \U$31271 ( \31586 , \22202 , \22596 );
nor \U$31272 ( \31587 , \31585 , \31586 );
xnor \U$31273 ( \31588 , \31587 , \22608 );
xor \U$31274 ( \31589 , \31584 , \31588 );
xor \U$31275 ( \31590 , \31575 , \31589 );
and \U$31276 ( \31591 , \31403 , \31407 );
and \U$31277 ( \31592 , \31407 , \31412 );
and \U$31278 ( \31593 , \31403 , \31412 );
or \U$31279 ( \31594 , \31591 , \31592 , \31593 );
and \U$31280 ( \31595 , \22397 , \22021 );
and \U$31281 ( \31596 , \22361 , \22019 );
nor \U$31282 ( \31597 , \31595 , \31596 );
xnor \U$31283 ( \31598 , \31597 , \21595 );
and \U$31284 ( \31599 , \22418 , \21983 );
and \U$31285 ( \31600 , \22386 , \21981 );
nor \U$31286 ( \31601 , \31599 , \31600 );
xnor \U$31287 ( \31602 , \31601 , \21995 );
xor \U$31288 ( \31603 , \31598 , \31602 );
and \U$31289 ( \31604 , \22407 , \21978 );
xor \U$31290 ( \31605 , \31603 , \31604 );
xnor \U$31291 ( \31606 , \31594 , \31605 );
xor \U$31292 ( \31607 , \31590 , \31606 );
and \U$31293 ( \31608 , \31359 , \31363 );
and \U$31294 ( \31609 , \31363 , \31368 );
and \U$31295 ( \31610 , \31359 , \31368 );
or \U$31296 ( \31611 , \31608 , \31609 , \31610 );
and \U$31297 ( \31612 , \31432 , \31436 );
and \U$31298 ( \31613 , \31436 , \31441 );
and \U$31299 ( \31614 , \31432 , \31441 );
or \U$31300 ( \31615 , \31612 , \31613 , \31614 );
xor \U$31301 ( \31616 , \31611 , \31615 );
and \U$31302 ( \31617 , \31417 , \31421 );
and \U$31303 ( \31618 , \31421 , \31426 );
and \U$31304 ( \31619 , \31417 , \31426 );
or \U$31305 ( \31620 , \31617 , \31618 , \31619 );
xor \U$31306 ( \31621 , \31616 , \31620 );
xor \U$31307 ( \31622 , \31607 , \31621 );
xor \U$31308 ( \31623 , \31546 , \31622 );
and \U$31309 ( \31624 , \31413 , \31427 );
and \U$31310 ( \31625 , \31427 , \31442 );
and \U$31311 ( \31626 , \31413 , \31442 );
or \U$31312 ( \31627 , \31624 , \31625 , \31626 );
and \U$31313 ( \31628 , \31369 , \31383 );
and \U$31314 ( \31629 , \31383 , \31398 );
and \U$31315 ( \31630 , \31369 , \31398 );
or \U$31316 ( \31631 , \31628 , \31629 , \31630 );
xor \U$31317 ( \31632 , \31627 , \31631 );
and \U$31318 ( \31633 , \22124 , \22484 );
and \U$31319 ( \31634 , \22089 , \22482 );
nor \U$31320 ( \31635 , \31633 , \31634 );
xnor \U$31321 ( \31636 , \31635 , \22494 );
and \U$31322 ( \31637 , \22145 , \22506 );
and \U$31323 ( \31638 , \22113 , \22504 );
nor \U$31324 ( \31639 , \31637 , \31638 );
xnor \U$31325 ( \31640 , \31639 , \22516 );
xor \U$31326 ( \31641 , \31636 , \31640 );
and \U$31327 ( \31642 , \22167 , \22530 );
and \U$31328 ( \31643 , \22134 , \22528 );
nor \U$31329 ( \31644 , \31642 , \31643 );
xnor \U$31330 ( \31645 , \31644 , \22540 );
xor \U$31331 ( \31646 , \31641 , \31645 );
and \U$31332 ( \31647 , \22894 , \22413 );
and \U$31333 ( \31648 , \23230 , \22411 );
nor \U$31334 ( \31649 , \31647 , \31648 );
xnor \U$31335 ( \31650 , \31649 , \22423 );
and \U$31336 ( \31651 , \22081 , \22435 );
and \U$31337 ( \31652 , \22858 , \22433 );
nor \U$31338 ( \31653 , \31651 , \31652 );
xnor \U$31339 ( \31654 , \31653 , \22445 );
xor \U$31340 ( \31655 , \31650 , \31654 );
and \U$31341 ( \31656 , \22100 , \22463 );
and \U$31342 ( \31657 , \22071 , \22461 );
nor \U$31343 ( \31658 , \31656 , \31657 );
xnor \U$31344 ( \31659 , \31658 , \22473 );
xor \U$31345 ( \31660 , \31655 , \31659 );
xor \U$31346 ( \31661 , \31646 , \31660 );
and \U$31347 ( \31662 , \21990 , \22345 );
not \U$31348 ( \31663 , \31662 );
xnor \U$31349 ( \31664 , \31663 , \22355 );
and \U$31350 ( \31665 , \22001 , \22367 );
and \U$31351 ( \31666 , \21977 , \22365 );
nor \U$31352 ( \31667 , \31665 , \31666 );
xnor \U$31353 ( \31668 , \31667 , \22377 );
xor \U$31354 ( \31669 , \31664 , \31668 );
and \U$31355 ( \31670 , \23329 , \22392 );
and \U$31356 ( \31671 , \22030 , \22390 );
nor \U$31357 ( \31672 , \31670 , \31671 );
xnor \U$31358 ( \31673 , \31672 , \22402 );
xor \U$31359 ( \31674 , \31669 , \31673 );
xor \U$31360 ( \31675 , \31661 , \31674 );
xor \U$31361 ( \31676 , \31632 , \31675 );
xor \U$31362 ( \31677 , \31623 , \31676 );
xor \U$31363 ( \31678 , \31532 , \31677 );
xor \U$31364 ( \31679 , \31523 , \31678 );
xor \U$31365 ( \31680 , \31479 , \31679 );
and \U$31366 ( \31681 , \31267 , \31471 );
nor \U$31367 ( \31682 , \31680 , \31681 );
and \U$31368 ( \31683 , \31483 , \31522 );
and \U$31369 ( \31684 , \31522 , \31678 );
and \U$31370 ( \31685 , \31483 , \31678 );
or \U$31371 ( \31686 , \31683 , \31684 , \31685 );
and \U$31372 ( \31687 , \31527 , \31531 );
and \U$31373 ( \31688 , \31531 , \31677 );
and \U$31374 ( \31689 , \31527 , \31677 );
or \U$31375 ( \31690 , \31687 , \31688 , \31689 );
and \U$31376 ( \31691 , \31497 , \31521 );
xor \U$31377 ( \31692 , \31690 , \31691 );
and \U$31378 ( \31693 , \31501 , \31505 );
and \U$31379 ( \31694 , \31505 , \31520 );
and \U$31380 ( \31695 , \31501 , \31520 );
or \U$31381 ( \31696 , \31693 , \31694 , \31695 );
and \U$31382 ( \31697 , \31536 , \31540 );
and \U$31383 ( \31698 , \31540 , \31545 );
and \U$31384 ( \31699 , \31536 , \31545 );
or \U$31385 ( \31700 , \31697 , \31698 , \31699 );
and \U$31386 ( \31701 , \31611 , \31615 );
and \U$31387 ( \31702 , \31615 , \31620 );
and \U$31388 ( \31703 , \31611 , \31620 );
or \U$31389 ( \31704 , \31701 , \31702 , \31703 );
xor \U$31390 ( \31705 , \31700 , \31704 );
or \U$31391 ( \31706 , \31594 , \31605 );
xor \U$31392 ( \31707 , \31705 , \31706 );
and \U$31393 ( \31708 , \31579 , \31583 );
and \U$31394 ( \31709 , \31583 , \31588 );
and \U$31395 ( \31710 , \31579 , \31588 );
or \U$31396 ( \31711 , \31708 , \31709 , \31710 );
and \U$31397 ( \31712 , \31564 , \31568 );
and \U$31398 ( \31713 , \31568 , \31573 );
and \U$31399 ( \31714 , \31564 , \31573 );
or \U$31400 ( \31715 , \31712 , \31713 , \31714 );
xor \U$31401 ( \31716 , \31711 , \31715 );
and \U$31402 ( \31717 , \31550 , \31554 );
and \U$31403 ( \31718 , \31554 , \31559 );
and \U$31404 ( \31719 , \31550 , \31559 );
or \U$31405 ( \31720 , \31717 , \31718 , \31719 );
xor \U$31406 ( \31721 , \31716 , \31720 );
and \U$31407 ( \31722 , \31664 , \31668 );
and \U$31408 ( \31723 , \31668 , \31673 );
and \U$31409 ( \31724 , \31664 , \31673 );
or \U$31410 ( \31725 , \31722 , \31723 , \31724 );
and \U$31411 ( \31726 , \31650 , \31654 );
and \U$31412 ( \31727 , \31654 , \31659 );
and \U$31413 ( \31728 , \31650 , \31659 );
or \U$31414 ( \31729 , \31726 , \31727 , \31728 );
xor \U$31415 ( \31730 , \31725 , \31729 );
and \U$31416 ( \31731 , \31636 , \31640 );
and \U$31417 ( \31732 , \31640 , \31645 );
and \U$31418 ( \31733 , \31636 , \31645 );
or \U$31419 ( \31734 , \31731 , \31732 , \31733 );
xor \U$31420 ( \31735 , \31730 , \31734 );
xor \U$31421 ( \31736 , \31721 , \31735 );
not \U$31422 ( \31737 , \22355 );
and \U$31423 ( \31738 , \21977 , \22367 );
and \U$31424 ( \31739 , \21990 , \22365 );
nor \U$31425 ( \31740 , \31738 , \31739 );
xnor \U$31426 ( \31741 , \31740 , \22377 );
xor \U$31427 ( \31742 , \31737 , \31741 );
and \U$31428 ( \31743 , \22030 , \22392 );
and \U$31429 ( \31744 , \22001 , \22390 );
nor \U$31430 ( \31745 , \31743 , \31744 );
xnor \U$31431 ( \31746 , \31745 , \22402 );
xor \U$31432 ( \31747 , \31742 , \31746 );
and \U$31433 ( \31748 , \22224 , \22619 );
and \U$31434 ( \31749 , \22235 , \22617 );
nor \U$31435 ( \31750 , \31748 , \31749 );
xnor \U$31436 ( \31751 , \31750 , \22629 );
and \U$31437 ( \31752 , \22251 , \22641 );
and \U$31438 ( \31753 , \22262 , \22639 );
nor \U$31439 ( \31754 , \31752 , \31753 );
xnor \U$31440 ( \31755 , \31754 , \22651 );
xor \U$31441 ( \31756 , \31751 , \31755 );
and \U$31442 ( \31757 , \22272 , \22671 );
and \U$31443 ( \31758 , \22283 , \22669 );
nor \U$31444 ( \31759 , \31757 , \31758 );
xnor \U$31445 ( \31760 , \31759 , \22681 );
xor \U$31446 ( \31761 , \31756 , \31760 );
and \U$31447 ( \31762 , \22156 , \22551 );
and \U$31448 ( \31763 , \22167 , \22549 );
nor \U$31449 ( \31764 , \31762 , \31763 );
xnor \U$31450 ( \31765 , \31764 , \22561 );
and \U$31451 ( \31766 , \22181 , \22573 );
and \U$31452 ( \31767 , \22192 , \22571 );
nor \U$31453 ( \31768 , \31766 , \31767 );
xnor \U$31454 ( \31769 , \31768 , \22583 );
xor \U$31455 ( \31770 , \31765 , \31769 );
and \U$31456 ( \31771 , \22202 , \22598 );
and \U$31457 ( \31772 , \22213 , \22596 );
nor \U$31458 ( \31773 , \31771 , \31772 );
xnor \U$31459 ( \31774 , \31773 , \22608 );
xor \U$31460 ( \31775 , \31770 , \31774 );
xor \U$31461 ( \31776 , \31761 , \31775 );
and \U$31462 ( \31777 , \22089 , \22484 );
and \U$31463 ( \31778 , \22100 , \22482 );
nor \U$31464 ( \31779 , \31777 , \31778 );
xnor \U$31465 ( \31780 , \31779 , \22494 );
and \U$31466 ( \31781 , \22113 , \22506 );
and \U$31467 ( \31782 , \22124 , \22504 );
nor \U$31468 ( \31783 , \31781 , \31782 );
xnor \U$31469 ( \31784 , \31783 , \22516 );
xor \U$31470 ( \31785 , \31780 , \31784 );
and \U$31471 ( \31786 , \22134 , \22530 );
and \U$31472 ( \31787 , \22145 , \22528 );
nor \U$31473 ( \31788 , \31786 , \31787 );
xnor \U$31474 ( \31789 , \31788 , \22540 );
xor \U$31475 ( \31790 , \31785 , \31789 );
xor \U$31476 ( \31791 , \31776 , \31790 );
xor \U$31477 ( \31792 , \31747 , \31791 );
and \U$31478 ( \31793 , \31598 , \31602 );
and \U$31479 ( \31794 , \31602 , \31604 );
and \U$31480 ( \31795 , \31598 , \31604 );
or \U$31481 ( \31796 , \31793 , \31794 , \31795 );
and \U$31482 ( \31797 , \22361 , \22021 );
and \U$31483 ( \31798 , \22372 , \22019 );
nor \U$31484 ( \31799 , \31797 , \31798 );
xnor \U$31485 ( \31800 , \31799 , \21595 );
and \U$31486 ( \31801 , \22386 , \21983 );
and \U$31487 ( \31802 , \22397 , \21981 );
nor \U$31488 ( \31803 , \31801 , \31802 );
xnor \U$31489 ( \31804 , \31803 , \21995 );
xor \U$31490 ( \31805 , \31800 , \31804 );
and \U$31491 ( \31806 , \22418 , \21978 );
xor \U$31492 ( \31807 , \31805 , \31806 );
xor \U$31493 ( \31808 , \31796 , \31807 );
and \U$31494 ( \31809 , \22294 , \22691 );
and \U$31495 ( \31810 , \22305 , \22689 );
nor \U$31496 ( \31811 , \31809 , \31810 );
xnor \U$31497 ( \31812 , \31811 , \22701 );
and \U$31498 ( \31813 , \22318 , \22720 );
and \U$31499 ( \31814 , \22329 , \22707 );
nor \U$31500 ( \31815 , \31813 , \31814 );
xnor \U$31501 ( \31816 , \31815 , \22067 );
xor \U$31502 ( \31817 , \31812 , \31816 );
and \U$31503 ( \31818 , \22339 , \23173 );
and \U$31504 ( \31819 , \22350 , \22999 );
nor \U$31505 ( \31820 , \31818 , \31819 );
xnor \U$31506 ( \31821 , \31820 , \22016 );
xor \U$31507 ( \31822 , \31817 , \31821 );
xor \U$31508 ( \31823 , \31808 , \31822 );
xor \U$31509 ( \31824 , \31792 , \31823 );
xor \U$31510 ( \31825 , \31736 , \31824 );
xor \U$31511 ( \31826 , \31707 , \31825 );
and \U$31512 ( \31827 , \31510 , \31514 );
and \U$31513 ( \31828 , \31514 , \31519 );
and \U$31514 ( \31829 , \31510 , \31519 );
or \U$31515 ( \31830 , \31827 , \31828 , \31829 );
and \U$31516 ( \31831 , \31627 , \31631 );
and \U$31517 ( \31832 , \31631 , \31675 );
and \U$31518 ( \31833 , \31627 , \31675 );
or \U$31519 ( \31834 , \31831 , \31832 , \31833 );
xor \U$31520 ( \31835 , \31830 , \31834 );
and \U$31521 ( \31836 , \31590 , \31606 );
and \U$31522 ( \31837 , \31606 , \31621 );
and \U$31523 ( \31838 , \31590 , \31621 );
or \U$31524 ( \31839 , \31836 , \31837 , \31838 );
xor \U$31525 ( \31840 , \31835 , \31839 );
xor \U$31526 ( \31841 , \31826 , \31840 );
xor \U$31527 ( \31842 , \31696 , \31841 );
and \U$31528 ( \31843 , \31487 , \31491 );
and \U$31529 ( \31844 , \31491 , \31496 );
and \U$31530 ( \31845 , \31487 , \31496 );
or \U$31531 ( \31846 , \31843 , \31844 , \31845 );
and \U$31532 ( \31847 , \31546 , \31622 );
and \U$31533 ( \31848 , \31622 , \31676 );
and \U$31534 ( \31849 , \31546 , \31676 );
or \U$31535 ( \31850 , \31847 , \31848 , \31849 );
xor \U$31536 ( \31851 , \31846 , \31850 );
and \U$31537 ( \31852 , \31560 , \31574 );
and \U$31538 ( \31853 , \31574 , \31589 );
and \U$31539 ( \31854 , \31560 , \31589 );
or \U$31540 ( \31855 , \31852 , \31853 , \31854 );
and \U$31541 ( \31856 , \31646 , \31660 );
and \U$31542 ( \31857 , \31660 , \31674 );
and \U$31543 ( \31858 , \31646 , \31674 );
or \U$31544 ( \31859 , \31856 , \31857 , \31858 );
xor \U$31545 ( \31860 , \31855 , \31859 );
and \U$31546 ( \31861 , \23230 , \22413 );
and \U$31547 ( \31862 , \23329 , \22411 );
nor \U$31548 ( \31863 , \31861 , \31862 );
xnor \U$31549 ( \31864 , \31863 , \22423 );
and \U$31550 ( \31865 , \22858 , \22435 );
and \U$31551 ( \31866 , \22894 , \22433 );
nor \U$31552 ( \31867 , \31865 , \31866 );
xnor \U$31553 ( \31868 , \31867 , \22445 );
xor \U$31554 ( \31869 , \31864 , \31868 );
and \U$31555 ( \31870 , \22071 , \22463 );
and \U$31556 ( \31871 , \22081 , \22461 );
nor \U$31557 ( \31872 , \31870 , \31871 );
xnor \U$31558 ( \31873 , \31872 , \22473 );
xor \U$31559 ( \31874 , \31869 , \31873 );
xor \U$31560 ( \31875 , \31860 , \31874 );
xor \U$31561 ( \31876 , \31851 , \31875 );
xor \U$31562 ( \31877 , \31842 , \31876 );
xor \U$31563 ( \31878 , \31692 , \31877 );
xor \U$31564 ( \31879 , \31686 , \31878 );
and \U$31565 ( \31880 , \31479 , \31679 );
nor \U$31566 ( \31881 , \31879 , \31880 );
nor \U$31567 ( \31882 , \31682 , \31881 );
nand \U$31568 ( \31883 , \31475 , \31882 );
and \U$31569 ( \31884 , \31690 , \31691 );
and \U$31570 ( \31885 , \31691 , \31877 );
and \U$31571 ( \31886 , \31690 , \31877 );
or \U$31572 ( \31887 , \31884 , \31885 , \31886 );
and \U$31573 ( \31888 , \31696 , \31841 );
and \U$31574 ( \31889 , \31841 , \31876 );
and \U$31575 ( \31890 , \31696 , \31876 );
or \U$31576 ( \31891 , \31888 , \31889 , \31890 );
and \U$31577 ( \31892 , \31830 , \31834 );
and \U$31578 ( \31893 , \31834 , \31839 );
and \U$31579 ( \31894 , \31830 , \31839 );
or \U$31580 ( \31895 , \31892 , \31893 , \31894 );
and \U$31581 ( \31896 , \31721 , \31735 );
and \U$31582 ( \31897 , \31735 , \31824 );
and \U$31583 ( \31898 , \31721 , \31824 );
or \U$31584 ( \31899 , \31896 , \31897 , \31898 );
xor \U$31585 ( \31900 , \31895 , \31899 );
and \U$31586 ( \31901 , \31800 , \31804 );
and \U$31587 ( \31902 , \31804 , \31806 );
and \U$31588 ( \31903 , \31800 , \31806 );
or \U$31589 ( \31904 , \31901 , \31902 , \31903 );
and \U$31590 ( \31905 , \22397 , \21983 );
and \U$31591 ( \31906 , \22361 , \21981 );
nor \U$31592 ( \31907 , \31905 , \31906 );
xnor \U$31593 ( \31908 , \31907 , \21995 );
and \U$31594 ( \31909 , \22386 , \21978 );
xnor \U$31595 ( \31910 , \31908 , \31909 );
xor \U$31596 ( \31911 , \31904 , \31910 );
and \U$31597 ( \31912 , \22329 , \22720 );
and \U$31598 ( \31913 , \22294 , \22707 );
nor \U$31599 ( \31914 , \31912 , \31913 );
xnor \U$31600 ( \31915 , \31914 , \22067 );
and \U$31601 ( \31916 , \22350 , \23173 );
and \U$31602 ( \31917 , \22318 , \22999 );
nor \U$31603 ( \31918 , \31916 , \31917 );
xnor \U$31604 ( \31919 , \31918 , \22016 );
xor \U$31605 ( \31920 , \31915 , \31919 );
and \U$31606 ( \31921 , \22372 , \22021 );
and \U$31607 ( \31922 , \22339 , \22019 );
nor \U$31608 ( \31923 , \31921 , \31922 );
xnor \U$31609 ( \31924 , \31923 , \21595 );
xor \U$31610 ( \31925 , \31920 , \31924 );
xor \U$31611 ( \31926 , \31911 , \31925 );
and \U$31612 ( \31927 , \31765 , \31769 );
and \U$31613 ( \31928 , \31769 , \31774 );
and \U$31614 ( \31929 , \31765 , \31774 );
or \U$31615 ( \31930 , \31927 , \31928 , \31929 );
and \U$31616 ( \31931 , \31751 , \31755 );
and \U$31617 ( \31932 , \31755 , \31760 );
and \U$31618 ( \31933 , \31751 , \31760 );
or \U$31619 ( \31934 , \31931 , \31932 , \31933 );
xor \U$31620 ( \31935 , \31930 , \31934 );
and \U$31621 ( \31936 , \31812 , \31816 );
and \U$31622 ( \31937 , \31816 , \31821 );
and \U$31623 ( \31938 , \31812 , \31821 );
or \U$31624 ( \31939 , \31936 , \31937 , \31938 );
xor \U$31625 ( \31940 , \31935 , \31939 );
xor \U$31626 ( \31941 , \31926 , \31940 );
and \U$31627 ( \31942 , \31737 , \31741 );
and \U$31628 ( \31943 , \31741 , \31746 );
and \U$31629 ( \31944 , \31737 , \31746 );
or \U$31630 ( \31945 , \31942 , \31943 , \31944 );
and \U$31631 ( \31946 , \31864 , \31868 );
and \U$31632 ( \31947 , \31868 , \31873 );
and \U$31633 ( \31948 , \31864 , \31873 );
or \U$31634 ( \31949 , \31946 , \31947 , \31948 );
xor \U$31635 ( \31950 , \31945 , \31949 );
and \U$31636 ( \31951 , \31780 , \31784 );
and \U$31637 ( \31952 , \31784 , \31789 );
and \U$31638 ( \31953 , \31780 , \31789 );
or \U$31639 ( \31954 , \31951 , \31952 , \31953 );
xor \U$31640 ( \31955 , \31950 , \31954 );
xor \U$31641 ( \31956 , \31941 , \31955 );
and \U$31642 ( \31957 , \31761 , \31775 );
and \U$31643 ( \31958 , \31775 , \31790 );
and \U$31644 ( \31959 , \31761 , \31790 );
or \U$31645 ( \31960 , \31957 , \31958 , \31959 );
and \U$31646 ( \31961 , \22894 , \22435 );
and \U$31647 ( \31962 , \23230 , \22433 );
nor \U$31648 ( \31963 , \31961 , \31962 );
xnor \U$31649 ( \31964 , \31963 , \22445 );
and \U$31650 ( \31965 , \22081 , \22463 );
and \U$31651 ( \31966 , \22858 , \22461 );
nor \U$31652 ( \31967 , \31965 , \31966 );
xnor \U$31653 ( \31968 , \31967 , \22473 );
xor \U$31654 ( \31969 , \31964 , \31968 );
and \U$31655 ( \31970 , \22100 , \22484 );
and \U$31656 ( \31971 , \22071 , \22482 );
nor \U$31657 ( \31972 , \31970 , \31971 );
xnor \U$31658 ( \31973 , \31972 , \22494 );
xor \U$31659 ( \31974 , \31969 , \31973 );
and \U$31660 ( \31975 , \21990 , \22367 );
not \U$31661 ( \31976 , \31975 );
xnor \U$31662 ( \31977 , \31976 , \22377 );
and \U$31663 ( \31978 , \22001 , \22392 );
and \U$31664 ( \31979 , \21977 , \22390 );
nor \U$31665 ( \31980 , \31978 , \31979 );
xnor \U$31666 ( \31981 , \31980 , \22402 );
xor \U$31667 ( \31982 , \31977 , \31981 );
and \U$31668 ( \31983 , \23329 , \22413 );
and \U$31669 ( \31984 , \22030 , \22411 );
nor \U$31670 ( \31985 , \31983 , \31984 );
xnor \U$31671 ( \31986 , \31985 , \22423 );
xor \U$31672 ( \31987 , \31982 , \31986 );
xor \U$31673 ( \31988 , \31974 , \31987 );
xor \U$31674 ( \31989 , \31960 , \31988 );
and \U$31675 ( \31990 , \22262 , \22641 );
and \U$31676 ( \31991 , \22224 , \22639 );
nor \U$31677 ( \31992 , \31990 , \31991 );
xnor \U$31678 ( \31993 , \31992 , \22651 );
and \U$31679 ( \31994 , \22283 , \22671 );
and \U$31680 ( \31995 , \22251 , \22669 );
nor \U$31681 ( \31996 , \31994 , \31995 );
xnor \U$31682 ( \31997 , \31996 , \22681 );
xor \U$31683 ( \31998 , \31993 , \31997 );
and \U$31684 ( \31999 , \22305 , \22691 );
and \U$31685 ( \32000 , \22272 , \22689 );
nor \U$31686 ( \32001 , \31999 , \32000 );
xnor \U$31687 ( \32002 , \32001 , \22701 );
xor \U$31688 ( \32003 , \31998 , \32002 );
and \U$31689 ( \32004 , \22192 , \22573 );
and \U$31690 ( \32005 , \22156 , \22571 );
nor \U$31691 ( \32006 , \32004 , \32005 );
xnor \U$31692 ( \32007 , \32006 , \22583 );
and \U$31693 ( \32008 , \22213 , \22598 );
and \U$31694 ( \32009 , \22181 , \22596 );
nor \U$31695 ( \32010 , \32008 , \32009 );
xnor \U$31696 ( \32011 , \32010 , \22608 );
xor \U$31697 ( \32012 , \32007 , \32011 );
and \U$31698 ( \32013 , \22235 , \22619 );
and \U$31699 ( \32014 , \22202 , \22617 );
nor \U$31700 ( \32015 , \32013 , \32014 );
xnor \U$31701 ( \32016 , \32015 , \22629 );
xor \U$31702 ( \32017 , \32012 , \32016 );
xor \U$31703 ( \32018 , \32003 , \32017 );
and \U$31704 ( \32019 , \22124 , \22506 );
and \U$31705 ( \32020 , \22089 , \22504 );
nor \U$31706 ( \32021 , \32019 , \32020 );
xnor \U$31707 ( \32022 , \32021 , \22516 );
and \U$31708 ( \32023 , \22145 , \22530 );
and \U$31709 ( \32024 , \22113 , \22528 );
nor \U$31710 ( \32025 , \32023 , \32024 );
xnor \U$31711 ( \32026 , \32025 , \22540 );
xor \U$31712 ( \32027 , \32022 , \32026 );
and \U$31713 ( \32028 , \22167 , \22551 );
and \U$31714 ( \32029 , \22134 , \22549 );
nor \U$31715 ( \32030 , \32028 , \32029 );
xnor \U$31716 ( \32031 , \32030 , \22561 );
xor \U$31717 ( \32032 , \32027 , \32031 );
xor \U$31718 ( \32033 , \32018 , \32032 );
xor \U$31719 ( \32034 , \31989 , \32033 );
xor \U$31720 ( \32035 , \31956 , \32034 );
and \U$31721 ( \32036 , \31725 , \31729 );
and \U$31722 ( \32037 , \31729 , \31734 );
and \U$31723 ( \32038 , \31725 , \31734 );
or \U$31724 ( \32039 , \32036 , \32037 , \32038 );
and \U$31725 ( \32040 , \31711 , \31715 );
and \U$31726 ( \32041 , \31715 , \31720 );
and \U$31727 ( \32042 , \31711 , \31720 );
or \U$31728 ( \32043 , \32040 , \32041 , \32042 );
xor \U$31729 ( \32044 , \32039 , \32043 );
and \U$31730 ( \32045 , \31796 , \31807 );
and \U$31731 ( \32046 , \31807 , \31822 );
and \U$31732 ( \32047 , \31796 , \31822 );
or \U$31733 ( \32048 , \32045 , \32046 , \32047 );
xor \U$31734 ( \32049 , \32044 , \32048 );
xor \U$31735 ( \32050 , \32035 , \32049 );
xor \U$31736 ( \32051 , \31900 , \32050 );
xor \U$31737 ( \32052 , \31891 , \32051 );
and \U$31738 ( \32053 , \31846 , \31850 );
and \U$31739 ( \32054 , \31850 , \31875 );
and \U$31740 ( \32055 , \31846 , \31875 );
or \U$31741 ( \32056 , \32053 , \32054 , \32055 );
and \U$31742 ( \32057 , \31707 , \31825 );
and \U$31743 ( \32058 , \31825 , \31840 );
and \U$31744 ( \32059 , \31707 , \31840 );
or \U$31745 ( \32060 , \32057 , \32058 , \32059 );
xor \U$31746 ( \32061 , \32056 , \32060 );
and \U$31747 ( \32062 , \31700 , \31704 );
and \U$31748 ( \32063 , \31704 , \31706 );
and \U$31749 ( \32064 , \31700 , \31706 );
or \U$31750 ( \32065 , \32062 , \32063 , \32064 );
and \U$31751 ( \32066 , \31855 , \31859 );
and \U$31752 ( \32067 , \31859 , \31874 );
and \U$31753 ( \32068 , \31855 , \31874 );
or \U$31754 ( \32069 , \32066 , \32067 , \32068 );
xor \U$31755 ( \32070 , \32065 , \32069 );
and \U$31756 ( \32071 , \31747 , \31791 );
and \U$31757 ( \32072 , \31791 , \31823 );
and \U$31758 ( \32073 , \31747 , \31823 );
or \U$31759 ( \32074 , \32071 , \32072 , \32073 );
xor \U$31760 ( \32075 , \32070 , \32074 );
xor \U$31761 ( \32076 , \32061 , \32075 );
xor \U$31762 ( \32077 , \32052 , \32076 );
xor \U$31763 ( \32078 , \31887 , \32077 );
and \U$31764 ( \32079 , \31686 , \31878 );
nor \U$31765 ( \32080 , \32078 , \32079 );
and \U$31766 ( \32081 , \31891 , \32051 );
and \U$31767 ( \32082 , \32051 , \32076 );
and \U$31768 ( \32083 , \31891 , \32076 );
or \U$31769 ( \32084 , \32081 , \32082 , \32083 );
and \U$31770 ( \32085 , \32056 , \32060 );
and \U$31771 ( \32086 , \32060 , \32075 );
and \U$31772 ( \32087 , \32056 , \32075 );
or \U$31773 ( \32088 , \32085 , \32086 , \32087 );
xor \U$31774 ( \32089 , \32084 , \32088 );
and \U$31775 ( \32090 , \31895 , \31899 );
and \U$31776 ( \32091 , \31899 , \32050 );
and \U$31777 ( \32092 , \31895 , \32050 );
or \U$31778 ( \32093 , \32090 , \32091 , \32092 );
and \U$31779 ( \32094 , \31977 , \31981 );
and \U$31780 ( \32095 , \31981 , \31986 );
and \U$31781 ( \32096 , \31977 , \31986 );
or \U$31782 ( \32097 , \32094 , \32095 , \32096 );
and \U$31783 ( \32098 , \31964 , \31968 );
and \U$31784 ( \32099 , \31968 , \31973 );
and \U$31785 ( \32100 , \31964 , \31973 );
or \U$31786 ( \32101 , \32098 , \32099 , \32100 );
xor \U$31787 ( \32102 , \32097 , \32101 );
and \U$31788 ( \32103 , \32022 , \32026 );
and \U$31789 ( \32104 , \32026 , \32031 );
and \U$31790 ( \32105 , \32022 , \32031 );
or \U$31791 ( \32106 , \32103 , \32104 , \32105 );
xor \U$31792 ( \32107 , \32102 , \32106 );
and \U$31793 ( \32108 , \22294 , \22720 );
and \U$31794 ( \32109 , \22305 , \22707 );
nor \U$31795 ( \32110 , \32108 , \32109 );
xnor \U$31796 ( \32111 , \32110 , \22067 );
and \U$31797 ( \32112 , \22318 , \23173 );
and \U$31798 ( \32113 , \22329 , \22999 );
nor \U$31799 ( \32114 , \32112 , \32113 );
xnor \U$31800 ( \32115 , \32114 , \22016 );
xor \U$31801 ( \32116 , \32111 , \32115 );
and \U$31802 ( \32117 , \22339 , \22021 );
and \U$31803 ( \32118 , \22350 , \22019 );
nor \U$31804 ( \32119 , \32117 , \32118 );
xnor \U$31805 ( \32120 , \32119 , \21595 );
xor \U$31806 ( \32121 , \32116 , \32120 );
and \U$31807 ( \32122 , \22224 , \22641 );
and \U$31808 ( \32123 , \22235 , \22639 );
nor \U$31809 ( \32124 , \32122 , \32123 );
xnor \U$31810 ( \32125 , \32124 , \22651 );
and \U$31811 ( \32126 , \22251 , \22671 );
and \U$31812 ( \32127 , \22262 , \22669 );
nor \U$31813 ( \32128 , \32126 , \32127 );
xnor \U$31814 ( \32129 , \32128 , \22681 );
xor \U$31815 ( \32130 , \32125 , \32129 );
and \U$31816 ( \32131 , \22272 , \22691 );
and \U$31817 ( \32132 , \22283 , \22689 );
nor \U$31818 ( \32133 , \32131 , \32132 );
xnor \U$31819 ( \32134 , \32133 , \22701 );
xor \U$31820 ( \32135 , \32130 , \32134 );
xor \U$31821 ( \32136 , \32121 , \32135 );
and \U$31822 ( \32137 , \22156 , \22573 );
and \U$31823 ( \32138 , \22167 , \22571 );
nor \U$31824 ( \32139 , \32137 , \32138 );
xnor \U$31825 ( \32140 , \32139 , \22583 );
and \U$31826 ( \32141 , \22181 , \22598 );
and \U$31827 ( \32142 , \22192 , \22596 );
nor \U$31828 ( \32143 , \32141 , \32142 );
xnor \U$31829 ( \32144 , \32143 , \22608 );
xor \U$31830 ( \32145 , \32140 , \32144 );
and \U$31831 ( \32146 , \22202 , \22619 );
and \U$31832 ( \32147 , \22213 , \22617 );
nor \U$31833 ( \32148 , \32146 , \32147 );
xnor \U$31834 ( \32149 , \32148 , \22629 );
xor \U$31835 ( \32150 , \32145 , \32149 );
xor \U$31836 ( \32151 , \32136 , \32150 );
or \U$31837 ( \32152 , \31908 , \31909 );
and \U$31838 ( \32153 , \22361 , \21983 );
and \U$31839 ( \32154 , \22372 , \21981 );
nor \U$31840 ( \32155 , \32153 , \32154 );
xnor \U$31841 ( \32156 , \32155 , \21995 );
xor \U$31842 ( \32157 , \32152 , \32156 );
and \U$31843 ( \32158 , \22397 , \21978 );
xor \U$31844 ( \32159 , \32157 , \32158 );
xor \U$31845 ( \32160 , \32151 , \32159 );
and \U$31846 ( \32161 , \32007 , \32011 );
and \U$31847 ( \32162 , \32011 , \32016 );
and \U$31848 ( \32163 , \32007 , \32016 );
or \U$31849 ( \32164 , \32161 , \32162 , \32163 );
and \U$31850 ( \32165 , \31993 , \31997 );
and \U$31851 ( \32166 , \31997 , \32002 );
and \U$31852 ( \32167 , \31993 , \32002 );
or \U$31853 ( \32168 , \32165 , \32166 , \32167 );
xor \U$31854 ( \32169 , \32164 , \32168 );
and \U$31855 ( \32170 , \31915 , \31919 );
and \U$31856 ( \32171 , \31919 , \31924 );
and \U$31857 ( \32172 , \31915 , \31924 );
or \U$31858 ( \32173 , \32170 , \32171 , \32172 );
xor \U$31859 ( \32174 , \32169 , \32173 );
xor \U$31860 ( \32175 , \32160 , \32174 );
xor \U$31861 ( \32176 , \32107 , \32175 );
and \U$31862 ( \32177 , \32003 , \32017 );
and \U$31863 ( \32178 , \32017 , \32032 );
and \U$31864 ( \32179 , \32003 , \32032 );
or \U$31865 ( \32180 , \32177 , \32178 , \32179 );
and \U$31866 ( \32181 , \31974 , \31987 );
xor \U$31867 ( \32182 , \32180 , \32181 );
and \U$31868 ( \32183 , \22089 , \22506 );
and \U$31869 ( \32184 , \22100 , \22504 );
nor \U$31870 ( \32185 , \32183 , \32184 );
xnor \U$31871 ( \32186 , \32185 , \22516 );
and \U$31872 ( \32187 , \22113 , \22530 );
and \U$31873 ( \32188 , \22124 , \22528 );
nor \U$31874 ( \32189 , \32187 , \32188 );
xnor \U$31875 ( \32190 , \32189 , \22540 );
xor \U$31876 ( \32191 , \32186 , \32190 );
and \U$31877 ( \32192 , \22134 , \22551 );
and \U$31878 ( \32193 , \22145 , \22549 );
nor \U$31879 ( \32194 , \32192 , \32193 );
xnor \U$31880 ( \32195 , \32194 , \22561 );
xor \U$31881 ( \32196 , \32191 , \32195 );
and \U$31882 ( \32197 , \23230 , \22435 );
and \U$31883 ( \32198 , \23329 , \22433 );
nor \U$31884 ( \32199 , \32197 , \32198 );
xnor \U$31885 ( \32200 , \32199 , \22445 );
and \U$31886 ( \32201 , \22858 , \22463 );
and \U$31887 ( \32202 , \22894 , \22461 );
nor \U$31888 ( \32203 , \32201 , \32202 );
xnor \U$31889 ( \32204 , \32203 , \22473 );
xor \U$31890 ( \32205 , \32200 , \32204 );
and \U$31891 ( \32206 , \22071 , \22484 );
and \U$31892 ( \32207 , \22081 , \22482 );
nor \U$31893 ( \32208 , \32206 , \32207 );
xnor \U$31894 ( \32209 , \32208 , \22494 );
xor \U$31895 ( \32210 , \32205 , \32209 );
xor \U$31896 ( \32211 , \32196 , \32210 );
not \U$31897 ( \32212 , \22377 );
and \U$31898 ( \32213 , \21977 , \22392 );
and \U$31899 ( \32214 , \21990 , \22390 );
nor \U$31900 ( \32215 , \32213 , \32214 );
xnor \U$31901 ( \32216 , \32215 , \22402 );
xor \U$31902 ( \32217 , \32212 , \32216 );
and \U$31903 ( \32218 , \22030 , \22413 );
and \U$31904 ( \32219 , \22001 , \22411 );
nor \U$31905 ( \32220 , \32218 , \32219 );
xnor \U$31906 ( \32221 , \32220 , \22423 );
xor \U$31907 ( \32222 , \32217 , \32221 );
xor \U$31908 ( \32223 , \32211 , \32222 );
xor \U$31909 ( \32224 , \32182 , \32223 );
xor \U$31910 ( \32225 , \32176 , \32224 );
and \U$31911 ( \32226 , \32039 , \32043 );
and \U$31912 ( \32227 , \32043 , \32048 );
and \U$31913 ( \32228 , \32039 , \32048 );
or \U$31914 ( \32229 , \32226 , \32227 , \32228 );
and \U$31915 ( \32230 , \31960 , \31988 );
and \U$31916 ( \32231 , \31988 , \32033 );
and \U$31917 ( \32232 , \31960 , \32033 );
or \U$31918 ( \32233 , \32230 , \32231 , \32232 );
xor \U$31919 ( \32234 , \32229 , \32233 );
and \U$31920 ( \32235 , \31926 , \31940 );
and \U$31921 ( \32236 , \31940 , \31955 );
and \U$31922 ( \32237 , \31926 , \31955 );
or \U$31923 ( \32238 , \32235 , \32236 , \32237 );
xor \U$31924 ( \32239 , \32234 , \32238 );
xor \U$31925 ( \32240 , \32225 , \32239 );
xor \U$31926 ( \32241 , \32093 , \32240 );
and \U$31927 ( \32242 , \32065 , \32069 );
and \U$31928 ( \32243 , \32069 , \32074 );
and \U$31929 ( \32244 , \32065 , \32074 );
or \U$31930 ( \32245 , \32242 , \32243 , \32244 );
and \U$31931 ( \32246 , \31956 , \32034 );
and \U$31932 ( \32247 , \32034 , \32049 );
and \U$31933 ( \32248 , \31956 , \32049 );
or \U$31934 ( \32249 , \32246 , \32247 , \32248 );
xor \U$31935 ( \32250 , \32245 , \32249 );
and \U$31936 ( \32251 , \31945 , \31949 );
and \U$31937 ( \32252 , \31949 , \31954 );
and \U$31938 ( \32253 , \31945 , \31954 );
or \U$31939 ( \32254 , \32251 , \32252 , \32253 );
and \U$31940 ( \32255 , \31930 , \31934 );
and \U$31941 ( \32256 , \31934 , \31939 );
and \U$31942 ( \32257 , \31930 , \31939 );
or \U$31943 ( \32258 , \32255 , \32256 , \32257 );
xor \U$31944 ( \32259 , \32254 , \32258 );
and \U$31945 ( \32260 , \31904 , \31910 );
and \U$31946 ( \32261 , \31910 , \31925 );
and \U$31947 ( \32262 , \31904 , \31925 );
or \U$31948 ( \32263 , \32260 , \32261 , \32262 );
xor \U$31949 ( \32264 , \32259 , \32263 );
xor \U$31950 ( \32265 , \32250 , \32264 );
xor \U$31951 ( \32266 , \32241 , \32265 );
xor \U$31952 ( \32267 , \32089 , \32266 );
and \U$31953 ( \32268 , \31887 , \32077 );
nor \U$31954 ( \32269 , \32267 , \32268 );
nor \U$31955 ( \32270 , \32080 , \32269 );
and \U$31956 ( \32271 , \32093 , \32240 );
and \U$31957 ( \32272 , \32240 , \32265 );
and \U$31958 ( \32273 , \32093 , \32265 );
or \U$31959 ( \32274 , \32271 , \32272 , \32273 );
and \U$31960 ( \32275 , \32229 , \32233 );
and \U$31961 ( \32276 , \32233 , \32238 );
and \U$31962 ( \32277 , \32229 , \32238 );
or \U$31963 ( \32278 , \32275 , \32276 , \32277 );
and \U$31964 ( \32279 , \32107 , \32175 );
and \U$31965 ( \32280 , \32175 , \32224 );
and \U$31966 ( \32281 , \32107 , \32224 );
or \U$31967 ( \32282 , \32279 , \32280 , \32281 );
xor \U$31968 ( \32283 , \32278 , \32282 );
and \U$31969 ( \32284 , \32121 , \32135 );
and \U$31970 ( \32285 , \32135 , \32150 );
and \U$31971 ( \32286 , \32121 , \32150 );
or \U$31972 ( \32287 , \32284 , \32285 , \32286 );
and \U$31973 ( \32288 , \32196 , \32210 );
and \U$31974 ( \32289 , \32210 , \32222 );
and \U$31975 ( \32290 , \32196 , \32222 );
or \U$31976 ( \32291 , \32288 , \32289 , \32290 );
xor \U$31977 ( \32292 , \32287 , \32291 );
and \U$31978 ( \32293 , \22894 , \22463 );
and \U$31979 ( \32294 , \23230 , \22461 );
nor \U$31980 ( \32295 , \32293 , \32294 );
xnor \U$31981 ( \32296 , \32295 , \22473 );
and \U$31982 ( \32297 , \22081 , \22484 );
and \U$31983 ( \32298 , \22858 , \22482 );
nor \U$31984 ( \32299 , \32297 , \32298 );
xnor \U$31985 ( \32300 , \32299 , \22494 );
xor \U$31986 ( \32301 , \32296 , \32300 );
and \U$31987 ( \32302 , \22100 , \22506 );
and \U$31988 ( \32303 , \22071 , \22504 );
nor \U$31989 ( \32304 , \32302 , \32303 );
xnor \U$31990 ( \32305 , \32304 , \22516 );
xor \U$31991 ( \32306 , \32301 , \32305 );
xor \U$31992 ( \32307 , \32292 , \32306 );
xor \U$31993 ( \32308 , \32283 , \32307 );
xor \U$31994 ( \32309 , \32274 , \32308 );
and \U$31995 ( \32310 , \32245 , \32249 );
and \U$31996 ( \32311 , \32249 , \32264 );
and \U$31997 ( \32312 , \32245 , \32264 );
or \U$31998 ( \32313 , \32310 , \32311 , \32312 );
and \U$31999 ( \32314 , \32225 , \32239 );
xor \U$32000 ( \32315 , \32313 , \32314 );
and \U$32001 ( \32316 , \32097 , \32101 );
and \U$32002 ( \32317 , \32101 , \32106 );
and \U$32003 ( \32318 , \32097 , \32106 );
or \U$32004 ( \32319 , \32316 , \32317 , \32318 );
and \U$32005 ( \32320 , \32164 , \32168 );
and \U$32006 ( \32321 , \32168 , \32173 );
and \U$32007 ( \32322 , \32164 , \32173 );
or \U$32008 ( \32323 , \32320 , \32321 , \32322 );
xor \U$32009 ( \32324 , \32319 , \32323 );
and \U$32010 ( \32325 , \32152 , \32156 );
and \U$32011 ( \32326 , \32156 , \32158 );
and \U$32012 ( \32327 , \32152 , \32158 );
or \U$32013 ( \32328 , \32325 , \32326 , \32327 );
xor \U$32014 ( \32329 , \32324 , \32328 );
and \U$32015 ( \32330 , \32140 , \32144 );
and \U$32016 ( \32331 , \32144 , \32149 );
and \U$32017 ( \32332 , \32140 , \32149 );
or \U$32018 ( \32333 , \32330 , \32331 , \32332 );
and \U$32019 ( \32334 , \32125 , \32129 );
and \U$32020 ( \32335 , \32129 , \32134 );
and \U$32021 ( \32336 , \32125 , \32134 );
or \U$32022 ( \32337 , \32334 , \32335 , \32336 );
xor \U$32023 ( \32338 , \32333 , \32337 );
and \U$32024 ( \32339 , \32111 , \32115 );
and \U$32025 ( \32340 , \32115 , \32120 );
and \U$32026 ( \32341 , \32111 , \32120 );
or \U$32027 ( \32342 , \32339 , \32340 , \32341 );
xor \U$32028 ( \32343 , \32338 , \32342 );
and \U$32029 ( \32344 , \32212 , \32216 );
and \U$32030 ( \32345 , \32216 , \32221 );
and \U$32031 ( \32346 , \32212 , \32221 );
or \U$32032 ( \32347 , \32344 , \32345 , \32346 );
and \U$32033 ( \32348 , \32200 , \32204 );
and \U$32034 ( \32349 , \32204 , \32209 );
and \U$32035 ( \32350 , \32200 , \32209 );
or \U$32036 ( \32351 , \32348 , \32349 , \32350 );
xor \U$32037 ( \32352 , \32347 , \32351 );
and \U$32038 ( \32353 , \32186 , \32190 );
and \U$32039 ( \32354 , \32190 , \32195 );
and \U$32040 ( \32355 , \32186 , \32195 );
or \U$32041 ( \32356 , \32353 , \32354 , \32355 );
xor \U$32042 ( \32357 , \32352 , \32356 );
xor \U$32043 ( \32358 , \32343 , \32357 );
and \U$32044 ( \32359 , \21990 , \22392 );
not \U$32045 ( \32360 , \32359 );
xnor \U$32046 ( \32361 , \32360 , \22402 );
and \U$32047 ( \32362 , \22001 , \22413 );
and \U$32048 ( \32363 , \21977 , \22411 );
nor \U$32049 ( \32364 , \32362 , \32363 );
xnor \U$32050 ( \32365 , \32364 , \22423 );
xor \U$32051 ( \32366 , \32361 , \32365 );
and \U$32052 ( \32367 , \23329 , \22435 );
and \U$32053 ( \32368 , \22030 , \22433 );
nor \U$32054 ( \32369 , \32367 , \32368 );
xnor \U$32055 ( \32370 , \32369 , \22445 );
xor \U$32056 ( \32371 , \32366 , \32370 );
and \U$32057 ( \32372 , \22262 , \22671 );
and \U$32058 ( \32373 , \22224 , \22669 );
nor \U$32059 ( \32374 , \32372 , \32373 );
xnor \U$32060 ( \32375 , \32374 , \22681 );
and \U$32061 ( \32376 , \22283 , \22691 );
and \U$32062 ( \32377 , \22251 , \22689 );
nor \U$32063 ( \32378 , \32376 , \32377 );
xnor \U$32064 ( \32379 , \32378 , \22701 );
xor \U$32065 ( \32380 , \32375 , \32379 );
and \U$32066 ( \32381 , \22305 , \22720 );
and \U$32067 ( \32382 , \22272 , \22707 );
nor \U$32068 ( \32383 , \32381 , \32382 );
xnor \U$32069 ( \32384 , \32383 , \22067 );
xor \U$32070 ( \32385 , \32380 , \32384 );
and \U$32071 ( \32386 , \22192 , \22598 );
and \U$32072 ( \32387 , \22156 , \22596 );
nor \U$32073 ( \32388 , \32386 , \32387 );
xnor \U$32074 ( \32389 , \32388 , \22608 );
and \U$32075 ( \32390 , \22213 , \22619 );
and \U$32076 ( \32391 , \22181 , \22617 );
nor \U$32077 ( \32392 , \32390 , \32391 );
xnor \U$32078 ( \32393 , \32392 , \22629 );
xor \U$32079 ( \32394 , \32389 , \32393 );
and \U$32080 ( \32395 , \22235 , \22641 );
and \U$32081 ( \32396 , \22202 , \22639 );
nor \U$32082 ( \32397 , \32395 , \32396 );
xnor \U$32083 ( \32398 , \32397 , \22651 );
xor \U$32084 ( \32399 , \32394 , \32398 );
xor \U$32085 ( \32400 , \32385 , \32399 );
and \U$32086 ( \32401 , \22124 , \22530 );
and \U$32087 ( \32402 , \22089 , \22528 );
nor \U$32088 ( \32403 , \32401 , \32402 );
xnor \U$32089 ( \32404 , \32403 , \22540 );
and \U$32090 ( \32405 , \22145 , \22551 );
and \U$32091 ( \32406 , \22113 , \22549 );
nor \U$32092 ( \32407 , \32405 , \32406 );
xnor \U$32093 ( \32408 , \32407 , \22561 );
xor \U$32094 ( \32409 , \32404 , \32408 );
and \U$32095 ( \32410 , \22167 , \22573 );
and \U$32096 ( \32411 , \22134 , \22571 );
nor \U$32097 ( \32412 , \32410 , \32411 );
xnor \U$32098 ( \32413 , \32412 , \22583 );
xor \U$32099 ( \32414 , \32409 , \32413 );
xor \U$32100 ( \32415 , \32400 , \32414 );
xor \U$32101 ( \32416 , \32371 , \32415 );
and \U$32102 ( \32417 , \22361 , \21978 );
and \U$32103 ( \32418 , \22329 , \23173 );
and \U$32104 ( \32419 , \22294 , \22999 );
nor \U$32105 ( \32420 , \32418 , \32419 );
xnor \U$32106 ( \32421 , \32420 , \22016 );
and \U$32107 ( \32422 , \22350 , \22021 );
and \U$32108 ( \32423 , \22318 , \22019 );
nor \U$32109 ( \32424 , \32422 , \32423 );
xnor \U$32110 ( \32425 , \32424 , \21595 );
xor \U$32111 ( \32426 , \32421 , \32425 );
and \U$32112 ( \32427 , \22372 , \21983 );
and \U$32113 ( \32428 , \22339 , \21981 );
nor \U$32114 ( \32429 , \32427 , \32428 );
xnor \U$32115 ( \32430 , \32429 , \21995 );
xor \U$32116 ( \32431 , \32426 , \32430 );
xnor \U$32117 ( \32432 , \32417 , \32431 );
xor \U$32118 ( \32433 , \32416 , \32432 );
xor \U$32119 ( \32434 , \32358 , \32433 );
xor \U$32120 ( \32435 , \32329 , \32434 );
and \U$32121 ( \32436 , \32254 , \32258 );
and \U$32122 ( \32437 , \32258 , \32263 );
and \U$32123 ( \32438 , \32254 , \32263 );
or \U$32124 ( \32439 , \32436 , \32437 , \32438 );
and \U$32125 ( \32440 , \32180 , \32181 );
and \U$32126 ( \32441 , \32181 , \32223 );
and \U$32127 ( \32442 , \32180 , \32223 );
or \U$32128 ( \32443 , \32440 , \32441 , \32442 );
xor \U$32129 ( \32444 , \32439 , \32443 );
and \U$32130 ( \32445 , \32151 , \32159 );
and \U$32131 ( \32446 , \32159 , \32174 );
and \U$32132 ( \32447 , \32151 , \32174 );
or \U$32133 ( \32448 , \32445 , \32446 , \32447 );
xor \U$32134 ( \32449 , \32444 , \32448 );
xor \U$32135 ( \32450 , \32435 , \32449 );
xor \U$32136 ( \32451 , \32315 , \32450 );
xor \U$32137 ( \32452 , \32309 , \32451 );
and \U$32138 ( \32453 , \32084 , \32088 );
and \U$32139 ( \32454 , \32088 , \32266 );
and \U$32140 ( \32455 , \32084 , \32266 );
or \U$32141 ( \32456 , \32453 , \32454 , \32455 );
nor \U$32142 ( \32457 , \32452 , \32456 );
and \U$32143 ( \32458 , \32313 , \32314 );
and \U$32144 ( \32459 , \32314 , \32450 );
and \U$32145 ( \32460 , \32313 , \32450 );
or \U$32146 ( \32461 , \32458 , \32459 , \32460 );
and \U$32147 ( \32462 , \32439 , \32443 );
and \U$32148 ( \32463 , \32443 , \32448 );
and \U$32149 ( \32464 , \32439 , \32448 );
or \U$32150 ( \32465 , \32462 , \32463 , \32464 );
and \U$32151 ( \32466 , \32343 , \32357 );
and \U$32152 ( \32467 , \32357 , \32433 );
and \U$32153 ( \32468 , \32343 , \32433 );
or \U$32154 ( \32469 , \32466 , \32467 , \32468 );
xor \U$32155 ( \32470 , \32465 , \32469 );
and \U$32156 ( \32471 , \22372 , \21978 );
and \U$32157 ( \32472 , \22294 , \23173 );
and \U$32158 ( \32473 , \22305 , \22999 );
nor \U$32159 ( \32474 , \32472 , \32473 );
xnor \U$32160 ( \32475 , \32474 , \22016 );
and \U$32161 ( \32476 , \22318 , \22021 );
and \U$32162 ( \32477 , \22329 , \22019 );
nor \U$32163 ( \32478 , \32476 , \32477 );
xnor \U$32164 ( \32479 , \32478 , \21595 );
xor \U$32165 ( \32480 , \32475 , \32479 );
and \U$32166 ( \32481 , \22339 , \21983 );
and \U$32167 ( \32482 , \22350 , \21981 );
nor \U$32168 ( \32483 , \32481 , \32482 );
xnor \U$32169 ( \32484 , \32483 , \21995 );
xor \U$32170 ( \32485 , \32480 , \32484 );
xor \U$32171 ( \32486 , \32471 , \32485 );
and \U$32172 ( \32487 , \22224 , \22671 );
and \U$32173 ( \32488 , \22235 , \22669 );
nor \U$32174 ( \32489 , \32487 , \32488 );
xnor \U$32175 ( \32490 , \32489 , \22681 );
and \U$32176 ( \32491 , \22251 , \22691 );
and \U$32177 ( \32492 , \22262 , \22689 );
nor \U$32178 ( \32493 , \32491 , \32492 );
xnor \U$32179 ( \32494 , \32493 , \22701 );
xor \U$32180 ( \32495 , \32490 , \32494 );
and \U$32181 ( \32496 , \22272 , \22720 );
and \U$32182 ( \32497 , \22283 , \22707 );
nor \U$32183 ( \32498 , \32496 , \32497 );
xnor \U$32184 ( \32499 , \32498 , \22067 );
xor \U$32185 ( \32500 , \32495 , \32499 );
xor \U$32186 ( \32501 , \32486 , \32500 );
and \U$32187 ( \32502 , \32389 , \32393 );
and \U$32188 ( \32503 , \32393 , \32398 );
and \U$32189 ( \32504 , \32389 , \32398 );
or \U$32190 ( \32505 , \32502 , \32503 , \32504 );
and \U$32191 ( \32506 , \32375 , \32379 );
and \U$32192 ( \32507 , \32379 , \32384 );
and \U$32193 ( \32508 , \32375 , \32384 );
or \U$32194 ( \32509 , \32506 , \32507 , \32508 );
xor \U$32195 ( \32510 , \32505 , \32509 );
and \U$32196 ( \32511 , \32421 , \32425 );
and \U$32197 ( \32512 , \32425 , \32430 );
and \U$32198 ( \32513 , \32421 , \32430 );
or \U$32199 ( \32514 , \32511 , \32512 , \32513 );
xor \U$32200 ( \32515 , \32510 , \32514 );
xor \U$32201 ( \32516 , \32501 , \32515 );
and \U$32202 ( \32517 , \32361 , \32365 );
and \U$32203 ( \32518 , \32365 , \32370 );
and \U$32204 ( \32519 , \32361 , \32370 );
or \U$32205 ( \32520 , \32517 , \32518 , \32519 );
and \U$32206 ( \32521 , \32296 , \32300 );
and \U$32207 ( \32522 , \32300 , \32305 );
and \U$32208 ( \32523 , \32296 , \32305 );
or \U$32209 ( \32524 , \32521 , \32522 , \32523 );
xor \U$32210 ( \32525 , \32520 , \32524 );
and \U$32211 ( \32526 , \32404 , \32408 );
and \U$32212 ( \32527 , \32408 , \32413 );
and \U$32213 ( \32528 , \32404 , \32413 );
or \U$32214 ( \32529 , \32526 , \32527 , \32528 );
xor \U$32215 ( \32530 , \32525 , \32529 );
xor \U$32216 ( \32531 , \32516 , \32530 );
and \U$32217 ( \32532 , \32385 , \32399 );
and \U$32218 ( \32533 , \32399 , \32414 );
and \U$32219 ( \32534 , \32385 , \32414 );
or \U$32220 ( \32535 , \32532 , \32533 , \32534 );
not \U$32221 ( \32536 , \22402 );
and \U$32222 ( \32537 , \21977 , \22413 );
and \U$32223 ( \32538 , \21990 , \22411 );
nor \U$32224 ( \32539 , \32537 , \32538 );
xnor \U$32225 ( \32540 , \32539 , \22423 );
xor \U$32226 ( \32541 , \32536 , \32540 );
and \U$32227 ( \32542 , \22030 , \22435 );
and \U$32228 ( \32543 , \22001 , \22433 );
nor \U$32229 ( \32544 , \32542 , \32543 );
xnor \U$32230 ( \32545 , \32544 , \22445 );
xor \U$32231 ( \32546 , \32541 , \32545 );
xor \U$32232 ( \32547 , \32535 , \32546 );
and \U$32233 ( \32548 , \22156 , \22598 );
and \U$32234 ( \32549 , \22167 , \22596 );
nor \U$32235 ( \32550 , \32548 , \32549 );
xnor \U$32236 ( \32551 , \32550 , \22608 );
and \U$32237 ( \32552 , \22181 , \22619 );
and \U$32238 ( \32553 , \22192 , \22617 );
nor \U$32239 ( \32554 , \32552 , \32553 );
xnor \U$32240 ( \32555 , \32554 , \22629 );
xor \U$32241 ( \32556 , \32551 , \32555 );
and \U$32242 ( \32557 , \22202 , \22641 );
and \U$32243 ( \32558 , \22213 , \22639 );
nor \U$32244 ( \32559 , \32557 , \32558 );
xnor \U$32245 ( \32560 , \32559 , \22651 );
xor \U$32246 ( \32561 , \32556 , \32560 );
and \U$32247 ( \32562 , \22089 , \22530 );
and \U$32248 ( \32563 , \22100 , \22528 );
nor \U$32249 ( \32564 , \32562 , \32563 );
xnor \U$32250 ( \32565 , \32564 , \22540 );
and \U$32251 ( \32566 , \22113 , \22551 );
and \U$32252 ( \32567 , \22124 , \22549 );
nor \U$32253 ( \32568 , \32566 , \32567 );
xnor \U$32254 ( \32569 , \32568 , \22561 );
xor \U$32255 ( \32570 , \32565 , \32569 );
and \U$32256 ( \32571 , \22134 , \22573 );
and \U$32257 ( \32572 , \22145 , \22571 );
nor \U$32258 ( \32573 , \32571 , \32572 );
xnor \U$32259 ( \32574 , \32573 , \22583 );
xor \U$32260 ( \32575 , \32570 , \32574 );
xor \U$32261 ( \32576 , \32561 , \32575 );
and \U$32262 ( \32577 , \23230 , \22463 );
and \U$32263 ( \32578 , \23329 , \22461 );
nor \U$32264 ( \32579 , \32577 , \32578 );
xnor \U$32265 ( \32580 , \32579 , \22473 );
and \U$32266 ( \32581 , \22858 , \22484 );
and \U$32267 ( \32582 , \22894 , \22482 );
nor \U$32268 ( \32583 , \32581 , \32582 );
xnor \U$32269 ( \32584 , \32583 , \22494 );
xor \U$32270 ( \32585 , \32580 , \32584 );
and \U$32271 ( \32586 , \22071 , \22506 );
and \U$32272 ( \32587 , \22081 , \22504 );
nor \U$32273 ( \32588 , \32586 , \32587 );
xnor \U$32274 ( \32589 , \32588 , \22516 );
xor \U$32275 ( \32590 , \32585 , \32589 );
xor \U$32276 ( \32591 , \32576 , \32590 );
xor \U$32277 ( \32592 , \32547 , \32591 );
xor \U$32278 ( \32593 , \32531 , \32592 );
and \U$32279 ( \32594 , \32347 , \32351 );
and \U$32280 ( \32595 , \32351 , \32356 );
and \U$32281 ( \32596 , \32347 , \32356 );
or \U$32282 ( \32597 , \32594 , \32595 , \32596 );
and \U$32283 ( \32598 , \32333 , \32337 );
and \U$32284 ( \32599 , \32337 , \32342 );
and \U$32285 ( \32600 , \32333 , \32342 );
or \U$32286 ( \32601 , \32598 , \32599 , \32600 );
xor \U$32287 ( \32602 , \32597 , \32601 );
or \U$32288 ( \32603 , \32417 , \32431 );
xor \U$32289 ( \32604 , \32602 , \32603 );
xor \U$32290 ( \32605 , \32593 , \32604 );
xor \U$32291 ( \32606 , \32470 , \32605 );
xor \U$32292 ( \32607 , \32461 , \32606 );
and \U$32293 ( \32608 , \32278 , \32282 );
and \U$32294 ( \32609 , \32282 , \32307 );
and \U$32295 ( \32610 , \32278 , \32307 );
or \U$32296 ( \32611 , \32608 , \32609 , \32610 );
and \U$32297 ( \32612 , \32329 , \32434 );
and \U$32298 ( \32613 , \32434 , \32449 );
and \U$32299 ( \32614 , \32329 , \32449 );
or \U$32300 ( \32615 , \32612 , \32613 , \32614 );
xor \U$32301 ( \32616 , \32611 , \32615 );
and \U$32302 ( \32617 , \32319 , \32323 );
and \U$32303 ( \32618 , \32323 , \32328 );
and \U$32304 ( \32619 , \32319 , \32328 );
or \U$32305 ( \32620 , \32617 , \32618 , \32619 );
and \U$32306 ( \32621 , \32287 , \32291 );
and \U$32307 ( \32622 , \32291 , \32306 );
and \U$32308 ( \32623 , \32287 , \32306 );
or \U$32309 ( \32624 , \32621 , \32622 , \32623 );
xor \U$32310 ( \32625 , \32620 , \32624 );
and \U$32311 ( \32626 , \32371 , \32415 );
and \U$32312 ( \32627 , \32415 , \32432 );
and \U$32313 ( \32628 , \32371 , \32432 );
or \U$32314 ( \32629 , \32626 , \32627 , \32628 );
xor \U$32315 ( \32630 , \32625 , \32629 );
xor \U$32316 ( \32631 , \32616 , \32630 );
xor \U$32317 ( \32632 , \32607 , \32631 );
and \U$32318 ( \32633 , \32274 , \32308 );
and \U$32319 ( \32634 , \32308 , \32451 );
and \U$32320 ( \32635 , \32274 , \32451 );
or \U$32321 ( \32636 , \32633 , \32634 , \32635 );
nor \U$32322 ( \32637 , \32632 , \32636 );
nor \U$32323 ( \32638 , \32457 , \32637 );
nand \U$32324 ( \32639 , \32270 , \32638 );
nor \U$32325 ( \32640 , \31883 , \32639 );
nand \U$32326 ( \32641 , \31045 , \32640 );
nor \U$32327 ( \32642 , \29124 , \32641 );
and \U$32328 ( \32643 , \32611 , \32615 );
and \U$32329 ( \32644 , \32615 , \32630 );
and \U$32330 ( \32645 , \32611 , \32630 );
or \U$32331 ( \32646 , \32643 , \32644 , \32645 );
and \U$32332 ( \32647 , \32465 , \32469 );
and \U$32333 ( \32648 , \32469 , \32605 );
and \U$32334 ( \32649 , \32465 , \32605 );
or \U$32335 ( \32650 , \32647 , \32648 , \32649 );
and \U$32336 ( \32651 , \32597 , \32601 );
and \U$32337 ( \32652 , \32601 , \32603 );
and \U$32338 ( \32653 , \32597 , \32603 );
or \U$32339 ( \32654 , \32651 , \32652 , \32653 );
and \U$32340 ( \32655 , \32535 , \32546 );
and \U$32341 ( \32656 , \32546 , \32591 );
and \U$32342 ( \32657 , \32535 , \32591 );
or \U$32343 ( \32658 , \32655 , \32656 , \32657 );
xor \U$32344 ( \32659 , \32654 , \32658 );
and \U$32345 ( \32660 , \32501 , \32515 );
and \U$32346 ( \32661 , \32515 , \32530 );
and \U$32347 ( \32662 , \32501 , \32530 );
or \U$32348 ( \32663 , \32660 , \32661 , \32662 );
xor \U$32349 ( \32664 , \32659 , \32663 );
xor \U$32350 ( \32665 , \32650 , \32664 );
and \U$32351 ( \32666 , \32620 , \32624 );
and \U$32352 ( \32667 , \32624 , \32629 );
and \U$32353 ( \32668 , \32620 , \32629 );
or \U$32354 ( \32669 , \32666 , \32667 , \32668 );
and \U$32355 ( \32670 , \32531 , \32592 );
and \U$32356 ( \32671 , \32592 , \32604 );
and \U$32357 ( \32672 , \32531 , \32604 );
or \U$32358 ( \32673 , \32670 , \32671 , \32672 );
xor \U$32359 ( \32674 , \32669 , \32673 );
and \U$32360 ( \32675 , \22329 , \22021 );
and \U$32361 ( \32676 , \22294 , \22019 );
nor \U$32362 ( \32677 , \32675 , \32676 );
xnor \U$32363 ( \32678 , \32677 , \21595 );
and \U$32364 ( \32679 , \22350 , \21983 );
and \U$32365 ( \32680 , \22318 , \21981 );
nor \U$32366 ( \32681 , \32679 , \32680 );
xnor \U$32367 ( \32682 , \32681 , \21995 );
xor \U$32368 ( \32683 , \32678 , \32682 );
and \U$32369 ( \32684 , \22339 , \21978 );
xor \U$32370 ( \32685 , \32683 , \32684 );
and \U$32371 ( \32686 , \22262 , \22691 );
and \U$32372 ( \32687 , \22224 , \22689 );
nor \U$32373 ( \32688 , \32686 , \32687 );
xnor \U$32374 ( \32689 , \32688 , \22701 );
and \U$32375 ( \32690 , \22283 , \22720 );
and \U$32376 ( \32691 , \22251 , \22707 );
nor \U$32377 ( \32692 , \32690 , \32691 );
xnor \U$32378 ( \32693 , \32692 , \22067 );
xor \U$32379 ( \32694 , \32689 , \32693 );
and \U$32380 ( \32695 , \22305 , \23173 );
and \U$32381 ( \32696 , \22272 , \22999 );
nor \U$32382 ( \32697 , \32695 , \32696 );
xnor \U$32383 ( \32698 , \32697 , \22016 );
xor \U$32384 ( \32699 , \32694 , \32698 );
xnor \U$32385 ( \32700 , \32685 , \32699 );
and \U$32386 ( \32701 , \32551 , \32555 );
and \U$32387 ( \32702 , \32555 , \32560 );
and \U$32388 ( \32703 , \32551 , \32560 );
or \U$32389 ( \32704 , \32701 , \32702 , \32703 );
and \U$32390 ( \32705 , \32490 , \32494 );
and \U$32391 ( \32706 , \32494 , \32499 );
and \U$32392 ( \32707 , \32490 , \32499 );
or \U$32393 ( \32708 , \32705 , \32706 , \32707 );
xor \U$32394 ( \32709 , \32704 , \32708 );
and \U$32395 ( \32710 , \32475 , \32479 );
and \U$32396 ( \32711 , \32479 , \32484 );
and \U$32397 ( \32712 , \32475 , \32484 );
or \U$32398 ( \32713 , \32710 , \32711 , \32712 );
xor \U$32399 ( \32714 , \32709 , \32713 );
xor \U$32400 ( \32715 , \32700 , \32714 );
and \U$32401 ( \32716 , \32536 , \32540 );
and \U$32402 ( \32717 , \32540 , \32545 );
and \U$32403 ( \32718 , \32536 , \32545 );
or \U$32404 ( \32719 , \32716 , \32717 , \32718 );
and \U$32405 ( \32720 , \32580 , \32584 );
and \U$32406 ( \32721 , \32584 , \32589 );
and \U$32407 ( \32722 , \32580 , \32589 );
or \U$32408 ( \32723 , \32720 , \32721 , \32722 );
xor \U$32409 ( \32724 , \32719 , \32723 );
and \U$32410 ( \32725 , \32565 , \32569 );
and \U$32411 ( \32726 , \32569 , \32574 );
and \U$32412 ( \32727 , \32565 , \32574 );
or \U$32413 ( \32728 , \32725 , \32726 , \32727 );
xor \U$32414 ( \32729 , \32724 , \32728 );
xor \U$32415 ( \32730 , \32715 , \32729 );
and \U$32416 ( \32731 , \32561 , \32575 );
and \U$32417 ( \32732 , \32575 , \32590 );
and \U$32418 ( \32733 , \32561 , \32590 );
or \U$32419 ( \32734 , \32731 , \32732 , \32733 );
and \U$32420 ( \32735 , \21990 , \22413 );
not \U$32421 ( \32736 , \32735 );
xnor \U$32422 ( \32737 , \32736 , \22423 );
and \U$32423 ( \32738 , \22001 , \22435 );
and \U$32424 ( \32739 , \21977 , \22433 );
nor \U$32425 ( \32740 , \32738 , \32739 );
xnor \U$32426 ( \32741 , \32740 , \22445 );
xor \U$32427 ( \32742 , \32737 , \32741 );
and \U$32428 ( \32743 , \23329 , \22463 );
and \U$32429 ( \32744 , \22030 , \22461 );
nor \U$32430 ( \32745 , \32743 , \32744 );
xnor \U$32431 ( \32746 , \32745 , \22473 );
xor \U$32432 ( \32747 , \32742 , \32746 );
xor \U$32433 ( \32748 , \32734 , \32747 );
and \U$32434 ( \32749 , \22192 , \22619 );
and \U$32435 ( \32750 , \22156 , \22617 );
nor \U$32436 ( \32751 , \32749 , \32750 );
xnor \U$32437 ( \32752 , \32751 , \22629 );
and \U$32438 ( \32753 , \22213 , \22641 );
and \U$32439 ( \32754 , \22181 , \22639 );
nor \U$32440 ( \32755 , \32753 , \32754 );
xnor \U$32441 ( \32756 , \32755 , \22651 );
xor \U$32442 ( \32757 , \32752 , \32756 );
and \U$32443 ( \32758 , \22235 , \22671 );
and \U$32444 ( \32759 , \22202 , \22669 );
nor \U$32445 ( \32760 , \32758 , \32759 );
xnor \U$32446 ( \32761 , \32760 , \22681 );
xor \U$32447 ( \32762 , \32757 , \32761 );
and \U$32448 ( \32763 , \22124 , \22551 );
and \U$32449 ( \32764 , \22089 , \22549 );
nor \U$32450 ( \32765 , \32763 , \32764 );
xnor \U$32451 ( \32766 , \32765 , \22561 );
and \U$32452 ( \32767 , \22145 , \22573 );
and \U$32453 ( \32768 , \22113 , \22571 );
nor \U$32454 ( \32769 , \32767 , \32768 );
xnor \U$32455 ( \32770 , \32769 , \22583 );
xor \U$32456 ( \32771 , \32766 , \32770 );
and \U$32457 ( \32772 , \22167 , \22598 );
and \U$32458 ( \32773 , \22134 , \22596 );
nor \U$32459 ( \32774 , \32772 , \32773 );
xnor \U$32460 ( \32775 , \32774 , \22608 );
xor \U$32461 ( \32776 , \32771 , \32775 );
xor \U$32462 ( \32777 , \32762 , \32776 );
and \U$32463 ( \32778 , \22894 , \22484 );
and \U$32464 ( \32779 , \23230 , \22482 );
nor \U$32465 ( \32780 , \32778 , \32779 );
xnor \U$32466 ( \32781 , \32780 , \22494 );
and \U$32467 ( \32782 , \22081 , \22506 );
and \U$32468 ( \32783 , \22858 , \22504 );
nor \U$32469 ( \32784 , \32782 , \32783 );
xnor \U$32470 ( \32785 , \32784 , \22516 );
xor \U$32471 ( \32786 , \32781 , \32785 );
and \U$32472 ( \32787 , \22100 , \22530 );
and \U$32473 ( \32788 , \22071 , \22528 );
nor \U$32474 ( \32789 , \32787 , \32788 );
xnor \U$32475 ( \32790 , \32789 , \22540 );
xor \U$32476 ( \32791 , \32786 , \32790 );
xor \U$32477 ( \32792 , \32777 , \32791 );
xor \U$32478 ( \32793 , \32748 , \32792 );
xor \U$32479 ( \32794 , \32730 , \32793 );
and \U$32480 ( \32795 , \32520 , \32524 );
and \U$32481 ( \32796 , \32524 , \32529 );
and \U$32482 ( \32797 , \32520 , \32529 );
or \U$32483 ( \32798 , \32795 , \32796 , \32797 );
and \U$32484 ( \32799 , \32505 , \32509 );
and \U$32485 ( \32800 , \32509 , \32514 );
and \U$32486 ( \32801 , \32505 , \32514 );
or \U$32487 ( \32802 , \32799 , \32800 , \32801 );
xor \U$32488 ( \32803 , \32798 , \32802 );
and \U$32489 ( \32804 , \32471 , \32485 );
and \U$32490 ( \32805 , \32485 , \32500 );
and \U$32491 ( \32806 , \32471 , \32500 );
or \U$32492 ( \32807 , \32804 , \32805 , \32806 );
xor \U$32493 ( \32808 , \32803 , \32807 );
xor \U$32494 ( \32809 , \32794 , \32808 );
xor \U$32495 ( \32810 , \32674 , \32809 );
xor \U$32496 ( \32811 , \32665 , \32810 );
xor \U$32497 ( \32812 , \32646 , \32811 );
and \U$32498 ( \32813 , \32461 , \32606 );
and \U$32499 ( \32814 , \32606 , \32631 );
and \U$32500 ( \32815 , \32461 , \32631 );
or \U$32501 ( \32816 , \32813 , \32814 , \32815 );
nor \U$32502 ( \32817 , \32812 , \32816 );
and \U$32503 ( \32818 , \32650 , \32664 );
and \U$32504 ( \32819 , \32664 , \32810 );
and \U$32505 ( \32820 , \32650 , \32810 );
or \U$32506 ( \32821 , \32818 , \32819 , \32820 );
and \U$32507 ( \32822 , \32669 , \32673 );
and \U$32508 ( \32823 , \32673 , \32809 );
and \U$32509 ( \32824 , \32669 , \32809 );
or \U$32510 ( \32825 , \32822 , \32823 , \32824 );
and \U$32511 ( \32826 , \32798 , \32802 );
and \U$32512 ( \32827 , \32802 , \32807 );
and \U$32513 ( \32828 , \32798 , \32807 );
or \U$32514 ( \32829 , \32826 , \32827 , \32828 );
and \U$32515 ( \32830 , \32734 , \32747 );
and \U$32516 ( \32831 , \32747 , \32792 );
and \U$32517 ( \32832 , \32734 , \32792 );
or \U$32518 ( \32833 , \32830 , \32831 , \32832 );
xor \U$32519 ( \32834 , \32829 , \32833 );
and \U$32520 ( \32835 , \32700 , \32714 );
and \U$32521 ( \32836 , \32714 , \32729 );
and \U$32522 ( \32837 , \32700 , \32729 );
or \U$32523 ( \32838 , \32835 , \32836 , \32837 );
xor \U$32524 ( \32839 , \32834 , \32838 );
xor \U$32525 ( \32840 , \32825 , \32839 );
and \U$32526 ( \32841 , \32654 , \32658 );
and \U$32527 ( \32842 , \32658 , \32663 );
and \U$32528 ( \32843 , \32654 , \32663 );
or \U$32529 ( \32844 , \32841 , \32842 , \32843 );
and \U$32530 ( \32845 , \32730 , \32793 );
and \U$32531 ( \32846 , \32793 , \32808 );
and \U$32532 ( \32847 , \32730 , \32808 );
or \U$32533 ( \32848 , \32845 , \32846 , \32847 );
xor \U$32534 ( \32849 , \32844 , \32848 );
and \U$32535 ( \32850 , \32752 , \32756 );
and \U$32536 ( \32851 , \32756 , \32761 );
and \U$32537 ( \32852 , \32752 , \32761 );
or \U$32538 ( \32853 , \32850 , \32851 , \32852 );
and \U$32539 ( \32854 , \32689 , \32693 );
and \U$32540 ( \32855 , \32693 , \32698 );
and \U$32541 ( \32856 , \32689 , \32698 );
or \U$32542 ( \32857 , \32854 , \32855 , \32856 );
xor \U$32543 ( \32858 , \32853 , \32857 );
and \U$32544 ( \32859 , \32678 , \32682 );
and \U$32545 ( \32860 , \32682 , \32684 );
and \U$32546 ( \32861 , \32678 , \32684 );
or \U$32547 ( \32862 , \32859 , \32860 , \32861 );
xor \U$32548 ( \32863 , \32858 , \32862 );
and \U$32549 ( \32864 , \32737 , \32741 );
and \U$32550 ( \32865 , \32741 , \32746 );
and \U$32551 ( \32866 , \32737 , \32746 );
or \U$32552 ( \32867 , \32864 , \32865 , \32866 );
and \U$32553 ( \32868 , \32781 , \32785 );
and \U$32554 ( \32869 , \32785 , \32790 );
and \U$32555 ( \32870 , \32781 , \32790 );
or \U$32556 ( \32871 , \32868 , \32869 , \32870 );
xor \U$32557 ( \32872 , \32867 , \32871 );
and \U$32558 ( \32873 , \32766 , \32770 );
and \U$32559 ( \32874 , \32770 , \32775 );
and \U$32560 ( \32875 , \32766 , \32775 );
or \U$32561 ( \32876 , \32873 , \32874 , \32875 );
xor \U$32562 ( \32877 , \32872 , \32876 );
xor \U$32563 ( \32878 , \32863 , \32877 );
and \U$32564 ( \32879 , \32762 , \32776 );
and \U$32565 ( \32880 , \32776 , \32791 );
and \U$32566 ( \32881 , \32762 , \32791 );
or \U$32567 ( \32882 , \32879 , \32880 , \32881 );
and \U$32568 ( \32883 , \22089 , \22551 );
and \U$32569 ( \32884 , \22100 , \22549 );
nor \U$32570 ( \32885 , \32883 , \32884 );
xnor \U$32571 ( \32886 , \32885 , \22561 );
and \U$32572 ( \32887 , \22113 , \22573 );
and \U$32573 ( \32888 , \22124 , \22571 );
nor \U$32574 ( \32889 , \32887 , \32888 );
xnor \U$32575 ( \32890 , \32889 , \22583 );
xor \U$32576 ( \32891 , \32886 , \32890 );
and \U$32577 ( \32892 , \22134 , \22598 );
and \U$32578 ( \32893 , \22145 , \22596 );
nor \U$32579 ( \32894 , \32892 , \32893 );
xnor \U$32580 ( \32895 , \32894 , \22608 );
xor \U$32581 ( \32896 , \32891 , \32895 );
and \U$32582 ( \32897 , \23230 , \22484 );
and \U$32583 ( \32898 , \23329 , \22482 );
nor \U$32584 ( \32899 , \32897 , \32898 );
xnor \U$32585 ( \32900 , \32899 , \22494 );
and \U$32586 ( \32901 , \22858 , \22506 );
and \U$32587 ( \32902 , \22894 , \22504 );
nor \U$32588 ( \32903 , \32901 , \32902 );
xnor \U$32589 ( \32904 , \32903 , \22516 );
xor \U$32590 ( \32905 , \32900 , \32904 );
and \U$32591 ( \32906 , \22071 , \22530 );
and \U$32592 ( \32907 , \22081 , \22528 );
nor \U$32593 ( \32908 , \32906 , \32907 );
xnor \U$32594 ( \32909 , \32908 , \22540 );
xor \U$32595 ( \32910 , \32905 , \32909 );
xor \U$32596 ( \32911 , \32896 , \32910 );
not \U$32597 ( \32912 , \22423 );
and \U$32598 ( \32913 , \21977 , \22435 );
and \U$32599 ( \32914 , \21990 , \22433 );
nor \U$32600 ( \32915 , \32913 , \32914 );
xnor \U$32601 ( \32916 , \32915 , \22445 );
xor \U$32602 ( \32917 , \32912 , \32916 );
and \U$32603 ( \32918 , \22030 , \22463 );
and \U$32604 ( \32919 , \22001 , \22461 );
nor \U$32605 ( \32920 , \32918 , \32919 );
xnor \U$32606 ( \32921 , \32920 , \22473 );
xor \U$32607 ( \32922 , \32917 , \32921 );
xor \U$32608 ( \32923 , \32911 , \32922 );
xor \U$32609 ( \32924 , \32882 , \32923 );
and \U$32610 ( \32925 , \22294 , \22021 );
and \U$32611 ( \32926 , \22305 , \22019 );
nor \U$32612 ( \32927 , \32925 , \32926 );
xnor \U$32613 ( \32928 , \32927 , \21595 );
and \U$32614 ( \32929 , \22318 , \21983 );
and \U$32615 ( \32930 , \22329 , \21981 );
nor \U$32616 ( \32931 , \32929 , \32930 );
xnor \U$32617 ( \32932 , \32931 , \21995 );
xor \U$32618 ( \32933 , \32928 , \32932 );
and \U$32619 ( \32934 , \22350 , \21978 );
xor \U$32620 ( \32935 , \32933 , \32934 );
and \U$32621 ( \32936 , \22224 , \22691 );
and \U$32622 ( \32937 , \22235 , \22689 );
nor \U$32623 ( \32938 , \32936 , \32937 );
xnor \U$32624 ( \32939 , \32938 , \22701 );
and \U$32625 ( \32940 , \22251 , \22720 );
and \U$32626 ( \32941 , \22262 , \22707 );
nor \U$32627 ( \32942 , \32940 , \32941 );
xnor \U$32628 ( \32943 , \32942 , \22067 );
xor \U$32629 ( \32944 , \32939 , \32943 );
and \U$32630 ( \32945 , \22272 , \23173 );
and \U$32631 ( \32946 , \22283 , \22999 );
nor \U$32632 ( \32947 , \32945 , \32946 );
xnor \U$32633 ( \32948 , \32947 , \22016 );
xor \U$32634 ( \32949 , \32944 , \32948 );
xor \U$32635 ( \32950 , \32935 , \32949 );
and \U$32636 ( \32951 , \22156 , \22619 );
and \U$32637 ( \32952 , \22167 , \22617 );
nor \U$32638 ( \32953 , \32951 , \32952 );
xnor \U$32639 ( \32954 , \32953 , \22629 );
and \U$32640 ( \32955 , \22181 , \22641 );
and \U$32641 ( \32956 , \22192 , \22639 );
nor \U$32642 ( \32957 , \32955 , \32956 );
xnor \U$32643 ( \32958 , \32957 , \22651 );
xor \U$32644 ( \32959 , \32954 , \32958 );
and \U$32645 ( \32960 , \22202 , \22671 );
and \U$32646 ( \32961 , \22213 , \22669 );
nor \U$32647 ( \32962 , \32960 , \32961 );
xnor \U$32648 ( \32963 , \32962 , \22681 );
xor \U$32649 ( \32964 , \32959 , \32963 );
xor \U$32650 ( \32965 , \32950 , \32964 );
xor \U$32651 ( \32966 , \32924 , \32965 );
xor \U$32652 ( \32967 , \32878 , \32966 );
and \U$32653 ( \32968 , \32719 , \32723 );
and \U$32654 ( \32969 , \32723 , \32728 );
and \U$32655 ( \32970 , \32719 , \32728 );
or \U$32656 ( \32971 , \32968 , \32969 , \32970 );
and \U$32657 ( \32972 , \32704 , \32708 );
and \U$32658 ( \32973 , \32708 , \32713 );
and \U$32659 ( \32974 , \32704 , \32713 );
or \U$32660 ( \32975 , \32972 , \32973 , \32974 );
xor \U$32661 ( \32976 , \32971 , \32975 );
or \U$32662 ( \32977 , \32685 , \32699 );
xor \U$32663 ( \32978 , \32976 , \32977 );
xor \U$32664 ( \32979 , \32967 , \32978 );
xor \U$32665 ( \32980 , \32849 , \32979 );
xor \U$32666 ( \32981 , \32840 , \32980 );
xor \U$32667 ( \32982 , \32821 , \32981 );
and \U$32668 ( \32983 , \32646 , \32811 );
nor \U$32669 ( \32984 , \32982 , \32983 );
nor \U$32670 ( \32985 , \32817 , \32984 );
and \U$32671 ( \32986 , \32825 , \32839 );
and \U$32672 ( \32987 , \32839 , \32980 );
and \U$32673 ( \32988 , \32825 , \32980 );
or \U$32674 ( \32989 , \32986 , \32987 , \32988 );
and \U$32675 ( \32990 , \32844 , \32848 );
and \U$32676 ( \32991 , \32848 , \32979 );
and \U$32677 ( \32992 , \32844 , \32979 );
or \U$32678 ( \32993 , \32990 , \32991 , \32992 );
and \U$32679 ( \32994 , \32971 , \32975 );
and \U$32680 ( \32995 , \32975 , \32977 );
and \U$32681 ( \32996 , \32971 , \32977 );
or \U$32682 ( \32997 , \32994 , \32995 , \32996 );
and \U$32683 ( \32998 , \32882 , \32923 );
and \U$32684 ( \32999 , \32923 , \32965 );
and \U$32685 ( \33000 , \32882 , \32965 );
or \U$32686 ( \33001 , \32998 , \32999 , \33000 );
xor \U$32687 ( \33002 , \32997 , \33001 );
and \U$32688 ( \33003 , \32863 , \32877 );
xor \U$32689 ( \33004 , \33002 , \33003 );
xor \U$32690 ( \33005 , \32993 , \33004 );
and \U$32691 ( \33006 , \32829 , \32833 );
and \U$32692 ( \33007 , \32833 , \32838 );
and \U$32693 ( \33008 , \32829 , \32838 );
or \U$32694 ( \33009 , \33006 , \33007 , \33008 );
and \U$32695 ( \33010 , \32878 , \32966 );
and \U$32696 ( \33011 , \32966 , \32978 );
and \U$32697 ( \33012 , \32878 , \32978 );
or \U$32698 ( \33013 , \33010 , \33011 , \33012 );
xor \U$32699 ( \33014 , \33009 , \33013 );
and \U$32700 ( \33015 , \32954 , \32958 );
and \U$32701 ( \33016 , \32958 , \32963 );
and \U$32702 ( \33017 , \32954 , \32963 );
or \U$32703 ( \33018 , \33015 , \33016 , \33017 );
and \U$32704 ( \33019 , \32939 , \32943 );
and \U$32705 ( \33020 , \32943 , \32948 );
and \U$32706 ( \33021 , \32939 , \32948 );
or \U$32707 ( \33022 , \33019 , \33020 , \33021 );
xor \U$32708 ( \33023 , \33018 , \33022 );
and \U$32709 ( \33024 , \32928 , \32932 );
and \U$32710 ( \33025 , \32932 , \32934 );
and \U$32711 ( \33026 , \32928 , \32934 );
or \U$32712 ( \33027 , \33024 , \33025 , \33026 );
xor \U$32713 ( \33028 , \33023 , \33027 );
and \U$32714 ( \33029 , \32912 , \32916 );
and \U$32715 ( \33030 , \32916 , \32921 );
and \U$32716 ( \33031 , \32912 , \32921 );
or \U$32717 ( \33032 , \33029 , \33030 , \33031 );
and \U$32718 ( \33033 , \32900 , \32904 );
and \U$32719 ( \33034 , \32904 , \32909 );
and \U$32720 ( \33035 , \32900 , \32909 );
or \U$32721 ( \33036 , \33033 , \33034 , \33035 );
xor \U$32722 ( \33037 , \33032 , \33036 );
and \U$32723 ( \33038 , \32886 , \32890 );
and \U$32724 ( \33039 , \32890 , \32895 );
and \U$32725 ( \33040 , \32886 , \32895 );
or \U$32726 ( \33041 , \33038 , \33039 , \33040 );
xor \U$32727 ( \33042 , \33037 , \33041 );
xor \U$32728 ( \33043 , \33028 , \33042 );
and \U$32729 ( \33044 , \32896 , \32910 );
and \U$32730 ( \33045 , \32910 , \32922 );
and \U$32731 ( \33046 , \32896 , \32922 );
or \U$32732 ( \33047 , \33044 , \33045 , \33046 );
and \U$32733 ( \33048 , \22124 , \22573 );
and \U$32734 ( \33049 , \22089 , \22571 );
nor \U$32735 ( \33050 , \33048 , \33049 );
xnor \U$32736 ( \33051 , \33050 , \22583 );
and \U$32737 ( \33052 , \22145 , \22598 );
and \U$32738 ( \33053 , \22113 , \22596 );
nor \U$32739 ( \33054 , \33052 , \33053 );
xnor \U$32740 ( \33055 , \33054 , \22608 );
xor \U$32741 ( \33056 , \33051 , \33055 );
and \U$32742 ( \33057 , \22167 , \22619 );
and \U$32743 ( \33058 , \22134 , \22617 );
nor \U$32744 ( \33059 , \33057 , \33058 );
xnor \U$32745 ( \33060 , \33059 , \22629 );
xor \U$32746 ( \33061 , \33056 , \33060 );
and \U$32747 ( \33062 , \22894 , \22506 );
and \U$32748 ( \33063 , \23230 , \22504 );
nor \U$32749 ( \33064 , \33062 , \33063 );
xnor \U$32750 ( \33065 , \33064 , \22516 );
and \U$32751 ( \33066 , \22081 , \22530 );
and \U$32752 ( \33067 , \22858 , \22528 );
nor \U$32753 ( \33068 , \33066 , \33067 );
xnor \U$32754 ( \33069 , \33068 , \22540 );
xor \U$32755 ( \33070 , \33065 , \33069 );
and \U$32756 ( \33071 , \22100 , \22551 );
and \U$32757 ( \33072 , \22071 , \22549 );
nor \U$32758 ( \33073 , \33071 , \33072 );
xnor \U$32759 ( \33074 , \33073 , \22561 );
xor \U$32760 ( \33075 , \33070 , \33074 );
xor \U$32761 ( \33076 , \33061 , \33075 );
and \U$32762 ( \33077 , \21990 , \22435 );
not \U$32763 ( \33078 , \33077 );
xnor \U$32764 ( \33079 , \33078 , \22445 );
and \U$32765 ( \33080 , \22001 , \22463 );
and \U$32766 ( \33081 , \21977 , \22461 );
nor \U$32767 ( \33082 , \33080 , \33081 );
xnor \U$32768 ( \33083 , \33082 , \22473 );
xor \U$32769 ( \33084 , \33079 , \33083 );
and \U$32770 ( \33085 , \23329 , \22484 );
and \U$32771 ( \33086 , \22030 , \22482 );
nor \U$32772 ( \33087 , \33085 , \33086 );
xnor \U$32773 ( \33088 , \33087 , \22494 );
xor \U$32774 ( \33089 , \33084 , \33088 );
xor \U$32775 ( \33090 , \33076 , \33089 );
xor \U$32776 ( \33091 , \33047 , \33090 );
and \U$32777 ( \33092 , \22329 , \21983 );
and \U$32778 ( \33093 , \22294 , \21981 );
nor \U$32779 ( \33094 , \33092 , \33093 );
xnor \U$32780 ( \33095 , \33094 , \21995 );
and \U$32781 ( \33096 , \22318 , \21978 );
xnor \U$32782 ( \33097 , \33095 , \33096 );
and \U$32783 ( \33098 , \22262 , \22720 );
and \U$32784 ( \33099 , \22224 , \22707 );
nor \U$32785 ( \33100 , \33098 , \33099 );
xnor \U$32786 ( \33101 , \33100 , \22067 );
and \U$32787 ( \33102 , \22283 , \23173 );
and \U$32788 ( \33103 , \22251 , \22999 );
nor \U$32789 ( \33104 , \33102 , \33103 );
xnor \U$32790 ( \33105 , \33104 , \22016 );
xor \U$32791 ( \33106 , \33101 , \33105 );
and \U$32792 ( \33107 , \22305 , \22021 );
and \U$32793 ( \33108 , \22272 , \22019 );
nor \U$32794 ( \33109 , \33107 , \33108 );
xnor \U$32795 ( \33110 , \33109 , \21595 );
xor \U$32796 ( \33111 , \33106 , \33110 );
xor \U$32797 ( \33112 , \33097 , \33111 );
and \U$32798 ( \33113 , \22192 , \22641 );
and \U$32799 ( \33114 , \22156 , \22639 );
nor \U$32800 ( \33115 , \33113 , \33114 );
xnor \U$32801 ( \33116 , \33115 , \22651 );
and \U$32802 ( \33117 , \22213 , \22671 );
and \U$32803 ( \33118 , \22181 , \22669 );
nor \U$32804 ( \33119 , \33117 , \33118 );
xnor \U$32805 ( \33120 , \33119 , \22681 );
xor \U$32806 ( \33121 , \33116 , \33120 );
and \U$32807 ( \33122 , \22235 , \22691 );
and \U$32808 ( \33123 , \22202 , \22689 );
nor \U$32809 ( \33124 , \33122 , \33123 );
xnor \U$32810 ( \33125 , \33124 , \22701 );
xor \U$32811 ( \33126 , \33121 , \33125 );
xor \U$32812 ( \33127 , \33112 , \33126 );
xor \U$32813 ( \33128 , \33091 , \33127 );
xor \U$32814 ( \33129 , \33043 , \33128 );
and \U$32815 ( \33130 , \32867 , \32871 );
and \U$32816 ( \33131 , \32871 , \32876 );
and \U$32817 ( \33132 , \32867 , \32876 );
or \U$32818 ( \33133 , \33130 , \33131 , \33132 );
and \U$32819 ( \33134 , \32853 , \32857 );
and \U$32820 ( \33135 , \32857 , \32862 );
and \U$32821 ( \33136 , \32853 , \32862 );
or \U$32822 ( \33137 , \33134 , \33135 , \33136 );
xor \U$32823 ( \33138 , \33133 , \33137 );
and \U$32824 ( \33139 , \32935 , \32949 );
and \U$32825 ( \33140 , \32949 , \32964 );
and \U$32826 ( \33141 , \32935 , \32964 );
or \U$32827 ( \33142 , \33139 , \33140 , \33141 );
xor \U$32828 ( \33143 , \33138 , \33142 );
xor \U$32829 ( \33144 , \33129 , \33143 );
xor \U$32830 ( \33145 , \33014 , \33144 );
xor \U$32831 ( \33146 , \33005 , \33145 );
xor \U$32832 ( \33147 , \32989 , \33146 );
and \U$32833 ( \33148 , \32821 , \32981 );
nor \U$32834 ( \33149 , \33147 , \33148 );
and \U$32835 ( \33150 , \32993 , \33004 );
and \U$32836 ( \33151 , \33004 , \33145 );
and \U$32837 ( \33152 , \32993 , \33145 );
or \U$32838 ( \33153 , \33150 , \33151 , \33152 );
and \U$32839 ( \33154 , \33009 , \33013 );
and \U$32840 ( \33155 , \33013 , \33144 );
and \U$32841 ( \33156 , \33009 , \33144 );
or \U$32842 ( \33157 , \33154 , \33155 , \33156 );
and \U$32843 ( \33158 , \33133 , \33137 );
and \U$32844 ( \33159 , \33137 , \33142 );
and \U$32845 ( \33160 , \33133 , \33142 );
or \U$32846 ( \33161 , \33158 , \33159 , \33160 );
and \U$32847 ( \33162 , \33047 , \33090 );
and \U$32848 ( \33163 , \33090 , \33127 );
and \U$32849 ( \33164 , \33047 , \33127 );
or \U$32850 ( \33165 , \33162 , \33163 , \33164 );
xor \U$32851 ( \33166 , \33161 , \33165 );
and \U$32852 ( \33167 , \33028 , \33042 );
xor \U$32853 ( \33168 , \33166 , \33167 );
xor \U$32854 ( \33169 , \33157 , \33168 );
and \U$32855 ( \33170 , \32997 , \33001 );
and \U$32856 ( \33171 , \33001 , \33003 );
and \U$32857 ( \33172 , \32997 , \33003 );
or \U$32858 ( \33173 , \33170 , \33171 , \33172 );
and \U$32859 ( \33174 , \33043 , \33128 );
and \U$32860 ( \33175 , \33128 , \33143 );
and \U$32861 ( \33176 , \33043 , \33143 );
or \U$32862 ( \33177 , \33174 , \33175 , \33176 );
xor \U$32863 ( \33178 , \33173 , \33177 );
and \U$32864 ( \33179 , \33116 , \33120 );
and \U$32865 ( \33180 , \33120 , \33125 );
and \U$32866 ( \33181 , \33116 , \33125 );
or \U$32867 ( \33182 , \33179 , \33180 , \33181 );
and \U$32868 ( \33183 , \33101 , \33105 );
and \U$32869 ( \33184 , \33105 , \33110 );
and \U$32870 ( \33185 , \33101 , \33110 );
or \U$32871 ( \33186 , \33183 , \33184 , \33185 );
xor \U$32872 ( \33187 , \33182 , \33186 );
or \U$32873 ( \33188 , \33095 , \33096 );
xor \U$32874 ( \33189 , \33187 , \33188 );
and \U$32875 ( \33190 , \33079 , \33083 );
and \U$32876 ( \33191 , \33083 , \33088 );
and \U$32877 ( \33192 , \33079 , \33088 );
or \U$32878 ( \33193 , \33190 , \33191 , \33192 );
and \U$32879 ( \33194 , \33065 , \33069 );
and \U$32880 ( \33195 , \33069 , \33074 );
and \U$32881 ( \33196 , \33065 , \33074 );
or \U$32882 ( \33197 , \33194 , \33195 , \33196 );
xor \U$32883 ( \33198 , \33193 , \33197 );
and \U$32884 ( \33199 , \33051 , \33055 );
and \U$32885 ( \33200 , \33055 , \33060 );
and \U$32886 ( \33201 , \33051 , \33060 );
or \U$32887 ( \33202 , \33199 , \33200 , \33201 );
xor \U$32888 ( \33203 , \33198 , \33202 );
xor \U$32889 ( \33204 , \33189 , \33203 );
and \U$32890 ( \33205 , \33061 , \33075 );
and \U$32891 ( \33206 , \33075 , \33089 );
and \U$32892 ( \33207 , \33061 , \33089 );
or \U$32893 ( \33208 , \33205 , \33206 , \33207 );
and \U$32894 ( \33209 , \22089 , \22573 );
and \U$32895 ( \33210 , \22100 , \22571 );
nor \U$32896 ( \33211 , \33209 , \33210 );
xnor \U$32897 ( \33212 , \33211 , \22583 );
and \U$32898 ( \33213 , \22113 , \22598 );
and \U$32899 ( \33214 , \22124 , \22596 );
nor \U$32900 ( \33215 , \33213 , \33214 );
xnor \U$32901 ( \33216 , \33215 , \22608 );
xor \U$32902 ( \33217 , \33212 , \33216 );
and \U$32903 ( \33218 , \22134 , \22619 );
and \U$32904 ( \33219 , \22145 , \22617 );
nor \U$32905 ( \33220 , \33218 , \33219 );
xnor \U$32906 ( \33221 , \33220 , \22629 );
xor \U$32907 ( \33222 , \33217 , \33221 );
and \U$32908 ( \33223 , \23230 , \22506 );
and \U$32909 ( \33224 , \23329 , \22504 );
nor \U$32910 ( \33225 , \33223 , \33224 );
xnor \U$32911 ( \33226 , \33225 , \22516 );
and \U$32912 ( \33227 , \22858 , \22530 );
and \U$32913 ( \33228 , \22894 , \22528 );
nor \U$32914 ( \33229 , \33227 , \33228 );
xnor \U$32915 ( \33230 , \33229 , \22540 );
xor \U$32916 ( \33231 , \33226 , \33230 );
and \U$32917 ( \33232 , \22071 , \22551 );
and \U$32918 ( \33233 , \22081 , \22549 );
nor \U$32919 ( \33234 , \33232 , \33233 );
xnor \U$32920 ( \33235 , \33234 , \22561 );
xor \U$32921 ( \33236 , \33231 , \33235 );
xor \U$32922 ( \33237 , \33222 , \33236 );
not \U$32923 ( \33238 , \22445 );
and \U$32924 ( \33239 , \21977 , \22463 );
and \U$32925 ( \33240 , \21990 , \22461 );
nor \U$32926 ( \33241 , \33239 , \33240 );
xnor \U$32927 ( \33242 , \33241 , \22473 );
xor \U$32928 ( \33243 , \33238 , \33242 );
and \U$32929 ( \33244 , \22030 , \22484 );
and \U$32930 ( \33245 , \22001 , \22482 );
nor \U$32931 ( \33246 , \33244 , \33245 );
xnor \U$32932 ( \33247 , \33246 , \22494 );
xor \U$32933 ( \33248 , \33243 , \33247 );
xor \U$32934 ( \33249 , \33237 , \33248 );
xor \U$32935 ( \33250 , \33208 , \33249 );
and \U$32936 ( \33251 , \22294 , \21983 );
and \U$32937 ( \33252 , \22305 , \21981 );
nor \U$32938 ( \33253 , \33251 , \33252 );
xnor \U$32939 ( \33254 , \33253 , \21995 );
and \U$32940 ( \33255 , \22329 , \21978 );
xor \U$32941 ( \33256 , \33254 , \33255 );
and \U$32942 ( \33257 , \22224 , \22720 );
and \U$32943 ( \33258 , \22235 , \22707 );
nor \U$32944 ( \33259 , \33257 , \33258 );
xnor \U$32945 ( \33260 , \33259 , \22067 );
and \U$32946 ( \33261 , \22251 , \23173 );
and \U$32947 ( \33262 , \22262 , \22999 );
nor \U$32948 ( \33263 , \33261 , \33262 );
xnor \U$32949 ( \33264 , \33263 , \22016 );
xor \U$32950 ( \33265 , \33260 , \33264 );
and \U$32951 ( \33266 , \22272 , \22021 );
and \U$32952 ( \33267 , \22283 , \22019 );
nor \U$32953 ( \33268 , \33266 , \33267 );
xnor \U$32954 ( \33269 , \33268 , \21595 );
xor \U$32955 ( \33270 , \33265 , \33269 );
xor \U$32956 ( \33271 , \33256 , \33270 );
and \U$32957 ( \33272 , \22156 , \22641 );
and \U$32958 ( \33273 , \22167 , \22639 );
nor \U$32959 ( \33274 , \33272 , \33273 );
xnor \U$32960 ( \33275 , \33274 , \22651 );
and \U$32961 ( \33276 , \22181 , \22671 );
and \U$32962 ( \33277 , \22192 , \22669 );
nor \U$32963 ( \33278 , \33276 , \33277 );
xnor \U$32964 ( \33279 , \33278 , \22681 );
xor \U$32965 ( \33280 , \33275 , \33279 );
and \U$32966 ( \33281 , \22202 , \22691 );
and \U$32967 ( \33282 , \22213 , \22689 );
nor \U$32968 ( \33283 , \33281 , \33282 );
xnor \U$32969 ( \33284 , \33283 , \22701 );
xor \U$32970 ( \33285 , \33280 , \33284 );
xor \U$32971 ( \33286 , \33271 , \33285 );
xor \U$32972 ( \33287 , \33250 , \33286 );
xor \U$32973 ( \33288 , \33204 , \33287 );
and \U$32974 ( \33289 , \33032 , \33036 );
and \U$32975 ( \33290 , \33036 , \33041 );
and \U$32976 ( \33291 , \33032 , \33041 );
or \U$32977 ( \33292 , \33289 , \33290 , \33291 );
and \U$32978 ( \33293 , \33018 , \33022 );
and \U$32979 ( \33294 , \33022 , \33027 );
and \U$32980 ( \33295 , \33018 , \33027 );
or \U$32981 ( \33296 , \33293 , \33294 , \33295 );
xor \U$32982 ( \33297 , \33292 , \33296 );
and \U$32983 ( \33298 , \33097 , \33111 );
and \U$32984 ( \33299 , \33111 , \33126 );
and \U$32985 ( \33300 , \33097 , \33126 );
or \U$32986 ( \33301 , \33298 , \33299 , \33300 );
xor \U$32987 ( \33302 , \33297 , \33301 );
xor \U$32988 ( \33303 , \33288 , \33302 );
xor \U$32989 ( \33304 , \33178 , \33303 );
xor \U$32990 ( \33305 , \33169 , \33304 );
xor \U$32991 ( \33306 , \33153 , \33305 );
and \U$32992 ( \33307 , \32989 , \33146 );
nor \U$32993 ( \33308 , \33306 , \33307 );
nor \U$32994 ( \33309 , \33149 , \33308 );
nand \U$32995 ( \33310 , \32985 , \33309 );
and \U$32996 ( \33311 , \33157 , \33168 );
and \U$32997 ( \33312 , \33168 , \33304 );
and \U$32998 ( \33313 , \33157 , \33304 );
or \U$32999 ( \33314 , \33311 , \33312 , \33313 );
and \U$33000 ( \33315 , \33173 , \33177 );
and \U$33001 ( \33316 , \33177 , \33303 );
and \U$33002 ( \33317 , \33173 , \33303 );
or \U$33003 ( \33318 , \33315 , \33316 , \33317 );
and \U$33004 ( \33319 , \33292 , \33296 );
and \U$33005 ( \33320 , \33296 , \33301 );
and \U$33006 ( \33321 , \33292 , \33301 );
or \U$33007 ( \33322 , \33319 , \33320 , \33321 );
and \U$33008 ( \33323 , \33208 , \33249 );
and \U$33009 ( \33324 , \33249 , \33286 );
and \U$33010 ( \33325 , \33208 , \33286 );
or \U$33011 ( \33326 , \33323 , \33324 , \33325 );
xor \U$33012 ( \33327 , \33322 , \33326 );
and \U$33013 ( \33328 , \33189 , \33203 );
xor \U$33014 ( \33329 , \33327 , \33328 );
xor \U$33015 ( \33330 , \33318 , \33329 );
and \U$33016 ( \33331 , \33161 , \33165 );
and \U$33017 ( \33332 , \33165 , \33167 );
and \U$33018 ( \33333 , \33161 , \33167 );
or \U$33019 ( \33334 , \33331 , \33332 , \33333 );
and \U$33020 ( \33335 , \33204 , \33287 );
and \U$33021 ( \33336 , \33287 , \33302 );
and \U$33022 ( \33337 , \33204 , \33302 );
or \U$33023 ( \33338 , \33335 , \33336 , \33337 );
xor \U$33024 ( \33339 , \33334 , \33338 );
and \U$33025 ( \33340 , \33275 , \33279 );
and \U$33026 ( \33341 , \33279 , \33284 );
and \U$33027 ( \33342 , \33275 , \33284 );
or \U$33028 ( \33343 , \33340 , \33341 , \33342 );
and \U$33029 ( \33344 , \33260 , \33264 );
and \U$33030 ( \33345 , \33264 , \33269 );
and \U$33031 ( \33346 , \33260 , \33269 );
or \U$33032 ( \33347 , \33344 , \33345 , \33346 );
xor \U$33033 ( \33348 , \33343 , \33347 );
and \U$33034 ( \33349 , \33254 , \33255 );
xor \U$33035 ( \33350 , \33348 , \33349 );
and \U$33036 ( \33351 , \33238 , \33242 );
and \U$33037 ( \33352 , \33242 , \33247 );
and \U$33038 ( \33353 , \33238 , \33247 );
or \U$33039 ( \33354 , \33351 , \33352 , \33353 );
and \U$33040 ( \33355 , \33226 , \33230 );
and \U$33041 ( \33356 , \33230 , \33235 );
and \U$33042 ( \33357 , \33226 , \33235 );
or \U$33043 ( \33358 , \33355 , \33356 , \33357 );
xor \U$33044 ( \33359 , \33354 , \33358 );
and \U$33045 ( \33360 , \33212 , \33216 );
and \U$33046 ( \33361 , \33216 , \33221 );
and \U$33047 ( \33362 , \33212 , \33221 );
or \U$33048 ( \33363 , \33360 , \33361 , \33362 );
xor \U$33049 ( \33364 , \33359 , \33363 );
xor \U$33050 ( \33365 , \33350 , \33364 );
and \U$33051 ( \33366 , \33222 , \33236 );
and \U$33052 ( \33367 , \33236 , \33248 );
and \U$33053 ( \33368 , \33222 , \33248 );
or \U$33054 ( \33369 , \33366 , \33367 , \33368 );
and \U$33055 ( \33370 , \22124 , \22598 );
and \U$33056 ( \33371 , \22089 , \22596 );
nor \U$33057 ( \33372 , \33370 , \33371 );
xnor \U$33058 ( \33373 , \33372 , \22608 );
and \U$33059 ( \33374 , \22145 , \22619 );
and \U$33060 ( \33375 , \22113 , \22617 );
nor \U$33061 ( \33376 , \33374 , \33375 );
xnor \U$33062 ( \33377 , \33376 , \22629 );
xor \U$33063 ( \33378 , \33373 , \33377 );
and \U$33064 ( \33379 , \22167 , \22641 );
and \U$33065 ( \33380 , \22134 , \22639 );
nor \U$33066 ( \33381 , \33379 , \33380 );
xnor \U$33067 ( \33382 , \33381 , \22651 );
xor \U$33068 ( \33383 , \33378 , \33382 );
and \U$33069 ( \33384 , \22894 , \22530 );
and \U$33070 ( \33385 , \23230 , \22528 );
nor \U$33071 ( \33386 , \33384 , \33385 );
xnor \U$33072 ( \33387 , \33386 , \22540 );
and \U$33073 ( \33388 , \22081 , \22551 );
and \U$33074 ( \33389 , \22858 , \22549 );
nor \U$33075 ( \33390 , \33388 , \33389 );
xnor \U$33076 ( \33391 , \33390 , \22561 );
xor \U$33077 ( \33392 , \33387 , \33391 );
and \U$33078 ( \33393 , \22100 , \22573 );
and \U$33079 ( \33394 , \22071 , \22571 );
nor \U$33080 ( \33395 , \33393 , \33394 );
xnor \U$33081 ( \33396 , \33395 , \22583 );
xor \U$33082 ( \33397 , \33392 , \33396 );
xor \U$33083 ( \33398 , \33383 , \33397 );
and \U$33084 ( \33399 , \21990 , \22463 );
not \U$33085 ( \33400 , \33399 );
xnor \U$33086 ( \33401 , \33400 , \22473 );
and \U$33087 ( \33402 , \22001 , \22484 );
and \U$33088 ( \33403 , \21977 , \22482 );
nor \U$33089 ( \33404 , \33402 , \33403 );
xnor \U$33090 ( \33405 , \33404 , \22494 );
xor \U$33091 ( \33406 , \33401 , \33405 );
and \U$33092 ( \33407 , \23329 , \22506 );
and \U$33093 ( \33408 , \22030 , \22504 );
nor \U$33094 ( \33409 , \33407 , \33408 );
xnor \U$33095 ( \33410 , \33409 , \22516 );
xor \U$33096 ( \33411 , \33406 , \33410 );
xor \U$33097 ( \33412 , \33398 , \33411 );
xor \U$33098 ( \33413 , \33369 , \33412 );
and \U$33099 ( \33414 , \22294 , \21978 );
not \U$33100 ( \33415 , \33414 );
and \U$33101 ( \33416 , \22262 , \23173 );
and \U$33102 ( \33417 , \22224 , \22999 );
nor \U$33103 ( \33418 , \33416 , \33417 );
xnor \U$33104 ( \33419 , \33418 , \22016 );
and \U$33105 ( \33420 , \22283 , \22021 );
and \U$33106 ( \33421 , \22251 , \22019 );
nor \U$33107 ( \33422 , \33420 , \33421 );
xnor \U$33108 ( \33423 , \33422 , \21595 );
xor \U$33109 ( \33424 , \33419 , \33423 );
and \U$33110 ( \33425 , \22305 , \21983 );
and \U$33111 ( \33426 , \22272 , \21981 );
nor \U$33112 ( \33427 , \33425 , \33426 );
xnor \U$33113 ( \33428 , \33427 , \21995 );
xor \U$33114 ( \33429 , \33424 , \33428 );
xor \U$33115 ( \33430 , \33415 , \33429 );
and \U$33116 ( \33431 , \22192 , \22671 );
and \U$33117 ( \33432 , \22156 , \22669 );
nor \U$33118 ( \33433 , \33431 , \33432 );
xnor \U$33119 ( \33434 , \33433 , \22681 );
and \U$33120 ( \33435 , \22213 , \22691 );
and \U$33121 ( \33436 , \22181 , \22689 );
nor \U$33122 ( \33437 , \33435 , \33436 );
xnor \U$33123 ( \33438 , \33437 , \22701 );
xor \U$33124 ( \33439 , \33434 , \33438 );
and \U$33125 ( \33440 , \22235 , \22720 );
and \U$33126 ( \33441 , \22202 , \22707 );
nor \U$33127 ( \33442 , \33440 , \33441 );
xnor \U$33128 ( \33443 , \33442 , \22067 );
xor \U$33129 ( \33444 , \33439 , \33443 );
xor \U$33130 ( \33445 , \33430 , \33444 );
xor \U$33131 ( \33446 , \33413 , \33445 );
xor \U$33132 ( \33447 , \33365 , \33446 );
and \U$33133 ( \33448 , \33193 , \33197 );
and \U$33134 ( \33449 , \33197 , \33202 );
and \U$33135 ( \33450 , \33193 , \33202 );
or \U$33136 ( \33451 , \33448 , \33449 , \33450 );
and \U$33137 ( \33452 , \33182 , \33186 );
and \U$33138 ( \33453 , \33186 , \33188 );
and \U$33139 ( \33454 , \33182 , \33188 );
or \U$33140 ( \33455 , \33452 , \33453 , \33454 );
xor \U$33141 ( \33456 , \33451 , \33455 );
and \U$33142 ( \33457 , \33256 , \33270 );
and \U$33143 ( \33458 , \33270 , \33285 );
and \U$33144 ( \33459 , \33256 , \33285 );
or \U$33145 ( \33460 , \33457 , \33458 , \33459 );
xor \U$33146 ( \33461 , \33456 , \33460 );
xor \U$33147 ( \33462 , \33447 , \33461 );
xor \U$33148 ( \33463 , \33339 , \33462 );
xor \U$33149 ( \33464 , \33330 , \33463 );
xor \U$33150 ( \33465 , \33314 , \33464 );
and \U$33151 ( \33466 , \33153 , \33305 );
nor \U$33152 ( \33467 , \33465 , \33466 );
and \U$33153 ( \33468 , \33318 , \33329 );
and \U$33154 ( \33469 , \33329 , \33463 );
and \U$33155 ( \33470 , \33318 , \33463 );
or \U$33156 ( \33471 , \33468 , \33469 , \33470 );
and \U$33157 ( \33472 , \33334 , \33338 );
and \U$33158 ( \33473 , \33338 , \33462 );
and \U$33159 ( \33474 , \33334 , \33462 );
or \U$33160 ( \33475 , \33472 , \33473 , \33474 );
and \U$33161 ( \33476 , \33451 , \33455 );
and \U$33162 ( \33477 , \33455 , \33460 );
and \U$33163 ( \33478 , \33451 , \33460 );
or \U$33164 ( \33479 , \33476 , \33477 , \33478 );
and \U$33165 ( \33480 , \33369 , \33412 );
and \U$33166 ( \33481 , \33412 , \33445 );
and \U$33167 ( \33482 , \33369 , \33445 );
or \U$33168 ( \33483 , \33480 , \33481 , \33482 );
xor \U$33169 ( \33484 , \33479 , \33483 );
and \U$33170 ( \33485 , \33350 , \33364 );
xor \U$33171 ( \33486 , \33484 , \33485 );
xor \U$33172 ( \33487 , \33475 , \33486 );
and \U$33173 ( \33488 , \33322 , \33326 );
and \U$33174 ( \33489 , \33326 , \33328 );
and \U$33175 ( \33490 , \33322 , \33328 );
or \U$33176 ( \33491 , \33488 , \33489 , \33490 );
and \U$33177 ( \33492 , \33365 , \33446 );
and \U$33178 ( \33493 , \33446 , \33461 );
and \U$33179 ( \33494 , \33365 , \33461 );
or \U$33180 ( \33495 , \33492 , \33493 , \33494 );
xor \U$33181 ( \33496 , \33491 , \33495 );
and \U$33182 ( \33497 , \33434 , \33438 );
and \U$33183 ( \33498 , \33438 , \33443 );
and \U$33184 ( \33499 , \33434 , \33443 );
or \U$33185 ( \33500 , \33497 , \33498 , \33499 );
and \U$33186 ( \33501 , \33419 , \33423 );
and \U$33187 ( \33502 , \33423 , \33428 );
and \U$33188 ( \33503 , \33419 , \33428 );
or \U$33189 ( \33504 , \33501 , \33502 , \33503 );
xor \U$33190 ( \33505 , \33500 , \33504 );
xor \U$33191 ( \33506 , \33505 , \33414 );
and \U$33192 ( \33507 , \33401 , \33405 );
and \U$33193 ( \33508 , \33405 , \33410 );
and \U$33194 ( \33509 , \33401 , \33410 );
or \U$33195 ( \33510 , \33507 , \33508 , \33509 );
and \U$33196 ( \33511 , \33387 , \33391 );
and \U$33197 ( \33512 , \33391 , \33396 );
and \U$33198 ( \33513 , \33387 , \33396 );
or \U$33199 ( \33514 , \33511 , \33512 , \33513 );
xor \U$33200 ( \33515 , \33510 , \33514 );
and \U$33201 ( \33516 , \33373 , \33377 );
and \U$33202 ( \33517 , \33377 , \33382 );
and \U$33203 ( \33518 , \33373 , \33382 );
or \U$33204 ( \33519 , \33516 , \33517 , \33518 );
xor \U$33205 ( \33520 , \33515 , \33519 );
xor \U$33206 ( \33521 , \33506 , \33520 );
and \U$33207 ( \33522 , \33383 , \33397 );
and \U$33208 ( \33523 , \33397 , \33411 );
and \U$33209 ( \33524 , \33383 , \33411 );
or \U$33210 ( \33525 , \33522 , \33523 , \33524 );
and \U$33211 ( \33526 , \22089 , \22598 );
and \U$33212 ( \33527 , \22100 , \22596 );
nor \U$33213 ( \33528 , \33526 , \33527 );
xnor \U$33214 ( \33529 , \33528 , \22608 );
and \U$33215 ( \33530 , \22113 , \22619 );
and \U$33216 ( \33531 , \22124 , \22617 );
nor \U$33217 ( \33532 , \33530 , \33531 );
xnor \U$33218 ( \33533 , \33532 , \22629 );
xor \U$33219 ( \33534 , \33529 , \33533 );
and \U$33220 ( \33535 , \22134 , \22641 );
and \U$33221 ( \33536 , \22145 , \22639 );
nor \U$33222 ( \33537 , \33535 , \33536 );
xnor \U$33223 ( \33538 , \33537 , \22651 );
xor \U$33224 ( \33539 , \33534 , \33538 );
and \U$33225 ( \33540 , \23230 , \22530 );
and \U$33226 ( \33541 , \23329 , \22528 );
nor \U$33227 ( \33542 , \33540 , \33541 );
xnor \U$33228 ( \33543 , \33542 , \22540 );
and \U$33229 ( \33544 , \22858 , \22551 );
and \U$33230 ( \33545 , \22894 , \22549 );
nor \U$33231 ( \33546 , \33544 , \33545 );
xnor \U$33232 ( \33547 , \33546 , \22561 );
xor \U$33233 ( \33548 , \33543 , \33547 );
and \U$33234 ( \33549 , \22071 , \22573 );
and \U$33235 ( \33550 , \22081 , \22571 );
nor \U$33236 ( \33551 , \33549 , \33550 );
xnor \U$33237 ( \33552 , \33551 , \22583 );
xor \U$33238 ( \33553 , \33548 , \33552 );
xor \U$33239 ( \33554 , \33539 , \33553 );
not \U$33240 ( \33555 , \22473 );
and \U$33241 ( \33556 , \21977 , \22484 );
and \U$33242 ( \33557 , \21990 , \22482 );
nor \U$33243 ( \33558 , \33556 , \33557 );
xnor \U$33244 ( \33559 , \33558 , \22494 );
xor \U$33245 ( \33560 , \33555 , \33559 );
and \U$33246 ( \33561 , \22030 , \22506 );
and \U$33247 ( \33562 , \22001 , \22504 );
nor \U$33248 ( \33563 , \33561 , \33562 );
xnor \U$33249 ( \33564 , \33563 , \22516 );
xor \U$33250 ( \33565 , \33560 , \33564 );
xor \U$33251 ( \33566 , \33554 , \33565 );
xor \U$33252 ( \33567 , \33525 , \33566 );
and \U$33253 ( \33568 , \22305 , \21978 );
and \U$33254 ( \33569 , \22224 , \23173 );
and \U$33255 ( \33570 , \22235 , \22999 );
nor \U$33256 ( \33571 , \33569 , \33570 );
xnor \U$33257 ( \33572 , \33571 , \22016 );
and \U$33258 ( \33573 , \22251 , \22021 );
and \U$33259 ( \33574 , \22262 , \22019 );
nor \U$33260 ( \33575 , \33573 , \33574 );
xnor \U$33261 ( \33576 , \33575 , \21595 );
xor \U$33262 ( \33577 , \33572 , \33576 );
and \U$33263 ( \33578 , \22272 , \21983 );
and \U$33264 ( \33579 , \22283 , \21981 );
nor \U$33265 ( \33580 , \33578 , \33579 );
xnor \U$33266 ( \33581 , \33580 , \21995 );
xor \U$33267 ( \33582 , \33577 , \33581 );
xor \U$33268 ( \33583 , \33568 , \33582 );
and \U$33269 ( \33584 , \22156 , \22671 );
and \U$33270 ( \33585 , \22167 , \22669 );
nor \U$33271 ( \33586 , \33584 , \33585 );
xnor \U$33272 ( \33587 , \33586 , \22681 );
and \U$33273 ( \33588 , \22181 , \22691 );
and \U$33274 ( \33589 , \22192 , \22689 );
nor \U$33275 ( \33590 , \33588 , \33589 );
xnor \U$33276 ( \33591 , \33590 , \22701 );
xor \U$33277 ( \33592 , \33587 , \33591 );
and \U$33278 ( \33593 , \22202 , \22720 );
and \U$33279 ( \33594 , \22213 , \22707 );
nor \U$33280 ( \33595 , \33593 , \33594 );
xnor \U$33281 ( \33596 , \33595 , \22067 );
xor \U$33282 ( \33597 , \33592 , \33596 );
xor \U$33283 ( \33598 , \33583 , \33597 );
xor \U$33284 ( \33599 , \33567 , \33598 );
xor \U$33285 ( \33600 , \33521 , \33599 );
and \U$33286 ( \33601 , \33354 , \33358 );
and \U$33287 ( \33602 , \33358 , \33363 );
and \U$33288 ( \33603 , \33354 , \33363 );
or \U$33289 ( \33604 , \33601 , \33602 , \33603 );
and \U$33290 ( \33605 , \33343 , \33347 );
and \U$33291 ( \33606 , \33347 , \33349 );
and \U$33292 ( \33607 , \33343 , \33349 );
or \U$33293 ( \33608 , \33605 , \33606 , \33607 );
xor \U$33294 ( \33609 , \33604 , \33608 );
and \U$33295 ( \33610 , \33415 , \33429 );
and \U$33296 ( \33611 , \33429 , \33444 );
and \U$33297 ( \33612 , \33415 , \33444 );
or \U$33298 ( \33613 , \33610 , \33611 , \33612 );
xor \U$33299 ( \33614 , \33609 , \33613 );
xor \U$33300 ( \33615 , \33600 , \33614 );
xor \U$33301 ( \33616 , \33496 , \33615 );
xor \U$33302 ( \33617 , \33487 , \33616 );
xor \U$33303 ( \33618 , \33471 , \33617 );
and \U$33304 ( \33619 , \33314 , \33464 );
nor \U$33305 ( \33620 , \33618 , \33619 );
nor \U$33306 ( \33621 , \33467 , \33620 );
and \U$33307 ( \33622 , \33475 , \33486 );
and \U$33308 ( \33623 , \33486 , \33616 );
and \U$33309 ( \33624 , \33475 , \33616 );
or \U$33310 ( \33625 , \33622 , \33623 , \33624 );
and \U$33311 ( \33626 , \33491 , \33495 );
and \U$33312 ( \33627 , \33495 , \33615 );
and \U$33313 ( \33628 , \33491 , \33615 );
or \U$33314 ( \33629 , \33626 , \33627 , \33628 );
and \U$33315 ( \33630 , \33604 , \33608 );
and \U$33316 ( \33631 , \33608 , \33613 );
and \U$33317 ( \33632 , \33604 , \33613 );
or \U$33318 ( \33633 , \33630 , \33631 , \33632 );
and \U$33319 ( \33634 , \33525 , \33566 );
and \U$33320 ( \33635 , \33566 , \33598 );
and \U$33321 ( \33636 , \33525 , \33598 );
or \U$33322 ( \33637 , \33634 , \33635 , \33636 );
xor \U$33323 ( \33638 , \33633 , \33637 );
and \U$33324 ( \33639 , \33506 , \33520 );
xor \U$33325 ( \33640 , \33638 , \33639 );
xor \U$33326 ( \33641 , \33629 , \33640 );
and \U$33327 ( \33642 , \33479 , \33483 );
and \U$33328 ( \33643 , \33483 , \33485 );
and \U$33329 ( \33644 , \33479 , \33485 );
or \U$33330 ( \33645 , \33642 , \33643 , \33644 );
and \U$33331 ( \33646 , \33521 , \33599 );
and \U$33332 ( \33647 , \33599 , \33614 );
and \U$33333 ( \33648 , \33521 , \33614 );
or \U$33334 ( \33649 , \33646 , \33647 , \33648 );
xor \U$33335 ( \33650 , \33645 , \33649 );
and \U$33336 ( \33651 , \22262 , \22021 );
and \U$33337 ( \33652 , \22224 , \22019 );
nor \U$33338 ( \33653 , \33651 , \33652 );
xnor \U$33339 ( \33654 , \33653 , \21595 );
and \U$33340 ( \33655 , \22283 , \21983 );
and \U$33341 ( \33656 , \22251 , \21981 );
nor \U$33342 ( \33657 , \33655 , \33656 );
xnor \U$33343 ( \33658 , \33657 , \21995 );
xor \U$33344 ( \33659 , \33654 , \33658 );
and \U$33345 ( \33660 , \22272 , \21978 );
xor \U$33346 ( \33661 , \33659 , \33660 );
and \U$33347 ( \33662 , \22192 , \22691 );
and \U$33348 ( \33663 , \22156 , \22689 );
nor \U$33349 ( \33664 , \33662 , \33663 );
xnor \U$33350 ( \33665 , \33664 , \22701 );
and \U$33351 ( \33666 , \22213 , \22720 );
and \U$33352 ( \33667 , \22181 , \22707 );
nor \U$33353 ( \33668 , \33666 , \33667 );
xnor \U$33354 ( \33669 , \33668 , \22067 );
xor \U$33355 ( \33670 , \33665 , \33669 );
and \U$33356 ( \33671 , \22235 , \23173 );
and \U$33357 ( \33672 , \22202 , \22999 );
nor \U$33358 ( \33673 , \33671 , \33672 );
xnor \U$33359 ( \33674 , \33673 , \22016 );
xor \U$33360 ( \33675 , \33670 , \33674 );
xor \U$33361 ( \33676 , \33661 , \33675 );
and \U$33362 ( \33677 , \22124 , \22619 );
and \U$33363 ( \33678 , \22089 , \22617 );
nor \U$33364 ( \33679 , \33677 , \33678 );
xnor \U$33365 ( \33680 , \33679 , \22629 );
and \U$33366 ( \33681 , \22145 , \22641 );
and \U$33367 ( \33682 , \22113 , \22639 );
nor \U$33368 ( \33683 , \33681 , \33682 );
xnor \U$33369 ( \33684 , \33683 , \22651 );
xor \U$33370 ( \33685 , \33680 , \33684 );
and \U$33371 ( \33686 , \22167 , \22671 );
and \U$33372 ( \33687 , \22134 , \22669 );
nor \U$33373 ( \33688 , \33686 , \33687 );
xnor \U$33374 ( \33689 , \33688 , \22681 );
xor \U$33375 ( \33690 , \33685 , \33689 );
xor \U$33376 ( \33691 , \33676 , \33690 );
and \U$33377 ( \33692 , \33587 , \33591 );
and \U$33378 ( \33693 , \33591 , \33596 );
and \U$33379 ( \33694 , \33587 , \33596 );
or \U$33380 ( \33695 , \33692 , \33693 , \33694 );
and \U$33381 ( \33696 , \33572 , \33576 );
and \U$33382 ( \33697 , \33576 , \33581 );
and \U$33383 ( \33698 , \33572 , \33581 );
or \U$33384 ( \33699 , \33696 , \33697 , \33698 );
xnor \U$33385 ( \33700 , \33695 , \33699 );
xor \U$33386 ( \33701 , \33691 , \33700 );
and \U$33387 ( \33702 , \33555 , \33559 );
and \U$33388 ( \33703 , \33559 , \33564 );
and \U$33389 ( \33704 , \33555 , \33564 );
or \U$33390 ( \33705 , \33702 , \33703 , \33704 );
and \U$33391 ( \33706 , \33543 , \33547 );
and \U$33392 ( \33707 , \33547 , \33552 );
and \U$33393 ( \33708 , \33543 , \33552 );
or \U$33394 ( \33709 , \33706 , \33707 , \33708 );
xor \U$33395 ( \33710 , \33705 , \33709 );
and \U$33396 ( \33711 , \33529 , \33533 );
and \U$33397 ( \33712 , \33533 , \33538 );
and \U$33398 ( \33713 , \33529 , \33538 );
or \U$33399 ( \33714 , \33711 , \33712 , \33713 );
xor \U$33400 ( \33715 , \33710 , \33714 );
xor \U$33401 ( \33716 , \33701 , \33715 );
and \U$33402 ( \33717 , \33539 , \33553 );
and \U$33403 ( \33718 , \33553 , \33565 );
and \U$33404 ( \33719 , \33539 , \33565 );
or \U$33405 ( \33720 , \33717 , \33718 , \33719 );
and \U$33406 ( \33721 , \22894 , \22551 );
and \U$33407 ( \33722 , \23230 , \22549 );
nor \U$33408 ( \33723 , \33721 , \33722 );
xnor \U$33409 ( \33724 , \33723 , \22561 );
and \U$33410 ( \33725 , \22081 , \22573 );
and \U$33411 ( \33726 , \22858 , \22571 );
nor \U$33412 ( \33727 , \33725 , \33726 );
xnor \U$33413 ( \33728 , \33727 , \22583 );
xor \U$33414 ( \33729 , \33724 , \33728 );
and \U$33415 ( \33730 , \22100 , \22598 );
and \U$33416 ( \33731 , \22071 , \22596 );
nor \U$33417 ( \33732 , \33730 , \33731 );
xnor \U$33418 ( \33733 , \33732 , \22608 );
xor \U$33419 ( \33734 , \33729 , \33733 );
xor \U$33420 ( \33735 , \33720 , \33734 );
and \U$33421 ( \33736 , \21990 , \22484 );
not \U$33422 ( \33737 , \33736 );
xnor \U$33423 ( \33738 , \33737 , \22494 );
and \U$33424 ( \33739 , \22001 , \22506 );
and \U$33425 ( \33740 , \21977 , \22504 );
nor \U$33426 ( \33741 , \33739 , \33740 );
xnor \U$33427 ( \33742 , \33741 , \22516 );
xor \U$33428 ( \33743 , \33738 , \33742 );
and \U$33429 ( \33744 , \23329 , \22530 );
and \U$33430 ( \33745 , \22030 , \22528 );
nor \U$33431 ( \33746 , \33744 , \33745 );
xnor \U$33432 ( \33747 , \33746 , \22540 );
xor \U$33433 ( \33748 , \33743 , \33747 );
xor \U$33434 ( \33749 , \33735 , \33748 );
xor \U$33435 ( \33750 , \33716 , \33749 );
and \U$33436 ( \33751 , \33510 , \33514 );
and \U$33437 ( \33752 , \33514 , \33519 );
and \U$33438 ( \33753 , \33510 , \33519 );
or \U$33439 ( \33754 , \33751 , \33752 , \33753 );
and \U$33440 ( \33755 , \33500 , \33504 );
and \U$33441 ( \33756 , \33504 , \33414 );
and \U$33442 ( \33757 , \33500 , \33414 );
or \U$33443 ( \33758 , \33755 , \33756 , \33757 );
xor \U$33444 ( \33759 , \33754 , \33758 );
and \U$33445 ( \33760 , \33568 , \33582 );
and \U$33446 ( \33761 , \33582 , \33597 );
and \U$33447 ( \33762 , \33568 , \33597 );
or \U$33448 ( \33763 , \33760 , \33761 , \33762 );
xor \U$33449 ( \33764 , \33759 , \33763 );
xor \U$33450 ( \33765 , \33750 , \33764 );
xor \U$33451 ( \33766 , \33650 , \33765 );
xor \U$33452 ( \33767 , \33641 , \33766 );
xor \U$33453 ( \33768 , \33625 , \33767 );
and \U$33454 ( \33769 , \33471 , \33617 );
nor \U$33455 ( \33770 , \33768 , \33769 );
and \U$33456 ( \33771 , \33629 , \33640 );
and \U$33457 ( \33772 , \33640 , \33766 );
and \U$33458 ( \33773 , \33629 , \33766 );
or \U$33459 ( \33774 , \33771 , \33772 , \33773 );
and \U$33460 ( \33775 , \33645 , \33649 );
and \U$33461 ( \33776 , \33649 , \33765 );
and \U$33462 ( \33777 , \33645 , \33765 );
or \U$33463 ( \33778 , \33775 , \33776 , \33777 );
and \U$33464 ( \33779 , \33754 , \33758 );
and \U$33465 ( \33780 , \33758 , \33763 );
and \U$33466 ( \33781 , \33754 , \33763 );
or \U$33467 ( \33782 , \33779 , \33780 , \33781 );
and \U$33468 ( \33783 , \33720 , \33734 );
and \U$33469 ( \33784 , \33734 , \33748 );
and \U$33470 ( \33785 , \33720 , \33748 );
or \U$33471 ( \33786 , \33783 , \33784 , \33785 );
xor \U$33472 ( \33787 , \33782 , \33786 );
and \U$33473 ( \33788 , \33691 , \33700 );
and \U$33474 ( \33789 , \33700 , \33715 );
and \U$33475 ( \33790 , \33691 , \33715 );
or \U$33476 ( \33791 , \33788 , \33789 , \33790 );
xor \U$33477 ( \33792 , \33787 , \33791 );
xor \U$33478 ( \33793 , \33778 , \33792 );
and \U$33479 ( \33794 , \33633 , \33637 );
and \U$33480 ( \33795 , \33637 , \33639 );
and \U$33481 ( \33796 , \33633 , \33639 );
or \U$33482 ( \33797 , \33794 , \33795 , \33796 );
and \U$33483 ( \33798 , \33716 , \33749 );
and \U$33484 ( \33799 , \33749 , \33764 );
and \U$33485 ( \33800 , \33716 , \33764 );
or \U$33486 ( \33801 , \33798 , \33799 , \33800 );
xor \U$33487 ( \33802 , \33797 , \33801 );
and \U$33488 ( \33803 , \33738 , \33742 );
and \U$33489 ( \33804 , \33742 , \33747 );
and \U$33490 ( \33805 , \33738 , \33747 );
or \U$33491 ( \33806 , \33803 , \33804 , \33805 );
and \U$33492 ( \33807 , \33724 , \33728 );
and \U$33493 ( \33808 , \33728 , \33733 );
and \U$33494 ( \33809 , \33724 , \33733 );
or \U$33495 ( \33810 , \33807 , \33808 , \33809 );
xor \U$33496 ( \33811 , \33806 , \33810 );
and \U$33497 ( \33812 , \33680 , \33684 );
and \U$33498 ( \33813 , \33684 , \33689 );
and \U$33499 ( \33814 , \33680 , \33689 );
or \U$33500 ( \33815 , \33812 , \33813 , \33814 );
xor \U$33501 ( \33816 , \33811 , \33815 );
not \U$33502 ( \33817 , \22494 );
and \U$33503 ( \33818 , \21977 , \22506 );
and \U$33504 ( \33819 , \21990 , \22504 );
nor \U$33505 ( \33820 , \33818 , \33819 );
xnor \U$33506 ( \33821 , \33820 , \22516 );
xor \U$33507 ( \33822 , \33817 , \33821 );
and \U$33508 ( \33823 , \22030 , \22530 );
and \U$33509 ( \33824 , \22001 , \22528 );
nor \U$33510 ( \33825 , \33823 , \33824 );
xnor \U$33511 ( \33826 , \33825 , \22540 );
xor \U$33512 ( \33827 , \33822 , \33826 );
and \U$33513 ( \33828 , \22156 , \22691 );
and \U$33514 ( \33829 , \22167 , \22689 );
nor \U$33515 ( \33830 , \33828 , \33829 );
xnor \U$33516 ( \33831 , \33830 , \22701 );
and \U$33517 ( \33832 , \22181 , \22720 );
and \U$33518 ( \33833 , \22192 , \22707 );
nor \U$33519 ( \33834 , \33832 , \33833 );
xnor \U$33520 ( \33835 , \33834 , \22067 );
xor \U$33521 ( \33836 , \33831 , \33835 );
and \U$33522 ( \33837 , \22202 , \23173 );
and \U$33523 ( \33838 , \22213 , \22999 );
nor \U$33524 ( \33839 , \33837 , \33838 );
xnor \U$33525 ( \33840 , \33839 , \22016 );
xor \U$33526 ( \33841 , \33836 , \33840 );
and \U$33527 ( \33842 , \22089 , \22619 );
and \U$33528 ( \33843 , \22100 , \22617 );
nor \U$33529 ( \33844 , \33842 , \33843 );
xnor \U$33530 ( \33845 , \33844 , \22629 );
and \U$33531 ( \33846 , \22113 , \22641 );
and \U$33532 ( \33847 , \22124 , \22639 );
nor \U$33533 ( \33848 , \33846 , \33847 );
xnor \U$33534 ( \33849 , \33848 , \22651 );
xor \U$33535 ( \33850 , \33845 , \33849 );
and \U$33536 ( \33851 , \22134 , \22671 );
and \U$33537 ( \33852 , \22145 , \22669 );
nor \U$33538 ( \33853 , \33851 , \33852 );
xnor \U$33539 ( \33854 , \33853 , \22681 );
xor \U$33540 ( \33855 , \33850 , \33854 );
xor \U$33541 ( \33856 , \33841 , \33855 );
and \U$33542 ( \33857 , \23230 , \22551 );
and \U$33543 ( \33858 , \23329 , \22549 );
nor \U$33544 ( \33859 , \33857 , \33858 );
xnor \U$33545 ( \33860 , \33859 , \22561 );
and \U$33546 ( \33861 , \22858 , \22573 );
and \U$33547 ( \33862 , \22894 , \22571 );
nor \U$33548 ( \33863 , \33861 , \33862 );
xnor \U$33549 ( \33864 , \33863 , \22583 );
xor \U$33550 ( \33865 , \33860 , \33864 );
and \U$33551 ( \33866 , \22071 , \22598 );
and \U$33552 ( \33867 , \22081 , \22596 );
nor \U$33553 ( \33868 , \33866 , \33867 );
xnor \U$33554 ( \33869 , \33868 , \22608 );
xor \U$33555 ( \33870 , \33865 , \33869 );
xor \U$33556 ( \33871 , \33856 , \33870 );
xor \U$33557 ( \33872 , \33827 , \33871 );
and \U$33558 ( \33873 , \33665 , \33669 );
and \U$33559 ( \33874 , \33669 , \33674 );
and \U$33560 ( \33875 , \33665 , \33674 );
or \U$33561 ( \33876 , \33873 , \33874 , \33875 );
and \U$33562 ( \33877 , \33654 , \33658 );
and \U$33563 ( \33878 , \33658 , \33660 );
and \U$33564 ( \33879 , \33654 , \33660 );
or \U$33565 ( \33880 , \33877 , \33878 , \33879 );
xor \U$33566 ( \33881 , \33876 , \33880 );
and \U$33567 ( \33882 , \22224 , \22021 );
and \U$33568 ( \33883 , \22235 , \22019 );
nor \U$33569 ( \33884 , \33882 , \33883 );
xnor \U$33570 ( \33885 , \33884 , \21595 );
and \U$33571 ( \33886 , \22251 , \21983 );
and \U$33572 ( \33887 , \22262 , \21981 );
nor \U$33573 ( \33888 , \33886 , \33887 );
xnor \U$33574 ( \33889 , \33888 , \21995 );
xor \U$33575 ( \33890 , \33885 , \33889 );
and \U$33576 ( \33891 , \22283 , \21978 );
xor \U$33577 ( \33892 , \33890 , \33891 );
xor \U$33578 ( \33893 , \33881 , \33892 );
xor \U$33579 ( \33894 , \33872 , \33893 );
xor \U$33580 ( \33895 , \33816 , \33894 );
and \U$33581 ( \33896 , \33705 , \33709 );
and \U$33582 ( \33897 , \33709 , \33714 );
and \U$33583 ( \33898 , \33705 , \33714 );
or \U$33584 ( \33899 , \33896 , \33897 , \33898 );
or \U$33585 ( \33900 , \33695 , \33699 );
xor \U$33586 ( \33901 , \33899 , \33900 );
and \U$33587 ( \33902 , \33661 , \33675 );
and \U$33588 ( \33903 , \33675 , \33690 );
and \U$33589 ( \33904 , \33661 , \33690 );
or \U$33590 ( \33905 , \33902 , \33903 , \33904 );
xor \U$33591 ( \33906 , \33901 , \33905 );
xor \U$33592 ( \33907 , \33895 , \33906 );
xor \U$33593 ( \33908 , \33802 , \33907 );
xor \U$33594 ( \33909 , \33793 , \33908 );
xor \U$33595 ( \33910 , \33774 , \33909 );
and \U$33596 ( \33911 , \33625 , \33767 );
nor \U$33597 ( \33912 , \33910 , \33911 );
nor \U$33598 ( \33913 , \33770 , \33912 );
nand \U$33599 ( \33914 , \33621 , \33913 );
nor \U$33600 ( \33915 , \33310 , \33914 );
and \U$33601 ( \33916 , \33778 , \33792 );
and \U$33602 ( \33917 , \33792 , \33908 );
and \U$33603 ( \33918 , \33778 , \33908 );
or \U$33604 ( \33919 , \33916 , \33917 , \33918 );
and \U$33605 ( \33920 , \33797 , \33801 );
and \U$33606 ( \33921 , \33801 , \33907 );
and \U$33607 ( \33922 , \33797 , \33907 );
or \U$33608 ( \33923 , \33920 , \33921 , \33922 );
and \U$33609 ( \33924 , \33806 , \33810 );
and \U$33610 ( \33925 , \33810 , \33815 );
and \U$33611 ( \33926 , \33806 , \33815 );
or \U$33612 ( \33927 , \33924 , \33925 , \33926 );
and \U$33613 ( \33928 , \33876 , \33880 );
and \U$33614 ( \33929 , \33880 , \33892 );
and \U$33615 ( \33930 , \33876 , \33892 );
or \U$33616 ( \33931 , \33928 , \33929 , \33930 );
xor \U$33617 ( \33932 , \33927 , \33931 );
and \U$33618 ( \33933 , \33841 , \33855 );
and \U$33619 ( \33934 , \33855 , \33870 );
and \U$33620 ( \33935 , \33841 , \33870 );
or \U$33621 ( \33936 , \33933 , \33934 , \33935 );
xor \U$33622 ( \33937 , \33932 , \33936 );
and \U$33623 ( \33938 , \33899 , \33900 );
and \U$33624 ( \33939 , \33900 , \33905 );
and \U$33625 ( \33940 , \33899 , \33905 );
or \U$33626 ( \33941 , \33938 , \33939 , \33940 );
and \U$33627 ( \33942 , \33827 , \33871 );
and \U$33628 ( \33943 , \33871 , \33893 );
and \U$33629 ( \33944 , \33827 , \33893 );
or \U$33630 ( \33945 , \33942 , \33943 , \33944 );
xor \U$33631 ( \33946 , \33941 , \33945 );
and \U$33632 ( \33947 , \33817 , \33821 );
and \U$33633 ( \33948 , \33821 , \33826 );
and \U$33634 ( \33949 , \33817 , \33826 );
or \U$33635 ( \33950 , \33947 , \33948 , \33949 );
and \U$33636 ( \33951 , \33860 , \33864 );
and \U$33637 ( \33952 , \33864 , \33869 );
and \U$33638 ( \33953 , \33860 , \33869 );
or \U$33639 ( \33954 , \33951 , \33952 , \33953 );
xor \U$33640 ( \33955 , \33950 , \33954 );
and \U$33641 ( \33956 , \33845 , \33849 );
and \U$33642 ( \33957 , \33849 , \33854 );
and \U$33643 ( \33958 , \33845 , \33854 );
or \U$33644 ( \33959 , \33956 , \33957 , \33958 );
xor \U$33645 ( \33960 , \33955 , \33959 );
xor \U$33646 ( \33961 , \33946 , \33960 );
xor \U$33647 ( \33962 , \33937 , \33961 );
xor \U$33648 ( \33963 , \33923 , \33962 );
and \U$33649 ( \33964 , \33782 , \33786 );
and \U$33650 ( \33965 , \33786 , \33791 );
and \U$33651 ( \33966 , \33782 , \33791 );
or \U$33652 ( \33967 , \33964 , \33965 , \33966 );
and \U$33653 ( \33968 , \33816 , \33894 );
and \U$33654 ( \33969 , \33894 , \33906 );
and \U$33655 ( \33970 , \33816 , \33906 );
or \U$33656 ( \33971 , \33968 , \33969 , \33970 );
xor \U$33657 ( \33972 , \33967 , \33971 );
and \U$33658 ( \33973 , \21990 , \22506 );
not \U$33659 ( \33974 , \33973 );
xnor \U$33660 ( \33975 , \33974 , \22516 );
and \U$33661 ( \33976 , \22001 , \22530 );
and \U$33662 ( \33977 , \21977 , \22528 );
nor \U$33663 ( \33978 , \33976 , \33977 );
xnor \U$33664 ( \33979 , \33978 , \22540 );
xor \U$33665 ( \33980 , \33975 , \33979 );
and \U$33666 ( \33981 , \23329 , \22551 );
and \U$33667 ( \33982 , \22030 , \22549 );
nor \U$33668 ( \33983 , \33981 , \33982 );
xnor \U$33669 ( \33984 , \33983 , \22561 );
xor \U$33670 ( \33985 , \33980 , \33984 );
and \U$33671 ( \33986 , \22192 , \22720 );
and \U$33672 ( \33987 , \22156 , \22707 );
nor \U$33673 ( \33988 , \33986 , \33987 );
xnor \U$33674 ( \33989 , \33988 , \22067 );
and \U$33675 ( \33990 , \22213 , \23173 );
and \U$33676 ( \33991 , \22181 , \22999 );
nor \U$33677 ( \33992 , \33990 , \33991 );
xnor \U$33678 ( \33993 , \33992 , \22016 );
xor \U$33679 ( \33994 , \33989 , \33993 );
and \U$33680 ( \33995 , \22235 , \22021 );
and \U$33681 ( \33996 , \22202 , \22019 );
nor \U$33682 ( \33997 , \33995 , \33996 );
xnor \U$33683 ( \33998 , \33997 , \21595 );
xor \U$33684 ( \33999 , \33994 , \33998 );
and \U$33685 ( \34000 , \22124 , \22641 );
and \U$33686 ( \34001 , \22089 , \22639 );
nor \U$33687 ( \34002 , \34000 , \34001 );
xnor \U$33688 ( \34003 , \34002 , \22651 );
and \U$33689 ( \34004 , \22145 , \22671 );
and \U$33690 ( \34005 , \22113 , \22669 );
nor \U$33691 ( \34006 , \34004 , \34005 );
xnor \U$33692 ( \34007 , \34006 , \22681 );
xor \U$33693 ( \34008 , \34003 , \34007 );
and \U$33694 ( \34009 , \22167 , \22691 );
and \U$33695 ( \34010 , \22134 , \22689 );
nor \U$33696 ( \34011 , \34009 , \34010 );
xnor \U$33697 ( \34012 , \34011 , \22701 );
xor \U$33698 ( \34013 , \34008 , \34012 );
xor \U$33699 ( \34014 , \33999 , \34013 );
and \U$33700 ( \34015 , \22894 , \22573 );
and \U$33701 ( \34016 , \23230 , \22571 );
nor \U$33702 ( \34017 , \34015 , \34016 );
xnor \U$33703 ( \34018 , \34017 , \22583 );
and \U$33704 ( \34019 , \22081 , \22598 );
and \U$33705 ( \34020 , \22858 , \22596 );
nor \U$33706 ( \34021 , \34019 , \34020 );
xnor \U$33707 ( \34022 , \34021 , \22608 );
xor \U$33708 ( \34023 , \34018 , \34022 );
and \U$33709 ( \34024 , \22100 , \22619 );
and \U$33710 ( \34025 , \22071 , \22617 );
nor \U$33711 ( \34026 , \34024 , \34025 );
xnor \U$33712 ( \34027 , \34026 , \22629 );
xor \U$33713 ( \34028 , \34023 , \34027 );
xor \U$33714 ( \34029 , \34014 , \34028 );
xor \U$33715 ( \34030 , \33985 , \34029 );
and \U$33716 ( \34031 , \33831 , \33835 );
and \U$33717 ( \34032 , \33835 , \33840 );
and \U$33718 ( \34033 , \33831 , \33840 );
or \U$33719 ( \34034 , \34031 , \34032 , \34033 );
and \U$33720 ( \34035 , \33885 , \33889 );
and \U$33721 ( \34036 , \33889 , \33891 );
and \U$33722 ( \34037 , \33885 , \33891 );
or \U$33723 ( \34038 , \34035 , \34036 , \34037 );
xor \U$33724 ( \34039 , \34034 , \34038 );
and \U$33725 ( \34040 , \22262 , \21983 );
and \U$33726 ( \34041 , \22224 , \21981 );
nor \U$33727 ( \34042 , \34040 , \34041 );
xnor \U$33728 ( \34043 , \34042 , \21995 );
and \U$33729 ( \34044 , \22251 , \21978 );
xnor \U$33730 ( \34045 , \34043 , \34044 );
xor \U$33731 ( \34046 , \34039 , \34045 );
xor \U$33732 ( \34047 , \34030 , \34046 );
xor \U$33733 ( \34048 , \33972 , \34047 );
xor \U$33734 ( \34049 , \33963 , \34048 );
xor \U$33735 ( \34050 , \33919 , \34049 );
and \U$33736 ( \34051 , \33774 , \33909 );
nor \U$33737 ( \34052 , \34050 , \34051 );
and \U$33738 ( \34053 , \33923 , \33962 );
and \U$33739 ( \34054 , \33962 , \34048 );
and \U$33740 ( \34055 , \33923 , \34048 );
or \U$33741 ( \34056 , \34053 , \34054 , \34055 );
and \U$33742 ( \34057 , \33967 , \33971 );
and \U$33743 ( \34058 , \33971 , \34047 );
and \U$33744 ( \34059 , \33967 , \34047 );
or \U$33745 ( \34060 , \34057 , \34058 , \34059 );
and \U$33746 ( \34061 , \33937 , \33961 );
xor \U$33747 ( \34062 , \34060 , \34061 );
and \U$33748 ( \34063 , \33941 , \33945 );
and \U$33749 ( \34064 , \33945 , \33960 );
and \U$33750 ( \34065 , \33941 , \33960 );
or \U$33751 ( \34066 , \34063 , \34064 , \34065 );
and \U$33752 ( \34067 , \33975 , \33979 );
and \U$33753 ( \34068 , \33979 , \33984 );
and \U$33754 ( \34069 , \33975 , \33984 );
or \U$33755 ( \34070 , \34067 , \34068 , \34069 );
and \U$33756 ( \34071 , \34018 , \34022 );
and \U$33757 ( \34072 , \34022 , \34027 );
and \U$33758 ( \34073 , \34018 , \34027 );
or \U$33759 ( \34074 , \34071 , \34072 , \34073 );
xor \U$33760 ( \34075 , \34070 , \34074 );
and \U$33761 ( \34076 , \34003 , \34007 );
and \U$33762 ( \34077 , \34007 , \34012 );
and \U$33763 ( \34078 , \34003 , \34012 );
or \U$33764 ( \34079 , \34076 , \34077 , \34078 );
xor \U$33765 ( \34080 , \34075 , \34079 );
and \U$33766 ( \34081 , \23230 , \22573 );
and \U$33767 ( \34082 , \23329 , \22571 );
nor \U$33768 ( \34083 , \34081 , \34082 );
xnor \U$33769 ( \34084 , \34083 , \22583 );
and \U$33770 ( \34085 , \22858 , \22598 );
and \U$33771 ( \34086 , \22894 , \22596 );
nor \U$33772 ( \34087 , \34085 , \34086 );
xnor \U$33773 ( \34088 , \34087 , \22608 );
xor \U$33774 ( \34089 , \34084 , \34088 );
and \U$33775 ( \34090 , \22071 , \22619 );
and \U$33776 ( \34091 , \22081 , \22617 );
nor \U$33777 ( \34092 , \34090 , \34091 );
xnor \U$33778 ( \34093 , \34092 , \22629 );
xor \U$33779 ( \34094 , \34089 , \34093 );
not \U$33780 ( \34095 , \22516 );
and \U$33781 ( \34096 , \21977 , \22530 );
and \U$33782 ( \34097 , \21990 , \22528 );
nor \U$33783 ( \34098 , \34096 , \34097 );
xnor \U$33784 ( \34099 , \34098 , \22540 );
xor \U$33785 ( \34100 , \34095 , \34099 );
and \U$33786 ( \34101 , \22030 , \22551 );
and \U$33787 ( \34102 , \22001 , \22549 );
nor \U$33788 ( \34103 , \34101 , \34102 );
xnor \U$33789 ( \34104 , \34103 , \22561 );
xor \U$33790 ( \34105 , \34100 , \34104 );
xor \U$33791 ( \34106 , \34094 , \34105 );
and \U$33792 ( \34107 , \22262 , \21978 );
and \U$33793 ( \34108 , \22156 , \22720 );
and \U$33794 ( \34109 , \22167 , \22707 );
nor \U$33795 ( \34110 , \34108 , \34109 );
xnor \U$33796 ( \34111 , \34110 , \22067 );
and \U$33797 ( \34112 , \22181 , \23173 );
and \U$33798 ( \34113 , \22192 , \22999 );
nor \U$33799 ( \34114 , \34112 , \34113 );
xnor \U$33800 ( \34115 , \34114 , \22016 );
xor \U$33801 ( \34116 , \34111 , \34115 );
and \U$33802 ( \34117 , \22202 , \22021 );
and \U$33803 ( \34118 , \22213 , \22019 );
nor \U$33804 ( \34119 , \34117 , \34118 );
xnor \U$33805 ( \34120 , \34119 , \21595 );
xor \U$33806 ( \34121 , \34116 , \34120 );
xor \U$33807 ( \34122 , \34107 , \34121 );
and \U$33808 ( \34123 , \22089 , \22641 );
and \U$33809 ( \34124 , \22100 , \22639 );
nor \U$33810 ( \34125 , \34123 , \34124 );
xnor \U$33811 ( \34126 , \34125 , \22651 );
and \U$33812 ( \34127 , \22113 , \22671 );
and \U$33813 ( \34128 , \22124 , \22669 );
nor \U$33814 ( \34129 , \34127 , \34128 );
xnor \U$33815 ( \34130 , \34129 , \22681 );
xor \U$33816 ( \34131 , \34126 , \34130 );
and \U$33817 ( \34132 , \22134 , \22691 );
and \U$33818 ( \34133 , \22145 , \22689 );
nor \U$33819 ( \34134 , \34132 , \34133 );
xnor \U$33820 ( \34135 , \34134 , \22701 );
xor \U$33821 ( \34136 , \34131 , \34135 );
xor \U$33822 ( \34137 , \34122 , \34136 );
xor \U$33823 ( \34138 , \34106 , \34137 );
xor \U$33824 ( \34139 , \34080 , \34138 );
and \U$33825 ( \34140 , \33950 , \33954 );
and \U$33826 ( \34141 , \33954 , \33959 );
and \U$33827 ( \34142 , \33950 , \33959 );
or \U$33828 ( \34143 , \34140 , \34141 , \34142 );
and \U$33829 ( \34144 , \34034 , \34038 );
and \U$33830 ( \34145 , \34038 , \34045 );
and \U$33831 ( \34146 , \34034 , \34045 );
or \U$33832 ( \34147 , \34144 , \34145 , \34146 );
xor \U$33833 ( \34148 , \34143 , \34147 );
and \U$33834 ( \34149 , \33999 , \34013 );
and \U$33835 ( \34150 , \34013 , \34028 );
and \U$33836 ( \34151 , \33999 , \34028 );
or \U$33837 ( \34152 , \34149 , \34150 , \34151 );
xor \U$33838 ( \34153 , \34148 , \34152 );
xor \U$33839 ( \34154 , \34139 , \34153 );
xor \U$33840 ( \34155 , \34066 , \34154 );
and \U$33841 ( \34156 , \33927 , \33931 );
and \U$33842 ( \34157 , \33931 , \33936 );
and \U$33843 ( \34158 , \33927 , \33936 );
or \U$33844 ( \34159 , \34156 , \34157 , \34158 );
and \U$33845 ( \34160 , \33985 , \34029 );
and \U$33846 ( \34161 , \34029 , \34046 );
and \U$33847 ( \34162 , \33985 , \34046 );
or \U$33848 ( \34163 , \34160 , \34161 , \34162 );
xor \U$33849 ( \34164 , \34159 , \34163 );
and \U$33850 ( \34165 , \33989 , \33993 );
and \U$33851 ( \34166 , \33993 , \33998 );
and \U$33852 ( \34167 , \33989 , \33998 );
or \U$33853 ( \34168 , \34165 , \34166 , \34167 );
or \U$33854 ( \34169 , \34043 , \34044 );
xor \U$33855 ( \34170 , \34168 , \34169 );
and \U$33856 ( \34171 , \22224 , \21983 );
and \U$33857 ( \34172 , \22235 , \21981 );
nor \U$33858 ( \34173 , \34171 , \34172 );
xnor \U$33859 ( \34174 , \34173 , \21995 );
xor \U$33860 ( \34175 , \34170 , \34174 );
xor \U$33861 ( \34176 , \34164 , \34175 );
xor \U$33862 ( \34177 , \34155 , \34176 );
xor \U$33863 ( \34178 , \34062 , \34177 );
xor \U$33864 ( \34179 , \34056 , \34178 );
and \U$33865 ( \34180 , \33919 , \34049 );
nor \U$33866 ( \34181 , \34179 , \34180 );
nor \U$33867 ( \34182 , \34052 , \34181 );
and \U$33868 ( \34183 , \34060 , \34061 );
and \U$33869 ( \34184 , \34061 , \34177 );
and \U$33870 ( \34185 , \34060 , \34177 );
or \U$33871 ( \34186 , \34183 , \34184 , \34185 );
and \U$33872 ( \34187 , \34066 , \34154 );
and \U$33873 ( \34188 , \34154 , \34176 );
and \U$33874 ( \34189 , \34066 , \34176 );
or \U$33875 ( \34190 , \34187 , \34188 , \34189 );
and \U$33876 ( \34191 , \34143 , \34147 );
and \U$33877 ( \34192 , \34147 , \34152 );
and \U$33878 ( \34193 , \34143 , \34152 );
or \U$33879 ( \34194 , \34191 , \34192 , \34193 );
and \U$33880 ( \34195 , \34094 , \34105 );
and \U$33881 ( \34196 , \34105 , \34137 );
and \U$33882 ( \34197 , \34094 , \34137 );
or \U$33883 ( \34198 , \34195 , \34196 , \34197 );
xor \U$33884 ( \34199 , \34194 , \34198 );
and \U$33885 ( \34200 , \22124 , \22671 );
and \U$33886 ( \34201 , \22089 , \22669 );
nor \U$33887 ( \34202 , \34200 , \34201 );
xnor \U$33888 ( \34203 , \34202 , \22681 );
and \U$33889 ( \34204 , \22145 , \22691 );
and \U$33890 ( \34205 , \22113 , \22689 );
nor \U$33891 ( \34206 , \34204 , \34205 );
xnor \U$33892 ( \34207 , \34206 , \22701 );
xor \U$33893 ( \34208 , \34203 , \34207 );
and \U$33894 ( \34209 , \22167 , \22720 );
and \U$33895 ( \34210 , \22134 , \22707 );
nor \U$33896 ( \34211 , \34209 , \34210 );
xnor \U$33897 ( \34212 , \34211 , \22067 );
xor \U$33898 ( \34213 , \34208 , \34212 );
and \U$33899 ( \34214 , \22894 , \22598 );
and \U$33900 ( \34215 , \23230 , \22596 );
nor \U$33901 ( \34216 , \34214 , \34215 );
xnor \U$33902 ( \34217 , \34216 , \22608 );
and \U$33903 ( \34218 , \22081 , \22619 );
and \U$33904 ( \34219 , \22858 , \22617 );
nor \U$33905 ( \34220 , \34218 , \34219 );
xnor \U$33906 ( \34221 , \34220 , \22629 );
xor \U$33907 ( \34222 , \34217 , \34221 );
and \U$33908 ( \34223 , \22100 , \22641 );
and \U$33909 ( \34224 , \22071 , \22639 );
nor \U$33910 ( \34225 , \34223 , \34224 );
xnor \U$33911 ( \34226 , \34225 , \22651 );
xor \U$33912 ( \34227 , \34222 , \34226 );
xor \U$33913 ( \34228 , \34213 , \34227 );
and \U$33914 ( \34229 , \21990 , \22530 );
not \U$33915 ( \34230 , \34229 );
xnor \U$33916 ( \34231 , \34230 , \22540 );
and \U$33917 ( \34232 , \22001 , \22551 );
and \U$33918 ( \34233 , \21977 , \22549 );
nor \U$33919 ( \34234 , \34232 , \34233 );
xnor \U$33920 ( \34235 , \34234 , \22561 );
xor \U$33921 ( \34236 , \34231 , \34235 );
and \U$33922 ( \34237 , \23329 , \22573 );
and \U$33923 ( \34238 , \22030 , \22571 );
nor \U$33924 ( \34239 , \34237 , \34238 );
xnor \U$33925 ( \34240 , \34239 , \22583 );
xor \U$33926 ( \34241 , \34236 , \34240 );
xor \U$33927 ( \34242 , \34228 , \34241 );
and \U$33928 ( \34243 , \34111 , \34115 );
and \U$33929 ( \34244 , \34115 , \34120 );
and \U$33930 ( \34245 , \34111 , \34120 );
or \U$33931 ( \34246 , \34243 , \34244 , \34245 );
and \U$33932 ( \34247 , \22224 , \21978 );
not \U$33933 ( \34248 , \34247 );
xor \U$33934 ( \34249 , \34246 , \34248 );
and \U$33935 ( \34250 , \22192 , \23173 );
and \U$33936 ( \34251 , \22156 , \22999 );
nor \U$33937 ( \34252 , \34250 , \34251 );
xnor \U$33938 ( \34253 , \34252 , \22016 );
and \U$33939 ( \34254 , \22213 , \22021 );
and \U$33940 ( \34255 , \22181 , \22019 );
nor \U$33941 ( \34256 , \34254 , \34255 );
xnor \U$33942 ( \34257 , \34256 , \21595 );
xor \U$33943 ( \34258 , \34253 , \34257 );
and \U$33944 ( \34259 , \22235 , \21983 );
and \U$33945 ( \34260 , \22202 , \21981 );
nor \U$33946 ( \34261 , \34259 , \34260 );
xnor \U$33947 ( \34262 , \34261 , \21995 );
xor \U$33948 ( \34263 , \34258 , \34262 );
xor \U$33949 ( \34264 , \34249 , \34263 );
xor \U$33950 ( \34265 , \34242 , \34264 );
and \U$33951 ( \34266 , \34095 , \34099 );
and \U$33952 ( \34267 , \34099 , \34104 );
and \U$33953 ( \34268 , \34095 , \34104 );
or \U$33954 ( \34269 , \34266 , \34267 , \34268 );
and \U$33955 ( \34270 , \34084 , \34088 );
and \U$33956 ( \34271 , \34088 , \34093 );
and \U$33957 ( \34272 , \34084 , \34093 );
or \U$33958 ( \34273 , \34270 , \34271 , \34272 );
xor \U$33959 ( \34274 , \34269 , \34273 );
and \U$33960 ( \34275 , \34126 , \34130 );
and \U$33961 ( \34276 , \34130 , \34135 );
and \U$33962 ( \34277 , \34126 , \34135 );
or \U$33963 ( \34278 , \34275 , \34276 , \34277 );
xor \U$33964 ( \34279 , \34274 , \34278 );
xor \U$33965 ( \34280 , \34265 , \34279 );
xor \U$33966 ( \34281 , \34199 , \34280 );
xor \U$33967 ( \34282 , \34190 , \34281 );
and \U$33968 ( \34283 , \34159 , \34163 );
and \U$33969 ( \34284 , \34163 , \34175 );
and \U$33970 ( \34285 , \34159 , \34175 );
or \U$33971 ( \34286 , \34283 , \34284 , \34285 );
and \U$33972 ( \34287 , \34080 , \34138 );
and \U$33973 ( \34288 , \34138 , \34153 );
and \U$33974 ( \34289 , \34080 , \34153 );
or \U$33975 ( \34290 , \34287 , \34288 , \34289 );
xor \U$33976 ( \34291 , \34286 , \34290 );
and \U$33977 ( \34292 , \34070 , \34074 );
and \U$33978 ( \34293 , \34074 , \34079 );
and \U$33979 ( \34294 , \34070 , \34079 );
or \U$33980 ( \34295 , \34292 , \34293 , \34294 );
and \U$33981 ( \34296 , \34168 , \34169 );
and \U$33982 ( \34297 , \34169 , \34174 );
and \U$33983 ( \34298 , \34168 , \34174 );
or \U$33984 ( \34299 , \34296 , \34297 , \34298 );
xor \U$33985 ( \34300 , \34295 , \34299 );
and \U$33986 ( \34301 , \34107 , \34121 );
and \U$33987 ( \34302 , \34121 , \34136 );
and \U$33988 ( \34303 , \34107 , \34136 );
or \U$33989 ( \34304 , \34301 , \34302 , \34303 );
xor \U$33990 ( \34305 , \34300 , \34304 );
xor \U$33991 ( \34306 , \34291 , \34305 );
xor \U$33992 ( \34307 , \34282 , \34306 );
xor \U$33993 ( \34308 , \34186 , \34307 );
and \U$33994 ( \34309 , \34056 , \34178 );
nor \U$33995 ( \34310 , \34308 , \34309 );
and \U$33996 ( \34311 , \34190 , \34281 );
and \U$33997 ( \34312 , \34281 , \34306 );
and \U$33998 ( \34313 , \34190 , \34306 );
or \U$33999 ( \34314 , \34311 , \34312 , \34313 );
and \U$34000 ( \34315 , \34286 , \34290 );
and \U$34001 ( \34316 , \34290 , \34305 );
and \U$34002 ( \34317 , \34286 , \34305 );
or \U$34003 ( \34318 , \34315 , \34316 , \34317 );
xor \U$34004 ( \34319 , \34314 , \34318 );
and \U$34005 ( \34320 , \34194 , \34198 );
and \U$34006 ( \34321 , \34198 , \34280 );
and \U$34007 ( \34322 , \34194 , \34280 );
or \U$34008 ( \34323 , \34320 , \34321 , \34322 );
not \U$34009 ( \34324 , \22540 );
and \U$34010 ( \34325 , \21977 , \22551 );
and \U$34011 ( \34326 , \21990 , \22549 );
nor \U$34012 ( \34327 , \34325 , \34326 );
xnor \U$34013 ( \34328 , \34327 , \22561 );
xor \U$34014 ( \34329 , \34324 , \34328 );
and \U$34015 ( \34330 , \22030 , \22573 );
and \U$34016 ( \34331 , \22001 , \22571 );
nor \U$34017 ( \34332 , \34330 , \34331 );
xnor \U$34018 ( \34333 , \34332 , \22583 );
xor \U$34019 ( \34334 , \34329 , \34333 );
and \U$34020 ( \34335 , \22156 , \23173 );
and \U$34021 ( \34336 , \22167 , \22999 );
nor \U$34022 ( \34337 , \34335 , \34336 );
xnor \U$34023 ( \34338 , \34337 , \22016 );
and \U$34024 ( \34339 , \22181 , \22021 );
and \U$34025 ( \34340 , \22192 , \22019 );
nor \U$34026 ( \34341 , \34339 , \34340 );
xnor \U$34027 ( \34342 , \34341 , \21595 );
xor \U$34028 ( \34343 , \34338 , \34342 );
and \U$34029 ( \34344 , \22202 , \21983 );
and \U$34030 ( \34345 , \22213 , \21981 );
nor \U$34031 ( \34346 , \34344 , \34345 );
xnor \U$34032 ( \34347 , \34346 , \21995 );
xor \U$34033 ( \34348 , \34343 , \34347 );
and \U$34034 ( \34349 , \22089 , \22671 );
and \U$34035 ( \34350 , \22100 , \22669 );
nor \U$34036 ( \34351 , \34349 , \34350 );
xnor \U$34037 ( \34352 , \34351 , \22681 );
and \U$34038 ( \34353 , \22113 , \22691 );
and \U$34039 ( \34354 , \22124 , \22689 );
nor \U$34040 ( \34355 , \34353 , \34354 );
xnor \U$34041 ( \34356 , \34355 , \22701 );
xor \U$34042 ( \34357 , \34352 , \34356 );
and \U$34043 ( \34358 , \22134 , \22720 );
and \U$34044 ( \34359 , \22145 , \22707 );
nor \U$34045 ( \34360 , \34358 , \34359 );
xnor \U$34046 ( \34361 , \34360 , \22067 );
xor \U$34047 ( \34362 , \34357 , \34361 );
xor \U$34048 ( \34363 , \34348 , \34362 );
and \U$34049 ( \34364 , \23230 , \22598 );
and \U$34050 ( \34365 , \23329 , \22596 );
nor \U$34051 ( \34366 , \34364 , \34365 );
xnor \U$34052 ( \34367 , \34366 , \22608 );
and \U$34053 ( \34368 , \22858 , \22619 );
and \U$34054 ( \34369 , \22894 , \22617 );
nor \U$34055 ( \34370 , \34368 , \34369 );
xnor \U$34056 ( \34371 , \34370 , \22629 );
xor \U$34057 ( \34372 , \34367 , \34371 );
and \U$34058 ( \34373 , \22071 , \22641 );
and \U$34059 ( \34374 , \22081 , \22639 );
nor \U$34060 ( \34375 , \34373 , \34374 );
xnor \U$34061 ( \34376 , \34375 , \22651 );
xor \U$34062 ( \34377 , \34372 , \34376 );
xor \U$34063 ( \34378 , \34363 , \34377 );
xor \U$34064 ( \34379 , \34334 , \34378 );
and \U$34065 ( \34380 , \34253 , \34257 );
and \U$34066 ( \34381 , \34257 , \34262 );
and \U$34067 ( \34382 , \34253 , \34262 );
or \U$34068 ( \34383 , \34380 , \34381 , \34382 );
xor \U$34069 ( \34384 , \34383 , \34247 );
and \U$34070 ( \34385 , \22235 , \21978 );
xor \U$34071 ( \34386 , \34384 , \34385 );
xor \U$34072 ( \34387 , \34379 , \34386 );
and \U$34073 ( \34388 , \34269 , \34273 );
and \U$34074 ( \34389 , \34273 , \34278 );
and \U$34075 ( \34390 , \34269 , \34278 );
or \U$34076 ( \34391 , \34388 , \34389 , \34390 );
and \U$34077 ( \34392 , \34246 , \34248 );
and \U$34078 ( \34393 , \34248 , \34263 );
and \U$34079 ( \34394 , \34246 , \34263 );
or \U$34080 ( \34395 , \34392 , \34393 , \34394 );
xor \U$34081 ( \34396 , \34391 , \34395 );
and \U$34082 ( \34397 , \34213 , \34227 );
and \U$34083 ( \34398 , \34227 , \34241 );
and \U$34084 ( \34399 , \34213 , \34241 );
or \U$34085 ( \34400 , \34397 , \34398 , \34399 );
xor \U$34086 ( \34401 , \34396 , \34400 );
xor \U$34087 ( \34402 , \34387 , \34401 );
xor \U$34088 ( \34403 , \34323 , \34402 );
and \U$34089 ( \34404 , \34295 , \34299 );
and \U$34090 ( \34405 , \34299 , \34304 );
and \U$34091 ( \34406 , \34295 , \34304 );
or \U$34092 ( \34407 , \34404 , \34405 , \34406 );
and \U$34093 ( \34408 , \34242 , \34264 );
and \U$34094 ( \34409 , \34264 , \34279 );
and \U$34095 ( \34410 , \34242 , \34279 );
or \U$34096 ( \34411 , \34408 , \34409 , \34410 );
xor \U$34097 ( \34412 , \34407 , \34411 );
and \U$34098 ( \34413 , \34231 , \34235 );
and \U$34099 ( \34414 , \34235 , \34240 );
and \U$34100 ( \34415 , \34231 , \34240 );
or \U$34101 ( \34416 , \34413 , \34414 , \34415 );
and \U$34102 ( \34417 , \34217 , \34221 );
and \U$34103 ( \34418 , \34221 , \34226 );
and \U$34104 ( \34419 , \34217 , \34226 );
or \U$34105 ( \34420 , \34417 , \34418 , \34419 );
xor \U$34106 ( \34421 , \34416 , \34420 );
and \U$34107 ( \34422 , \34203 , \34207 );
and \U$34108 ( \34423 , \34207 , \34212 );
and \U$34109 ( \34424 , \34203 , \34212 );
or \U$34110 ( \34425 , \34422 , \34423 , \34424 );
xor \U$34111 ( \34426 , \34421 , \34425 );
xor \U$34112 ( \34427 , \34412 , \34426 );
xor \U$34113 ( \34428 , \34403 , \34427 );
xor \U$34114 ( \34429 , \34319 , \34428 );
and \U$34115 ( \34430 , \34186 , \34307 );
nor \U$34116 ( \34431 , \34429 , \34430 );
nor \U$34117 ( \34432 , \34310 , \34431 );
nand \U$34118 ( \34433 , \34182 , \34432 );
and \U$34119 ( \34434 , \34323 , \34402 );
and \U$34120 ( \34435 , \34402 , \34427 );
and \U$34121 ( \34436 , \34323 , \34427 );
or \U$34122 ( \34437 , \34434 , \34435 , \34436 );
and \U$34123 ( \34438 , \34391 , \34395 );
and \U$34124 ( \34439 , \34395 , \34400 );
and \U$34125 ( \34440 , \34391 , \34400 );
or \U$34126 ( \34441 , \34438 , \34439 , \34440 );
and \U$34127 ( \34442 , \34334 , \34378 );
and \U$34128 ( \34443 , \34378 , \34386 );
and \U$34129 ( \34444 , \34334 , \34386 );
or \U$34130 ( \34445 , \34442 , \34443 , \34444 );
xor \U$34131 ( \34446 , \34441 , \34445 );
and \U$34132 ( \34447 , \22124 , \22691 );
and \U$34133 ( \34448 , \22089 , \22689 );
nor \U$34134 ( \34449 , \34447 , \34448 );
xnor \U$34135 ( \34450 , \34449 , \22701 );
and \U$34136 ( \34451 , \22145 , \22720 );
and \U$34137 ( \34452 , \22113 , \22707 );
nor \U$34138 ( \34453 , \34451 , \34452 );
xnor \U$34139 ( \34454 , \34453 , \22067 );
xor \U$34140 ( \34455 , \34450 , \34454 );
and \U$34141 ( \34456 , \22167 , \23173 );
and \U$34142 ( \34457 , \22134 , \22999 );
nor \U$34143 ( \34458 , \34456 , \34457 );
xnor \U$34144 ( \34459 , \34458 , \22016 );
xor \U$34145 ( \34460 , \34455 , \34459 );
and \U$34146 ( \34461 , \22894 , \22619 );
and \U$34147 ( \34462 , \23230 , \22617 );
nor \U$34148 ( \34463 , \34461 , \34462 );
xnor \U$34149 ( \34464 , \34463 , \22629 );
and \U$34150 ( \34465 , \22081 , \22641 );
and \U$34151 ( \34466 , \22858 , \22639 );
nor \U$34152 ( \34467 , \34465 , \34466 );
xnor \U$34153 ( \34468 , \34467 , \22651 );
xor \U$34154 ( \34469 , \34464 , \34468 );
and \U$34155 ( \34470 , \22100 , \22671 );
and \U$34156 ( \34471 , \22071 , \22669 );
nor \U$34157 ( \34472 , \34470 , \34471 );
xnor \U$34158 ( \34473 , \34472 , \22681 );
xor \U$34159 ( \34474 , \34469 , \34473 );
xor \U$34160 ( \34475 , \34460 , \34474 );
and \U$34161 ( \34476 , \21990 , \22551 );
not \U$34162 ( \34477 , \34476 );
xnor \U$34163 ( \34478 , \34477 , \22561 );
and \U$34164 ( \34479 , \22001 , \22573 );
and \U$34165 ( \34480 , \21977 , \22571 );
nor \U$34166 ( \34481 , \34479 , \34480 );
xnor \U$34167 ( \34482 , \34481 , \22583 );
xor \U$34168 ( \34483 , \34478 , \34482 );
and \U$34169 ( \34484 , \23329 , \22598 );
and \U$34170 ( \34485 , \22030 , \22596 );
nor \U$34171 ( \34486 , \34484 , \34485 );
xnor \U$34172 ( \34487 , \34486 , \22608 );
xor \U$34173 ( \34488 , \34483 , \34487 );
xor \U$34174 ( \34489 , \34475 , \34488 );
and \U$34175 ( \34490 , \34338 , \34342 );
and \U$34176 ( \34491 , \34342 , \34347 );
and \U$34177 ( \34492 , \34338 , \34347 );
or \U$34178 ( \34493 , \34490 , \34491 , \34492 );
and \U$34179 ( \34494 , \22192 , \22021 );
and \U$34180 ( \34495 , \22156 , \22019 );
nor \U$34181 ( \34496 , \34494 , \34495 );
xnor \U$34182 ( \34497 , \34496 , \21595 );
and \U$34183 ( \34498 , \22213 , \21983 );
and \U$34184 ( \34499 , \22181 , \21981 );
nor \U$34185 ( \34500 , \34498 , \34499 );
xnor \U$34186 ( \34501 , \34500 , \21995 );
xor \U$34187 ( \34502 , \34497 , \34501 );
and \U$34188 ( \34503 , \22202 , \21978 );
xor \U$34189 ( \34504 , \34502 , \34503 );
xnor \U$34190 ( \34505 , \34493 , \34504 );
xor \U$34191 ( \34506 , \34489 , \34505 );
and \U$34192 ( \34507 , \34324 , \34328 );
and \U$34193 ( \34508 , \34328 , \34333 );
and \U$34194 ( \34509 , \34324 , \34333 );
or \U$34195 ( \34510 , \34507 , \34508 , \34509 );
and \U$34196 ( \34511 , \34367 , \34371 );
and \U$34197 ( \34512 , \34371 , \34376 );
and \U$34198 ( \34513 , \34367 , \34376 );
or \U$34199 ( \34514 , \34511 , \34512 , \34513 );
xor \U$34200 ( \34515 , \34510 , \34514 );
and \U$34201 ( \34516 , \34352 , \34356 );
and \U$34202 ( \34517 , \34356 , \34361 );
and \U$34203 ( \34518 , \34352 , \34361 );
or \U$34204 ( \34519 , \34516 , \34517 , \34518 );
xor \U$34205 ( \34520 , \34515 , \34519 );
xor \U$34206 ( \34521 , \34506 , \34520 );
xor \U$34207 ( \34522 , \34446 , \34521 );
xor \U$34208 ( \34523 , \34437 , \34522 );
and \U$34209 ( \34524 , \34407 , \34411 );
and \U$34210 ( \34525 , \34411 , \34426 );
and \U$34211 ( \34526 , \34407 , \34426 );
or \U$34212 ( \34527 , \34524 , \34525 , \34526 );
and \U$34213 ( \34528 , \34387 , \34401 );
xor \U$34214 ( \34529 , \34527 , \34528 );
and \U$34215 ( \34530 , \34416 , \34420 );
and \U$34216 ( \34531 , \34420 , \34425 );
and \U$34217 ( \34532 , \34416 , \34425 );
or \U$34218 ( \34533 , \34530 , \34531 , \34532 );
and \U$34219 ( \34534 , \34383 , \34247 );
and \U$34220 ( \34535 , \34247 , \34385 );
and \U$34221 ( \34536 , \34383 , \34385 );
or \U$34222 ( \34537 , \34534 , \34535 , \34536 );
xor \U$34223 ( \34538 , \34533 , \34537 );
and \U$34224 ( \34539 , \34348 , \34362 );
and \U$34225 ( \34540 , \34362 , \34377 );
and \U$34226 ( \34541 , \34348 , \34377 );
or \U$34227 ( \34542 , \34539 , \34540 , \34541 );
xor \U$34228 ( \34543 , \34538 , \34542 );
xor \U$34229 ( \34544 , \34529 , \34543 );
xor \U$34230 ( \34545 , \34523 , \34544 );
and \U$34231 ( \34546 , \34314 , \34318 );
and \U$34232 ( \34547 , \34318 , \34428 );
and \U$34233 ( \34548 , \34314 , \34428 );
or \U$34234 ( \34549 , \34546 , \34547 , \34548 );
nor \U$34235 ( \34550 , \34545 , \34549 );
and \U$34236 ( \34551 , \34527 , \34528 );
and \U$34237 ( \34552 , \34528 , \34543 );
and \U$34238 ( \34553 , \34527 , \34543 );
or \U$34239 ( \34554 , \34551 , \34552 , \34553 );
and \U$34240 ( \34555 , \34441 , \34445 );
and \U$34241 ( \34556 , \34445 , \34521 );
and \U$34242 ( \34557 , \34441 , \34521 );
or \U$34243 ( \34558 , \34555 , \34556 , \34557 );
and \U$34244 ( \34559 , \34510 , \34514 );
and \U$34245 ( \34560 , \34514 , \34519 );
and \U$34246 ( \34561 , \34510 , \34519 );
or \U$34247 ( \34562 , \34559 , \34560 , \34561 );
or \U$34248 ( \34563 , \34493 , \34504 );
xor \U$34249 ( \34564 , \34562 , \34563 );
and \U$34250 ( \34565 , \34460 , \34474 );
and \U$34251 ( \34566 , \34474 , \34488 );
and \U$34252 ( \34567 , \34460 , \34488 );
or \U$34253 ( \34568 , \34565 , \34566 , \34567 );
xor \U$34254 ( \34569 , \34564 , \34568 );
xor \U$34255 ( \34570 , \34558 , \34569 );
and \U$34256 ( \34571 , \34533 , \34537 );
and \U$34257 ( \34572 , \34537 , \34542 );
and \U$34258 ( \34573 , \34533 , \34542 );
or \U$34259 ( \34574 , \34571 , \34572 , \34573 );
and \U$34260 ( \34575 , \34489 , \34505 );
and \U$34261 ( \34576 , \34505 , \34520 );
and \U$34262 ( \34577 , \34489 , \34520 );
or \U$34263 ( \34578 , \34575 , \34576 , \34577 );
xor \U$34264 ( \34579 , \34574 , \34578 );
and \U$34265 ( \34580 , \23230 , \22619 );
and \U$34266 ( \34581 , \23329 , \22617 );
nor \U$34267 ( \34582 , \34580 , \34581 );
xnor \U$34268 ( \34583 , \34582 , \22629 );
and \U$34269 ( \34584 , \22858 , \22641 );
and \U$34270 ( \34585 , \22894 , \22639 );
nor \U$34271 ( \34586 , \34584 , \34585 );
xnor \U$34272 ( \34587 , \34586 , \22651 );
xor \U$34273 ( \34588 , \34583 , \34587 );
and \U$34274 ( \34589 , \22071 , \22671 );
and \U$34275 ( \34590 , \22081 , \22669 );
nor \U$34276 ( \34591 , \34589 , \34590 );
xnor \U$34277 ( \34592 , \34591 , \22681 );
xor \U$34278 ( \34593 , \34588 , \34592 );
not \U$34279 ( \34594 , \22561 );
and \U$34280 ( \34595 , \21977 , \22573 );
and \U$34281 ( \34596 , \21990 , \22571 );
nor \U$34282 ( \34597 , \34595 , \34596 );
xnor \U$34283 ( \34598 , \34597 , \22583 );
xor \U$34284 ( \34599 , \34594 , \34598 );
and \U$34285 ( \34600 , \22030 , \22598 );
and \U$34286 ( \34601 , \22001 , \22596 );
nor \U$34287 ( \34602 , \34600 , \34601 );
xnor \U$34288 ( \34603 , \34602 , \22608 );
xor \U$34289 ( \34604 , \34599 , \34603 );
xor \U$34290 ( \34605 , \34593 , \34604 );
and \U$34291 ( \34606 , \34497 , \34501 );
and \U$34292 ( \34607 , \34501 , \34503 );
and \U$34293 ( \34608 , \34497 , \34503 );
or \U$34294 ( \34609 , \34606 , \34607 , \34608 );
and \U$34295 ( \34610 , \22156 , \22021 );
and \U$34296 ( \34611 , \22167 , \22019 );
nor \U$34297 ( \34612 , \34610 , \34611 );
xnor \U$34298 ( \34613 , \34612 , \21595 );
and \U$34299 ( \34614 , \22181 , \21983 );
and \U$34300 ( \34615 , \22192 , \21981 );
nor \U$34301 ( \34616 , \34614 , \34615 );
xnor \U$34302 ( \34617 , \34616 , \21995 );
xor \U$34303 ( \34618 , \34613 , \34617 );
and \U$34304 ( \34619 , \22213 , \21978 );
xor \U$34305 ( \34620 , \34618 , \34619 );
xor \U$34306 ( \34621 , \34609 , \34620 );
and \U$34307 ( \34622 , \22089 , \22691 );
and \U$34308 ( \34623 , \22100 , \22689 );
nor \U$34309 ( \34624 , \34622 , \34623 );
xnor \U$34310 ( \34625 , \34624 , \22701 );
and \U$34311 ( \34626 , \22113 , \22720 );
and \U$34312 ( \34627 , \22124 , \22707 );
nor \U$34313 ( \34628 , \34626 , \34627 );
xnor \U$34314 ( \34629 , \34628 , \22067 );
xor \U$34315 ( \34630 , \34625 , \34629 );
and \U$34316 ( \34631 , \22134 , \23173 );
and \U$34317 ( \34632 , \22145 , \22999 );
nor \U$34318 ( \34633 , \34631 , \34632 );
xnor \U$34319 ( \34634 , \34633 , \22016 );
xor \U$34320 ( \34635 , \34630 , \34634 );
xor \U$34321 ( \34636 , \34621 , \34635 );
xor \U$34322 ( \34637 , \34605 , \34636 );
and \U$34323 ( \34638 , \34478 , \34482 );
and \U$34324 ( \34639 , \34482 , \34487 );
and \U$34325 ( \34640 , \34478 , \34487 );
or \U$34326 ( \34641 , \34638 , \34639 , \34640 );
and \U$34327 ( \34642 , \34464 , \34468 );
and \U$34328 ( \34643 , \34468 , \34473 );
and \U$34329 ( \34644 , \34464 , \34473 );
or \U$34330 ( \34645 , \34642 , \34643 , \34644 );
xor \U$34331 ( \34646 , \34641 , \34645 );
and \U$34332 ( \34647 , \34450 , \34454 );
and \U$34333 ( \34648 , \34454 , \34459 );
and \U$34334 ( \34649 , \34450 , \34459 );
or \U$34335 ( \34650 , \34647 , \34648 , \34649 );
xor \U$34336 ( \34651 , \34646 , \34650 );
xor \U$34337 ( \34652 , \34637 , \34651 );
xor \U$34338 ( \34653 , \34579 , \34652 );
xor \U$34339 ( \34654 , \34570 , \34653 );
xor \U$34340 ( \34655 , \34554 , \34654 );
and \U$34341 ( \34656 , \34437 , \34522 );
and \U$34342 ( \34657 , \34522 , \34544 );
and \U$34343 ( \34658 , \34437 , \34544 );
or \U$34344 ( \34659 , \34656 , \34657 , \34658 );
nor \U$34345 ( \34660 , \34655 , \34659 );
nor \U$34346 ( \34661 , \34550 , \34660 );
and \U$34347 ( \34662 , \34558 , \34569 );
and \U$34348 ( \34663 , \34569 , \34653 );
and \U$34349 ( \34664 , \34558 , \34653 );
or \U$34350 ( \34665 , \34662 , \34663 , \34664 );
and \U$34351 ( \34666 , \34574 , \34578 );
and \U$34352 ( \34667 , \34578 , \34652 );
and \U$34353 ( \34668 , \34574 , \34652 );
or \U$34354 ( \34669 , \34666 , \34667 , \34668 );
and \U$34355 ( \34670 , \34641 , \34645 );
and \U$34356 ( \34671 , \34645 , \34650 );
and \U$34357 ( \34672 , \34641 , \34650 );
or \U$34358 ( \34673 , \34670 , \34671 , \34672 );
and \U$34359 ( \34674 , \34609 , \34620 );
and \U$34360 ( \34675 , \34620 , \34635 );
and \U$34361 ( \34676 , \34609 , \34635 );
or \U$34362 ( \34677 , \34674 , \34675 , \34676 );
xor \U$34363 ( \34678 , \34673 , \34677 );
and \U$34364 ( \34679 , \34593 , \34604 );
xor \U$34365 ( \34680 , \34678 , \34679 );
xor \U$34366 ( \34681 , \34669 , \34680 );
and \U$34367 ( \34682 , \34562 , \34563 );
and \U$34368 ( \34683 , \34563 , \34568 );
and \U$34369 ( \34684 , \34562 , \34568 );
or \U$34370 ( \34685 , \34682 , \34683 , \34684 );
and \U$34371 ( \34686 , \34605 , \34636 );
and \U$34372 ( \34687 , \34636 , \34651 );
and \U$34373 ( \34688 , \34605 , \34651 );
or \U$34374 ( \34689 , \34686 , \34687 , \34688 );
xor \U$34375 ( \34690 , \34685 , \34689 );
and \U$34376 ( \34691 , \22894 , \22641 );
and \U$34377 ( \34692 , \23230 , \22639 );
nor \U$34378 ( \34693 , \34691 , \34692 );
xnor \U$34379 ( \34694 , \34693 , \22651 );
and \U$34380 ( \34695 , \22081 , \22671 );
and \U$34381 ( \34696 , \22858 , \22669 );
nor \U$34382 ( \34697 , \34695 , \34696 );
xnor \U$34383 ( \34698 , \34697 , \22681 );
xor \U$34384 ( \34699 , \34694 , \34698 );
and \U$34385 ( \34700 , \22100 , \22691 );
and \U$34386 ( \34701 , \22071 , \22689 );
nor \U$34387 ( \34702 , \34700 , \34701 );
xnor \U$34388 ( \34703 , \34702 , \22701 );
xor \U$34389 ( \34704 , \34699 , \34703 );
and \U$34390 ( \34705 , \21990 , \22573 );
not \U$34391 ( \34706 , \34705 );
xnor \U$34392 ( \34707 , \34706 , \22583 );
and \U$34393 ( \34708 , \22001 , \22598 );
and \U$34394 ( \34709 , \21977 , \22596 );
nor \U$34395 ( \34710 , \34708 , \34709 );
xnor \U$34396 ( \34711 , \34710 , \22608 );
xor \U$34397 ( \34712 , \34707 , \34711 );
and \U$34398 ( \34713 , \23329 , \22619 );
and \U$34399 ( \34714 , \22030 , \22617 );
nor \U$34400 ( \34715 , \34713 , \34714 );
xnor \U$34401 ( \34716 , \34715 , \22629 );
xor \U$34402 ( \34717 , \34712 , \34716 );
xor \U$34403 ( \34718 , \34704 , \34717 );
and \U$34404 ( \34719 , \34613 , \34617 );
and \U$34405 ( \34720 , \34617 , \34619 );
and \U$34406 ( \34721 , \34613 , \34619 );
or \U$34407 ( \34722 , \34719 , \34720 , \34721 );
and \U$34408 ( \34723 , \22192 , \21983 );
and \U$34409 ( \34724 , \22156 , \21981 );
nor \U$34410 ( \34725 , \34723 , \34724 );
xnor \U$34411 ( \34726 , \34725 , \21995 );
and \U$34412 ( \34727 , \22181 , \21978 );
xnor \U$34413 ( \34728 , \34726 , \34727 );
xor \U$34414 ( \34729 , \34722 , \34728 );
and \U$34415 ( \34730 , \22124 , \22720 );
and \U$34416 ( \34731 , \22089 , \22707 );
nor \U$34417 ( \34732 , \34730 , \34731 );
xnor \U$34418 ( \34733 , \34732 , \22067 );
and \U$34419 ( \34734 , \22145 , \23173 );
and \U$34420 ( \34735 , \22113 , \22999 );
nor \U$34421 ( \34736 , \34734 , \34735 );
xnor \U$34422 ( \34737 , \34736 , \22016 );
xor \U$34423 ( \34738 , \34733 , \34737 );
and \U$34424 ( \34739 , \22167 , \22021 );
and \U$34425 ( \34740 , \22134 , \22019 );
nor \U$34426 ( \34741 , \34739 , \34740 );
xnor \U$34427 ( \34742 , \34741 , \21595 );
xor \U$34428 ( \34743 , \34738 , \34742 );
xor \U$34429 ( \34744 , \34729 , \34743 );
xor \U$34430 ( \34745 , \34718 , \34744 );
and \U$34431 ( \34746 , \34594 , \34598 );
and \U$34432 ( \34747 , \34598 , \34603 );
and \U$34433 ( \34748 , \34594 , \34603 );
or \U$34434 ( \34749 , \34746 , \34747 , \34748 );
and \U$34435 ( \34750 , \34583 , \34587 );
and \U$34436 ( \34751 , \34587 , \34592 );
and \U$34437 ( \34752 , \34583 , \34592 );
or \U$34438 ( \34753 , \34750 , \34751 , \34752 );
xor \U$34439 ( \34754 , \34749 , \34753 );
and \U$34440 ( \34755 , \34625 , \34629 );
and \U$34441 ( \34756 , \34629 , \34634 );
and \U$34442 ( \34757 , \34625 , \34634 );
or \U$34443 ( \34758 , \34755 , \34756 , \34757 );
xor \U$34444 ( \34759 , \34754 , \34758 );
xor \U$34445 ( \34760 , \34745 , \34759 );
xor \U$34446 ( \34761 , \34690 , \34760 );
xor \U$34447 ( \34762 , \34681 , \34761 );
xor \U$34448 ( \34763 , \34665 , \34762 );
and \U$34449 ( \34764 , \34554 , \34654 );
nor \U$34450 ( \34765 , \34763 , \34764 );
and \U$34451 ( \34766 , \34669 , \34680 );
and \U$34452 ( \34767 , \34680 , \34761 );
and \U$34453 ( \34768 , \34669 , \34761 );
or \U$34454 ( \34769 , \34766 , \34767 , \34768 );
and \U$34455 ( \34770 , \34685 , \34689 );
and \U$34456 ( \34771 , \34689 , \34760 );
and \U$34457 ( \34772 , \34685 , \34760 );
or \U$34458 ( \34773 , \34770 , \34771 , \34772 );
and \U$34459 ( \34774 , \34749 , \34753 );
and \U$34460 ( \34775 , \34753 , \34758 );
and \U$34461 ( \34776 , \34749 , \34758 );
or \U$34462 ( \34777 , \34774 , \34775 , \34776 );
and \U$34463 ( \34778 , \34722 , \34728 );
and \U$34464 ( \34779 , \34728 , \34743 );
and \U$34465 ( \34780 , \34722 , \34743 );
or \U$34466 ( \34781 , \34778 , \34779 , \34780 );
xor \U$34467 ( \34782 , \34777 , \34781 );
and \U$34468 ( \34783 , \34704 , \34717 );
xor \U$34469 ( \34784 , \34782 , \34783 );
xor \U$34470 ( \34785 , \34773 , \34784 );
and \U$34471 ( \34786 , \34673 , \34677 );
and \U$34472 ( \34787 , \34677 , \34679 );
and \U$34473 ( \34788 , \34673 , \34679 );
or \U$34474 ( \34789 , \34786 , \34787 , \34788 );
and \U$34475 ( \34790 , \34718 , \34744 );
and \U$34476 ( \34791 , \34744 , \34759 );
and \U$34477 ( \34792 , \34718 , \34759 );
or \U$34478 ( \34793 , \34790 , \34791 , \34792 );
xor \U$34479 ( \34794 , \34789 , \34793 );
and \U$34480 ( \34795 , \22089 , \22720 );
and \U$34481 ( \34796 , \22100 , \22707 );
nor \U$34482 ( \34797 , \34795 , \34796 );
xnor \U$34483 ( \34798 , \34797 , \22067 );
and \U$34484 ( \34799 , \22113 , \23173 );
and \U$34485 ( \34800 , \22124 , \22999 );
nor \U$34486 ( \34801 , \34799 , \34800 );
xnor \U$34487 ( \34802 , \34801 , \22016 );
xor \U$34488 ( \34803 , \34798 , \34802 );
and \U$34489 ( \34804 , \22134 , \22021 );
and \U$34490 ( \34805 , \22145 , \22019 );
nor \U$34491 ( \34806 , \34804 , \34805 );
xnor \U$34492 ( \34807 , \34806 , \21595 );
xor \U$34493 ( \34808 , \34803 , \34807 );
and \U$34494 ( \34809 , \23230 , \22641 );
and \U$34495 ( \34810 , \23329 , \22639 );
nor \U$34496 ( \34811 , \34809 , \34810 );
xnor \U$34497 ( \34812 , \34811 , \22651 );
and \U$34498 ( \34813 , \22858 , \22671 );
and \U$34499 ( \34814 , \22894 , \22669 );
nor \U$34500 ( \34815 , \34813 , \34814 );
xnor \U$34501 ( \34816 , \34815 , \22681 );
xor \U$34502 ( \34817 , \34812 , \34816 );
and \U$34503 ( \34818 , \22071 , \22691 );
and \U$34504 ( \34819 , \22081 , \22689 );
nor \U$34505 ( \34820 , \34818 , \34819 );
xnor \U$34506 ( \34821 , \34820 , \22701 );
xor \U$34507 ( \34822 , \34817 , \34821 );
xor \U$34508 ( \34823 , \34808 , \34822 );
not \U$34509 ( \34824 , \22583 );
and \U$34510 ( \34825 , \21977 , \22598 );
and \U$34511 ( \34826 , \21990 , \22596 );
nor \U$34512 ( \34827 , \34825 , \34826 );
xnor \U$34513 ( \34828 , \34827 , \22608 );
xor \U$34514 ( \34829 , \34824 , \34828 );
and \U$34515 ( \34830 , \22030 , \22619 );
and \U$34516 ( \34831 , \22001 , \22617 );
nor \U$34517 ( \34832 , \34830 , \34831 );
xnor \U$34518 ( \34833 , \34832 , \22629 );
xor \U$34519 ( \34834 , \34829 , \34833 );
xor \U$34520 ( \34835 , \34823 , \34834 );
or \U$34521 ( \34836 , \34726 , \34727 );
and \U$34522 ( \34837 , \22156 , \21983 );
and \U$34523 ( \34838 , \22167 , \21981 );
nor \U$34524 ( \34839 , \34837 , \34838 );
xnor \U$34525 ( \34840 , \34839 , \21995 );
xor \U$34526 ( \34841 , \34836 , \34840 );
and \U$34527 ( \34842 , \22192 , \21978 );
xor \U$34528 ( \34843 , \34841 , \34842 );
xor \U$34529 ( \34844 , \34835 , \34843 );
and \U$34530 ( \34845 , \34707 , \34711 );
and \U$34531 ( \34846 , \34711 , \34716 );
and \U$34532 ( \34847 , \34707 , \34716 );
or \U$34533 ( \34848 , \34845 , \34846 , \34847 );
and \U$34534 ( \34849 , \34694 , \34698 );
and \U$34535 ( \34850 , \34698 , \34703 );
and \U$34536 ( \34851 , \34694 , \34703 );
or \U$34537 ( \34852 , \34849 , \34850 , \34851 );
xor \U$34538 ( \34853 , \34848 , \34852 );
and \U$34539 ( \34854 , \34733 , \34737 );
and \U$34540 ( \34855 , \34737 , \34742 );
and \U$34541 ( \34856 , \34733 , \34742 );
or \U$34542 ( \34857 , \34854 , \34855 , \34856 );
xor \U$34543 ( \34858 , \34853 , \34857 );
xor \U$34544 ( \34859 , \34844 , \34858 );
xor \U$34545 ( \34860 , \34794 , \34859 );
xor \U$34546 ( \34861 , \34785 , \34860 );
xor \U$34547 ( \34862 , \34769 , \34861 );
and \U$34548 ( \34863 , \34665 , \34762 );
nor \U$34549 ( \34864 , \34862 , \34863 );
nor \U$34550 ( \34865 , \34765 , \34864 );
nand \U$34551 ( \34866 , \34661 , \34865 );
nor \U$34552 ( \34867 , \34433 , \34866 );
nand \U$34553 ( \34868 , \33915 , \34867 );
and \U$34554 ( \34869 , \34773 , \34784 );
and \U$34555 ( \34870 , \34784 , \34860 );
and \U$34556 ( \34871 , \34773 , \34860 );
or \U$34557 ( \34872 , \34869 , \34870 , \34871 );
and \U$34558 ( \34873 , \34789 , \34793 );
and \U$34559 ( \34874 , \34793 , \34859 );
and \U$34560 ( \34875 , \34789 , \34859 );
or \U$34561 ( \34876 , \34873 , \34874 , \34875 );
and \U$34562 ( \34877 , \34848 , \34852 );
and \U$34563 ( \34878 , \34852 , \34857 );
and \U$34564 ( \34879 , \34848 , \34857 );
or \U$34565 ( \34880 , \34877 , \34878 , \34879 );
and \U$34566 ( \34881 , \34836 , \34840 );
and \U$34567 ( \34882 , \34840 , \34842 );
and \U$34568 ( \34883 , \34836 , \34842 );
or \U$34569 ( \34884 , \34881 , \34882 , \34883 );
xor \U$34570 ( \34885 , \34880 , \34884 );
and \U$34571 ( \34886 , \34808 , \34822 );
and \U$34572 ( \34887 , \34822 , \34834 );
and \U$34573 ( \34888 , \34808 , \34834 );
or \U$34574 ( \34889 , \34886 , \34887 , \34888 );
xor \U$34575 ( \34890 , \34885 , \34889 );
xor \U$34576 ( \34891 , \34876 , \34890 );
and \U$34577 ( \34892 , \34777 , \34781 );
and \U$34578 ( \34893 , \34781 , \34783 );
and \U$34579 ( \34894 , \34777 , \34783 );
or \U$34580 ( \34895 , \34892 , \34893 , \34894 );
and \U$34581 ( \34896 , \34835 , \34843 );
and \U$34582 ( \34897 , \34843 , \34858 );
and \U$34583 ( \34898 , \34835 , \34858 );
or \U$34584 ( \34899 , \34896 , \34897 , \34898 );
xor \U$34585 ( \34900 , \34895 , \34899 );
and \U$34586 ( \34901 , \22894 , \22671 );
and \U$34587 ( \34902 , \23230 , \22669 );
nor \U$34588 ( \34903 , \34901 , \34902 );
xnor \U$34589 ( \34904 , \34903 , \22681 );
and \U$34590 ( \34905 , \22081 , \22691 );
and \U$34591 ( \34906 , \22858 , \22689 );
nor \U$34592 ( \34907 , \34905 , \34906 );
xnor \U$34593 ( \34908 , \34907 , \22701 );
xor \U$34594 ( \34909 , \34904 , \34908 );
and \U$34595 ( \34910 , \22100 , \22720 );
and \U$34596 ( \34911 , \22071 , \22707 );
nor \U$34597 ( \34912 , \34910 , \34911 );
xnor \U$34598 ( \34913 , \34912 , \22067 );
xor \U$34599 ( \34914 , \34909 , \34913 );
and \U$34600 ( \34915 , \21990 , \22598 );
not \U$34601 ( \34916 , \34915 );
xnor \U$34602 ( \34917 , \34916 , \22608 );
and \U$34603 ( \34918 , \22001 , \22619 );
and \U$34604 ( \34919 , \21977 , \22617 );
nor \U$34605 ( \34920 , \34918 , \34919 );
xnor \U$34606 ( \34921 , \34920 , \22629 );
xor \U$34607 ( \34922 , \34917 , \34921 );
and \U$34608 ( \34923 , \23329 , \22641 );
and \U$34609 ( \34924 , \22030 , \22639 );
nor \U$34610 ( \34925 , \34923 , \34924 );
xnor \U$34611 ( \34926 , \34925 , \22651 );
xor \U$34612 ( \34927 , \34922 , \34926 );
xor \U$34613 ( \34928 , \34914 , \34927 );
and \U$34614 ( \34929 , \22156 , \21978 );
and \U$34615 ( \34930 , \22124 , \23173 );
and \U$34616 ( \34931 , \22089 , \22999 );
nor \U$34617 ( \34932 , \34930 , \34931 );
xnor \U$34618 ( \34933 , \34932 , \22016 );
and \U$34619 ( \34934 , \22145 , \22021 );
and \U$34620 ( \34935 , \22113 , \22019 );
nor \U$34621 ( \34936 , \34934 , \34935 );
xnor \U$34622 ( \34937 , \34936 , \21595 );
xor \U$34623 ( \34938 , \34933 , \34937 );
and \U$34624 ( \34939 , \22167 , \21983 );
and \U$34625 ( \34940 , \22134 , \21981 );
nor \U$34626 ( \34941 , \34939 , \34940 );
xnor \U$34627 ( \34942 , \34941 , \21995 );
xor \U$34628 ( \34943 , \34938 , \34942 );
xnor \U$34629 ( \34944 , \34929 , \34943 );
xor \U$34630 ( \34945 , \34928 , \34944 );
and \U$34631 ( \34946 , \34824 , \34828 );
and \U$34632 ( \34947 , \34828 , \34833 );
and \U$34633 ( \34948 , \34824 , \34833 );
or \U$34634 ( \34949 , \34946 , \34947 , \34948 );
and \U$34635 ( \34950 , \34812 , \34816 );
and \U$34636 ( \34951 , \34816 , \34821 );
and \U$34637 ( \34952 , \34812 , \34821 );
or \U$34638 ( \34953 , \34950 , \34951 , \34952 );
xor \U$34639 ( \34954 , \34949 , \34953 );
and \U$34640 ( \34955 , \34798 , \34802 );
and \U$34641 ( \34956 , \34802 , \34807 );
and \U$34642 ( \34957 , \34798 , \34807 );
or \U$34643 ( \34958 , \34955 , \34956 , \34957 );
xor \U$34644 ( \34959 , \34954 , \34958 );
xor \U$34645 ( \34960 , \34945 , \34959 );
xor \U$34646 ( \34961 , \34900 , \34960 );
xor \U$34647 ( \34962 , \34891 , \34961 );
xor \U$34648 ( \34963 , \34872 , \34962 );
and \U$34649 ( \34964 , \34769 , \34861 );
nor \U$34650 ( \34965 , \34963 , \34964 );
and \U$34651 ( \34966 , \34876 , \34890 );
and \U$34652 ( \34967 , \34890 , \34961 );
and \U$34653 ( \34968 , \34876 , \34961 );
or \U$34654 ( \34969 , \34966 , \34967 , \34968 );
and \U$34655 ( \34970 , \34895 , \34899 );
and \U$34656 ( \34971 , \34899 , \34960 );
and \U$34657 ( \34972 , \34895 , \34960 );
or \U$34658 ( \34973 , \34970 , \34971 , \34972 );
and \U$34659 ( \34974 , \34949 , \34953 );
and \U$34660 ( \34975 , \34953 , \34958 );
and \U$34661 ( \34976 , \34949 , \34958 );
or \U$34662 ( \34977 , \34974 , \34975 , \34976 );
or \U$34663 ( \34978 , \34929 , \34943 );
xor \U$34664 ( \34979 , \34977 , \34978 );
and \U$34665 ( \34980 , \34914 , \34927 );
xor \U$34666 ( \34981 , \34979 , \34980 );
xor \U$34667 ( \34982 , \34973 , \34981 );
and \U$34668 ( \34983 , \34880 , \34884 );
and \U$34669 ( \34984 , \34884 , \34889 );
and \U$34670 ( \34985 , \34880 , \34889 );
or \U$34671 ( \34986 , \34983 , \34984 , \34985 );
and \U$34672 ( \34987 , \34928 , \34944 );
and \U$34673 ( \34988 , \34944 , \34959 );
and \U$34674 ( \34989 , \34928 , \34959 );
or \U$34675 ( \34990 , \34987 , \34988 , \34989 );
xor \U$34676 ( \34991 , \34986 , \34990 );
not \U$34677 ( \34992 , \22608 );
and \U$34678 ( \34993 , \21977 , \22619 );
and \U$34679 ( \34994 , \21990 , \22617 );
nor \U$34680 ( \34995 , \34993 , \34994 );
xnor \U$34681 ( \34996 , \34995 , \22629 );
xor \U$34682 ( \34997 , \34992 , \34996 );
and \U$34683 ( \34998 , \22030 , \22641 );
and \U$34684 ( \34999 , \22001 , \22639 );
nor \U$34685 ( \35000 , \34998 , \34999 );
xnor \U$34686 ( \35001 , \35000 , \22651 );
xor \U$34687 ( \35002 , \34997 , \35001 );
and \U$34688 ( \35003 , \22167 , \21978 );
and \U$34689 ( \35004 , \22089 , \23173 );
and \U$34690 ( \35005 , \22100 , \22999 );
nor \U$34691 ( \35006 , \35004 , \35005 );
xnor \U$34692 ( \35007 , \35006 , \22016 );
and \U$34693 ( \35008 , \22113 , \22021 );
and \U$34694 ( \35009 , \22124 , \22019 );
nor \U$34695 ( \35010 , \35008 , \35009 );
xnor \U$34696 ( \35011 , \35010 , \21595 );
xor \U$34697 ( \35012 , \35007 , \35011 );
and \U$34698 ( \35013 , \22134 , \21983 );
and \U$34699 ( \35014 , \22145 , \21981 );
nor \U$34700 ( \35015 , \35013 , \35014 );
xnor \U$34701 ( \35016 , \35015 , \21995 );
xor \U$34702 ( \35017 , \35012 , \35016 );
xor \U$34703 ( \35018 , \35003 , \35017 );
and \U$34704 ( \35019 , \23230 , \22671 );
and \U$34705 ( \35020 , \23329 , \22669 );
nor \U$34706 ( \35021 , \35019 , \35020 );
xnor \U$34707 ( \35022 , \35021 , \22681 );
and \U$34708 ( \35023 , \22858 , \22691 );
and \U$34709 ( \35024 , \22894 , \22689 );
nor \U$34710 ( \35025 , \35023 , \35024 );
xnor \U$34711 ( \35026 , \35025 , \22701 );
xor \U$34712 ( \35027 , \35022 , \35026 );
and \U$34713 ( \35028 , \22071 , \22720 );
and \U$34714 ( \35029 , \22081 , \22707 );
nor \U$34715 ( \35030 , \35028 , \35029 );
xnor \U$34716 ( \35031 , \35030 , \22067 );
xor \U$34717 ( \35032 , \35027 , \35031 );
xor \U$34718 ( \35033 , \35018 , \35032 );
xor \U$34719 ( \35034 , \35002 , \35033 );
and \U$34720 ( \35035 , \34917 , \34921 );
and \U$34721 ( \35036 , \34921 , \34926 );
and \U$34722 ( \35037 , \34917 , \34926 );
or \U$34723 ( \35038 , \35035 , \35036 , \35037 );
and \U$34724 ( \35039 , \34904 , \34908 );
and \U$34725 ( \35040 , \34908 , \34913 );
and \U$34726 ( \35041 , \34904 , \34913 );
or \U$34727 ( \35042 , \35039 , \35040 , \35041 );
xor \U$34728 ( \35043 , \35038 , \35042 );
and \U$34729 ( \35044 , \34933 , \34937 );
and \U$34730 ( \35045 , \34937 , \34942 );
and \U$34731 ( \35046 , \34933 , \34942 );
or \U$34732 ( \35047 , \35044 , \35045 , \35046 );
xor \U$34733 ( \35048 , \35043 , \35047 );
xor \U$34734 ( \35049 , \35034 , \35048 );
xor \U$34735 ( \35050 , \34991 , \35049 );
xor \U$34736 ( \35051 , \34982 , \35050 );
xor \U$34737 ( \35052 , \34969 , \35051 );
and \U$34738 ( \35053 , \34872 , \34962 );
nor \U$34739 ( \35054 , \35052 , \35053 );
nor \U$34740 ( \35055 , \34965 , \35054 );
and \U$34741 ( \35056 , \34973 , \34981 );
and \U$34742 ( \35057 , \34981 , \35050 );
and \U$34743 ( \35058 , \34973 , \35050 );
or \U$34744 ( \35059 , \35056 , \35057 , \35058 );
and \U$34745 ( \35060 , \34986 , \34990 );
and \U$34746 ( \35061 , \34990 , \35049 );
and \U$34747 ( \35062 , \34986 , \35049 );
or \U$34748 ( \35063 , \35060 , \35061 , \35062 );
and \U$34749 ( \35064 , \34992 , \34996 );
and \U$34750 ( \35065 , \34996 , \35001 );
and \U$34751 ( \35066 , \34992 , \35001 );
or \U$34752 ( \35067 , \35064 , \35065 , \35066 );
and \U$34753 ( \35068 , \35022 , \35026 );
and \U$34754 ( \35069 , \35026 , \35031 );
and \U$34755 ( \35070 , \35022 , \35031 );
or \U$34756 ( \35071 , \35068 , \35069 , \35070 );
xor \U$34757 ( \35072 , \35067 , \35071 );
and \U$34758 ( \35073 , \35007 , \35011 );
and \U$34759 ( \35074 , \35011 , \35016 );
and \U$34760 ( \35075 , \35007 , \35016 );
or \U$34761 ( \35076 , \35073 , \35074 , \35075 );
xor \U$34762 ( \35077 , \35072 , \35076 );
and \U$34763 ( \35078 , \35038 , \35042 );
and \U$34764 ( \35079 , \35042 , \35047 );
and \U$34765 ( \35080 , \35038 , \35047 );
or \U$34766 ( \35081 , \35078 , \35079 , \35080 );
and \U$34767 ( \35082 , \35003 , \35017 );
and \U$34768 ( \35083 , \35017 , \35032 );
and \U$34769 ( \35084 , \35003 , \35032 );
or \U$34770 ( \35085 , \35082 , \35083 , \35084 );
xor \U$34771 ( \35086 , \35081 , \35085 );
and \U$34772 ( \35087 , \21990 , \22619 );
not \U$34773 ( \35088 , \35087 );
xnor \U$34774 ( \35089 , \35088 , \22629 );
and \U$34775 ( \35090 , \22001 , \22641 );
and \U$34776 ( \35091 , \21977 , \22639 );
nor \U$34777 ( \35092 , \35090 , \35091 );
xnor \U$34778 ( \35093 , \35092 , \22651 );
xor \U$34779 ( \35094 , \35089 , \35093 );
and \U$34780 ( \35095 , \23329 , \22671 );
and \U$34781 ( \35096 , \22030 , \22669 );
nor \U$34782 ( \35097 , \35095 , \35096 );
xnor \U$34783 ( \35098 , \35097 , \22681 );
xor \U$34784 ( \35099 , \35094 , \35098 );
xor \U$34785 ( \35100 , \35086 , \35099 );
xor \U$34786 ( \35101 , \35077 , \35100 );
xor \U$34787 ( \35102 , \35063 , \35101 );
and \U$34788 ( \35103 , \34977 , \34978 );
and \U$34789 ( \35104 , \34978 , \34980 );
and \U$34790 ( \35105 , \34977 , \34980 );
or \U$34791 ( \35106 , \35103 , \35104 , \35105 );
and \U$34792 ( \35107 , \35002 , \35033 );
and \U$34793 ( \35108 , \35033 , \35048 );
and \U$34794 ( \35109 , \35002 , \35048 );
or \U$34795 ( \35110 , \35107 , \35108 , \35109 );
xor \U$34796 ( \35111 , \35106 , \35110 );
and \U$34797 ( \35112 , \22124 , \22021 );
and \U$34798 ( \35113 , \22089 , \22019 );
nor \U$34799 ( \35114 , \35112 , \35113 );
xnor \U$34800 ( \35115 , \35114 , \21595 );
and \U$34801 ( \35116 , \22145 , \21983 );
and \U$34802 ( \35117 , \22113 , \21981 );
nor \U$34803 ( \35118 , \35116 , \35117 );
xnor \U$34804 ( \35119 , \35118 , \21995 );
xor \U$34805 ( \35120 , \35115 , \35119 );
and \U$34806 ( \35121 , \22134 , \21978 );
xor \U$34807 ( \35122 , \35120 , \35121 );
and \U$34808 ( \35123 , \22894 , \22691 );
and \U$34809 ( \35124 , \23230 , \22689 );
nor \U$34810 ( \35125 , \35123 , \35124 );
xnor \U$34811 ( \35126 , \35125 , \22701 );
and \U$34812 ( \35127 , \22081 , \22720 );
and \U$34813 ( \35128 , \22858 , \22707 );
nor \U$34814 ( \35129 , \35127 , \35128 );
xnor \U$34815 ( \35130 , \35129 , \22067 );
xor \U$34816 ( \35131 , \35126 , \35130 );
and \U$34817 ( \35132 , \22100 , \23173 );
and \U$34818 ( \35133 , \22071 , \22999 );
nor \U$34819 ( \35134 , \35132 , \35133 );
xnor \U$34820 ( \35135 , \35134 , \22016 );
xor \U$34821 ( \35136 , \35131 , \35135 );
xnor \U$34822 ( \35137 , \35122 , \35136 );
xor \U$34823 ( \35138 , \35111 , \35137 );
xor \U$34824 ( \35139 , \35102 , \35138 );
xor \U$34825 ( \35140 , \35059 , \35139 );
and \U$34826 ( \35141 , \34969 , \35051 );
nor \U$34827 ( \35142 , \35140 , \35141 );
and \U$34828 ( \35143 , \35063 , \35101 );
and \U$34829 ( \35144 , \35101 , \35138 );
and \U$34830 ( \35145 , \35063 , \35138 );
or \U$34831 ( \35146 , \35143 , \35144 , \35145 );
and \U$34832 ( \35147 , \35106 , \35110 );
and \U$34833 ( \35148 , \35110 , \35137 );
and \U$34834 ( \35149 , \35106 , \35137 );
or \U$34835 ( \35150 , \35147 , \35148 , \35149 );
and \U$34836 ( \35151 , \35077 , \35100 );
xor \U$34837 ( \35152 , \35150 , \35151 );
and \U$34838 ( \35153 , \35081 , \35085 );
and \U$34839 ( \35154 , \35085 , \35099 );
and \U$34840 ( \35155 , \35081 , \35099 );
or \U$34841 ( \35156 , \35153 , \35154 , \35155 );
and \U$34842 ( \35157 , \35089 , \35093 );
and \U$34843 ( \35158 , \35093 , \35098 );
and \U$34844 ( \35159 , \35089 , \35098 );
or \U$34845 ( \35160 , \35157 , \35158 , \35159 );
and \U$34846 ( \35161 , \35126 , \35130 );
and \U$34847 ( \35162 , \35130 , \35135 );
and \U$34848 ( \35163 , \35126 , \35135 );
or \U$34849 ( \35164 , \35161 , \35162 , \35163 );
xor \U$34850 ( \35165 , \35160 , \35164 );
and \U$34851 ( \35166 , \35115 , \35119 );
and \U$34852 ( \35167 , \35119 , \35121 );
and \U$34853 ( \35168 , \35115 , \35121 );
or \U$34854 ( \35169 , \35166 , \35167 , \35168 );
xor \U$34855 ( \35170 , \35165 , \35169 );
xor \U$34856 ( \35171 , \35156 , \35170 );
and \U$34857 ( \35172 , \35067 , \35071 );
and \U$34858 ( \35173 , \35071 , \35076 );
and \U$34859 ( \35174 , \35067 , \35076 );
or \U$34860 ( \35175 , \35172 , \35173 , \35174 );
or \U$34861 ( \35176 , \35122 , \35136 );
xor \U$34862 ( \35177 , \35175 , \35176 );
and \U$34863 ( \35178 , \22089 , \22021 );
and \U$34864 ( \35179 , \22100 , \22019 );
nor \U$34865 ( \35180 , \35178 , \35179 );
xnor \U$34866 ( \35181 , \35180 , \21595 );
and \U$34867 ( \35182 , \22113 , \21983 );
and \U$34868 ( \35183 , \22124 , \21981 );
nor \U$34869 ( \35184 , \35182 , \35183 );
xnor \U$34870 ( \35185 , \35184 , \21995 );
xor \U$34871 ( \35186 , \35181 , \35185 );
and \U$34872 ( \35187 , \22145 , \21978 );
xor \U$34873 ( \35188 , \35186 , \35187 );
and \U$34874 ( \35189 , \23230 , \22691 );
and \U$34875 ( \35190 , \23329 , \22689 );
nor \U$34876 ( \35191 , \35189 , \35190 );
xnor \U$34877 ( \35192 , \35191 , \22701 );
and \U$34878 ( \35193 , \22858 , \22720 );
and \U$34879 ( \35194 , \22894 , \22707 );
nor \U$34880 ( \35195 , \35193 , \35194 );
xnor \U$34881 ( \35196 , \35195 , \22067 );
xor \U$34882 ( \35197 , \35192 , \35196 );
and \U$34883 ( \35198 , \22071 , \23173 );
and \U$34884 ( \35199 , \22081 , \22999 );
nor \U$34885 ( \35200 , \35198 , \35199 );
xnor \U$34886 ( \35201 , \35200 , \22016 );
xor \U$34887 ( \35202 , \35197 , \35201 );
xor \U$34888 ( \35203 , \35188 , \35202 );
not \U$34889 ( \35204 , \22629 );
and \U$34890 ( \35205 , \21977 , \22641 );
and \U$34891 ( \35206 , \21990 , \22639 );
nor \U$34892 ( \35207 , \35205 , \35206 );
xnor \U$34893 ( \35208 , \35207 , \22651 );
xor \U$34894 ( \35209 , \35204 , \35208 );
and \U$34895 ( \35210 , \22030 , \22671 );
and \U$34896 ( \35211 , \22001 , \22669 );
nor \U$34897 ( \35212 , \35210 , \35211 );
xnor \U$34898 ( \35213 , \35212 , \22681 );
xor \U$34899 ( \35214 , \35209 , \35213 );
xor \U$34900 ( \35215 , \35203 , \35214 );
xor \U$34901 ( \35216 , \35177 , \35215 );
xor \U$34902 ( \35217 , \35171 , \35216 );
xor \U$34903 ( \35218 , \35152 , \35217 );
xor \U$34904 ( \35219 , \35146 , \35218 );
and \U$34905 ( \35220 , \35059 , \35139 );
nor \U$34906 ( \35221 , \35219 , \35220 );
nor \U$34907 ( \35222 , \35142 , \35221 );
nand \U$34908 ( \35223 , \35055 , \35222 );
and \U$34909 ( \35224 , \35150 , \35151 );
and \U$34910 ( \35225 , \35151 , \35217 );
and \U$34911 ( \35226 , \35150 , \35217 );
or \U$34912 ( \35227 , \35224 , \35225 , \35226 );
and \U$34913 ( \35228 , \35156 , \35170 );
and \U$34914 ( \35229 , \35170 , \35216 );
and \U$34915 ( \35230 , \35156 , \35216 );
or \U$34916 ( \35231 , \35228 , \35229 , \35230 );
xor \U$34917 ( \35232 , \35227 , \35231 );
and \U$34918 ( \35233 , \35175 , \35176 );
and \U$34919 ( \35234 , \35176 , \35215 );
and \U$34920 ( \35235 , \35175 , \35215 );
or \U$34921 ( \35236 , \35233 , \35234 , \35235 );
and \U$34922 ( \35237 , \35204 , \35208 );
and \U$34923 ( \35238 , \35208 , \35213 );
and \U$34924 ( \35239 , \35204 , \35213 );
or \U$34925 ( \35240 , \35237 , \35238 , \35239 );
and \U$34926 ( \35241 , \35192 , \35196 );
and \U$34927 ( \35242 , \35196 , \35201 );
and \U$34928 ( \35243 , \35192 , \35201 );
or \U$34929 ( \35244 , \35241 , \35242 , \35243 );
xor \U$34930 ( \35245 , \35240 , \35244 );
and \U$34931 ( \35246 , \35181 , \35185 );
and \U$34932 ( \35247 , \35185 , \35187 );
and \U$34933 ( \35248 , \35181 , \35187 );
or \U$34934 ( \35249 , \35246 , \35247 , \35248 );
xor \U$34935 ( \35250 , \35245 , \35249 );
xor \U$34936 ( \35251 , \35236 , \35250 );
and \U$34937 ( \35252 , \35160 , \35164 );
and \U$34938 ( \35253 , \35164 , \35169 );
and \U$34939 ( \35254 , \35160 , \35169 );
or \U$34940 ( \35255 , \35252 , \35253 , \35254 );
and \U$34941 ( \35256 , \35188 , \35202 );
and \U$34942 ( \35257 , \35202 , \35214 );
and \U$34943 ( \35258 , \35188 , \35214 );
or \U$34944 ( \35259 , \35256 , \35257 , \35258 );
xor \U$34945 ( \35260 , \35255 , \35259 );
and \U$34946 ( \35261 , \22124 , \21983 );
and \U$34947 ( \35262 , \22089 , \21981 );
nor \U$34948 ( \35263 , \35261 , \35262 );
xnor \U$34949 ( \35264 , \35263 , \21995 );
and \U$34950 ( \35265 , \22113 , \21978 );
xnor \U$34951 ( \35266 , \35264 , \35265 );
and \U$34952 ( \35267 , \22894 , \22720 );
and \U$34953 ( \35268 , \23230 , \22707 );
nor \U$34954 ( \35269 , \35267 , \35268 );
xnor \U$34955 ( \35270 , \35269 , \22067 );
and \U$34956 ( \35271 , \22081 , \23173 );
and \U$34957 ( \35272 , \22858 , \22999 );
nor \U$34958 ( \35273 , \35271 , \35272 );
xnor \U$34959 ( \35274 , \35273 , \22016 );
xor \U$34960 ( \35275 , \35270 , \35274 );
and \U$34961 ( \35276 , \22100 , \22021 );
and \U$34962 ( \35277 , \22071 , \22019 );
nor \U$34963 ( \35278 , \35276 , \35277 );
xnor \U$34964 ( \35279 , \35278 , \21595 );
xor \U$34965 ( \35280 , \35275 , \35279 );
xor \U$34966 ( \35281 , \35266 , \35280 );
and \U$34967 ( \35282 , \21990 , \22641 );
not \U$34968 ( \35283 , \35282 );
xnor \U$34969 ( \35284 , \35283 , \22651 );
and \U$34970 ( \35285 , \22001 , \22671 );
and \U$34971 ( \35286 , \21977 , \22669 );
nor \U$34972 ( \35287 , \35285 , \35286 );
xnor \U$34973 ( \35288 , \35287 , \22681 );
xor \U$34974 ( \35289 , \35284 , \35288 );
and \U$34975 ( \35290 , \23329 , \22691 );
and \U$34976 ( \35291 , \22030 , \22689 );
nor \U$34977 ( \35292 , \35290 , \35291 );
xnor \U$34978 ( \35293 , \35292 , \22701 );
xor \U$34979 ( \35294 , \35289 , \35293 );
xor \U$34980 ( \35295 , \35281 , \35294 );
xor \U$34981 ( \35296 , \35260 , \35295 );
xor \U$34982 ( \35297 , \35251 , \35296 );
xor \U$34983 ( \35298 , \35232 , \35297 );
and \U$34984 ( \35299 , \35146 , \35218 );
nor \U$34985 ( \35300 , \35298 , \35299 );
and \U$34986 ( \35301 , \35236 , \35250 );
and \U$34987 ( \35302 , \35250 , \35296 );
and \U$34988 ( \35303 , \35236 , \35296 );
or \U$34989 ( \35304 , \35301 , \35302 , \35303 );
and \U$34990 ( \35305 , \35255 , \35259 );
and \U$34991 ( \35306 , \35259 , \35295 );
and \U$34992 ( \35307 , \35255 , \35295 );
or \U$34993 ( \35308 , \35305 , \35306 , \35307 );
and \U$34994 ( \35309 , \35284 , \35288 );
and \U$34995 ( \35310 , \35288 , \35293 );
and \U$34996 ( \35311 , \35284 , \35293 );
or \U$34997 ( \35312 , \35309 , \35310 , \35311 );
and \U$34998 ( \35313 , \35270 , \35274 );
and \U$34999 ( \35314 , \35274 , \35279 );
and \U$35000 ( \35315 , \35270 , \35279 );
or \U$35001 ( \35316 , \35313 , \35314 , \35315 );
xor \U$35002 ( \35317 , \35312 , \35316 );
or \U$35003 ( \35318 , \35264 , \35265 );
xor \U$35004 ( \35319 , \35317 , \35318 );
xor \U$35005 ( \35320 , \35308 , \35319 );
and \U$35006 ( \35321 , \35240 , \35244 );
and \U$35007 ( \35322 , \35244 , \35249 );
and \U$35008 ( \35323 , \35240 , \35249 );
or \U$35009 ( \35324 , \35321 , \35322 , \35323 );
and \U$35010 ( \35325 , \35266 , \35280 );
and \U$35011 ( \35326 , \35280 , \35294 );
and \U$35012 ( \35327 , \35266 , \35294 );
or \U$35013 ( \35328 , \35325 , \35326 , \35327 );
xor \U$35014 ( \35329 , \35324 , \35328 );
and \U$35015 ( \35330 , \22089 , \21983 );
and \U$35016 ( \35331 , \22100 , \21981 );
nor \U$35017 ( \35332 , \35330 , \35331 );
xnor \U$35018 ( \35333 , \35332 , \21995 );
and \U$35019 ( \35334 , \22124 , \21978 );
xor \U$35020 ( \35335 , \35333 , \35334 );
and \U$35021 ( \35336 , \23230 , \22720 );
and \U$35022 ( \35337 , \23329 , \22707 );
nor \U$35023 ( \35338 , \35336 , \35337 );
xnor \U$35024 ( \35339 , \35338 , \22067 );
and \U$35025 ( \35340 , \22858 , \23173 );
and \U$35026 ( \35341 , \22894 , \22999 );
nor \U$35027 ( \35342 , \35340 , \35341 );
xnor \U$35028 ( \35343 , \35342 , \22016 );
xor \U$35029 ( \35344 , \35339 , \35343 );
and \U$35030 ( \35345 , \22071 , \22021 );
and \U$35031 ( \35346 , \22081 , \22019 );
nor \U$35032 ( \35347 , \35345 , \35346 );
xnor \U$35033 ( \35348 , \35347 , \21595 );
xor \U$35034 ( \35349 , \35344 , \35348 );
xor \U$35035 ( \35350 , \35335 , \35349 );
not \U$35036 ( \35351 , \22651 );
and \U$35037 ( \35352 , \21977 , \22671 );
and \U$35038 ( \35353 , \21990 , \22669 );
nor \U$35039 ( \35354 , \35352 , \35353 );
xnor \U$35040 ( \35355 , \35354 , \22681 );
xor \U$35041 ( \35356 , \35351 , \35355 );
and \U$35042 ( \35357 , \22030 , \22691 );
and \U$35043 ( \35358 , \22001 , \22689 );
nor \U$35044 ( \35359 , \35357 , \35358 );
xnor \U$35045 ( \35360 , \35359 , \22701 );
xor \U$35046 ( \35361 , \35356 , \35360 );
xor \U$35047 ( \35362 , \35350 , \35361 );
xor \U$35048 ( \35363 , \35329 , \35362 );
xor \U$35049 ( \35364 , \35320 , \35363 );
xor \U$35050 ( \35365 , \35304 , \35364 );
and \U$35051 ( \35366 , \35227 , \35231 );
and \U$35052 ( \35367 , \35231 , \35297 );
and \U$35053 ( \35368 , \35227 , \35297 );
or \U$35054 ( \35369 , \35366 , \35367 , \35368 );
nor \U$35055 ( \35370 , \35365 , \35369 );
nor \U$35056 ( \35371 , \35300 , \35370 );
and \U$35057 ( \35372 , \35308 , \35319 );
and \U$35058 ( \35373 , \35319 , \35363 );
and \U$35059 ( \35374 , \35308 , \35363 );
or \U$35060 ( \35375 , \35372 , \35373 , \35374 );
and \U$35061 ( \35376 , \35324 , \35328 );
and \U$35062 ( \35377 , \35328 , \35362 );
and \U$35063 ( \35378 , \35324 , \35362 );
or \U$35064 ( \35379 , \35376 , \35377 , \35378 );
and \U$35065 ( \35380 , \35351 , \35355 );
and \U$35066 ( \35381 , \35355 , \35360 );
and \U$35067 ( \35382 , \35351 , \35360 );
or \U$35068 ( \35383 , \35380 , \35381 , \35382 );
and \U$35069 ( \35384 , \35339 , \35343 );
and \U$35070 ( \35385 , \35343 , \35348 );
and \U$35071 ( \35386 , \35339 , \35348 );
or \U$35072 ( \35387 , \35384 , \35385 , \35386 );
xor \U$35073 ( \35388 , \35383 , \35387 );
and \U$35074 ( \35389 , \35333 , \35334 );
xor \U$35075 ( \35390 , \35388 , \35389 );
xor \U$35076 ( \35391 , \35379 , \35390 );
and \U$35077 ( \35392 , \35312 , \35316 );
and \U$35078 ( \35393 , \35316 , \35318 );
and \U$35079 ( \35394 , \35312 , \35318 );
or \U$35080 ( \35395 , \35392 , \35393 , \35394 );
and \U$35081 ( \35396 , \35335 , \35349 );
and \U$35082 ( \35397 , \35349 , \35361 );
and \U$35083 ( \35398 , \35335 , \35361 );
or \U$35084 ( \35399 , \35396 , \35397 , \35398 );
xor \U$35085 ( \35400 , \35395 , \35399 );
and \U$35086 ( \35401 , \22089 , \21978 );
not \U$35087 ( \35402 , \35401 );
and \U$35088 ( \35403 , \22894 , \23173 );
and \U$35089 ( \35404 , \23230 , \22999 );
nor \U$35090 ( \35405 , \35403 , \35404 );
xnor \U$35091 ( \35406 , \35405 , \22016 );
and \U$35092 ( \35407 , \22081 , \22021 );
and \U$35093 ( \35408 , \22858 , \22019 );
nor \U$35094 ( \35409 , \35407 , \35408 );
xnor \U$35095 ( \35410 , \35409 , \21595 );
xor \U$35096 ( \35411 , \35406 , \35410 );
and \U$35097 ( \35412 , \22100 , \21983 );
and \U$35098 ( \35413 , \22071 , \21981 );
nor \U$35099 ( \35414 , \35412 , \35413 );
xnor \U$35100 ( \35415 , \35414 , \21995 );
xor \U$35101 ( \35416 , \35411 , \35415 );
xor \U$35102 ( \35417 , \35402 , \35416 );
and \U$35103 ( \35418 , \21990 , \22671 );
not \U$35104 ( \35419 , \35418 );
xnor \U$35105 ( \35420 , \35419 , \22681 );
and \U$35106 ( \35421 , \22001 , \22691 );
and \U$35107 ( \35422 , \21977 , \22689 );
nor \U$35108 ( \35423 , \35421 , \35422 );
xnor \U$35109 ( \35424 , \35423 , \22701 );
xor \U$35110 ( \35425 , \35420 , \35424 );
and \U$35111 ( \35426 , \23329 , \22720 );
and \U$35112 ( \35427 , \22030 , \22707 );
nor \U$35113 ( \35428 , \35426 , \35427 );
xnor \U$35114 ( \35429 , \35428 , \22067 );
xor \U$35115 ( \35430 , \35425 , \35429 );
xor \U$35116 ( \35431 , \35417 , \35430 );
xor \U$35117 ( \35432 , \35400 , \35431 );
xor \U$35118 ( \35433 , \35391 , \35432 );
xor \U$35119 ( \35434 , \35375 , \35433 );
and \U$35120 ( \35435 , \35304 , \35364 );
nor \U$35121 ( \35436 , \35434 , \35435 );
and \U$35122 ( \35437 , \35379 , \35390 );
and \U$35123 ( \35438 , \35390 , \35432 );
and \U$35124 ( \35439 , \35379 , \35432 );
or \U$35125 ( \35440 , \35437 , \35438 , \35439 );
and \U$35126 ( \35441 , \35395 , \35399 );
and \U$35127 ( \35442 , \35399 , \35431 );
and \U$35128 ( \35443 , \35395 , \35431 );
or \U$35129 ( \35444 , \35441 , \35442 , \35443 );
and \U$35130 ( \35445 , \35420 , \35424 );
and \U$35131 ( \35446 , \35424 , \35429 );
and \U$35132 ( \35447 , \35420 , \35429 );
or \U$35133 ( \35448 , \35445 , \35446 , \35447 );
and \U$35134 ( \35449 , \35406 , \35410 );
and \U$35135 ( \35450 , \35410 , \35415 );
and \U$35136 ( \35451 , \35406 , \35415 );
or \U$35137 ( \35452 , \35449 , \35450 , \35451 );
xor \U$35138 ( \35453 , \35448 , \35452 );
xor \U$35139 ( \35454 , \35453 , \35401 );
xor \U$35140 ( \35455 , \35444 , \35454 );
and \U$35141 ( \35456 , \35383 , \35387 );
and \U$35142 ( \35457 , \35387 , \35389 );
and \U$35143 ( \35458 , \35383 , \35389 );
or \U$35144 ( \35459 , \35456 , \35457 , \35458 );
and \U$35145 ( \35460 , \35402 , \35416 );
and \U$35146 ( \35461 , \35416 , \35430 );
and \U$35147 ( \35462 , \35402 , \35430 );
or \U$35148 ( \35463 , \35460 , \35461 , \35462 );
xor \U$35149 ( \35464 , \35459 , \35463 );
and \U$35150 ( \35465 , \22100 , \21978 );
and \U$35151 ( \35466 , \23230 , \23173 );
and \U$35152 ( \35467 , \23329 , \22999 );
nor \U$35153 ( \35468 , \35466 , \35467 );
xnor \U$35154 ( \35469 , \35468 , \22016 );
and \U$35155 ( \35470 , \22858 , \22021 );
and \U$35156 ( \35471 , \22894 , \22019 );
nor \U$35157 ( \35472 , \35470 , \35471 );
xnor \U$35158 ( \35473 , \35472 , \21595 );
xor \U$35159 ( \35474 , \35469 , \35473 );
and \U$35160 ( \35475 , \22071 , \21983 );
and \U$35161 ( \35476 , \22081 , \21981 );
nor \U$35162 ( \35477 , \35475 , \35476 );
xnor \U$35163 ( \35478 , \35477 , \21995 );
xor \U$35164 ( \35479 , \35474 , \35478 );
xor \U$35165 ( \35480 , \35465 , \35479 );
not \U$35166 ( \35481 , \22681 );
and \U$35167 ( \35482 , \21977 , \22691 );
and \U$35168 ( \35483 , \21990 , \22689 );
nor \U$35169 ( \35484 , \35482 , \35483 );
xnor \U$35170 ( \35485 , \35484 , \22701 );
xor \U$35171 ( \35486 , \35481 , \35485 );
and \U$35172 ( \35487 , \22030 , \22720 );
and \U$35173 ( \35488 , \22001 , \22707 );
nor \U$35174 ( \35489 , \35487 , \35488 );
xnor \U$35175 ( \35490 , \35489 , \22067 );
xor \U$35176 ( \35491 , \35486 , \35490 );
xor \U$35177 ( \35492 , \35480 , \35491 );
xor \U$35178 ( \35493 , \35464 , \35492 );
xor \U$35179 ( \35494 , \35455 , \35493 );
xor \U$35180 ( \35495 , \35440 , \35494 );
and \U$35181 ( \35496 , \35375 , \35433 );
nor \U$35182 ( \35497 , \35495 , \35496 );
nor \U$35183 ( \35498 , \35436 , \35497 );
nand \U$35184 ( \35499 , \35371 , \35498 );
nor \U$35185 ( \35500 , \35223 , \35499 );
and \U$35186 ( \35501 , \35444 , \35454 );
and \U$35187 ( \35502 , \35454 , \35493 );
and \U$35188 ( \35503 , \35444 , \35493 );
or \U$35189 ( \35504 , \35501 , \35502 , \35503 );
and \U$35190 ( \35505 , \35459 , \35463 );
and \U$35191 ( \35506 , \35463 , \35492 );
and \U$35192 ( \35507 , \35459 , \35492 );
or \U$35193 ( \35508 , \35505 , \35506 , \35507 );
and \U$35194 ( \35509 , \21990 , \22691 );
not \U$35195 ( \35510 , \35509 );
xnor \U$35196 ( \35511 , \35510 , \22701 );
and \U$35197 ( \35512 , \22001 , \22720 );
and \U$35198 ( \35513 , \21977 , \22707 );
nor \U$35199 ( \35514 , \35512 , \35513 );
xnor \U$35200 ( \35515 , \35514 , \22067 );
xor \U$35201 ( \35516 , \35511 , \35515 );
and \U$35202 ( \35517 , \23329 , \23173 );
and \U$35203 ( \35518 , \22030 , \22999 );
nor \U$35204 ( \35519 , \35517 , \35518 );
xnor \U$35205 ( \35520 , \35519 , \22016 );
xor \U$35206 ( \35521 , \35516 , \35520 );
and \U$35207 ( \35522 , \35481 , \35485 );
and \U$35208 ( \35523 , \35485 , \35490 );
and \U$35209 ( \35524 , \35481 , \35490 );
or \U$35210 ( \35525 , \35522 , \35523 , \35524 );
and \U$35211 ( \35526 , \35469 , \35473 );
and \U$35212 ( \35527 , \35473 , \35478 );
and \U$35213 ( \35528 , \35469 , \35478 );
or \U$35214 ( \35529 , \35526 , \35527 , \35528 );
xnor \U$35215 ( \35530 , \35525 , \35529 );
xor \U$35216 ( \35531 , \35521 , \35530 );
xor \U$35217 ( \35532 , \35508 , \35531 );
and \U$35218 ( \35533 , \35448 , \35452 );
and \U$35219 ( \35534 , \35452 , \35401 );
and \U$35220 ( \35535 , \35448 , \35401 );
or \U$35221 ( \35536 , \35533 , \35534 , \35535 );
and \U$35222 ( \35537 , \35465 , \35479 );
and \U$35223 ( \35538 , \35479 , \35491 );
and \U$35224 ( \35539 , \35465 , \35491 );
or \U$35225 ( \35540 , \35537 , \35538 , \35539 );
xor \U$35226 ( \35541 , \35536 , \35540 );
and \U$35227 ( \35542 , \22894 , \22021 );
and \U$35228 ( \35543 , \23230 , \22019 );
nor \U$35229 ( \35544 , \35542 , \35543 );
xnor \U$35230 ( \35545 , \35544 , \21595 );
and \U$35231 ( \35546 , \22081 , \21983 );
and \U$35232 ( \35547 , \22858 , \21981 );
nor \U$35233 ( \35548 , \35546 , \35547 );
xnor \U$35234 ( \35549 , \35548 , \21995 );
xor \U$35235 ( \35550 , \35545 , \35549 );
and \U$35236 ( \35551 , \22071 , \21978 );
xor \U$35237 ( \35552 , \35550 , \35551 );
xor \U$35238 ( \35553 , \35541 , \35552 );
xor \U$35239 ( \35554 , \35532 , \35553 );
xor \U$35240 ( \35555 , \35504 , \35554 );
and \U$35241 ( \35556 , \35440 , \35494 );
nor \U$35242 ( \35557 , \35555 , \35556 );
and \U$35243 ( \35558 , \35508 , \35531 );
and \U$35244 ( \35559 , \35531 , \35553 );
and \U$35245 ( \35560 , \35508 , \35553 );
or \U$35246 ( \35561 , \35558 , \35559 , \35560 );
and \U$35247 ( \35562 , \35536 , \35540 );
and \U$35248 ( \35563 , \35540 , \35552 );
and \U$35249 ( \35564 , \35536 , \35552 );
or \U$35250 ( \35565 , \35562 , \35563 , \35564 );
and \U$35251 ( \35566 , \35521 , \35530 );
xor \U$35252 ( \35567 , \35565 , \35566 );
or \U$35253 ( \35568 , \35525 , \35529 );
not \U$35254 ( \35569 , \22701 );
and \U$35255 ( \35570 , \21977 , \22720 );
and \U$35256 ( \35571 , \21990 , \22707 );
nor \U$35257 ( \35572 , \35570 , \35571 );
xnor \U$35258 ( \35573 , \35572 , \22067 );
xor \U$35259 ( \35574 , \35569 , \35573 );
and \U$35260 ( \35575 , \22030 , \23173 );
and \U$35261 ( \35576 , \22001 , \22999 );
nor \U$35262 ( \35577 , \35575 , \35576 );
xnor \U$35263 ( \35578 , \35577 , \22016 );
xor \U$35264 ( \35579 , \35574 , \35578 );
xor \U$35265 ( \35580 , \35568 , \35579 );
and \U$35266 ( \35581 , \35511 , \35515 );
and \U$35267 ( \35582 , \35515 , \35520 );
and \U$35268 ( \35583 , \35511 , \35520 );
or \U$35269 ( \35584 , \35581 , \35582 , \35583 );
and \U$35270 ( \35585 , \35545 , \35549 );
and \U$35271 ( \35586 , \35549 , \35551 );
and \U$35272 ( \35587 , \35545 , \35551 );
or \U$35273 ( \35588 , \35585 , \35586 , \35587 );
xor \U$35274 ( \35589 , \35584 , \35588 );
and \U$35275 ( \35590 , \23230 , \22021 );
and \U$35276 ( \35591 , \23329 , \22019 );
nor \U$35277 ( \35592 , \35590 , \35591 );
xnor \U$35278 ( \35593 , \35592 , \21595 );
and \U$35279 ( \35594 , \22858 , \21983 );
and \U$35280 ( \35595 , \22894 , \21981 );
nor \U$35281 ( \35596 , \35594 , \35595 );
xnor \U$35282 ( \35597 , \35596 , \21995 );
xor \U$35283 ( \35598 , \35593 , \35597 );
and \U$35284 ( \35599 , \22081 , \21978 );
xor \U$35285 ( \35600 , \35598 , \35599 );
xor \U$35286 ( \35601 , \35589 , \35600 );
xor \U$35287 ( \35602 , \35580 , \35601 );
xor \U$35288 ( \35603 , \35567 , \35602 );
xor \U$35289 ( \35604 , \35561 , \35603 );
and \U$35290 ( \35605 , \35504 , \35554 );
nor \U$35291 ( \35606 , \35604 , \35605 );
nor \U$35292 ( \35607 , \35557 , \35606 );
and \U$35293 ( \35608 , \35565 , \35566 );
and \U$35294 ( \35609 , \35566 , \35602 );
and \U$35295 ( \35610 , \35565 , \35602 );
or \U$35296 ( \35611 , \35608 , \35609 , \35610 );
and \U$35297 ( \35612 , \35568 , \35579 );
and \U$35298 ( \35613 , \35579 , \35601 );
and \U$35299 ( \35614 , \35568 , \35601 );
or \U$35300 ( \35615 , \35612 , \35613 , \35614 );
xor \U$35301 ( \35616 , \35611 , \35615 );
and \U$35302 ( \35617 , \35584 , \35588 );
and \U$35303 ( \35618 , \35588 , \35600 );
and \U$35304 ( \35619 , \35584 , \35600 );
or \U$35305 ( \35620 , \35617 , \35618 , \35619 );
and \U$35306 ( \35621 , \21990 , \22720 );
not \U$35307 ( \35622 , \35621 );
xnor \U$35308 ( \35623 , \35622 , \22067 );
and \U$35309 ( \35624 , \22001 , \23173 );
and \U$35310 ( \35625 , \21977 , \22999 );
nor \U$35311 ( \35626 , \35624 , \35625 );
xnor \U$35312 ( \35627 , \35626 , \22016 );
xor \U$35313 ( \35628 , \35623 , \35627 );
and \U$35314 ( \35629 , \23329 , \22021 );
and \U$35315 ( \35630 , \22030 , \22019 );
nor \U$35316 ( \35631 , \35629 , \35630 );
xnor \U$35317 ( \35632 , \35631 , \21595 );
xor \U$35318 ( \35633 , \35628 , \35632 );
xor \U$35319 ( \35634 , \35620 , \35633 );
and \U$35320 ( \35635 , \35569 , \35573 );
and \U$35321 ( \35636 , \35573 , \35578 );
and \U$35322 ( \35637 , \35569 , \35578 );
or \U$35323 ( \35638 , \35635 , \35636 , \35637 );
and \U$35324 ( \35639 , \35593 , \35597 );
and \U$35325 ( \35640 , \35597 , \35599 );
and \U$35326 ( \35641 , \35593 , \35599 );
or \U$35327 ( \35642 , \35639 , \35640 , \35641 );
xor \U$35328 ( \35643 , \35638 , \35642 );
and \U$35329 ( \35644 , \22894 , \21983 );
and \U$35330 ( \35645 , \23230 , \21981 );
nor \U$35331 ( \35646 , \35644 , \35645 );
xnor \U$35332 ( \35647 , \35646 , \21995 );
and \U$35333 ( \35648 , \22858 , \21978 );
xnor \U$35334 ( \35649 , \35647 , \35648 );
xor \U$35335 ( \35650 , \35643 , \35649 );
xor \U$35336 ( \35651 , \35634 , \35650 );
xor \U$35337 ( \35652 , \35616 , \35651 );
and \U$35338 ( \35653 , \35561 , \35603 );
nor \U$35339 ( \35654 , \35652 , \35653 );
and \U$35340 ( \35655 , \35620 , \35633 );
and \U$35341 ( \35656 , \35633 , \35650 );
and \U$35342 ( \35657 , \35620 , \35650 );
or \U$35343 ( \35658 , \35655 , \35656 , \35657 );
and \U$35344 ( \35659 , \35638 , \35642 );
and \U$35345 ( \35660 , \35642 , \35649 );
and \U$35346 ( \35661 , \35638 , \35649 );
or \U$35347 ( \35662 , \35659 , \35660 , \35661 );
and \U$35348 ( \35663 , \22894 , \21978 );
not \U$35349 ( \35664 , \22067 );
and \U$35350 ( \35665 , \21977 , \23173 );
and \U$35351 ( \35666 , \21990 , \22999 );
nor \U$35352 ( \35667 , \35665 , \35666 );
xnor \U$35353 ( \35668 , \35667 , \22016 );
xor \U$35354 ( \35669 , \35664 , \35668 );
and \U$35355 ( \35670 , \22030 , \22021 );
and \U$35356 ( \35671 , \22001 , \22019 );
nor \U$35357 ( \35672 , \35670 , \35671 );
xnor \U$35358 ( \35673 , \35672 , \21595 );
xor \U$35359 ( \35674 , \35669 , \35673 );
xor \U$35360 ( \35675 , \35663 , \35674 );
xor \U$35361 ( \35676 , \35662 , \35675 );
and \U$35362 ( \35677 , \35623 , \35627 );
and \U$35363 ( \35678 , \35627 , \35632 );
and \U$35364 ( \35679 , \35623 , \35632 );
or \U$35365 ( \35680 , \35677 , \35678 , \35679 );
or \U$35366 ( \35681 , \35647 , \35648 );
xor \U$35367 ( \35682 , \35680 , \35681 );
and \U$35368 ( \35683 , \23230 , \21983 );
and \U$35369 ( \35684 , \23329 , \21981 );
nor \U$35370 ( \35685 , \35683 , \35684 );
xnor \U$35371 ( \35686 , \35685 , \21995 );
xor \U$35372 ( \35687 , \35682 , \35686 );
xor \U$35373 ( \35688 , \35676 , \35687 );
xor \U$35374 ( \35689 , \35658 , \35688 );
and \U$35375 ( \35690 , \35611 , \35615 );
and \U$35376 ( \35691 , \35615 , \35651 );
and \U$35377 ( \35692 , \35611 , \35651 );
or \U$35378 ( \35693 , \35690 , \35691 , \35692 );
nor \U$35379 ( \35694 , \35689 , \35693 );
nor \U$35380 ( \35695 , \35654 , \35694 );
nand \U$35381 ( \35696 , \35607 , \35695 );
and \U$35382 ( \35697 , \35662 , \35675 );
and \U$35383 ( \35698 , \35675 , \35687 );
and \U$35384 ( \35699 , \35662 , \35687 );
or \U$35385 ( \35700 , \35697 , \35698 , \35699 );
and \U$35386 ( \35701 , \35680 , \35681 );
and \U$35387 ( \35702 , \35681 , \35686 );
and \U$35388 ( \35703 , \35680 , \35686 );
or \U$35389 ( \35704 , \35701 , \35702 , \35703 );
and \U$35390 ( \35705 , \35663 , \35674 );
xor \U$35391 ( \35706 , \35704 , \35705 );
and \U$35392 ( \35707 , \35664 , \35668 );
and \U$35393 ( \35708 , \35668 , \35673 );
and \U$35394 ( \35709 , \35664 , \35673 );
or \U$35395 ( \35710 , \35707 , \35708 , \35709 );
and \U$35396 ( \35711 , \23230 , \21978 );
not \U$35397 ( \35712 , \35711 );
xor \U$35398 ( \35713 , \35710 , \35712 );
and \U$35399 ( \35714 , \21990 , \23173 );
not \U$35400 ( \35715 , \35714 );
xnor \U$35401 ( \35716 , \35715 , \22016 );
and \U$35402 ( \35717 , \22001 , \22021 );
and \U$35403 ( \35718 , \21977 , \22019 );
nor \U$35404 ( \35719 , \35717 , \35718 );
xnor \U$35405 ( \35720 , \35719 , \21595 );
xor \U$35406 ( \35721 , \35716 , \35720 );
and \U$35407 ( \35722 , \23329 , \21983 );
and \U$35408 ( \35723 , \22030 , \21981 );
nor \U$35409 ( \35724 , \35722 , \35723 );
xnor \U$35410 ( \35725 , \35724 , \21995 );
xor \U$35411 ( \35726 , \35721 , \35725 );
xor \U$35412 ( \35727 , \35713 , \35726 );
xor \U$35413 ( \35728 , \35706 , \35727 );
xor \U$35414 ( \35729 , \35700 , \35728 );
and \U$35415 ( \35730 , \35658 , \35688 );
nor \U$35416 ( \35731 , \35729 , \35730 );
and \U$35417 ( \35732 , \35704 , \35705 );
and \U$35418 ( \35733 , \35705 , \35727 );
and \U$35419 ( \35734 , \35704 , \35727 );
or \U$35420 ( \35735 , \35732 , \35733 , \35734 );
and \U$35421 ( \35736 , \35710 , \35712 );
and \U$35422 ( \35737 , \35712 , \35726 );
and \U$35423 ( \35738 , \35710 , \35726 );
or \U$35424 ( \35739 , \35736 , \35737 , \35738 );
xor \U$35425 ( \35740 , \22017 , \22025 );
xor \U$35426 ( \35741 , \35740 , \22034 );
xor \U$35427 ( \35742 , \35739 , \35741 );
and \U$35428 ( \35743 , \35716 , \35720 );
and \U$35429 ( \35744 , \35720 , \35725 );
and \U$35430 ( \35745 , \35716 , \35725 );
or \U$35431 ( \35746 , \35743 , \35744 , \35745 );
xor \U$35432 ( \35747 , \35746 , \35711 );
and \U$35433 ( \35748 , \23329 , \21978 );
xor \U$35434 ( \35749 , \35747 , \35748 );
xor \U$35435 ( \35750 , \35742 , \35749 );
xor \U$35436 ( \35751 , \35735 , \35750 );
and \U$35437 ( \35752 , \35700 , \35728 );
nor \U$35438 ( \35753 , \35751 , \35752 );
nor \U$35439 ( \35754 , \35731 , \35753 );
and \U$35440 ( \35755 , \35739 , \35741 );
and \U$35441 ( \35756 , \35741 , \35749 );
and \U$35442 ( \35757 , \35739 , \35749 );
or \U$35443 ( \35758 , \35755 , \35756 , \35757 );
and \U$35444 ( \35759 , \35746 , \35711 );
and \U$35445 ( \35760 , \35711 , \35748 );
and \U$35446 ( \35761 , \35746 , \35748 );
or \U$35447 ( \35762 , \35759 , \35760 , \35761 );
xor \U$35448 ( \35763 , \35758 , \35762 );
xnor \U$35449 ( \35764 , \22037 , \22047 );
xor \U$35450 ( \35765 , \35763 , \35764 );
and \U$35451 ( \35766 , \35735 , \35750 );
nor \U$35452 ( \35767 , \35765 , \35766 );
xor \U$35453 ( \35768 , \22048 , \22052 );
xor \U$35454 ( \35769 , \35768 , \22055 );
and \U$35455 ( \35770 , \35758 , \35762 );
and \U$35456 ( \35771 , \35762 , \35764 );
and \U$35457 ( \35772 , \35758 , \35764 );
or \U$35458 ( \35773 , \35770 , \35771 , \35772 );
nor \U$35459 ( \35774 , \35769 , \35773 );
nor \U$35460 ( \35775 , \35767 , \35774 );
nand \U$35461 ( \35776 , \35754 , \35775 );
nor \U$35462 ( \35777 , \35696 , \35776 );
nand \U$35463 ( \35778 , \35500 , \35777 );
nor \U$35464 ( \35779 , \34868 , \35778 );
nand \U$35465 ( \35780 , \32642 , \35779 );
and \U$35466 ( \35781 , \22407 , \22076 );
and \U$35467 ( \35782 , \22418 , \22073 );
nor \U$35468 ( \35783 , \35781 , \35782 );
xnor \U$35469 ( \35784 , \35783 , \22072 );
and \U$35470 ( \35785 , \22377 , \35784 );
and \U$35471 ( \35786 , \22429 , \22095 );
and \U$35472 ( \35787 , \22440 , \22093 );
nor \U$35473 ( \35788 , \35786 , \35787 );
xnor \U$35474 ( \35789 , \35788 , \22105 );
and \U$35475 ( \35790 , \35784 , \35789 );
and \U$35476 ( \35791 , \22377 , \35789 );
or \U$35477 ( \35792 , \35785 , \35790 , \35791 );
and \U$35478 ( \35793 , \22457 , \22119 );
and \U$35479 ( \35794 , \22468 , \22117 );
nor \U$35480 ( \35795 , \35793 , \35794 );
xnor \U$35481 ( \35796 , \35795 , \22129 );
and \U$35482 ( \35797 , \22478 , \22140 );
and \U$35483 ( \35798 , \22489 , \22138 );
nor \U$35484 ( \35799 , \35797 , \35798 );
xnor \U$35485 ( \35800 , \35799 , \22150 );
and \U$35486 ( \35801 , \35796 , \35800 );
and \U$35487 ( \35802 , \22500 , \22162 );
and \U$35488 ( \35803 , \22511 , \22160 );
nor \U$35489 ( \35804 , \35802 , \35803 );
xnor \U$35490 ( \35805 , \35804 , \22172 );
and \U$35491 ( \35806 , \35800 , \35805 );
and \U$35492 ( \35807 , \35796 , \35805 );
or \U$35493 ( \35808 , \35801 , \35806 , \35807 );
and \U$35494 ( \35809 , \35792 , \35808 );
and \U$35495 ( \35810 , \22524 , \22187 );
and \U$35496 ( \35811 , \22535 , \22185 );
nor \U$35497 ( \35812 , \35810 , \35811 );
xnor \U$35498 ( \35813 , \35812 , \22197 );
and \U$35499 ( \35814 , \22545 , \22208 );
and \U$35500 ( \35815 , \22556 , \22206 );
nor \U$35501 ( \35816 , \35814 , \35815 );
xnor \U$35502 ( \35817 , \35816 , \22218 );
and \U$35503 ( \35818 , \35813 , \35817 );
and \U$35504 ( \35819 , \22567 , \22230 );
and \U$35505 ( \35820 , \22578 , \22228 );
nor \U$35506 ( \35821 , \35819 , \35820 );
xnor \U$35507 ( \35822 , \35821 , \22240 );
and \U$35508 ( \35823 , \35817 , \35822 );
and \U$35509 ( \35824 , \35813 , \35822 );
or \U$35510 ( \35825 , \35818 , \35823 , \35824 );
and \U$35511 ( \35826 , \35808 , \35825 );
and \U$35512 ( \35827 , \35792 , \35825 );
or \U$35513 ( \35828 , \35809 , \35826 , \35827 );
and \U$35514 ( \35829 , \22592 , \22257 );
and \U$35515 ( \35830 , \22603 , \22255 );
nor \U$35516 ( \35831 , \35829 , \35830 );
xnor \U$35517 ( \35832 , \35831 , \22267 );
and \U$35518 ( \35833 , \22613 , \22278 );
and \U$35519 ( \35834 , \22624 , \22276 );
nor \U$35520 ( \35835 , \35833 , \35834 );
xnor \U$35521 ( \35836 , \35835 , \22288 );
and \U$35522 ( \35837 , \35832 , \35836 );
and \U$35523 ( \35838 , \22635 , \22300 );
and \U$35524 ( \35839 , \22646 , \22298 );
nor \U$35525 ( \35840 , \35838 , \35839 );
xnor \U$35526 ( \35841 , \35840 , \22310 );
and \U$35527 ( \35842 , \35836 , \35841 );
and \U$35528 ( \35843 , \35832 , \35841 );
or \U$35529 ( \35844 , \35837 , \35842 , \35843 );
and \U$35530 ( \35845 , \22665 , \22324 );
and \U$35531 ( \35846 , \22676 , \22322 );
nor \U$35532 ( \35847 , \35845 , \35846 );
xnor \U$35533 ( \35848 , \35847 , \22334 );
and \U$35534 ( \35849 , \22686 , \22345 );
and \U$35535 ( \35850 , \22696 , \22343 );
nor \U$35536 ( \35851 , \35849 , \35850 );
xnor \U$35537 ( \35852 , \35851 , \22355 );
and \U$35538 ( \35853 , \35848 , \35852 );
nand \U$35539 ( \35854 , \22706 , \22365 );
xnor \U$35540 ( \35855 , \35854 , \22377 );
and \U$35541 ( \35856 , \35852 , \35855 );
and \U$35542 ( \35857 , \35848 , \35855 );
or \U$35543 ( \35858 , \35853 , \35856 , \35857 );
and \U$35544 ( \35859 , \35844 , \35858 );
and \U$35545 ( \35860 , \22696 , \22345 );
and \U$35546 ( \35861 , \22665 , \22343 );
nor \U$35547 ( \35862 , \35860 , \35861 );
xnor \U$35548 ( \35863 , \35862 , \22355 );
and \U$35549 ( \35864 , \35858 , \35863 );
and \U$35550 ( \35865 , \35844 , \35863 );
or \U$35551 ( \35866 , \35859 , \35864 , \35865 );
and \U$35552 ( \35867 , \35828 , \35866 );
and \U$35553 ( \35868 , \22706 , \22367 );
and \U$35554 ( \35869 , \22686 , \22365 );
nor \U$35555 ( \35870 , \35868 , \35869 );
xnor \U$35556 ( \35871 , \35870 , \22377 );
and \U$35557 ( \35872 , \22624 , \22278 );
and \U$35558 ( \35873 , \22592 , \22276 );
nor \U$35559 ( \35874 , \35872 , \35873 );
xnor \U$35560 ( \35875 , \35874 , \22288 );
and \U$35561 ( \35876 , \22646 , \22300 );
and \U$35562 ( \35877 , \22613 , \22298 );
nor \U$35563 ( \35878 , \35876 , \35877 );
xnor \U$35564 ( \35879 , \35878 , \22310 );
xor \U$35565 ( \35880 , \35875 , \35879 );
and \U$35566 ( \35881 , \22676 , \22324 );
and \U$35567 ( \35882 , \22635 , \22322 );
nor \U$35568 ( \35883 , \35881 , \35882 );
xnor \U$35569 ( \35884 , \35883 , \22334 );
xor \U$35570 ( \35885 , \35880 , \35884 );
and \U$35571 ( \35886 , \35871 , \35885 );
and \U$35572 ( \35887 , \22556 , \22208 );
and \U$35573 ( \35888 , \22524 , \22206 );
nor \U$35574 ( \35889 , \35887 , \35888 );
xnor \U$35575 ( \35890 , \35889 , \22218 );
and \U$35576 ( \35891 , \22578 , \22230 );
and \U$35577 ( \35892 , \22545 , \22228 );
nor \U$35578 ( \35893 , \35891 , \35892 );
xnor \U$35579 ( \35894 , \35893 , \22240 );
xor \U$35580 ( \35895 , \35890 , \35894 );
and \U$35581 ( \35896 , \22603 , \22257 );
and \U$35582 ( \35897 , \22567 , \22255 );
nor \U$35583 ( \35898 , \35896 , \35897 );
xnor \U$35584 ( \35899 , \35898 , \22267 );
xor \U$35585 ( \35900 , \35895 , \35899 );
and \U$35586 ( \35901 , \35885 , \35900 );
and \U$35587 ( \35902 , \35871 , \35900 );
or \U$35588 ( \35903 , \35886 , \35901 , \35902 );
and \U$35589 ( \35904 , \35866 , \35903 );
and \U$35590 ( \35905 , \35828 , \35903 );
or \U$35591 ( \35906 , \35867 , \35904 , \35905 );
and \U$35592 ( \35907 , \22386 , \22076 );
and \U$35593 ( \35908 , \22397 , \22073 );
nor \U$35594 ( \35909 , \35907 , \35908 );
xnor \U$35595 ( \35910 , \35909 , \22072 );
xor \U$35596 ( \35911 , \22402 , \35910 );
and \U$35597 ( \35912 , \22407 , \22095 );
and \U$35598 ( \35913 , \22418 , \22093 );
nor \U$35599 ( \35914 , \35912 , \35913 );
xnor \U$35600 ( \35915 , \35914 , \22105 );
xor \U$35601 ( \35916 , \35911 , \35915 );
and \U$35602 ( \35917 , \22567 , \22257 );
and \U$35603 ( \35918 , \22578 , \22255 );
nor \U$35604 ( \35919 , \35917 , \35918 );
xnor \U$35605 ( \35920 , \35919 , \22267 );
and \U$35606 ( \35921 , \22592 , \22278 );
and \U$35607 ( \35922 , \22603 , \22276 );
nor \U$35608 ( \35923 , \35921 , \35922 );
xnor \U$35609 ( \35924 , \35923 , \22288 );
xor \U$35610 ( \35925 , \35920 , \35924 );
and \U$35611 ( \35926 , \22613 , \22300 );
and \U$35612 ( \35927 , \22624 , \22298 );
nor \U$35613 ( \35928 , \35926 , \35927 );
xnor \U$35614 ( \35929 , \35928 , \22310 );
xor \U$35615 ( \35930 , \35925 , \35929 );
and \U$35616 ( \35931 , \22500 , \22187 );
and \U$35617 ( \35932 , \22511 , \22185 );
nor \U$35618 ( \35933 , \35931 , \35932 );
xnor \U$35619 ( \35934 , \35933 , \22197 );
and \U$35620 ( \35935 , \22524 , \22208 );
and \U$35621 ( \35936 , \22535 , \22206 );
nor \U$35622 ( \35937 , \35935 , \35936 );
xnor \U$35623 ( \35938 , \35937 , \22218 );
xor \U$35624 ( \35939 , \35934 , \35938 );
and \U$35625 ( \35940 , \22545 , \22230 );
and \U$35626 ( \35941 , \22556 , \22228 );
nor \U$35627 ( \35942 , \35940 , \35941 );
xnor \U$35628 ( \35943 , \35942 , \22240 );
xor \U$35629 ( \35944 , \35939 , \35943 );
xor \U$35630 ( \35945 , \35930 , \35944 );
and \U$35631 ( \35946 , \22429 , \22119 );
and \U$35632 ( \35947 , \22440 , \22117 );
nor \U$35633 ( \35948 , \35946 , \35947 );
xnor \U$35634 ( \35949 , \35948 , \22129 );
and \U$35635 ( \35950 , \22457 , \22140 );
and \U$35636 ( \35951 , \22468 , \22138 );
nor \U$35637 ( \35952 , \35950 , \35951 );
xnor \U$35638 ( \35953 , \35952 , \22150 );
xor \U$35639 ( \35954 , \35949 , \35953 );
and \U$35640 ( \35955 , \22478 , \22162 );
and \U$35641 ( \35956 , \22489 , \22160 );
nor \U$35642 ( \35957 , \35955 , \35956 );
xnor \U$35643 ( \35958 , \35957 , \22172 );
xor \U$35644 ( \35959 , \35954 , \35958 );
xor \U$35645 ( \35960 , \35945 , \35959 );
and \U$35646 ( \35961 , \35916 , \35960 );
and \U$35647 ( \35962 , \35875 , \35879 );
and \U$35648 ( \35963 , \35879 , \35884 );
and \U$35649 ( \35964 , \35875 , \35884 );
or \U$35650 ( \35965 , \35962 , \35963 , \35964 );
nand \U$35651 ( \35966 , \22706 , \22390 );
xnor \U$35652 ( \35967 , \35966 , \22402 );
xor \U$35653 ( \35968 , \35965 , \35967 );
and \U$35654 ( \35969 , \22635 , \22324 );
and \U$35655 ( \35970 , \22646 , \22322 );
nor \U$35656 ( \35971 , \35969 , \35970 );
xnor \U$35657 ( \35972 , \35971 , \22334 );
and \U$35658 ( \35973 , \22665 , \22345 );
and \U$35659 ( \35974 , \22676 , \22343 );
nor \U$35660 ( \35975 , \35973 , \35974 );
xnor \U$35661 ( \35976 , \35975 , \22355 );
xor \U$35662 ( \35977 , \35972 , \35976 );
and \U$35663 ( \35978 , \22686 , \22367 );
and \U$35664 ( \35979 , \22696 , \22365 );
nor \U$35665 ( \35980 , \35978 , \35979 );
xnor \U$35666 ( \35981 , \35980 , \22377 );
xor \U$35667 ( \35982 , \35977 , \35981 );
xor \U$35668 ( \35983 , \35968 , \35982 );
and \U$35669 ( \35984 , \35960 , \35983 );
and \U$35670 ( \35985 , \35916 , \35983 );
or \U$35671 ( \35986 , \35961 , \35984 , \35985 );
and \U$35672 ( \35987 , \35906 , \35986 );
and \U$35673 ( \35988 , \22402 , \35910 );
and \U$35674 ( \35989 , \35910 , \35915 );
and \U$35675 ( \35990 , \22402 , \35915 );
or \U$35676 ( \35991 , \35988 , \35989 , \35990 );
and \U$35677 ( \35992 , \35949 , \35953 );
and \U$35678 ( \35993 , \35953 , \35958 );
and \U$35679 ( \35994 , \35949 , \35958 );
or \U$35680 ( \35995 , \35992 , \35993 , \35994 );
xor \U$35681 ( \35996 , \35991 , \35995 );
and \U$35682 ( \35997 , \35934 , \35938 );
and \U$35683 ( \35998 , \35938 , \35943 );
and \U$35684 ( \35999 , \35934 , \35943 );
or \U$35685 ( \36000 , \35997 , \35998 , \35999 );
xor \U$35686 ( \36001 , \35996 , \36000 );
and \U$35687 ( \36002 , \35986 , \36001 );
and \U$35688 ( \36003 , \35906 , \36001 );
or \U$35689 ( \36004 , \35987 , \36002 , \36003 );
and \U$35690 ( \36005 , \22397 , \22076 );
and \U$35691 ( \36006 , \22361 , \22073 );
nor \U$35692 ( \36007 , \36005 , \36006 );
xnor \U$35693 ( \36008 , \36007 , \22072 );
and \U$35694 ( \36009 , \22418 , \22095 );
and \U$35695 ( \36010 , \22386 , \22093 );
nor \U$35696 ( \36011 , \36009 , \36010 );
xnor \U$35697 ( \36012 , \36011 , \22105 );
xor \U$35698 ( \36013 , \36008 , \36012 );
and \U$35699 ( \36014 , \22440 , \22119 );
and \U$35700 ( \36015 , \22407 , \22117 );
nor \U$35701 ( \36016 , \36014 , \36015 );
xnor \U$35702 ( \36017 , \36016 , \22129 );
xor \U$35703 ( \36018 , \36013 , \36017 );
and \U$35704 ( \36019 , \22603 , \22278 );
and \U$35705 ( \36020 , \22567 , \22276 );
nor \U$35706 ( \36021 , \36019 , \36020 );
xnor \U$35707 ( \36022 , \36021 , \22288 );
and \U$35708 ( \36023 , \22624 , \22300 );
and \U$35709 ( \36024 , \22592 , \22298 );
nor \U$35710 ( \36025 , \36023 , \36024 );
xnor \U$35711 ( \36026 , \36025 , \22310 );
xor \U$35712 ( \36027 , \36022 , \36026 );
and \U$35713 ( \36028 , \22646 , \22324 );
and \U$35714 ( \36029 , \22613 , \22322 );
nor \U$35715 ( \36030 , \36028 , \36029 );
xnor \U$35716 ( \36031 , \36030 , \22334 );
xor \U$35717 ( \36032 , \36027 , \36031 );
and \U$35718 ( \36033 , \22535 , \22208 );
and \U$35719 ( \36034 , \22500 , \22206 );
nor \U$35720 ( \36035 , \36033 , \36034 );
xnor \U$35721 ( \36036 , \36035 , \22218 );
and \U$35722 ( \36037 , \22556 , \22230 );
and \U$35723 ( \36038 , \22524 , \22228 );
nor \U$35724 ( \36039 , \36037 , \36038 );
xnor \U$35725 ( \36040 , \36039 , \22240 );
xor \U$35726 ( \36041 , \36036 , \36040 );
and \U$35727 ( \36042 , \22578 , \22257 );
and \U$35728 ( \36043 , \22545 , \22255 );
nor \U$35729 ( \36044 , \36042 , \36043 );
xnor \U$35730 ( \36045 , \36044 , \22267 );
xor \U$35731 ( \36046 , \36041 , \36045 );
xor \U$35732 ( \36047 , \36032 , \36046 );
and \U$35733 ( \36048 , \22468 , \22140 );
and \U$35734 ( \36049 , \22429 , \22138 );
nor \U$35735 ( \36050 , \36048 , \36049 );
xnor \U$35736 ( \36051 , \36050 , \22150 );
and \U$35737 ( \36052 , \22489 , \22162 );
and \U$35738 ( \36053 , \22457 , \22160 );
nor \U$35739 ( \36054 , \36052 , \36053 );
xnor \U$35740 ( \36055 , \36054 , \22172 );
xor \U$35741 ( \36056 , \36051 , \36055 );
and \U$35742 ( \36057 , \22511 , \22187 );
and \U$35743 ( \36058 , \22478 , \22185 );
nor \U$35744 ( \36059 , \36057 , \36058 );
xnor \U$35745 ( \36060 , \36059 , \22197 );
xor \U$35746 ( \36061 , \36056 , \36060 );
xor \U$35747 ( \36062 , \36047 , \36061 );
xor \U$35748 ( \36063 , \36018 , \36062 );
and \U$35749 ( \36064 , \35920 , \35924 );
and \U$35750 ( \36065 , \35924 , \35929 );
and \U$35751 ( \36066 , \35920 , \35929 );
or \U$35752 ( \36067 , \36064 , \36065 , \36066 );
and \U$35753 ( \36068 , \35972 , \35976 );
and \U$35754 ( \36069 , \35976 , \35981 );
and \U$35755 ( \36070 , \35972 , \35981 );
or \U$35756 ( \36071 , \36068 , \36069 , \36070 );
xor \U$35757 ( \36072 , \36067 , \36071 );
and \U$35758 ( \36073 , \22676 , \22345 );
and \U$35759 ( \36074 , \22635 , \22343 );
nor \U$35760 ( \36075 , \36073 , \36074 );
xnor \U$35761 ( \36076 , \36075 , \22355 );
and \U$35762 ( \36077 , \22696 , \22367 );
and \U$35763 ( \36078 , \22665 , \22365 );
nor \U$35764 ( \36079 , \36077 , \36078 );
xnor \U$35765 ( \36080 , \36079 , \22377 );
xor \U$35766 ( \36081 , \36076 , \36080 );
and \U$35767 ( \36082 , \22706 , \22392 );
and \U$35768 ( \36083 , \22686 , \22390 );
nor \U$35769 ( \36084 , \36082 , \36083 );
xnor \U$35770 ( \36085 , \36084 , \22402 );
xor \U$35771 ( \36086 , \36081 , \36085 );
xor \U$35772 ( \36087 , \36072 , \36086 );
xor \U$35773 ( \36088 , \36063 , \36087 );
and \U$35774 ( \36089 , \22418 , \22076 );
and \U$35775 ( \36090 , \22386 , \22073 );
nor \U$35776 ( \36091 , \36089 , \36090 );
xnor \U$35777 ( \36092 , \36091 , \22072 );
and \U$35778 ( \36093 , \22440 , \22095 );
and \U$35779 ( \36094 , \22407 , \22093 );
nor \U$35780 ( \36095 , \36093 , \36094 );
xnor \U$35781 ( \36096 , \36095 , \22105 );
and \U$35782 ( \36097 , \36092 , \36096 );
and \U$35783 ( \36098 , \22468 , \22119 );
and \U$35784 ( \36099 , \22429 , \22117 );
nor \U$35785 ( \36100 , \36098 , \36099 );
xnor \U$35786 ( \36101 , \36100 , \22129 );
and \U$35787 ( \36102 , \36096 , \36101 );
and \U$35788 ( \36103 , \36092 , \36101 );
or \U$35789 ( \36104 , \36097 , \36102 , \36103 );
and \U$35790 ( \36105 , \22489 , \22140 );
and \U$35791 ( \36106 , \22457 , \22138 );
nor \U$35792 ( \36107 , \36105 , \36106 );
xnor \U$35793 ( \36108 , \36107 , \22150 );
and \U$35794 ( \36109 , \22511 , \22162 );
and \U$35795 ( \36110 , \22478 , \22160 );
nor \U$35796 ( \36111 , \36109 , \36110 );
xnor \U$35797 ( \36112 , \36111 , \22172 );
and \U$35798 ( \36113 , \36108 , \36112 );
and \U$35799 ( \36114 , \22535 , \22187 );
and \U$35800 ( \36115 , \22500 , \22185 );
nor \U$35801 ( \36116 , \36114 , \36115 );
xnor \U$35802 ( \36117 , \36116 , \22197 );
and \U$35803 ( \36118 , \36112 , \36117 );
and \U$35804 ( \36119 , \36108 , \36117 );
or \U$35805 ( \36120 , \36113 , \36118 , \36119 );
and \U$35806 ( \36121 , \36104 , \36120 );
and \U$35807 ( \36122 , \35890 , \35894 );
and \U$35808 ( \36123 , \35894 , \35899 );
and \U$35809 ( \36124 , \35890 , \35899 );
or \U$35810 ( \36125 , \36122 , \36123 , \36124 );
and \U$35811 ( \36126 , \36120 , \36125 );
and \U$35812 ( \36127 , \36104 , \36125 );
or \U$35813 ( \36128 , \36121 , \36126 , \36127 );
and \U$35814 ( \36129 , \35965 , \35967 );
and \U$35815 ( \36130 , \35967 , \35982 );
and \U$35816 ( \36131 , \35965 , \35982 );
or \U$35817 ( \36132 , \36129 , \36130 , \36131 );
xor \U$35818 ( \36133 , \36128 , \36132 );
and \U$35819 ( \36134 , \35930 , \35944 );
and \U$35820 ( \36135 , \35944 , \35959 );
and \U$35821 ( \36136 , \35930 , \35959 );
or \U$35822 ( \36137 , \36134 , \36135 , \36136 );
xor \U$35823 ( \36138 , \36133 , \36137 );
and \U$35824 ( \36139 , \36088 , \36138 );
and \U$35825 ( \36140 , \36004 , \36139 );
and \U$35826 ( \36141 , \22478 , \22187 );
and \U$35827 ( \36142 , \22489 , \22185 );
nor \U$35828 ( \36143 , \36141 , \36142 );
xnor \U$35829 ( \36144 , \36143 , \22197 );
and \U$35830 ( \36145 , \22500 , \22208 );
and \U$35831 ( \36146 , \22511 , \22206 );
nor \U$35832 ( \36147 , \36145 , \36146 );
xnor \U$35833 ( \36148 , \36147 , \22218 );
xor \U$35834 ( \36149 , \36144 , \36148 );
and \U$35835 ( \36150 , \22524 , \22230 );
and \U$35836 ( \36151 , \22535 , \22228 );
nor \U$35837 ( \36152 , \36150 , \36151 );
xnor \U$35838 ( \36153 , \36152 , \22240 );
xor \U$35839 ( \36154 , \36149 , \36153 );
and \U$35840 ( \36155 , \22407 , \22119 );
and \U$35841 ( \36156 , \22418 , \22117 );
nor \U$35842 ( \36157 , \36155 , \36156 );
xnor \U$35843 ( \36158 , \36157 , \22129 );
and \U$35844 ( \36159 , \22429 , \22140 );
and \U$35845 ( \36160 , \22440 , \22138 );
nor \U$35846 ( \36161 , \36159 , \36160 );
xnor \U$35847 ( \36162 , \36161 , \22150 );
xor \U$35848 ( \36163 , \36158 , \36162 );
and \U$35849 ( \36164 , \22457 , \22162 );
and \U$35850 ( \36165 , \22468 , \22160 );
nor \U$35851 ( \36166 , \36164 , \36165 );
xnor \U$35852 ( \36167 , \36166 , \22172 );
xor \U$35853 ( \36168 , \36163 , \36167 );
xor \U$35854 ( \36169 , \36154 , \36168 );
and \U$35855 ( \36170 , \22361 , \22076 );
and \U$35856 ( \36171 , \22372 , \22073 );
nor \U$35857 ( \36172 , \36170 , \36171 );
xnor \U$35858 ( \36173 , \36172 , \22072 );
xor \U$35859 ( \36174 , \22423 , \36173 );
and \U$35860 ( \36175 , \22386 , \22095 );
and \U$35861 ( \36176 , \22397 , \22093 );
nor \U$35862 ( \36177 , \36175 , \36176 );
xnor \U$35863 ( \36178 , \36177 , \22105 );
xor \U$35864 ( \36179 , \36174 , \36178 );
xor \U$35865 ( \36180 , \36169 , \36179 );
nand \U$35866 ( \36181 , \22706 , \22411 );
xnor \U$35867 ( \36182 , \36181 , \22423 );
and \U$35868 ( \36183 , \22613 , \22324 );
and \U$35869 ( \36184 , \22624 , \22322 );
nor \U$35870 ( \36185 , \36183 , \36184 );
xnor \U$35871 ( \36186 , \36185 , \22334 );
and \U$35872 ( \36187 , \22635 , \22345 );
and \U$35873 ( \36188 , \22646 , \22343 );
nor \U$35874 ( \36189 , \36187 , \36188 );
xnor \U$35875 ( \36190 , \36189 , \22355 );
xor \U$35876 ( \36191 , \36186 , \36190 );
and \U$35877 ( \36192 , \22665 , \22367 );
and \U$35878 ( \36193 , \22676 , \22365 );
nor \U$35879 ( \36194 , \36192 , \36193 );
xnor \U$35880 ( \36195 , \36194 , \22377 );
xor \U$35881 ( \36196 , \36191 , \36195 );
xor \U$35882 ( \36197 , \36182 , \36196 );
and \U$35883 ( \36198 , \22545 , \22257 );
and \U$35884 ( \36199 , \22556 , \22255 );
nor \U$35885 ( \36200 , \36198 , \36199 );
xnor \U$35886 ( \36201 , \36200 , \22267 );
and \U$35887 ( \36202 , \22567 , \22278 );
and \U$35888 ( \36203 , \22578 , \22276 );
nor \U$35889 ( \36204 , \36202 , \36203 );
xnor \U$35890 ( \36205 , \36204 , \22288 );
xor \U$35891 ( \36206 , \36201 , \36205 );
and \U$35892 ( \36207 , \22592 , \22300 );
and \U$35893 ( \36208 , \22603 , \22298 );
nor \U$35894 ( \36209 , \36207 , \36208 );
xnor \U$35895 ( \36210 , \36209 , \22310 );
xor \U$35896 ( \36211 , \36206 , \36210 );
xor \U$35897 ( \36212 , \36197 , \36211 );
xor \U$35898 ( \36213 , \36180 , \36212 );
and \U$35899 ( \36214 , \36022 , \36026 );
and \U$35900 ( \36215 , \36026 , \36031 );
and \U$35901 ( \36216 , \36022 , \36031 );
or \U$35902 ( \36217 , \36214 , \36215 , \36216 );
and \U$35903 ( \36218 , \36076 , \36080 );
and \U$35904 ( \36219 , \36080 , \36085 );
and \U$35905 ( \36220 , \36076 , \36085 );
or \U$35906 ( \36221 , \36218 , \36219 , \36220 );
xor \U$35907 ( \36222 , \36217 , \36221 );
and \U$35908 ( \36223 , \22686 , \22392 );
and \U$35909 ( \36224 , \22696 , \22390 );
nor \U$35910 ( \36225 , \36223 , \36224 );
xnor \U$35911 ( \36226 , \36225 , \22402 );
xor \U$35912 ( \36227 , \36222 , \36226 );
xor \U$35913 ( \36228 , \36213 , \36227 );
and \U$35914 ( \36229 , \36139 , \36228 );
and \U$35915 ( \36230 , \36004 , \36228 );
or \U$35916 ( \36231 , \36140 , \36229 , \36230 );
and \U$35917 ( \36232 , \35991 , \35995 );
and \U$35918 ( \36233 , \35995 , \36000 );
and \U$35919 ( \36234 , \35991 , \36000 );
or \U$35920 ( \36235 , \36232 , \36233 , \36234 );
and \U$35921 ( \36236 , \36067 , \36071 );
and \U$35922 ( \36237 , \36071 , \36086 );
and \U$35923 ( \36238 , \36067 , \36086 );
or \U$35924 ( \36239 , \36236 , \36237 , \36238 );
xor \U$35925 ( \36240 , \36235 , \36239 );
and \U$35926 ( \36241 , \36032 , \36046 );
and \U$35927 ( \36242 , \36046 , \36061 );
and \U$35928 ( \36243 , \36032 , \36061 );
or \U$35929 ( \36244 , \36241 , \36242 , \36243 );
xor \U$35930 ( \36245 , \36240 , \36244 );
and \U$35931 ( \36246 , \36128 , \36132 );
and \U$35932 ( \36247 , \36132 , \36137 );
and \U$35933 ( \36248 , \36128 , \36137 );
or \U$35934 ( \36249 , \36246 , \36247 , \36248 );
and \U$35935 ( \36250 , \36018 , \36062 );
and \U$35936 ( \36251 , \36062 , \36087 );
and \U$35937 ( \36252 , \36018 , \36087 );
or \U$35938 ( \36253 , \36250 , \36251 , \36252 );
xor \U$35939 ( \36254 , \36249 , \36253 );
and \U$35940 ( \36255 , \36008 , \36012 );
and \U$35941 ( \36256 , \36012 , \36017 );
and \U$35942 ( \36257 , \36008 , \36017 );
or \U$35943 ( \36258 , \36255 , \36256 , \36257 );
and \U$35944 ( \36259 , \36051 , \36055 );
and \U$35945 ( \36260 , \36055 , \36060 );
and \U$35946 ( \36261 , \36051 , \36060 );
or \U$35947 ( \36262 , \36259 , \36260 , \36261 );
xor \U$35948 ( \36263 , \36258 , \36262 );
and \U$35949 ( \36264 , \36036 , \36040 );
and \U$35950 ( \36265 , \36040 , \36045 );
and \U$35951 ( \36266 , \36036 , \36045 );
or \U$35952 ( \36267 , \36264 , \36265 , \36266 );
xor \U$35953 ( \36268 , \36263 , \36267 );
xor \U$35954 ( \36269 , \36254 , \36268 );
and \U$35955 ( \36270 , \36245 , \36269 );
xor \U$35956 ( \36271 , \36231 , \36270 );
and \U$35957 ( \36272 , \36249 , \36253 );
and \U$35958 ( \36273 , \36253 , \36268 );
and \U$35959 ( \36274 , \36249 , \36268 );
or \U$35960 ( \36275 , \36272 , \36273 , \36274 );
and \U$35961 ( \36276 , \36154 , \36168 );
and \U$35962 ( \36277 , \36168 , \36179 );
and \U$35963 ( \36278 , \36154 , \36179 );
or \U$35964 ( \36279 , \36276 , \36277 , \36278 );
and \U$35965 ( \36280 , \22440 , \22140 );
and \U$35966 ( \36281 , \22407 , \22138 );
nor \U$35967 ( \36282 , \36280 , \36281 );
xnor \U$35968 ( \36283 , \36282 , \22150 );
and \U$35969 ( \36284 , \22468 , \22162 );
and \U$35970 ( \36285 , \22429 , \22160 );
nor \U$35971 ( \36286 , \36284 , \36285 );
xnor \U$35972 ( \36287 , \36286 , \22172 );
xor \U$35973 ( \36288 , \36283 , \36287 );
and \U$35974 ( \36289 , \22489 , \22187 );
and \U$35975 ( \36290 , \22457 , \22185 );
nor \U$35976 ( \36291 , \36289 , \36290 );
xnor \U$35977 ( \36292 , \36291 , \22197 );
xor \U$35978 ( \36293 , \36288 , \36292 );
xor \U$35979 ( \36294 , \36279 , \36293 );
and \U$35980 ( \36295 , \22372 , \22076 );
and \U$35981 ( \36296 , \22339 , \22073 );
nor \U$35982 ( \36297 , \36295 , \36296 );
xnor \U$35983 ( \36298 , \36297 , \22072 );
and \U$35984 ( \36299 , \22397 , \22095 );
and \U$35985 ( \36300 , \22361 , \22093 );
nor \U$35986 ( \36301 , \36299 , \36300 );
xnor \U$35987 ( \36302 , \36301 , \22105 );
xor \U$35988 ( \36303 , \36298 , \36302 );
and \U$35989 ( \36304 , \22418 , \22119 );
and \U$35990 ( \36305 , \22386 , \22117 );
nor \U$35991 ( \36306 , \36304 , \36305 );
xnor \U$35992 ( \36307 , \36306 , \22129 );
xor \U$35993 ( \36308 , \36303 , \36307 );
xor \U$35994 ( \36309 , \36294 , \36308 );
and \U$35995 ( \36310 , \36258 , \36262 );
and \U$35996 ( \36311 , \36262 , \36267 );
and \U$35997 ( \36312 , \36258 , \36267 );
or \U$35998 ( \36313 , \36310 , \36311 , \36312 );
and \U$35999 ( \36314 , \36217 , \36221 );
and \U$36000 ( \36315 , \36221 , \36226 );
and \U$36001 ( \36316 , \36217 , \36226 );
or \U$36002 ( \36317 , \36314 , \36315 , \36316 );
xor \U$36003 ( \36318 , \36313 , \36317 );
and \U$36004 ( \36319 , \36182 , \36196 );
and \U$36005 ( \36320 , \36196 , \36211 );
and \U$36006 ( \36321 , \36182 , \36211 );
or \U$36007 ( \36322 , \36319 , \36320 , \36321 );
xor \U$36008 ( \36323 , \36318 , \36322 );
xor \U$36009 ( \36324 , \36309 , \36323 );
xor \U$36010 ( \36325 , \36275 , \36324 );
and \U$36011 ( \36326 , \36235 , \36239 );
and \U$36012 ( \36327 , \36239 , \36244 );
and \U$36013 ( \36328 , \36235 , \36244 );
or \U$36014 ( \36329 , \36326 , \36327 , \36328 );
and \U$36015 ( \36330 , \36180 , \36212 );
and \U$36016 ( \36331 , \36212 , \36227 );
and \U$36017 ( \36332 , \36180 , \36227 );
or \U$36018 ( \36333 , \36330 , \36331 , \36332 );
xor \U$36019 ( \36334 , \36329 , \36333 );
and \U$36020 ( \36335 , \22646 , \22345 );
and \U$36021 ( \36336 , \22613 , \22343 );
nor \U$36022 ( \36337 , \36335 , \36336 );
xnor \U$36023 ( \36338 , \36337 , \22355 );
and \U$36024 ( \36339 , \22676 , \22367 );
and \U$36025 ( \36340 , \22635 , \22365 );
nor \U$36026 ( \36341 , \36339 , \36340 );
xnor \U$36027 ( \36342 , \36341 , \22377 );
xor \U$36028 ( \36343 , \36338 , \36342 );
and \U$36029 ( \36344 , \22696 , \22392 );
and \U$36030 ( \36345 , \22665 , \22390 );
nor \U$36031 ( \36346 , \36344 , \36345 );
xnor \U$36032 ( \36347 , \36346 , \22402 );
xor \U$36033 ( \36348 , \36343 , \36347 );
and \U$36034 ( \36349 , \22578 , \22278 );
and \U$36035 ( \36350 , \22545 , \22276 );
nor \U$36036 ( \36351 , \36349 , \36350 );
xnor \U$36037 ( \36352 , \36351 , \22288 );
and \U$36038 ( \36353 , \22603 , \22300 );
and \U$36039 ( \36354 , \22567 , \22298 );
nor \U$36040 ( \36355 , \36353 , \36354 );
xnor \U$36041 ( \36356 , \36355 , \22310 );
xor \U$36042 ( \36357 , \36352 , \36356 );
and \U$36043 ( \36358 , \22624 , \22324 );
and \U$36044 ( \36359 , \22592 , \22322 );
nor \U$36045 ( \36360 , \36358 , \36359 );
xnor \U$36046 ( \36361 , \36360 , \22334 );
xor \U$36047 ( \36362 , \36357 , \36361 );
xor \U$36048 ( \36363 , \36348 , \36362 );
and \U$36049 ( \36364 , \22511 , \22208 );
and \U$36050 ( \36365 , \22478 , \22206 );
nor \U$36051 ( \36366 , \36364 , \36365 );
xnor \U$36052 ( \36367 , \36366 , \22218 );
and \U$36053 ( \36368 , \22535 , \22230 );
and \U$36054 ( \36369 , \22500 , \22228 );
nor \U$36055 ( \36370 , \36368 , \36369 );
xnor \U$36056 ( \36371 , \36370 , \22240 );
xor \U$36057 ( \36372 , \36367 , \36371 );
and \U$36058 ( \36373 , \22556 , \22257 );
and \U$36059 ( \36374 , \22524 , \22255 );
nor \U$36060 ( \36375 , \36373 , \36374 );
xnor \U$36061 ( \36376 , \36375 , \22267 );
xor \U$36062 ( \36377 , \36372 , \36376 );
xor \U$36063 ( \36378 , \36363 , \36377 );
and \U$36064 ( \36379 , \36201 , \36205 );
and \U$36065 ( \36380 , \36205 , \36210 );
and \U$36066 ( \36381 , \36201 , \36210 );
or \U$36067 ( \36382 , \36379 , \36380 , \36381 );
and \U$36068 ( \36383 , \36186 , \36190 );
and \U$36069 ( \36384 , \36190 , \36195 );
and \U$36070 ( \36385 , \36186 , \36195 );
or \U$36071 ( \36386 , \36383 , \36384 , \36385 );
xor \U$36072 ( \36387 , \36382 , \36386 );
and \U$36073 ( \36388 , \22706 , \22413 );
and \U$36074 ( \36389 , \22686 , \22411 );
nor \U$36075 ( \36390 , \36388 , \36389 );
xnor \U$36076 ( \36391 , \36390 , \22423 );
xor \U$36077 ( \36392 , \36387 , \36391 );
xor \U$36078 ( \36393 , \36378 , \36392 );
and \U$36079 ( \36394 , \22423 , \36173 );
and \U$36080 ( \36395 , \36173 , \36178 );
and \U$36081 ( \36396 , \22423 , \36178 );
or \U$36082 ( \36397 , \36394 , \36395 , \36396 );
and \U$36083 ( \36398 , \36158 , \36162 );
and \U$36084 ( \36399 , \36162 , \36167 );
and \U$36085 ( \36400 , \36158 , \36167 );
or \U$36086 ( \36401 , \36398 , \36399 , \36400 );
xor \U$36087 ( \36402 , \36397 , \36401 );
and \U$36088 ( \36403 , \36144 , \36148 );
and \U$36089 ( \36404 , \36148 , \36153 );
and \U$36090 ( \36405 , \36144 , \36153 );
or \U$36091 ( \36406 , \36403 , \36404 , \36405 );
xor \U$36092 ( \36407 , \36402 , \36406 );
xor \U$36093 ( \36408 , \36393 , \36407 );
xor \U$36094 ( \36409 , \36334 , \36408 );
xor \U$36095 ( \36410 , \36325 , \36409 );
xor \U$36096 ( \36411 , \36271 , \36410 );
and \U$36097 ( \36412 , \22440 , \22076 );
and \U$36098 ( \36413 , \22407 , \22073 );
nor \U$36099 ( \36414 , \36412 , \36413 );
xnor \U$36100 ( \36415 , \36414 , \22072 );
and \U$36101 ( \36416 , \22468 , \22095 );
and \U$36102 ( \36417 , \22429 , \22093 );
nor \U$36103 ( \36418 , \36416 , \36417 );
xnor \U$36104 ( \36419 , \36418 , \22105 );
and \U$36105 ( \36420 , \36415 , \36419 );
and \U$36106 ( \36421 , \22489 , \22119 );
and \U$36107 ( \36422 , \22457 , \22117 );
nor \U$36108 ( \36423 , \36421 , \36422 );
xnor \U$36109 ( \36424 , \36423 , \22129 );
and \U$36110 ( \36425 , \36419 , \36424 );
and \U$36111 ( \36426 , \36415 , \36424 );
or \U$36112 ( \36427 , \36420 , \36425 , \36426 );
and \U$36113 ( \36428 , \22511 , \22140 );
and \U$36114 ( \36429 , \22478 , \22138 );
nor \U$36115 ( \36430 , \36428 , \36429 );
xnor \U$36116 ( \36431 , \36430 , \22150 );
and \U$36117 ( \36432 , \22535 , \22162 );
and \U$36118 ( \36433 , \22500 , \22160 );
nor \U$36119 ( \36434 , \36432 , \36433 );
xnor \U$36120 ( \36435 , \36434 , \22172 );
and \U$36121 ( \36436 , \36431 , \36435 );
and \U$36122 ( \36437 , \22556 , \22187 );
and \U$36123 ( \36438 , \22524 , \22185 );
nor \U$36124 ( \36439 , \36437 , \36438 );
xnor \U$36125 ( \36440 , \36439 , \22197 );
and \U$36126 ( \36441 , \36435 , \36440 );
and \U$36127 ( \36442 , \36431 , \36440 );
or \U$36128 ( \36443 , \36436 , \36441 , \36442 );
and \U$36129 ( \36444 , \36427 , \36443 );
and \U$36130 ( \36445 , \22578 , \22208 );
and \U$36131 ( \36446 , \22545 , \22206 );
nor \U$36132 ( \36447 , \36445 , \36446 );
xnor \U$36133 ( \36448 , \36447 , \22218 );
and \U$36134 ( \36449 , \22603 , \22230 );
and \U$36135 ( \36450 , \22567 , \22228 );
nor \U$36136 ( \36451 , \36449 , \36450 );
xnor \U$36137 ( \36452 , \36451 , \22240 );
and \U$36138 ( \36453 , \36448 , \36452 );
and \U$36139 ( \36454 , \22624 , \22257 );
and \U$36140 ( \36455 , \22592 , \22255 );
nor \U$36141 ( \36456 , \36454 , \36455 );
xnor \U$36142 ( \36457 , \36456 , \22267 );
and \U$36143 ( \36458 , \36452 , \36457 );
and \U$36144 ( \36459 , \36448 , \36457 );
or \U$36145 ( \36460 , \36453 , \36458 , \36459 );
and \U$36146 ( \36461 , \36443 , \36460 );
and \U$36147 ( \36462 , \36427 , \36460 );
or \U$36148 ( \36463 , \36444 , \36461 , \36462 );
and \U$36149 ( \36464 , \22646 , \22278 );
and \U$36150 ( \36465 , \22613 , \22276 );
nor \U$36151 ( \36466 , \36464 , \36465 );
xnor \U$36152 ( \36467 , \36466 , \22288 );
and \U$36153 ( \36468 , \22676 , \22300 );
and \U$36154 ( \36469 , \22635 , \22298 );
nor \U$36155 ( \36470 , \36468 , \36469 );
xnor \U$36156 ( \36471 , \36470 , \22310 );
and \U$36157 ( \36472 , \36467 , \36471 );
and \U$36158 ( \36473 , \22696 , \22324 );
and \U$36159 ( \36474 , \22665 , \22322 );
nor \U$36160 ( \36475 , \36473 , \36474 );
xnor \U$36161 ( \36476 , \36475 , \22334 );
and \U$36162 ( \36477 , \36471 , \36476 );
and \U$36163 ( \36478 , \36467 , \36476 );
or \U$36164 ( \36479 , \36472 , \36477 , \36478 );
xor \U$36165 ( \36480 , \35848 , \35852 );
xor \U$36166 ( \36481 , \36480 , \35855 );
and \U$36167 ( \36482 , \36479 , \36481 );
xor \U$36168 ( \36483 , \35832 , \35836 );
xor \U$36169 ( \36484 , \36483 , \35841 );
and \U$36170 ( \36485 , \36481 , \36484 );
and \U$36171 ( \36486 , \36479 , \36484 );
or \U$36172 ( \36487 , \36482 , \36485 , \36486 );
and \U$36173 ( \36488 , \36463 , \36487 );
xor \U$36174 ( \36489 , \35813 , \35817 );
xor \U$36175 ( \36490 , \36489 , \35822 );
xor \U$36176 ( \36491 , \35796 , \35800 );
xor \U$36177 ( \36492 , \36491 , \35805 );
and \U$36178 ( \36493 , \36490 , \36492 );
xor \U$36179 ( \36494 , \22377 , \35784 );
xor \U$36180 ( \36495 , \36494 , \35789 );
and \U$36181 ( \36496 , \36492 , \36495 );
and \U$36182 ( \36497 , \36490 , \36495 );
or \U$36183 ( \36498 , \36493 , \36496 , \36497 );
and \U$36184 ( \36499 , \36487 , \36498 );
and \U$36185 ( \36500 , \36463 , \36498 );
or \U$36186 ( \36501 , \36488 , \36499 , \36500 );
xor \U$36187 ( \36502 , \36108 , \36112 );
xor \U$36188 ( \36503 , \36502 , \36117 );
xor \U$36189 ( \36504 , \36092 , \36096 );
xor \U$36190 ( \36505 , \36504 , \36101 );
and \U$36191 ( \36506 , \36503 , \36505 );
xor \U$36192 ( \36507 , \35871 , \35885 );
xor \U$36193 ( \36508 , \36507 , \35900 );
and \U$36194 ( \36509 , \36505 , \36508 );
and \U$36195 ( \36510 , \36503 , \36508 );
or \U$36196 ( \36511 , \36506 , \36509 , \36510 );
and \U$36197 ( \36512 , \36501 , \36511 );
xor \U$36198 ( \36513 , \36104 , \36120 );
xor \U$36199 ( \36514 , \36513 , \36125 );
and \U$36200 ( \36515 , \36511 , \36514 );
and \U$36201 ( \36516 , \36501 , \36514 );
or \U$36202 ( \36517 , \36512 , \36515 , \36516 );
xor \U$36203 ( \36518 , \36088 , \36138 );
and \U$36204 ( \36519 , \36517 , \36518 );
xor \U$36205 ( \36520 , \35906 , \35986 );
xor \U$36206 ( \36521 , \36520 , \36001 );
and \U$36207 ( \36522 , \36518 , \36521 );
and \U$36208 ( \36523 , \36517 , \36521 );
or \U$36209 ( \36524 , \36519 , \36522 , \36523 );
xor \U$36210 ( \36525 , \36245 , \36269 );
and \U$36211 ( \36526 , \36524 , \36525 );
xor \U$36212 ( \36527 , \36004 , \36139 );
xor \U$36213 ( \36528 , \36527 , \36228 );
and \U$36214 ( \36529 , \36525 , \36528 );
and \U$36215 ( \36530 , \36524 , \36528 );
or \U$36216 ( \36531 , \36526 , \36529 , \36530 );
nor \U$36217 ( \36532 , \36411 , \36531 );
and \U$36218 ( \36533 , \36275 , \36324 );
and \U$36219 ( \36534 , \36324 , \36409 );
and \U$36220 ( \36535 , \36275 , \36409 );
or \U$36221 ( \36536 , \36533 , \36534 , \36535 );
and \U$36222 ( \36537 , \36313 , \36317 );
and \U$36223 ( \36538 , \36317 , \36322 );
and \U$36224 ( \36539 , \36313 , \36322 );
or \U$36225 ( \36540 , \36537 , \36538 , \36539 );
and \U$36226 ( \36541 , \36279 , \36293 );
and \U$36227 ( \36542 , \36293 , \36308 );
and \U$36228 ( \36543 , \36279 , \36308 );
or \U$36229 ( \36544 , \36541 , \36542 , \36543 );
xor \U$36230 ( \36545 , \36540 , \36544 );
and \U$36231 ( \36546 , \36378 , \36392 );
and \U$36232 ( \36547 , \36392 , \36407 );
and \U$36233 ( \36548 , \36378 , \36407 );
or \U$36234 ( \36549 , \36546 , \36547 , \36548 );
xor \U$36235 ( \36550 , \36545 , \36549 );
xor \U$36236 ( \36551 , \36536 , \36550 );
and \U$36237 ( \36552 , \36329 , \36333 );
and \U$36238 ( \36553 , \36333 , \36408 );
and \U$36239 ( \36554 , \36329 , \36408 );
or \U$36240 ( \36555 , \36552 , \36553 , \36554 );
and \U$36241 ( \36556 , \36309 , \36323 );
xor \U$36242 ( \36557 , \36555 , \36556 );
and \U$36243 ( \36558 , \36352 , \36356 );
and \U$36244 ( \36559 , \36356 , \36361 );
and \U$36245 ( \36560 , \36352 , \36361 );
or \U$36246 ( \36561 , \36558 , \36559 , \36560 );
and \U$36247 ( \36562 , \36338 , \36342 );
and \U$36248 ( \36563 , \36342 , \36347 );
and \U$36249 ( \36564 , \36338 , \36347 );
or \U$36250 ( \36565 , \36562 , \36563 , \36564 );
xor \U$36251 ( \36566 , \36561 , \36565 );
and \U$36252 ( \36567 , \22665 , \22392 );
and \U$36253 ( \36568 , \22676 , \22390 );
nor \U$36254 ( \36569 , \36567 , \36568 );
xnor \U$36255 ( \36570 , \36569 , \22402 );
and \U$36256 ( \36571 , \22686 , \22413 );
and \U$36257 ( \36572 , \22696 , \22411 );
nor \U$36258 ( \36573 , \36571 , \36572 );
xnor \U$36259 ( \36574 , \36573 , \22423 );
xor \U$36260 ( \36575 , \36570 , \36574 );
nand \U$36261 ( \36576 , \22706 , \22433 );
xnor \U$36262 ( \36577 , \36576 , \22445 );
xor \U$36263 ( \36578 , \36575 , \36577 );
xor \U$36264 ( \36579 , \36566 , \36578 );
and \U$36265 ( \36580 , \36298 , \36302 );
and \U$36266 ( \36581 , \36302 , \36307 );
and \U$36267 ( \36582 , \36298 , \36307 );
or \U$36268 ( \36583 , \36580 , \36581 , \36582 );
and \U$36269 ( \36584 , \36283 , \36287 );
and \U$36270 ( \36585 , \36287 , \36292 );
and \U$36271 ( \36586 , \36283 , \36292 );
or \U$36272 ( \36587 , \36584 , \36585 , \36586 );
xor \U$36273 ( \36588 , \36583 , \36587 );
and \U$36274 ( \36589 , \36367 , \36371 );
and \U$36275 ( \36590 , \36371 , \36376 );
and \U$36276 ( \36591 , \36367 , \36376 );
or \U$36277 ( \36592 , \36589 , \36590 , \36591 );
xor \U$36278 ( \36593 , \36588 , \36592 );
xor \U$36279 ( \36594 , \36579 , \36593 );
and \U$36280 ( \36595 , \22386 , \22119 );
and \U$36281 ( \36596 , \22397 , \22117 );
nor \U$36282 ( \36597 , \36595 , \36596 );
xnor \U$36283 ( \36598 , \36597 , \22129 );
and \U$36284 ( \36599 , \22407 , \22140 );
and \U$36285 ( \36600 , \22418 , \22138 );
nor \U$36286 ( \36601 , \36599 , \36600 );
xnor \U$36287 ( \36602 , \36601 , \22150 );
xor \U$36288 ( \36603 , \36598 , \36602 );
and \U$36289 ( \36604 , \22429 , \22162 );
and \U$36290 ( \36605 , \22440 , \22160 );
nor \U$36291 ( \36606 , \36604 , \36605 );
xnor \U$36292 ( \36607 , \36606 , \22172 );
xor \U$36293 ( \36608 , \36603 , \36607 );
and \U$36294 ( \36609 , \22339 , \22076 );
and \U$36295 ( \36610 , \22350 , \22073 );
nor \U$36296 ( \36611 , \36609 , \36610 );
xnor \U$36297 ( \36612 , \36611 , \22072 );
xor \U$36298 ( \36613 , \22445 , \36612 );
and \U$36299 ( \36614 , \22361 , \22095 );
and \U$36300 ( \36615 , \22372 , \22093 );
nor \U$36301 ( \36616 , \36614 , \36615 );
xnor \U$36302 ( \36617 , \36616 , \22105 );
xor \U$36303 ( \36618 , \36613 , \36617 );
xor \U$36304 ( \36619 , \36608 , \36618 );
and \U$36305 ( \36620 , \22592 , \22324 );
and \U$36306 ( \36621 , \22603 , \22322 );
nor \U$36307 ( \36622 , \36620 , \36621 );
xnor \U$36308 ( \36623 , \36622 , \22334 );
and \U$36309 ( \36624 , \22613 , \22345 );
and \U$36310 ( \36625 , \22624 , \22343 );
nor \U$36311 ( \36626 , \36624 , \36625 );
xnor \U$36312 ( \36627 , \36626 , \22355 );
xor \U$36313 ( \36628 , \36623 , \36627 );
and \U$36314 ( \36629 , \22635 , \22367 );
and \U$36315 ( \36630 , \22646 , \22365 );
nor \U$36316 ( \36631 , \36629 , \36630 );
xnor \U$36317 ( \36632 , \36631 , \22377 );
xor \U$36318 ( \36633 , \36628 , \36632 );
and \U$36319 ( \36634 , \22524 , \22257 );
and \U$36320 ( \36635 , \22535 , \22255 );
nor \U$36321 ( \36636 , \36634 , \36635 );
xnor \U$36322 ( \36637 , \36636 , \22267 );
and \U$36323 ( \36638 , \22545 , \22278 );
and \U$36324 ( \36639 , \22556 , \22276 );
nor \U$36325 ( \36640 , \36638 , \36639 );
xnor \U$36326 ( \36641 , \36640 , \22288 );
xor \U$36327 ( \36642 , \36637 , \36641 );
and \U$36328 ( \36643 , \22567 , \22300 );
and \U$36329 ( \36644 , \22578 , \22298 );
nor \U$36330 ( \36645 , \36643 , \36644 );
xnor \U$36331 ( \36646 , \36645 , \22310 );
xor \U$36332 ( \36647 , \36642 , \36646 );
xor \U$36333 ( \36648 , \36633 , \36647 );
and \U$36334 ( \36649 , \22457 , \22187 );
and \U$36335 ( \36650 , \22468 , \22185 );
nor \U$36336 ( \36651 , \36649 , \36650 );
xnor \U$36337 ( \36652 , \36651 , \22197 );
and \U$36338 ( \36653 , \22478 , \22208 );
and \U$36339 ( \36654 , \22489 , \22206 );
nor \U$36340 ( \36655 , \36653 , \36654 );
xnor \U$36341 ( \36656 , \36655 , \22218 );
xor \U$36342 ( \36657 , \36652 , \36656 );
and \U$36343 ( \36658 , \22500 , \22230 );
and \U$36344 ( \36659 , \22511 , \22228 );
nor \U$36345 ( \36660 , \36658 , \36659 );
xnor \U$36346 ( \36661 , \36660 , \22240 );
xor \U$36347 ( \36662 , \36657 , \36661 );
xor \U$36348 ( \36663 , \36648 , \36662 );
xor \U$36349 ( \36664 , \36619 , \36663 );
xor \U$36350 ( \36665 , \36594 , \36664 );
and \U$36351 ( \36666 , \36397 , \36401 );
and \U$36352 ( \36667 , \36401 , \36406 );
and \U$36353 ( \36668 , \36397 , \36406 );
or \U$36354 ( \36669 , \36666 , \36667 , \36668 );
and \U$36355 ( \36670 , \36382 , \36386 );
and \U$36356 ( \36671 , \36386 , \36391 );
and \U$36357 ( \36672 , \36382 , \36391 );
or \U$36358 ( \36673 , \36670 , \36671 , \36672 );
xor \U$36359 ( \36674 , \36669 , \36673 );
and \U$36360 ( \36675 , \36348 , \36362 );
and \U$36361 ( \36676 , \36362 , \36377 );
and \U$36362 ( \36677 , \36348 , \36377 );
or \U$36363 ( \36678 , \36675 , \36676 , \36677 );
xor \U$36364 ( \36679 , \36674 , \36678 );
xor \U$36365 ( \36680 , \36665 , \36679 );
xor \U$36366 ( \36681 , \36557 , \36680 );
xor \U$36367 ( \36682 , \36551 , \36681 );
and \U$36368 ( \36683 , \36231 , \36270 );
and \U$36369 ( \36684 , \36270 , \36410 );
and \U$36370 ( \36685 , \36231 , \36410 );
or \U$36371 ( \36686 , \36683 , \36684 , \36685 );
nor \U$36372 ( \36687 , \36682 , \36686 );
nor \U$36373 ( \36688 , \36532 , \36687 );
and \U$36374 ( \36689 , \36555 , \36556 );
and \U$36375 ( \36690 , \36556 , \36680 );
and \U$36376 ( \36691 , \36555 , \36680 );
or \U$36377 ( \36692 , \36689 , \36690 , \36691 );
and \U$36378 ( \36693 , \36669 , \36673 );
and \U$36379 ( \36694 , \36673 , \36678 );
and \U$36380 ( \36695 , \36669 , \36678 );
or \U$36381 ( \36696 , \36693 , \36694 , \36695 );
and \U$36382 ( \36697 , \36608 , \36618 );
and \U$36383 ( \36698 , \36618 , \36663 );
and \U$36384 ( \36699 , \36608 , \36663 );
or \U$36385 ( \36700 , \36697 , \36698 , \36699 );
xor \U$36386 ( \36701 , \36696 , \36700 );
and \U$36387 ( \36702 , \36579 , \36593 );
xor \U$36388 ( \36703 , \36701 , \36702 );
xor \U$36389 ( \36704 , \36692 , \36703 );
and \U$36390 ( \36705 , \36540 , \36544 );
and \U$36391 ( \36706 , \36544 , \36549 );
and \U$36392 ( \36707 , \36540 , \36549 );
or \U$36393 ( \36708 , \36705 , \36706 , \36707 );
and \U$36394 ( \36709 , \36594 , \36664 );
and \U$36395 ( \36710 , \36664 , \36679 );
and \U$36396 ( \36711 , \36594 , \36679 );
or \U$36397 ( \36712 , \36709 , \36710 , \36711 );
xor \U$36398 ( \36713 , \36708 , \36712 );
and \U$36399 ( \36714 , \22445 , \36612 );
and \U$36400 ( \36715 , \36612 , \36617 );
and \U$36401 ( \36716 , \22445 , \36617 );
or \U$36402 ( \36717 , \36714 , \36715 , \36716 );
and \U$36403 ( \36718 , \36598 , \36602 );
and \U$36404 ( \36719 , \36602 , \36607 );
and \U$36405 ( \36720 , \36598 , \36607 );
or \U$36406 ( \36721 , \36718 , \36719 , \36720 );
xor \U$36407 ( \36722 , \36717 , \36721 );
and \U$36408 ( \36723 , \36652 , \36656 );
and \U$36409 ( \36724 , \36656 , \36661 );
and \U$36410 ( \36725 , \36652 , \36661 );
or \U$36411 ( \36726 , \36723 , \36724 , \36725 );
xor \U$36412 ( \36727 , \36722 , \36726 );
and \U$36413 ( \36728 , \22489 , \22208 );
and \U$36414 ( \36729 , \22457 , \22206 );
nor \U$36415 ( \36730 , \36728 , \36729 );
xnor \U$36416 ( \36731 , \36730 , \22218 );
and \U$36417 ( \36732 , \22511 , \22230 );
and \U$36418 ( \36733 , \22478 , \22228 );
nor \U$36419 ( \36734 , \36732 , \36733 );
xnor \U$36420 ( \36735 , \36734 , \22240 );
xor \U$36421 ( \36736 , \36731 , \36735 );
and \U$36422 ( \36737 , \22535 , \22257 );
and \U$36423 ( \36738 , \22500 , \22255 );
nor \U$36424 ( \36739 , \36737 , \36738 );
xnor \U$36425 ( \36740 , \36739 , \22267 );
xor \U$36426 ( \36741 , \36736 , \36740 );
and \U$36427 ( \36742 , \22418 , \22140 );
and \U$36428 ( \36743 , \22386 , \22138 );
nor \U$36429 ( \36744 , \36742 , \36743 );
xnor \U$36430 ( \36745 , \36744 , \22150 );
and \U$36431 ( \36746 , \22440 , \22162 );
and \U$36432 ( \36747 , \22407 , \22160 );
nor \U$36433 ( \36748 , \36746 , \36747 );
xnor \U$36434 ( \36749 , \36748 , \22172 );
xor \U$36435 ( \36750 , \36745 , \36749 );
and \U$36436 ( \36751 , \22468 , \22187 );
and \U$36437 ( \36752 , \22429 , \22185 );
nor \U$36438 ( \36753 , \36751 , \36752 );
xnor \U$36439 ( \36754 , \36753 , \22197 );
xor \U$36440 ( \36755 , \36750 , \36754 );
xor \U$36441 ( \36756 , \36741 , \36755 );
and \U$36442 ( \36757 , \22350 , \22076 );
and \U$36443 ( \36758 , \22318 , \22073 );
nor \U$36444 ( \36759 , \36757 , \36758 );
xnor \U$36445 ( \36760 , \36759 , \22072 );
and \U$36446 ( \36761 , \22372 , \22095 );
and \U$36447 ( \36762 , \22339 , \22093 );
nor \U$36448 ( \36763 , \36761 , \36762 );
xnor \U$36449 ( \36764 , \36763 , \22105 );
xor \U$36450 ( \36765 , \36760 , \36764 );
and \U$36451 ( \36766 , \22397 , \22119 );
and \U$36452 ( \36767 , \22361 , \22117 );
nor \U$36453 ( \36768 , \36766 , \36767 );
xnor \U$36454 ( \36769 , \36768 , \22129 );
xor \U$36455 ( \36770 , \36765 , \36769 );
xor \U$36456 ( \36771 , \36756 , \36770 );
and \U$36457 ( \36772 , \22696 , \22413 );
and \U$36458 ( \36773 , \22665 , \22411 );
nor \U$36459 ( \36774 , \36772 , \36773 );
xnor \U$36460 ( \36775 , \36774 , \22423 );
and \U$36461 ( \36776 , \22706 , \22435 );
and \U$36462 ( \36777 , \22686 , \22433 );
nor \U$36463 ( \36778 , \36776 , \36777 );
xnor \U$36464 ( \36779 , \36778 , \22445 );
xor \U$36465 ( \36780 , \36775 , \36779 );
and \U$36466 ( \36781 , \22624 , \22345 );
and \U$36467 ( \36782 , \22592 , \22343 );
nor \U$36468 ( \36783 , \36781 , \36782 );
xnor \U$36469 ( \36784 , \36783 , \22355 );
and \U$36470 ( \36785 , \22646 , \22367 );
and \U$36471 ( \36786 , \22613 , \22365 );
nor \U$36472 ( \36787 , \36785 , \36786 );
xnor \U$36473 ( \36788 , \36787 , \22377 );
xor \U$36474 ( \36789 , \36784 , \36788 );
and \U$36475 ( \36790 , \22676 , \22392 );
and \U$36476 ( \36791 , \22635 , \22390 );
nor \U$36477 ( \36792 , \36790 , \36791 );
xnor \U$36478 ( \36793 , \36792 , \22402 );
xor \U$36479 ( \36794 , \36789 , \36793 );
xor \U$36480 ( \36795 , \36780 , \36794 );
and \U$36481 ( \36796 , \22556 , \22278 );
and \U$36482 ( \36797 , \22524 , \22276 );
nor \U$36483 ( \36798 , \36796 , \36797 );
xnor \U$36484 ( \36799 , \36798 , \22288 );
and \U$36485 ( \36800 , \22578 , \22300 );
and \U$36486 ( \36801 , \22545 , \22298 );
nor \U$36487 ( \36802 , \36800 , \36801 );
xnor \U$36488 ( \36803 , \36802 , \22310 );
xor \U$36489 ( \36804 , \36799 , \36803 );
and \U$36490 ( \36805 , \22603 , \22324 );
and \U$36491 ( \36806 , \22567 , \22322 );
nor \U$36492 ( \36807 , \36805 , \36806 );
xnor \U$36493 ( \36808 , \36807 , \22334 );
xor \U$36494 ( \36809 , \36804 , \36808 );
xor \U$36495 ( \36810 , \36795 , \36809 );
xor \U$36496 ( \36811 , \36771 , \36810 );
and \U$36497 ( \36812 , \36637 , \36641 );
and \U$36498 ( \36813 , \36641 , \36646 );
and \U$36499 ( \36814 , \36637 , \36646 );
or \U$36500 ( \36815 , \36812 , \36813 , \36814 );
and \U$36501 ( \36816 , \36623 , \36627 );
and \U$36502 ( \36817 , \36627 , \36632 );
and \U$36503 ( \36818 , \36623 , \36632 );
or \U$36504 ( \36819 , \36816 , \36817 , \36818 );
xor \U$36505 ( \36820 , \36815 , \36819 );
and \U$36506 ( \36821 , \36570 , \36574 );
and \U$36507 ( \36822 , \36574 , \36577 );
and \U$36508 ( \36823 , \36570 , \36577 );
or \U$36509 ( \36824 , \36821 , \36822 , \36823 );
xor \U$36510 ( \36825 , \36820 , \36824 );
xor \U$36511 ( \36826 , \36811 , \36825 );
xor \U$36512 ( \36827 , \36727 , \36826 );
and \U$36513 ( \36828 , \36583 , \36587 );
and \U$36514 ( \36829 , \36587 , \36592 );
and \U$36515 ( \36830 , \36583 , \36592 );
or \U$36516 ( \36831 , \36828 , \36829 , \36830 );
and \U$36517 ( \36832 , \36561 , \36565 );
and \U$36518 ( \36833 , \36565 , \36578 );
and \U$36519 ( \36834 , \36561 , \36578 );
or \U$36520 ( \36835 , \36832 , \36833 , \36834 );
xor \U$36521 ( \36836 , \36831 , \36835 );
and \U$36522 ( \36837 , \36633 , \36647 );
and \U$36523 ( \36838 , \36647 , \36662 );
and \U$36524 ( \36839 , \36633 , \36662 );
or \U$36525 ( \36840 , \36837 , \36838 , \36839 );
xor \U$36526 ( \36841 , \36836 , \36840 );
xor \U$36527 ( \36842 , \36827 , \36841 );
xor \U$36528 ( \36843 , \36713 , \36842 );
xor \U$36529 ( \36844 , \36704 , \36843 );
and \U$36530 ( \36845 , \36536 , \36550 );
and \U$36531 ( \36846 , \36550 , \36681 );
and \U$36532 ( \36847 , \36536 , \36681 );
or \U$36533 ( \36848 , \36845 , \36846 , \36847 );
nor \U$36534 ( \36849 , \36844 , \36848 );
and \U$36535 ( \36850 , \36708 , \36712 );
and \U$36536 ( \36851 , \36712 , \36842 );
and \U$36537 ( \36852 , \36708 , \36842 );
or \U$36538 ( \36853 , \36850 , \36851 , \36852 );
and \U$36539 ( \36854 , \36717 , \36721 );
and \U$36540 ( \36855 , \36721 , \36726 );
and \U$36541 ( \36856 , \36717 , \36726 );
or \U$36542 ( \36857 , \36854 , \36855 , \36856 );
and \U$36543 ( \36858 , \36815 , \36819 );
and \U$36544 ( \36859 , \36819 , \36824 );
and \U$36545 ( \36860 , \36815 , \36824 );
or \U$36546 ( \36861 , \36858 , \36859 , \36860 );
xor \U$36547 ( \36862 , \36857 , \36861 );
and \U$36548 ( \36863 , \36780 , \36794 );
and \U$36549 ( \36864 , \36794 , \36809 );
and \U$36550 ( \36865 , \36780 , \36809 );
or \U$36551 ( \36866 , \36863 , \36864 , \36865 );
xor \U$36552 ( \36867 , \36862 , \36866 );
and \U$36553 ( \36868 , \36831 , \36835 );
and \U$36554 ( \36869 , \36835 , \36840 );
and \U$36555 ( \36870 , \36831 , \36840 );
or \U$36556 ( \36871 , \36868 , \36869 , \36870 );
and \U$36557 ( \36872 , \36771 , \36810 );
and \U$36558 ( \36873 , \36810 , \36825 );
and \U$36559 ( \36874 , \36771 , \36825 );
or \U$36560 ( \36875 , \36872 , \36873 , \36874 );
xor \U$36561 ( \36876 , \36871 , \36875 );
nand \U$36562 ( \36877 , \22706 , \22461 );
xnor \U$36563 ( \36878 , \36877 , \22473 );
and \U$36564 ( \36879 , \22635 , \22392 );
and \U$36565 ( \36880 , \22646 , \22390 );
nor \U$36566 ( \36881 , \36879 , \36880 );
xnor \U$36567 ( \36882 , \36881 , \22402 );
and \U$36568 ( \36883 , \22665 , \22413 );
and \U$36569 ( \36884 , \22676 , \22411 );
nor \U$36570 ( \36885 , \36883 , \36884 );
xnor \U$36571 ( \36886 , \36885 , \22423 );
xor \U$36572 ( \36887 , \36882 , \36886 );
and \U$36573 ( \36888 , \22686 , \22435 );
and \U$36574 ( \36889 , \22696 , \22433 );
nor \U$36575 ( \36890 , \36888 , \36889 );
xnor \U$36576 ( \36891 , \36890 , \22445 );
xor \U$36577 ( \36892 , \36887 , \36891 );
xor \U$36578 ( \36893 , \36878 , \36892 );
and \U$36579 ( \36894 , \22567 , \22324 );
and \U$36580 ( \36895 , \22578 , \22322 );
nor \U$36581 ( \36896 , \36894 , \36895 );
xnor \U$36582 ( \36897 , \36896 , \22334 );
and \U$36583 ( \36898 , \22592 , \22345 );
and \U$36584 ( \36899 , \22603 , \22343 );
nor \U$36585 ( \36900 , \36898 , \36899 );
xnor \U$36586 ( \36901 , \36900 , \22355 );
xor \U$36587 ( \36902 , \36897 , \36901 );
and \U$36588 ( \36903 , \22613 , \22367 );
and \U$36589 ( \36904 , \22624 , \22365 );
nor \U$36590 ( \36905 , \36903 , \36904 );
xnor \U$36591 ( \36906 , \36905 , \22377 );
xor \U$36592 ( \36907 , \36902 , \36906 );
xor \U$36593 ( \36908 , \36893 , \36907 );
and \U$36594 ( \36909 , \36799 , \36803 );
and \U$36595 ( \36910 , \36803 , \36808 );
and \U$36596 ( \36911 , \36799 , \36808 );
or \U$36597 ( \36912 , \36909 , \36910 , \36911 );
and \U$36598 ( \36913 , \36784 , \36788 );
and \U$36599 ( \36914 , \36788 , \36793 );
and \U$36600 ( \36915 , \36784 , \36793 );
or \U$36601 ( \36916 , \36913 , \36914 , \36915 );
xor \U$36602 ( \36917 , \36912 , \36916 );
and \U$36603 ( \36918 , \36775 , \36779 );
xor \U$36604 ( \36919 , \36917 , \36918 );
xor \U$36605 ( \36920 , \36908 , \36919 );
and \U$36606 ( \36921 , \36760 , \36764 );
and \U$36607 ( \36922 , \36764 , \36769 );
and \U$36608 ( \36923 , \36760 , \36769 );
or \U$36609 ( \36924 , \36921 , \36922 , \36923 );
and \U$36610 ( \36925 , \36745 , \36749 );
and \U$36611 ( \36926 , \36749 , \36754 );
and \U$36612 ( \36927 , \36745 , \36754 );
or \U$36613 ( \36928 , \36925 , \36926 , \36927 );
xor \U$36614 ( \36929 , \36924 , \36928 );
and \U$36615 ( \36930 , \36731 , \36735 );
and \U$36616 ( \36931 , \36735 , \36740 );
and \U$36617 ( \36932 , \36731 , \36740 );
or \U$36618 ( \36933 , \36930 , \36931 , \36932 );
xor \U$36619 ( \36934 , \36929 , \36933 );
xor \U$36620 ( \36935 , \36920 , \36934 );
xor \U$36621 ( \36936 , \36876 , \36935 );
xor \U$36622 ( \36937 , \36867 , \36936 );
xor \U$36623 ( \36938 , \36853 , \36937 );
and \U$36624 ( \36939 , \36696 , \36700 );
and \U$36625 ( \36940 , \36700 , \36702 );
and \U$36626 ( \36941 , \36696 , \36702 );
or \U$36627 ( \36942 , \36939 , \36940 , \36941 );
and \U$36628 ( \36943 , \36727 , \36826 );
and \U$36629 ( \36944 , \36826 , \36841 );
and \U$36630 ( \36945 , \36727 , \36841 );
or \U$36631 ( \36946 , \36943 , \36944 , \36945 );
xor \U$36632 ( \36947 , \36942 , \36946 );
and \U$36633 ( \36948 , \36741 , \36755 );
and \U$36634 ( \36949 , \36755 , \36770 );
and \U$36635 ( \36950 , \36741 , \36770 );
or \U$36636 ( \36951 , \36948 , \36949 , \36950 );
and \U$36637 ( \36952 , \22318 , \22076 );
and \U$36638 ( \36953 , \22329 , \22073 );
nor \U$36639 ( \36954 , \36952 , \36953 );
xnor \U$36640 ( \36955 , \36954 , \22072 );
xor \U$36641 ( \36956 , \22473 , \36955 );
and \U$36642 ( \36957 , \22339 , \22095 );
and \U$36643 ( \36958 , \22350 , \22093 );
nor \U$36644 ( \36959 , \36957 , \36958 );
xnor \U$36645 ( \36960 , \36959 , \22105 );
xor \U$36646 ( \36961 , \36956 , \36960 );
xor \U$36647 ( \36962 , \36951 , \36961 );
and \U$36648 ( \36963 , \22500 , \22257 );
and \U$36649 ( \36964 , \22511 , \22255 );
nor \U$36650 ( \36965 , \36963 , \36964 );
xnor \U$36651 ( \36966 , \36965 , \22267 );
and \U$36652 ( \36967 , \22524 , \22278 );
and \U$36653 ( \36968 , \22535 , \22276 );
nor \U$36654 ( \36969 , \36967 , \36968 );
xnor \U$36655 ( \36970 , \36969 , \22288 );
xor \U$36656 ( \36971 , \36966 , \36970 );
and \U$36657 ( \36972 , \22545 , \22300 );
and \U$36658 ( \36973 , \22556 , \22298 );
nor \U$36659 ( \36974 , \36972 , \36973 );
xnor \U$36660 ( \36975 , \36974 , \22310 );
xor \U$36661 ( \36976 , \36971 , \36975 );
and \U$36662 ( \36977 , \22429 , \22187 );
and \U$36663 ( \36978 , \22440 , \22185 );
nor \U$36664 ( \36979 , \36977 , \36978 );
xnor \U$36665 ( \36980 , \36979 , \22197 );
and \U$36666 ( \36981 , \22457 , \22208 );
and \U$36667 ( \36982 , \22468 , \22206 );
nor \U$36668 ( \36983 , \36981 , \36982 );
xnor \U$36669 ( \36984 , \36983 , \22218 );
xor \U$36670 ( \36985 , \36980 , \36984 );
and \U$36671 ( \36986 , \22478 , \22230 );
and \U$36672 ( \36987 , \22489 , \22228 );
nor \U$36673 ( \36988 , \36986 , \36987 );
xnor \U$36674 ( \36989 , \36988 , \22240 );
xor \U$36675 ( \36990 , \36985 , \36989 );
xor \U$36676 ( \36991 , \36976 , \36990 );
and \U$36677 ( \36992 , \22361 , \22119 );
and \U$36678 ( \36993 , \22372 , \22117 );
nor \U$36679 ( \36994 , \36992 , \36993 );
xnor \U$36680 ( \36995 , \36994 , \22129 );
and \U$36681 ( \36996 , \22386 , \22140 );
and \U$36682 ( \36997 , \22397 , \22138 );
nor \U$36683 ( \36998 , \36996 , \36997 );
xnor \U$36684 ( \36999 , \36998 , \22150 );
xor \U$36685 ( \37000 , \36995 , \36999 );
and \U$36686 ( \37001 , \22407 , \22162 );
and \U$36687 ( \37002 , \22418 , \22160 );
nor \U$36688 ( \37003 , \37001 , \37002 );
xnor \U$36689 ( \37004 , \37003 , \22172 );
xor \U$36690 ( \37005 , \37000 , \37004 );
xor \U$36691 ( \37006 , \36991 , \37005 );
xor \U$36692 ( \37007 , \36962 , \37006 );
xor \U$36693 ( \37008 , \36947 , \37007 );
xor \U$36694 ( \37009 , \36938 , \37008 );
and \U$36695 ( \37010 , \36692 , \36703 );
and \U$36696 ( \37011 , \36703 , \36843 );
and \U$36697 ( \37012 , \36692 , \36843 );
or \U$36698 ( \37013 , \37010 , \37011 , \37012 );
nor \U$36699 ( \37014 , \37009 , \37013 );
nor \U$36700 ( \37015 , \36849 , \37014 );
nand \U$36701 ( \37016 , \36688 , \37015 );
and \U$36702 ( \37017 , \36942 , \36946 );
and \U$36703 ( \37018 , \36946 , \37007 );
and \U$36704 ( \37019 , \36942 , \37007 );
or \U$36705 ( \37020 , \37017 , \37018 , \37019 );
and \U$36706 ( \37021 , \36867 , \36936 );
xor \U$36707 ( \37022 , \37020 , \37021 );
and \U$36708 ( \37023 , \36871 , \36875 );
and \U$36709 ( \37024 , \36875 , \36935 );
and \U$36710 ( \37025 , \36871 , \36935 );
or \U$36711 ( \37026 , \37023 , \37024 , \37025 );
and \U$36712 ( \37027 , \36966 , \36970 );
and \U$36713 ( \37028 , \36970 , \36975 );
and \U$36714 ( \37029 , \36966 , \36975 );
or \U$36715 ( \37030 , \37027 , \37028 , \37029 );
and \U$36716 ( \37031 , \36897 , \36901 );
and \U$36717 ( \37032 , \36901 , \36906 );
and \U$36718 ( \37033 , \36897 , \36906 );
or \U$36719 ( \37034 , \37031 , \37032 , \37033 );
xor \U$36720 ( \37035 , \37030 , \37034 );
and \U$36721 ( \37036 , \36882 , \36886 );
and \U$36722 ( \37037 , \36886 , \36891 );
and \U$36723 ( \37038 , \36882 , \36891 );
or \U$36724 ( \37039 , \37036 , \37037 , \37038 );
xor \U$36725 ( \37040 , \37035 , \37039 );
and \U$36726 ( \37041 , \22473 , \36955 );
and \U$36727 ( \37042 , \36955 , \36960 );
and \U$36728 ( \37043 , \22473 , \36960 );
or \U$36729 ( \37044 , \37041 , \37042 , \37043 );
and \U$36730 ( \37045 , \36995 , \36999 );
and \U$36731 ( \37046 , \36999 , \37004 );
and \U$36732 ( \37047 , \36995 , \37004 );
or \U$36733 ( \37048 , \37045 , \37046 , \37047 );
xor \U$36734 ( \37049 , \37044 , \37048 );
and \U$36735 ( \37050 , \36980 , \36984 );
and \U$36736 ( \37051 , \36984 , \36989 );
and \U$36737 ( \37052 , \36980 , \36989 );
or \U$36738 ( \37053 , \37050 , \37051 , \37052 );
xor \U$36739 ( \37054 , \37049 , \37053 );
xor \U$36740 ( \37055 , \37040 , \37054 );
and \U$36741 ( \37056 , \36976 , \36990 );
and \U$36742 ( \37057 , \36990 , \37005 );
and \U$36743 ( \37058 , \36976 , \37005 );
or \U$36744 ( \37059 , \37056 , \37057 , \37058 );
and \U$36745 ( \37060 , \22468 , \22208 );
and \U$36746 ( \37061 , \22429 , \22206 );
nor \U$36747 ( \37062 , \37060 , \37061 );
xnor \U$36748 ( \37063 , \37062 , \22218 );
and \U$36749 ( \37064 , \22489 , \22230 );
and \U$36750 ( \37065 , \22457 , \22228 );
nor \U$36751 ( \37066 , \37064 , \37065 );
xnor \U$36752 ( \37067 , \37066 , \22240 );
xor \U$36753 ( \37068 , \37063 , \37067 );
and \U$36754 ( \37069 , \22511 , \22257 );
and \U$36755 ( \37070 , \22478 , \22255 );
nor \U$36756 ( \37071 , \37069 , \37070 );
xnor \U$36757 ( \37072 , \37071 , \22267 );
xor \U$36758 ( \37073 , \37068 , \37072 );
and \U$36759 ( \37074 , \22397 , \22140 );
and \U$36760 ( \37075 , \22361 , \22138 );
nor \U$36761 ( \37076 , \37074 , \37075 );
xnor \U$36762 ( \37077 , \37076 , \22150 );
and \U$36763 ( \37078 , \22418 , \22162 );
and \U$36764 ( \37079 , \22386 , \22160 );
nor \U$36765 ( \37080 , \37078 , \37079 );
xnor \U$36766 ( \37081 , \37080 , \22172 );
xor \U$36767 ( \37082 , \37077 , \37081 );
and \U$36768 ( \37083 , \22440 , \22187 );
and \U$36769 ( \37084 , \22407 , \22185 );
nor \U$36770 ( \37085 , \37083 , \37084 );
xnor \U$36771 ( \37086 , \37085 , \22197 );
xor \U$36772 ( \37087 , \37082 , \37086 );
xor \U$36773 ( \37088 , \37073 , \37087 );
and \U$36774 ( \37089 , \22329 , \22076 );
and \U$36775 ( \37090 , \22294 , \22073 );
nor \U$36776 ( \37091 , \37089 , \37090 );
xnor \U$36777 ( \37092 , \37091 , \22072 );
and \U$36778 ( \37093 , \22350 , \22095 );
and \U$36779 ( \37094 , \22318 , \22093 );
nor \U$36780 ( \37095 , \37093 , \37094 );
xnor \U$36781 ( \37096 , \37095 , \22105 );
xor \U$36782 ( \37097 , \37092 , \37096 );
and \U$36783 ( \37098 , \22372 , \22119 );
and \U$36784 ( \37099 , \22339 , \22117 );
nor \U$36785 ( \37100 , \37098 , \37099 );
xnor \U$36786 ( \37101 , \37100 , \22129 );
xor \U$36787 ( \37102 , \37097 , \37101 );
xor \U$36788 ( \37103 , \37088 , \37102 );
xor \U$36789 ( \37104 , \37059 , \37103 );
and \U$36790 ( \37105 , \22676 , \22413 );
and \U$36791 ( \37106 , \22635 , \22411 );
nor \U$36792 ( \37107 , \37105 , \37106 );
xnor \U$36793 ( \37108 , \37107 , \22423 );
and \U$36794 ( \37109 , \22696 , \22435 );
and \U$36795 ( \37110 , \22665 , \22433 );
nor \U$36796 ( \37111 , \37109 , \37110 );
xnor \U$36797 ( \37112 , \37111 , \22445 );
xor \U$36798 ( \37113 , \37108 , \37112 );
and \U$36799 ( \37114 , \22706 , \22463 );
and \U$36800 ( \37115 , \22686 , \22461 );
nor \U$36801 ( \37116 , \37114 , \37115 );
xnor \U$36802 ( \37117 , \37116 , \22473 );
xor \U$36803 ( \37118 , \37113 , \37117 );
and \U$36804 ( \37119 , \22603 , \22345 );
and \U$36805 ( \37120 , \22567 , \22343 );
nor \U$36806 ( \37121 , \37119 , \37120 );
xnor \U$36807 ( \37122 , \37121 , \22355 );
and \U$36808 ( \37123 , \22624 , \22367 );
and \U$36809 ( \37124 , \22592 , \22365 );
nor \U$36810 ( \37125 , \37123 , \37124 );
xnor \U$36811 ( \37126 , \37125 , \22377 );
xor \U$36812 ( \37127 , \37122 , \37126 );
and \U$36813 ( \37128 , \22646 , \22392 );
and \U$36814 ( \37129 , \22613 , \22390 );
nor \U$36815 ( \37130 , \37128 , \37129 );
xnor \U$36816 ( \37131 , \37130 , \22402 );
xor \U$36817 ( \37132 , \37127 , \37131 );
xor \U$36818 ( \37133 , \37118 , \37132 );
and \U$36819 ( \37134 , \22535 , \22278 );
and \U$36820 ( \37135 , \22500 , \22276 );
nor \U$36821 ( \37136 , \37134 , \37135 );
xnor \U$36822 ( \37137 , \37136 , \22288 );
and \U$36823 ( \37138 , \22556 , \22300 );
and \U$36824 ( \37139 , \22524 , \22298 );
nor \U$36825 ( \37140 , \37138 , \37139 );
xnor \U$36826 ( \37141 , \37140 , \22310 );
xor \U$36827 ( \37142 , \37137 , \37141 );
and \U$36828 ( \37143 , \22578 , \22324 );
and \U$36829 ( \37144 , \22545 , \22322 );
nor \U$36830 ( \37145 , \37143 , \37144 );
xnor \U$36831 ( \37146 , \37145 , \22334 );
xor \U$36832 ( \37147 , \37142 , \37146 );
xor \U$36833 ( \37148 , \37133 , \37147 );
xor \U$36834 ( \37149 , \37104 , \37148 );
xor \U$36835 ( \37150 , \37055 , \37149 );
and \U$36836 ( \37151 , \36924 , \36928 );
and \U$36837 ( \37152 , \36928 , \36933 );
and \U$36838 ( \37153 , \36924 , \36933 );
or \U$36839 ( \37154 , \37151 , \37152 , \37153 );
and \U$36840 ( \37155 , \36912 , \36916 );
and \U$36841 ( \37156 , \36916 , \36918 );
and \U$36842 ( \37157 , \36912 , \36918 );
or \U$36843 ( \37158 , \37155 , \37156 , \37157 );
xor \U$36844 ( \37159 , \37154 , \37158 );
and \U$36845 ( \37160 , \36878 , \36892 );
and \U$36846 ( \37161 , \36892 , \36907 );
and \U$36847 ( \37162 , \36878 , \36907 );
or \U$36848 ( \37163 , \37160 , \37161 , \37162 );
xor \U$36849 ( \37164 , \37159 , \37163 );
xor \U$36850 ( \37165 , \37150 , \37164 );
xor \U$36851 ( \37166 , \37026 , \37165 );
and \U$36852 ( \37167 , \36857 , \36861 );
and \U$36853 ( \37168 , \36861 , \36866 );
and \U$36854 ( \37169 , \36857 , \36866 );
or \U$36855 ( \37170 , \37167 , \37168 , \37169 );
and \U$36856 ( \37171 , \36951 , \36961 );
and \U$36857 ( \37172 , \36961 , \37006 );
and \U$36858 ( \37173 , \36951 , \37006 );
or \U$36859 ( \37174 , \37171 , \37172 , \37173 );
xor \U$36860 ( \37175 , \37170 , \37174 );
and \U$36861 ( \37176 , \36908 , \36919 );
and \U$36862 ( \37177 , \36919 , \36934 );
and \U$36863 ( \37178 , \36908 , \36934 );
or \U$36864 ( \37179 , \37176 , \37177 , \37178 );
xor \U$36865 ( \37180 , \37175 , \37179 );
xor \U$36866 ( \37181 , \37166 , \37180 );
xor \U$36867 ( \37182 , \37022 , \37181 );
and \U$36868 ( \37183 , \36853 , \36937 );
and \U$36869 ( \37184 , \36937 , \37008 );
and \U$36870 ( \37185 , \36853 , \37008 );
or \U$36871 ( \37186 , \37183 , \37184 , \37185 );
nor \U$36872 ( \37187 , \37182 , \37186 );
and \U$36873 ( \37188 , \37026 , \37165 );
and \U$36874 ( \37189 , \37165 , \37180 );
and \U$36875 ( \37190 , \37026 , \37180 );
or \U$36876 ( \37191 , \37188 , \37189 , \37190 );
and \U$36877 ( \37192 , \37154 , \37158 );
and \U$36878 ( \37193 , \37158 , \37163 );
and \U$36879 ( \37194 , \37154 , \37163 );
or \U$36880 ( \37195 , \37192 , \37193 , \37194 );
and \U$36881 ( \37196 , \37059 , \37103 );
and \U$36882 ( \37197 , \37103 , \37148 );
and \U$36883 ( \37198 , \37059 , \37148 );
or \U$36884 ( \37199 , \37196 , \37197 , \37198 );
xor \U$36885 ( \37200 , \37195 , \37199 );
and \U$36886 ( \37201 , \37040 , \37054 );
xor \U$36887 ( \37202 , \37200 , \37201 );
xor \U$36888 ( \37203 , \37191 , \37202 );
and \U$36889 ( \37204 , \37170 , \37174 );
and \U$36890 ( \37205 , \37174 , \37179 );
and \U$36891 ( \37206 , \37170 , \37179 );
or \U$36892 ( \37207 , \37204 , \37205 , \37206 );
and \U$36893 ( \37208 , \37055 , \37149 );
and \U$36894 ( \37209 , \37149 , \37164 );
and \U$36895 ( \37210 , \37055 , \37164 );
or \U$36896 ( \37211 , \37208 , \37209 , \37210 );
xor \U$36897 ( \37212 , \37207 , \37211 );
and \U$36898 ( \37213 , \22686 , \22463 );
and \U$36899 ( \37214 , \22696 , \22461 );
nor \U$36900 ( \37215 , \37213 , \37214 );
xnor \U$36901 ( \37216 , \37215 , \22473 );
nand \U$36902 ( \37217 , \22706 , \22482 );
xnor \U$36903 ( \37218 , \37217 , \22494 );
xor \U$36904 ( \37219 , \37216 , \37218 );
and \U$36905 ( \37220 , \22613 , \22392 );
and \U$36906 ( \37221 , \22624 , \22390 );
nor \U$36907 ( \37222 , \37220 , \37221 );
xnor \U$36908 ( \37223 , \37222 , \22402 );
and \U$36909 ( \37224 , \22635 , \22413 );
and \U$36910 ( \37225 , \22646 , \22411 );
nor \U$36911 ( \37226 , \37224 , \37225 );
xnor \U$36912 ( \37227 , \37226 , \22423 );
xor \U$36913 ( \37228 , \37223 , \37227 );
and \U$36914 ( \37229 , \22665 , \22435 );
and \U$36915 ( \37230 , \22676 , \22433 );
nor \U$36916 ( \37231 , \37229 , \37230 );
xnor \U$36917 ( \37232 , \37231 , \22445 );
xor \U$36918 ( \37233 , \37228 , \37232 );
xor \U$36919 ( \37234 , \37219 , \37233 );
and \U$36920 ( \37235 , \37137 , \37141 );
and \U$36921 ( \37236 , \37141 , \37146 );
and \U$36922 ( \37237 , \37137 , \37146 );
or \U$36923 ( \37238 , \37235 , \37236 , \37237 );
and \U$36924 ( \37239 , \37122 , \37126 );
and \U$36925 ( \37240 , \37126 , \37131 );
and \U$36926 ( \37241 , \37122 , \37131 );
or \U$36927 ( \37242 , \37239 , \37240 , \37241 );
xor \U$36928 ( \37243 , \37238 , \37242 );
and \U$36929 ( \37244 , \37108 , \37112 );
and \U$36930 ( \37245 , \37112 , \37117 );
and \U$36931 ( \37246 , \37108 , \37117 );
or \U$36932 ( \37247 , \37244 , \37245 , \37246 );
xor \U$36933 ( \37248 , \37243 , \37247 );
xor \U$36934 ( \37249 , \37234 , \37248 );
and \U$36935 ( \37250 , \37092 , \37096 );
and \U$36936 ( \37251 , \37096 , \37101 );
and \U$36937 ( \37252 , \37092 , \37101 );
or \U$36938 ( \37253 , \37250 , \37251 , \37252 );
and \U$36939 ( \37254 , \37077 , \37081 );
and \U$36940 ( \37255 , \37081 , \37086 );
and \U$36941 ( \37256 , \37077 , \37086 );
or \U$36942 ( \37257 , \37254 , \37255 , \37256 );
xor \U$36943 ( \37258 , \37253 , \37257 );
and \U$36944 ( \37259 , \37063 , \37067 );
and \U$36945 ( \37260 , \37067 , \37072 );
and \U$36946 ( \37261 , \37063 , \37072 );
or \U$36947 ( \37262 , \37259 , \37260 , \37261 );
xor \U$36948 ( \37263 , \37258 , \37262 );
xor \U$36949 ( \37264 , \37249 , \37263 );
and \U$36950 ( \37265 , \37073 , \37087 );
and \U$36951 ( \37266 , \37087 , \37102 );
and \U$36952 ( \37267 , \37073 , \37102 );
or \U$36953 ( \37268 , \37265 , \37266 , \37267 );
and \U$36954 ( \37269 , \22339 , \22119 );
and \U$36955 ( \37270 , \22350 , \22117 );
nor \U$36956 ( \37271 , \37269 , \37270 );
xnor \U$36957 ( \37272 , \37271 , \22129 );
and \U$36958 ( \37273 , \22361 , \22140 );
and \U$36959 ( \37274 , \22372 , \22138 );
nor \U$36960 ( \37275 , \37273 , \37274 );
xnor \U$36961 ( \37276 , \37275 , \22150 );
xor \U$36962 ( \37277 , \37272 , \37276 );
and \U$36963 ( \37278 , \22386 , \22162 );
and \U$36964 ( \37279 , \22397 , \22160 );
nor \U$36965 ( \37280 , \37278 , \37279 );
xnor \U$36966 ( \37281 , \37280 , \22172 );
xor \U$36967 ( \37282 , \37277 , \37281 );
and \U$36968 ( \37283 , \22294 , \22076 );
and \U$36969 ( \37284 , \22305 , \22073 );
nor \U$36970 ( \37285 , \37283 , \37284 );
xnor \U$36971 ( \37286 , \37285 , \22072 );
xor \U$36972 ( \37287 , \22494 , \37286 );
and \U$36973 ( \37288 , \22318 , \22095 );
and \U$36974 ( \37289 , \22329 , \22093 );
nor \U$36975 ( \37290 , \37288 , \37289 );
xnor \U$36976 ( \37291 , \37290 , \22105 );
xor \U$36977 ( \37292 , \37287 , \37291 );
xor \U$36978 ( \37293 , \37282 , \37292 );
xor \U$36979 ( \37294 , \37268 , \37293 );
and \U$36980 ( \37295 , \22545 , \22324 );
and \U$36981 ( \37296 , \22556 , \22322 );
nor \U$36982 ( \37297 , \37295 , \37296 );
xnor \U$36983 ( \37298 , \37297 , \22334 );
and \U$36984 ( \37299 , \22567 , \22345 );
and \U$36985 ( \37300 , \22578 , \22343 );
nor \U$36986 ( \37301 , \37299 , \37300 );
xnor \U$36987 ( \37302 , \37301 , \22355 );
xor \U$36988 ( \37303 , \37298 , \37302 );
and \U$36989 ( \37304 , \22592 , \22367 );
and \U$36990 ( \37305 , \22603 , \22365 );
nor \U$36991 ( \37306 , \37304 , \37305 );
xnor \U$36992 ( \37307 , \37306 , \22377 );
xor \U$36993 ( \37308 , \37303 , \37307 );
and \U$36994 ( \37309 , \22478 , \22257 );
and \U$36995 ( \37310 , \22489 , \22255 );
nor \U$36996 ( \37311 , \37309 , \37310 );
xnor \U$36997 ( \37312 , \37311 , \22267 );
and \U$36998 ( \37313 , \22500 , \22278 );
and \U$36999 ( \37314 , \22511 , \22276 );
nor \U$37000 ( \37315 , \37313 , \37314 );
xnor \U$37001 ( \37316 , \37315 , \22288 );
xor \U$37002 ( \37317 , \37312 , \37316 );
and \U$37003 ( \37318 , \22524 , \22300 );
and \U$37004 ( \37319 , \22535 , \22298 );
nor \U$37005 ( \37320 , \37318 , \37319 );
xnor \U$37006 ( \37321 , \37320 , \22310 );
xor \U$37007 ( \37322 , \37317 , \37321 );
xor \U$37008 ( \37323 , \37308 , \37322 );
and \U$37009 ( \37324 , \22407 , \22187 );
and \U$37010 ( \37325 , \22418 , \22185 );
nor \U$37011 ( \37326 , \37324 , \37325 );
xnor \U$37012 ( \37327 , \37326 , \22197 );
and \U$37013 ( \37328 , \22429 , \22208 );
and \U$37014 ( \37329 , \22440 , \22206 );
nor \U$37015 ( \37330 , \37328 , \37329 );
xnor \U$37016 ( \37331 , \37330 , \22218 );
xor \U$37017 ( \37332 , \37327 , \37331 );
and \U$37018 ( \37333 , \22457 , \22230 );
and \U$37019 ( \37334 , \22468 , \22228 );
nor \U$37020 ( \37335 , \37333 , \37334 );
xnor \U$37021 ( \37336 , \37335 , \22240 );
xor \U$37022 ( \37337 , \37332 , \37336 );
xor \U$37023 ( \37338 , \37323 , \37337 );
xor \U$37024 ( \37339 , \37294 , \37338 );
xor \U$37025 ( \37340 , \37264 , \37339 );
and \U$37026 ( \37341 , \37044 , \37048 );
and \U$37027 ( \37342 , \37048 , \37053 );
and \U$37028 ( \37343 , \37044 , \37053 );
or \U$37029 ( \37344 , \37341 , \37342 , \37343 );
and \U$37030 ( \37345 , \37030 , \37034 );
and \U$37031 ( \37346 , \37034 , \37039 );
and \U$37032 ( \37347 , \37030 , \37039 );
or \U$37033 ( \37348 , \37345 , \37346 , \37347 );
xor \U$37034 ( \37349 , \37344 , \37348 );
and \U$37035 ( \37350 , \37118 , \37132 );
and \U$37036 ( \37351 , \37132 , \37147 );
and \U$37037 ( \37352 , \37118 , \37147 );
or \U$37038 ( \37353 , \37350 , \37351 , \37352 );
xor \U$37039 ( \37354 , \37349 , \37353 );
xor \U$37040 ( \37355 , \37340 , \37354 );
xor \U$37041 ( \37356 , \37212 , \37355 );
xor \U$37042 ( \37357 , \37203 , \37356 );
and \U$37043 ( \37358 , \37020 , \37021 );
and \U$37044 ( \37359 , \37021 , \37181 );
and \U$37045 ( \37360 , \37020 , \37181 );
or \U$37046 ( \37361 , \37358 , \37359 , \37360 );
nor \U$37047 ( \37362 , \37357 , \37361 );
nor \U$37048 ( \37363 , \37187 , \37362 );
and \U$37049 ( \37364 , \37207 , \37211 );
and \U$37050 ( \37365 , \37211 , \37355 );
and \U$37051 ( \37366 , \37207 , \37355 );
or \U$37052 ( \37367 , \37364 , \37365 , \37366 );
and \U$37053 ( \37368 , \22494 , \37286 );
and \U$37054 ( \37369 , \37286 , \37291 );
and \U$37055 ( \37370 , \22494 , \37291 );
or \U$37056 ( \37371 , \37368 , \37369 , \37370 );
and \U$37057 ( \37372 , \37272 , \37276 );
and \U$37058 ( \37373 , \37276 , \37281 );
and \U$37059 ( \37374 , \37272 , \37281 );
or \U$37060 ( \37375 , \37372 , \37373 , \37374 );
xor \U$37061 ( \37376 , \37371 , \37375 );
and \U$37062 ( \37377 , \37327 , \37331 );
and \U$37063 ( \37378 , \37331 , \37336 );
and \U$37064 ( \37379 , \37327 , \37336 );
or \U$37065 ( \37380 , \37377 , \37378 , \37379 );
xor \U$37066 ( \37381 , \37376 , \37380 );
and \U$37067 ( \37382 , \22511 , \22278 );
and \U$37068 ( \37383 , \22478 , \22276 );
nor \U$37069 ( \37384 , \37382 , \37383 );
xnor \U$37070 ( \37385 , \37384 , \22288 );
and \U$37071 ( \37386 , \22535 , \22300 );
and \U$37072 ( \37387 , \22500 , \22298 );
nor \U$37073 ( \37388 , \37386 , \37387 );
xnor \U$37074 ( \37389 , \37388 , \22310 );
xor \U$37075 ( \37390 , \37385 , \37389 );
and \U$37076 ( \37391 , \22556 , \22324 );
and \U$37077 ( \37392 , \22524 , \22322 );
nor \U$37078 ( \37393 , \37391 , \37392 );
xnor \U$37079 ( \37394 , \37393 , \22334 );
xor \U$37080 ( \37395 , \37390 , \37394 );
and \U$37081 ( \37396 , \22440 , \22208 );
and \U$37082 ( \37397 , \22407 , \22206 );
nor \U$37083 ( \37398 , \37396 , \37397 );
xnor \U$37084 ( \37399 , \37398 , \22218 );
and \U$37085 ( \37400 , \22468 , \22230 );
and \U$37086 ( \37401 , \22429 , \22228 );
nor \U$37087 ( \37402 , \37400 , \37401 );
xnor \U$37088 ( \37403 , \37402 , \22240 );
xor \U$37089 ( \37404 , \37399 , \37403 );
and \U$37090 ( \37405 , \22489 , \22257 );
and \U$37091 ( \37406 , \22457 , \22255 );
nor \U$37092 ( \37407 , \37405 , \37406 );
xnor \U$37093 ( \37408 , \37407 , \22267 );
xor \U$37094 ( \37409 , \37404 , \37408 );
xor \U$37095 ( \37410 , \37395 , \37409 );
and \U$37096 ( \37411 , \22372 , \22140 );
and \U$37097 ( \37412 , \22339 , \22138 );
nor \U$37098 ( \37413 , \37411 , \37412 );
xnor \U$37099 ( \37414 , \37413 , \22150 );
and \U$37100 ( \37415 , \22397 , \22162 );
and \U$37101 ( \37416 , \22361 , \22160 );
nor \U$37102 ( \37417 , \37415 , \37416 );
xnor \U$37103 ( \37418 , \37417 , \22172 );
xor \U$37104 ( \37419 , \37414 , \37418 );
and \U$37105 ( \37420 , \22418 , \22187 );
and \U$37106 ( \37421 , \22386 , \22185 );
nor \U$37107 ( \37422 , \37420 , \37421 );
xnor \U$37108 ( \37423 , \37422 , \22197 );
xor \U$37109 ( \37424 , \37419 , \37423 );
xor \U$37110 ( \37425 , \37410 , \37424 );
and \U$37111 ( \37426 , \22706 , \22484 );
and \U$37112 ( \37427 , \22686 , \22482 );
nor \U$37113 ( \37428 , \37426 , \37427 );
xnor \U$37114 ( \37429 , \37428 , \22494 );
and \U$37115 ( \37430 , \22646 , \22413 );
and \U$37116 ( \37431 , \22613 , \22411 );
nor \U$37117 ( \37432 , \37430 , \37431 );
xnor \U$37118 ( \37433 , \37432 , \22423 );
and \U$37119 ( \37434 , \22676 , \22435 );
and \U$37120 ( \37435 , \22635 , \22433 );
nor \U$37121 ( \37436 , \37434 , \37435 );
xnor \U$37122 ( \37437 , \37436 , \22445 );
xor \U$37123 ( \37438 , \37433 , \37437 );
and \U$37124 ( \37439 , \22696 , \22463 );
and \U$37125 ( \37440 , \22665 , \22461 );
nor \U$37126 ( \37441 , \37439 , \37440 );
xnor \U$37127 ( \37442 , \37441 , \22473 );
xor \U$37128 ( \37443 , \37438 , \37442 );
xor \U$37129 ( \37444 , \37429 , \37443 );
and \U$37130 ( \37445 , \22578 , \22345 );
and \U$37131 ( \37446 , \22545 , \22343 );
nor \U$37132 ( \37447 , \37445 , \37446 );
xnor \U$37133 ( \37448 , \37447 , \22355 );
and \U$37134 ( \37449 , \22603 , \22367 );
and \U$37135 ( \37450 , \22567 , \22365 );
nor \U$37136 ( \37451 , \37449 , \37450 );
xnor \U$37137 ( \37452 , \37451 , \22377 );
xor \U$37138 ( \37453 , \37448 , \37452 );
and \U$37139 ( \37454 , \22624 , \22392 );
and \U$37140 ( \37455 , \22592 , \22390 );
nor \U$37141 ( \37456 , \37454 , \37455 );
xnor \U$37142 ( \37457 , \37456 , \22402 );
xor \U$37143 ( \37458 , \37453 , \37457 );
xor \U$37144 ( \37459 , \37444 , \37458 );
xor \U$37145 ( \37460 , \37425 , \37459 );
and \U$37146 ( \37461 , \37312 , \37316 );
and \U$37147 ( \37462 , \37316 , \37321 );
and \U$37148 ( \37463 , \37312 , \37321 );
or \U$37149 ( \37464 , \37461 , \37462 , \37463 );
and \U$37150 ( \37465 , \37298 , \37302 );
and \U$37151 ( \37466 , \37302 , \37307 );
and \U$37152 ( \37467 , \37298 , \37307 );
or \U$37153 ( \37468 , \37465 , \37466 , \37467 );
xor \U$37154 ( \37469 , \37464 , \37468 );
and \U$37155 ( \37470 , \37223 , \37227 );
and \U$37156 ( \37471 , \37227 , \37232 );
and \U$37157 ( \37472 , \37223 , \37232 );
or \U$37158 ( \37473 , \37470 , \37471 , \37472 );
xor \U$37159 ( \37474 , \37469 , \37473 );
xor \U$37160 ( \37475 , \37460 , \37474 );
xor \U$37161 ( \37476 , \37381 , \37475 );
and \U$37162 ( \37477 , \37308 , \37322 );
and \U$37163 ( \37478 , \37322 , \37337 );
and \U$37164 ( \37479 , \37308 , \37337 );
or \U$37165 ( \37480 , \37477 , \37478 , \37479 );
and \U$37166 ( \37481 , \37282 , \37292 );
xor \U$37167 ( \37482 , \37480 , \37481 );
and \U$37168 ( \37483 , \22305 , \22076 );
and \U$37169 ( \37484 , \22272 , \22073 );
nor \U$37170 ( \37485 , \37483 , \37484 );
xnor \U$37171 ( \37486 , \37485 , \22072 );
and \U$37172 ( \37487 , \22329 , \22095 );
and \U$37173 ( \37488 , \22294 , \22093 );
nor \U$37174 ( \37489 , \37487 , \37488 );
xnor \U$37175 ( \37490 , \37489 , \22105 );
xor \U$37176 ( \37491 , \37486 , \37490 );
and \U$37177 ( \37492 , \22350 , \22119 );
and \U$37178 ( \37493 , \22318 , \22117 );
nor \U$37179 ( \37494 , \37492 , \37493 );
xnor \U$37180 ( \37495 , \37494 , \22129 );
xor \U$37181 ( \37496 , \37491 , \37495 );
xor \U$37182 ( \37497 , \37482 , \37496 );
xor \U$37183 ( \37498 , \37476 , \37497 );
and \U$37184 ( \37499 , \37344 , \37348 );
and \U$37185 ( \37500 , \37348 , \37353 );
and \U$37186 ( \37501 , \37344 , \37353 );
or \U$37187 ( \37502 , \37499 , \37500 , \37501 );
and \U$37188 ( \37503 , \37268 , \37293 );
and \U$37189 ( \37504 , \37293 , \37338 );
and \U$37190 ( \37505 , \37268 , \37338 );
or \U$37191 ( \37506 , \37503 , \37504 , \37505 );
xor \U$37192 ( \37507 , \37502 , \37506 );
and \U$37193 ( \37508 , \37234 , \37248 );
and \U$37194 ( \37509 , \37248 , \37263 );
and \U$37195 ( \37510 , \37234 , \37263 );
or \U$37196 ( \37511 , \37508 , \37509 , \37510 );
xor \U$37197 ( \37512 , \37507 , \37511 );
xor \U$37198 ( \37513 , \37498 , \37512 );
xor \U$37199 ( \37514 , \37367 , \37513 );
and \U$37200 ( \37515 , \37195 , \37199 );
and \U$37201 ( \37516 , \37199 , \37201 );
and \U$37202 ( \37517 , \37195 , \37201 );
or \U$37203 ( \37518 , \37515 , \37516 , \37517 );
and \U$37204 ( \37519 , \37264 , \37339 );
and \U$37205 ( \37520 , \37339 , \37354 );
and \U$37206 ( \37521 , \37264 , \37354 );
or \U$37207 ( \37522 , \37519 , \37520 , \37521 );
xor \U$37208 ( \37523 , \37518 , \37522 );
and \U$37209 ( \37524 , \37253 , \37257 );
and \U$37210 ( \37525 , \37257 , \37262 );
and \U$37211 ( \37526 , \37253 , \37262 );
or \U$37212 ( \37527 , \37524 , \37525 , \37526 );
and \U$37213 ( \37528 , \37238 , \37242 );
and \U$37214 ( \37529 , \37242 , \37247 );
and \U$37215 ( \37530 , \37238 , \37247 );
or \U$37216 ( \37531 , \37528 , \37529 , \37530 );
xor \U$37217 ( \37532 , \37527 , \37531 );
and \U$37218 ( \37533 , \37216 , \37218 );
and \U$37219 ( \37534 , \37218 , \37233 );
and \U$37220 ( \37535 , \37216 , \37233 );
or \U$37221 ( \37536 , \37533 , \37534 , \37535 );
xor \U$37222 ( \37537 , \37532 , \37536 );
xor \U$37223 ( \37538 , \37523 , \37537 );
xor \U$37224 ( \37539 , \37514 , \37538 );
and \U$37225 ( \37540 , \37191 , \37202 );
and \U$37226 ( \37541 , \37202 , \37356 );
and \U$37227 ( \37542 , \37191 , \37356 );
or \U$37228 ( \37543 , \37540 , \37541 , \37542 );
nor \U$37229 ( \37544 , \37539 , \37543 );
and \U$37230 ( \37545 , \37502 , \37506 );
and \U$37231 ( \37546 , \37506 , \37511 );
and \U$37232 ( \37547 , \37502 , \37511 );
or \U$37233 ( \37548 , \37545 , \37546 , \37547 );
and \U$37234 ( \37549 , \37381 , \37475 );
and \U$37235 ( \37550 , \37475 , \37497 );
and \U$37236 ( \37551 , \37381 , \37497 );
or \U$37237 ( \37552 , \37549 , \37550 , \37551 );
xor \U$37238 ( \37553 , \37548 , \37552 );
and \U$37239 ( \37554 , \22665 , \22463 );
and \U$37240 ( \37555 , \22676 , \22461 );
nor \U$37241 ( \37556 , \37554 , \37555 );
xnor \U$37242 ( \37557 , \37556 , \22473 );
and \U$37243 ( \37558 , \22686 , \22484 );
and \U$37244 ( \37559 , \22696 , \22482 );
nor \U$37245 ( \37560 , \37558 , \37559 );
xnor \U$37246 ( \37561 , \37560 , \22494 );
xor \U$37247 ( \37562 , \37557 , \37561 );
nand \U$37248 ( \37563 , \22706 , \22504 );
xnor \U$37249 ( \37564 , \37563 , \22516 );
xor \U$37250 ( \37565 , \37562 , \37564 );
and \U$37251 ( \37566 , \22592 , \22392 );
and \U$37252 ( \37567 , \22603 , \22390 );
nor \U$37253 ( \37568 , \37566 , \37567 );
xnor \U$37254 ( \37569 , \37568 , \22402 );
and \U$37255 ( \37570 , \22613 , \22413 );
and \U$37256 ( \37571 , \22624 , \22411 );
nor \U$37257 ( \37572 , \37570 , \37571 );
xnor \U$37258 ( \37573 , \37572 , \22423 );
xor \U$37259 ( \37574 , \37569 , \37573 );
and \U$37260 ( \37575 , \22635 , \22435 );
and \U$37261 ( \37576 , \22646 , \22433 );
nor \U$37262 ( \37577 , \37575 , \37576 );
xnor \U$37263 ( \37578 , \37577 , \22445 );
xor \U$37264 ( \37579 , \37574 , \37578 );
xor \U$37265 ( \37580 , \37565 , \37579 );
and \U$37266 ( \37581 , \22524 , \22324 );
and \U$37267 ( \37582 , \22535 , \22322 );
nor \U$37268 ( \37583 , \37581 , \37582 );
xnor \U$37269 ( \37584 , \37583 , \22334 );
and \U$37270 ( \37585 , \22545 , \22345 );
and \U$37271 ( \37586 , \22556 , \22343 );
nor \U$37272 ( \37587 , \37585 , \37586 );
xnor \U$37273 ( \37588 , \37587 , \22355 );
xor \U$37274 ( \37589 , \37584 , \37588 );
and \U$37275 ( \37590 , \22567 , \22367 );
and \U$37276 ( \37591 , \22578 , \22365 );
nor \U$37277 ( \37592 , \37590 , \37591 );
xnor \U$37278 ( \37593 , \37592 , \22377 );
xor \U$37279 ( \37594 , \37589 , \37593 );
xor \U$37280 ( \37595 , \37580 , \37594 );
and \U$37281 ( \37596 , \37385 , \37389 );
and \U$37282 ( \37597 , \37389 , \37394 );
and \U$37283 ( \37598 , \37385 , \37394 );
or \U$37284 ( \37599 , \37596 , \37597 , \37598 );
and \U$37285 ( \37600 , \37448 , \37452 );
and \U$37286 ( \37601 , \37452 , \37457 );
and \U$37287 ( \37602 , \37448 , \37457 );
or \U$37288 ( \37603 , \37600 , \37601 , \37602 );
xor \U$37289 ( \37604 , \37599 , \37603 );
and \U$37290 ( \37605 , \37433 , \37437 );
and \U$37291 ( \37606 , \37437 , \37442 );
and \U$37292 ( \37607 , \37433 , \37442 );
or \U$37293 ( \37608 , \37605 , \37606 , \37607 );
xor \U$37294 ( \37609 , \37604 , \37608 );
xor \U$37295 ( \37610 , \37595 , \37609 );
and \U$37296 ( \37611 , \37486 , \37490 );
and \U$37297 ( \37612 , \37490 , \37495 );
and \U$37298 ( \37613 , \37486 , \37495 );
or \U$37299 ( \37614 , \37611 , \37612 , \37613 );
and \U$37300 ( \37615 , \37414 , \37418 );
and \U$37301 ( \37616 , \37418 , \37423 );
and \U$37302 ( \37617 , \37414 , \37423 );
or \U$37303 ( \37618 , \37615 , \37616 , \37617 );
xor \U$37304 ( \37619 , \37614 , \37618 );
and \U$37305 ( \37620 , \37399 , \37403 );
and \U$37306 ( \37621 , \37403 , \37408 );
and \U$37307 ( \37622 , \37399 , \37408 );
or \U$37308 ( \37623 , \37620 , \37621 , \37622 );
xor \U$37309 ( \37624 , \37619 , \37623 );
xor \U$37310 ( \37625 , \37610 , \37624 );
and \U$37311 ( \37626 , \37395 , \37409 );
and \U$37312 ( \37627 , \37409 , \37424 );
and \U$37313 ( \37628 , \37395 , \37424 );
or \U$37314 ( \37629 , \37626 , \37627 , \37628 );
and \U$37315 ( \37630 , \22272 , \22076 );
and \U$37316 ( \37631 , \22283 , \22073 );
nor \U$37317 ( \37632 , \37630 , \37631 );
xnor \U$37318 ( \37633 , \37632 , \22072 );
xor \U$37319 ( \37634 , \22516 , \37633 );
and \U$37320 ( \37635 , \22294 , \22095 );
and \U$37321 ( \37636 , \22305 , \22093 );
nor \U$37322 ( \37637 , \37635 , \37636 );
xnor \U$37323 ( \37638 , \37637 , \22105 );
xor \U$37324 ( \37639 , \37634 , \37638 );
xor \U$37325 ( \37640 , \37629 , \37639 );
and \U$37326 ( \37641 , \22457 , \22257 );
and \U$37327 ( \37642 , \22468 , \22255 );
nor \U$37328 ( \37643 , \37641 , \37642 );
xnor \U$37329 ( \37644 , \37643 , \22267 );
and \U$37330 ( \37645 , \22478 , \22278 );
and \U$37331 ( \37646 , \22489 , \22276 );
nor \U$37332 ( \37647 , \37645 , \37646 );
xnor \U$37333 ( \37648 , \37647 , \22288 );
xor \U$37334 ( \37649 , \37644 , \37648 );
and \U$37335 ( \37650 , \22500 , \22300 );
and \U$37336 ( \37651 , \22511 , \22298 );
nor \U$37337 ( \37652 , \37650 , \37651 );
xnor \U$37338 ( \37653 , \37652 , \22310 );
xor \U$37339 ( \37654 , \37649 , \37653 );
and \U$37340 ( \37655 , \22386 , \22187 );
and \U$37341 ( \37656 , \22397 , \22185 );
nor \U$37342 ( \37657 , \37655 , \37656 );
xnor \U$37343 ( \37658 , \37657 , \22197 );
and \U$37344 ( \37659 , \22407 , \22208 );
and \U$37345 ( \37660 , \22418 , \22206 );
nor \U$37346 ( \37661 , \37659 , \37660 );
xnor \U$37347 ( \37662 , \37661 , \22218 );
xor \U$37348 ( \37663 , \37658 , \37662 );
and \U$37349 ( \37664 , \22429 , \22230 );
and \U$37350 ( \37665 , \22440 , \22228 );
nor \U$37351 ( \37666 , \37664 , \37665 );
xnor \U$37352 ( \37667 , \37666 , \22240 );
xor \U$37353 ( \37668 , \37663 , \37667 );
xor \U$37354 ( \37669 , \37654 , \37668 );
and \U$37355 ( \37670 , \22318 , \22119 );
and \U$37356 ( \37671 , \22329 , \22117 );
nor \U$37357 ( \37672 , \37670 , \37671 );
xnor \U$37358 ( \37673 , \37672 , \22129 );
and \U$37359 ( \37674 , \22339 , \22140 );
and \U$37360 ( \37675 , \22350 , \22138 );
nor \U$37361 ( \37676 , \37674 , \37675 );
xnor \U$37362 ( \37677 , \37676 , \22150 );
xor \U$37363 ( \37678 , \37673 , \37677 );
and \U$37364 ( \37679 , \22361 , \22162 );
and \U$37365 ( \37680 , \22372 , \22160 );
nor \U$37366 ( \37681 , \37679 , \37680 );
xnor \U$37367 ( \37682 , \37681 , \22172 );
xor \U$37368 ( \37683 , \37678 , \37682 );
xor \U$37369 ( \37684 , \37669 , \37683 );
xor \U$37370 ( \37685 , \37640 , \37684 );
xor \U$37371 ( \37686 , \37625 , \37685 );
and \U$37372 ( \37687 , \37371 , \37375 );
and \U$37373 ( \37688 , \37375 , \37380 );
and \U$37374 ( \37689 , \37371 , \37380 );
or \U$37375 ( \37690 , \37687 , \37688 , \37689 );
and \U$37376 ( \37691 , \37464 , \37468 );
and \U$37377 ( \37692 , \37468 , \37473 );
and \U$37378 ( \37693 , \37464 , \37473 );
or \U$37379 ( \37694 , \37691 , \37692 , \37693 );
xor \U$37380 ( \37695 , \37690 , \37694 );
and \U$37381 ( \37696 , \37429 , \37443 );
and \U$37382 ( \37697 , \37443 , \37458 );
and \U$37383 ( \37698 , \37429 , \37458 );
or \U$37384 ( \37699 , \37696 , \37697 , \37698 );
xor \U$37385 ( \37700 , \37695 , \37699 );
xor \U$37386 ( \37701 , \37686 , \37700 );
xor \U$37387 ( \37702 , \37553 , \37701 );
and \U$37388 ( \37703 , \37518 , \37522 );
and \U$37389 ( \37704 , \37522 , \37537 );
and \U$37390 ( \37705 , \37518 , \37537 );
or \U$37391 ( \37706 , \37703 , \37704 , \37705 );
and \U$37392 ( \37707 , \37498 , \37512 );
xor \U$37393 ( \37708 , \37706 , \37707 );
and \U$37394 ( \37709 , \37527 , \37531 );
and \U$37395 ( \37710 , \37531 , \37536 );
and \U$37396 ( \37711 , \37527 , \37536 );
or \U$37397 ( \37712 , \37709 , \37710 , \37711 );
and \U$37398 ( \37713 , \37480 , \37481 );
and \U$37399 ( \37714 , \37481 , \37496 );
and \U$37400 ( \37715 , \37480 , \37496 );
or \U$37401 ( \37716 , \37713 , \37714 , \37715 );
xor \U$37402 ( \37717 , \37712 , \37716 );
and \U$37403 ( \37718 , \37425 , \37459 );
and \U$37404 ( \37719 , \37459 , \37474 );
and \U$37405 ( \37720 , \37425 , \37474 );
or \U$37406 ( \37721 , \37718 , \37719 , \37720 );
xor \U$37407 ( \37722 , \37717 , \37721 );
xor \U$37408 ( \37723 , \37708 , \37722 );
xor \U$37409 ( \37724 , \37702 , \37723 );
and \U$37410 ( \37725 , \37367 , \37513 );
and \U$37411 ( \37726 , \37513 , \37538 );
and \U$37412 ( \37727 , \37367 , \37538 );
or \U$37413 ( \37728 , \37725 , \37726 , \37727 );
nor \U$37414 ( \37729 , \37724 , \37728 );
nor \U$37415 ( \37730 , \37544 , \37729 );
nand \U$37416 ( \37731 , \37363 , \37730 );
nor \U$37417 ( \37732 , \37016 , \37731 );
and \U$37418 ( \37733 , \37706 , \37707 );
and \U$37419 ( \37734 , \37707 , \37722 );
and \U$37420 ( \37735 , \37706 , \37722 );
or \U$37421 ( \37736 , \37733 , \37734 , \37735 );
and \U$37422 ( \37737 , \37548 , \37552 );
and \U$37423 ( \37738 , \37552 , \37701 );
and \U$37424 ( \37739 , \37548 , \37701 );
or \U$37425 ( \37740 , \37737 , \37738 , \37739 );
and \U$37426 ( \37741 , \37690 , \37694 );
and \U$37427 ( \37742 , \37694 , \37699 );
and \U$37428 ( \37743 , \37690 , \37699 );
or \U$37429 ( \37744 , \37741 , \37742 , \37743 );
and \U$37430 ( \37745 , \37629 , \37639 );
and \U$37431 ( \37746 , \37639 , \37684 );
and \U$37432 ( \37747 , \37629 , \37684 );
or \U$37433 ( \37748 , \37745 , \37746 , \37747 );
xor \U$37434 ( \37749 , \37744 , \37748 );
and \U$37435 ( \37750 , \37595 , \37609 );
and \U$37436 ( \37751 , \37609 , \37624 );
and \U$37437 ( \37752 , \37595 , \37624 );
or \U$37438 ( \37753 , \37750 , \37751 , \37752 );
xor \U$37439 ( \37754 , \37749 , \37753 );
xor \U$37440 ( \37755 , \37740 , \37754 );
and \U$37441 ( \37756 , \37712 , \37716 );
and \U$37442 ( \37757 , \37716 , \37721 );
and \U$37443 ( \37758 , \37712 , \37721 );
or \U$37444 ( \37759 , \37756 , \37757 , \37758 );
and \U$37445 ( \37760 , \37625 , \37685 );
and \U$37446 ( \37761 , \37685 , \37700 );
and \U$37447 ( \37762 , \37625 , \37700 );
or \U$37448 ( \37763 , \37760 , \37761 , \37762 );
xor \U$37449 ( \37764 , \37759 , \37763 );
and \U$37450 ( \37765 , \37557 , \37561 );
and \U$37451 ( \37766 , \37561 , \37564 );
and \U$37452 ( \37767 , \37557 , \37564 );
or \U$37453 ( \37768 , \37765 , \37766 , \37767 );
and \U$37454 ( \37769 , \22696 , \22484 );
and \U$37455 ( \37770 , \22665 , \22482 );
nor \U$37456 ( \37771 , \37769 , \37770 );
xnor \U$37457 ( \37772 , \37771 , \22494 );
xor \U$37458 ( \37773 , \37768 , \37772 );
and \U$37459 ( \37774 , \22706 , \22506 );
and \U$37460 ( \37775 , \22686 , \22504 );
nor \U$37461 ( \37776 , \37774 , \37775 );
xnor \U$37462 ( \37777 , \37776 , \22516 );
xor \U$37463 ( \37778 , \37773 , \37777 );
and \U$37464 ( \37779 , \37644 , \37648 );
and \U$37465 ( \37780 , \37648 , \37653 );
and \U$37466 ( \37781 , \37644 , \37653 );
or \U$37467 ( \37782 , \37779 , \37780 , \37781 );
and \U$37468 ( \37783 , \37584 , \37588 );
and \U$37469 ( \37784 , \37588 , \37593 );
and \U$37470 ( \37785 , \37584 , \37593 );
or \U$37471 ( \37786 , \37783 , \37784 , \37785 );
xor \U$37472 ( \37787 , \37782 , \37786 );
and \U$37473 ( \37788 , \37569 , \37573 );
and \U$37474 ( \37789 , \37573 , \37578 );
and \U$37475 ( \37790 , \37569 , \37578 );
or \U$37476 ( \37791 , \37788 , \37789 , \37790 );
xor \U$37477 ( \37792 , \37787 , \37791 );
xor \U$37478 ( \37793 , \37778 , \37792 );
and \U$37479 ( \37794 , \22516 , \37633 );
and \U$37480 ( \37795 , \37633 , \37638 );
and \U$37481 ( \37796 , \22516 , \37638 );
or \U$37482 ( \37797 , \37794 , \37795 , \37796 );
and \U$37483 ( \37798 , \37673 , \37677 );
and \U$37484 ( \37799 , \37677 , \37682 );
and \U$37485 ( \37800 , \37673 , \37682 );
or \U$37486 ( \37801 , \37798 , \37799 , \37800 );
xor \U$37487 ( \37802 , \37797 , \37801 );
and \U$37488 ( \37803 , \37658 , \37662 );
and \U$37489 ( \37804 , \37662 , \37667 );
and \U$37490 ( \37805 , \37658 , \37667 );
or \U$37491 ( \37806 , \37803 , \37804 , \37805 );
xor \U$37492 ( \37807 , \37802 , \37806 );
xor \U$37493 ( \37808 , \37793 , \37807 );
and \U$37494 ( \37809 , \37654 , \37668 );
and \U$37495 ( \37810 , \37668 , \37683 );
and \U$37496 ( \37811 , \37654 , \37683 );
or \U$37497 ( \37812 , \37809 , \37810 , \37811 );
and \U$37498 ( \37813 , \22418 , \22208 );
and \U$37499 ( \37814 , \22386 , \22206 );
nor \U$37500 ( \37815 , \37813 , \37814 );
xnor \U$37501 ( \37816 , \37815 , \22218 );
and \U$37502 ( \37817 , \22440 , \22230 );
and \U$37503 ( \37818 , \22407 , \22228 );
nor \U$37504 ( \37819 , \37817 , \37818 );
xnor \U$37505 ( \37820 , \37819 , \22240 );
xor \U$37506 ( \37821 , \37816 , \37820 );
and \U$37507 ( \37822 , \22468 , \22257 );
and \U$37508 ( \37823 , \22429 , \22255 );
nor \U$37509 ( \37824 , \37822 , \37823 );
xnor \U$37510 ( \37825 , \37824 , \22267 );
xor \U$37511 ( \37826 , \37821 , \37825 );
and \U$37512 ( \37827 , \22350 , \22140 );
and \U$37513 ( \37828 , \22318 , \22138 );
nor \U$37514 ( \37829 , \37827 , \37828 );
xnor \U$37515 ( \37830 , \37829 , \22150 );
and \U$37516 ( \37831 , \22372 , \22162 );
and \U$37517 ( \37832 , \22339 , \22160 );
nor \U$37518 ( \37833 , \37831 , \37832 );
xnor \U$37519 ( \37834 , \37833 , \22172 );
xor \U$37520 ( \37835 , \37830 , \37834 );
and \U$37521 ( \37836 , \22397 , \22187 );
and \U$37522 ( \37837 , \22361 , \22185 );
nor \U$37523 ( \37838 , \37836 , \37837 );
xnor \U$37524 ( \37839 , \37838 , \22197 );
xor \U$37525 ( \37840 , \37835 , \37839 );
xor \U$37526 ( \37841 , \37826 , \37840 );
and \U$37527 ( \37842 , \22283 , \22076 );
and \U$37528 ( \37843 , \22251 , \22073 );
nor \U$37529 ( \37844 , \37842 , \37843 );
xnor \U$37530 ( \37845 , \37844 , \22072 );
and \U$37531 ( \37846 , \22305 , \22095 );
and \U$37532 ( \37847 , \22272 , \22093 );
nor \U$37533 ( \37848 , \37846 , \37847 );
xnor \U$37534 ( \37849 , \37848 , \22105 );
xor \U$37535 ( \37850 , \37845 , \37849 );
and \U$37536 ( \37851 , \22329 , \22119 );
and \U$37537 ( \37852 , \22294 , \22117 );
nor \U$37538 ( \37853 , \37851 , \37852 );
xnor \U$37539 ( \37854 , \37853 , \22129 );
xor \U$37540 ( \37855 , \37850 , \37854 );
xor \U$37541 ( \37856 , \37841 , \37855 );
xor \U$37542 ( \37857 , \37812 , \37856 );
and \U$37543 ( \37858 , \22624 , \22413 );
and \U$37544 ( \37859 , \22592 , \22411 );
nor \U$37545 ( \37860 , \37858 , \37859 );
xnor \U$37546 ( \37861 , \37860 , \22423 );
and \U$37547 ( \37862 , \22646 , \22435 );
and \U$37548 ( \37863 , \22613 , \22433 );
nor \U$37549 ( \37864 , \37862 , \37863 );
xnor \U$37550 ( \37865 , \37864 , \22445 );
xor \U$37551 ( \37866 , \37861 , \37865 );
and \U$37552 ( \37867 , \22676 , \22463 );
and \U$37553 ( \37868 , \22635 , \22461 );
nor \U$37554 ( \37869 , \37867 , \37868 );
xnor \U$37555 ( \37870 , \37869 , \22473 );
xor \U$37556 ( \37871 , \37866 , \37870 );
and \U$37557 ( \37872 , \22556 , \22345 );
and \U$37558 ( \37873 , \22524 , \22343 );
nor \U$37559 ( \37874 , \37872 , \37873 );
xnor \U$37560 ( \37875 , \37874 , \22355 );
and \U$37561 ( \37876 , \22578 , \22367 );
and \U$37562 ( \37877 , \22545 , \22365 );
nor \U$37563 ( \37878 , \37876 , \37877 );
xnor \U$37564 ( \37879 , \37878 , \22377 );
xor \U$37565 ( \37880 , \37875 , \37879 );
and \U$37566 ( \37881 , \22603 , \22392 );
and \U$37567 ( \37882 , \22567 , \22390 );
nor \U$37568 ( \37883 , \37881 , \37882 );
xnor \U$37569 ( \37884 , \37883 , \22402 );
xor \U$37570 ( \37885 , \37880 , \37884 );
xor \U$37571 ( \37886 , \37871 , \37885 );
and \U$37572 ( \37887 , \22489 , \22278 );
and \U$37573 ( \37888 , \22457 , \22276 );
nor \U$37574 ( \37889 , \37887 , \37888 );
xnor \U$37575 ( \37890 , \37889 , \22288 );
and \U$37576 ( \37891 , \22511 , \22300 );
and \U$37577 ( \37892 , \22478 , \22298 );
nor \U$37578 ( \37893 , \37891 , \37892 );
xnor \U$37579 ( \37894 , \37893 , \22310 );
xor \U$37580 ( \37895 , \37890 , \37894 );
and \U$37581 ( \37896 , \22535 , \22324 );
and \U$37582 ( \37897 , \22500 , \22322 );
nor \U$37583 ( \37898 , \37896 , \37897 );
xnor \U$37584 ( \37899 , \37898 , \22334 );
xor \U$37585 ( \37900 , \37895 , \37899 );
xor \U$37586 ( \37901 , \37886 , \37900 );
xor \U$37587 ( \37902 , \37857 , \37901 );
xor \U$37588 ( \37903 , \37808 , \37902 );
and \U$37589 ( \37904 , \37614 , \37618 );
and \U$37590 ( \37905 , \37618 , \37623 );
and \U$37591 ( \37906 , \37614 , \37623 );
or \U$37592 ( \37907 , \37904 , \37905 , \37906 );
and \U$37593 ( \37908 , \37599 , \37603 );
and \U$37594 ( \37909 , \37603 , \37608 );
and \U$37595 ( \37910 , \37599 , \37608 );
or \U$37596 ( \37911 , \37908 , \37909 , \37910 );
xor \U$37597 ( \37912 , \37907 , \37911 );
and \U$37598 ( \37913 , \37565 , \37579 );
and \U$37599 ( \37914 , \37579 , \37594 );
and \U$37600 ( \37915 , \37565 , \37594 );
or \U$37601 ( \37916 , \37913 , \37914 , \37915 );
xor \U$37602 ( \37917 , \37912 , \37916 );
xor \U$37603 ( \37918 , \37903 , \37917 );
xor \U$37604 ( \37919 , \37764 , \37918 );
xor \U$37605 ( \37920 , \37755 , \37919 );
xor \U$37606 ( \37921 , \37736 , \37920 );
and \U$37607 ( \37922 , \37702 , \37723 );
nor \U$37608 ( \37923 , \37921 , \37922 );
and \U$37609 ( \37924 , \37740 , \37754 );
and \U$37610 ( \37925 , \37754 , \37919 );
and \U$37611 ( \37926 , \37740 , \37919 );
or \U$37612 ( \37927 , \37924 , \37925 , \37926 );
and \U$37613 ( \37928 , \37759 , \37763 );
and \U$37614 ( \37929 , \37763 , \37918 );
and \U$37615 ( \37930 , \37759 , \37918 );
or \U$37616 ( \37931 , \37928 , \37929 , \37930 );
and \U$37617 ( \37932 , \37797 , \37801 );
and \U$37618 ( \37933 , \37801 , \37806 );
and \U$37619 ( \37934 , \37797 , \37806 );
or \U$37620 ( \37935 , \37932 , \37933 , \37934 );
and \U$37621 ( \37936 , \37782 , \37786 );
and \U$37622 ( \37937 , \37786 , \37791 );
and \U$37623 ( \37938 , \37782 , \37791 );
or \U$37624 ( \37939 , \37936 , \37937 , \37938 );
xor \U$37625 ( \37940 , \37935 , \37939 );
and \U$37626 ( \37941 , \37768 , \37772 );
and \U$37627 ( \37942 , \37772 , \37777 );
and \U$37628 ( \37943 , \37768 , \37777 );
or \U$37629 ( \37944 , \37941 , \37942 , \37943 );
xor \U$37630 ( \37945 , \37940 , \37944 );
and \U$37631 ( \37946 , \37890 , \37894 );
and \U$37632 ( \37947 , \37894 , \37899 );
and \U$37633 ( \37948 , \37890 , \37899 );
or \U$37634 ( \37949 , \37946 , \37947 , \37948 );
and \U$37635 ( \37950 , \37875 , \37879 );
and \U$37636 ( \37951 , \37879 , \37884 );
and \U$37637 ( \37952 , \37875 , \37884 );
or \U$37638 ( \37953 , \37950 , \37951 , \37952 );
xor \U$37639 ( \37954 , \37949 , \37953 );
and \U$37640 ( \37955 , \37861 , \37865 );
and \U$37641 ( \37956 , \37865 , \37870 );
and \U$37642 ( \37957 , \37861 , \37870 );
or \U$37643 ( \37958 , \37955 , \37956 , \37957 );
xor \U$37644 ( \37959 , \37954 , \37958 );
and \U$37645 ( \37960 , \37845 , \37849 );
and \U$37646 ( \37961 , \37849 , \37854 );
and \U$37647 ( \37962 , \37845 , \37854 );
or \U$37648 ( \37963 , \37960 , \37961 , \37962 );
and \U$37649 ( \37964 , \37830 , \37834 );
and \U$37650 ( \37965 , \37834 , \37839 );
and \U$37651 ( \37966 , \37830 , \37839 );
or \U$37652 ( \37967 , \37964 , \37965 , \37966 );
xor \U$37653 ( \37968 , \37963 , \37967 );
and \U$37654 ( \37969 , \37816 , \37820 );
and \U$37655 ( \37970 , \37820 , \37825 );
and \U$37656 ( \37971 , \37816 , \37825 );
or \U$37657 ( \37972 , \37969 , \37970 , \37971 );
xor \U$37658 ( \37973 , \37968 , \37972 );
xor \U$37659 ( \37974 , \37959 , \37973 );
and \U$37660 ( \37975 , \22251 , \22076 );
and \U$37661 ( \37976 , \22262 , \22073 );
nor \U$37662 ( \37977 , \37975 , \37976 );
xnor \U$37663 ( \37978 , \37977 , \22072 );
xor \U$37664 ( \37979 , \22540 , \37978 );
and \U$37665 ( \37980 , \22272 , \22095 );
and \U$37666 ( \37981 , \22283 , \22093 );
nor \U$37667 ( \37982 , \37980 , \37981 );
xnor \U$37668 ( \37983 , \37982 , \22105 );
xor \U$37669 ( \37984 , \37979 , \37983 );
and \U$37670 ( \37985 , \22500 , \22324 );
and \U$37671 ( \37986 , \22511 , \22322 );
nor \U$37672 ( \37987 , \37985 , \37986 );
xnor \U$37673 ( \37988 , \37987 , \22334 );
and \U$37674 ( \37989 , \22524 , \22345 );
and \U$37675 ( \37990 , \22535 , \22343 );
nor \U$37676 ( \37991 , \37989 , \37990 );
xnor \U$37677 ( \37992 , \37991 , \22355 );
xor \U$37678 ( \37993 , \37988 , \37992 );
and \U$37679 ( \37994 , \22545 , \22367 );
and \U$37680 ( \37995 , \22556 , \22365 );
nor \U$37681 ( \37996 , \37994 , \37995 );
xnor \U$37682 ( \37997 , \37996 , \22377 );
xor \U$37683 ( \37998 , \37993 , \37997 );
and \U$37684 ( \37999 , \22429 , \22257 );
and \U$37685 ( \38000 , \22440 , \22255 );
nor \U$37686 ( \38001 , \37999 , \38000 );
xnor \U$37687 ( \38002 , \38001 , \22267 );
and \U$37688 ( \38003 , \22457 , \22278 );
and \U$37689 ( \38004 , \22468 , \22276 );
nor \U$37690 ( \38005 , \38003 , \38004 );
xnor \U$37691 ( \38006 , \38005 , \22288 );
xor \U$37692 ( \38007 , \38002 , \38006 );
and \U$37693 ( \38008 , \22478 , \22300 );
and \U$37694 ( \38009 , \22489 , \22298 );
nor \U$37695 ( \38010 , \38008 , \38009 );
xnor \U$37696 ( \38011 , \38010 , \22310 );
xor \U$37697 ( \38012 , \38007 , \38011 );
xor \U$37698 ( \38013 , \37998 , \38012 );
and \U$37699 ( \38014 , \22361 , \22187 );
and \U$37700 ( \38015 , \22372 , \22185 );
nor \U$37701 ( \38016 , \38014 , \38015 );
xnor \U$37702 ( \38017 , \38016 , \22197 );
and \U$37703 ( \38018 , \22386 , \22208 );
and \U$37704 ( \38019 , \22397 , \22206 );
nor \U$37705 ( \38020 , \38018 , \38019 );
xnor \U$37706 ( \38021 , \38020 , \22218 );
xor \U$37707 ( \38022 , \38017 , \38021 );
and \U$37708 ( \38023 , \22407 , \22230 );
and \U$37709 ( \38024 , \22418 , \22228 );
nor \U$37710 ( \38025 , \38023 , \38024 );
xnor \U$37711 ( \38026 , \38025 , \22240 );
xor \U$37712 ( \38027 , \38022 , \38026 );
xor \U$37713 ( \38028 , \38013 , \38027 );
xor \U$37714 ( \38029 , \37984 , \38028 );
nand \U$37715 ( \38030 , \22706 , \22528 );
xnor \U$37716 ( \38031 , \38030 , \22540 );
and \U$37717 ( \38032 , \22635 , \22463 );
and \U$37718 ( \38033 , \22646 , \22461 );
nor \U$37719 ( \38034 , \38032 , \38033 );
xnor \U$37720 ( \38035 , \38034 , \22473 );
and \U$37721 ( \38036 , \22665 , \22484 );
and \U$37722 ( \38037 , \22676 , \22482 );
nor \U$37723 ( \38038 , \38036 , \38037 );
xnor \U$37724 ( \38039 , \38038 , \22494 );
xor \U$37725 ( \38040 , \38035 , \38039 );
and \U$37726 ( \38041 , \22686 , \22506 );
and \U$37727 ( \38042 , \22696 , \22504 );
nor \U$37728 ( \38043 , \38041 , \38042 );
xnor \U$37729 ( \38044 , \38043 , \22516 );
xor \U$37730 ( \38045 , \38040 , \38044 );
xor \U$37731 ( \38046 , \38031 , \38045 );
and \U$37732 ( \38047 , \22567 , \22392 );
and \U$37733 ( \38048 , \22578 , \22390 );
nor \U$37734 ( \38049 , \38047 , \38048 );
xnor \U$37735 ( \38050 , \38049 , \22402 );
and \U$37736 ( \38051 , \22592 , \22413 );
and \U$37737 ( \38052 , \22603 , \22411 );
nor \U$37738 ( \38053 , \38051 , \38052 );
xnor \U$37739 ( \38054 , \38053 , \22423 );
xor \U$37740 ( \38055 , \38050 , \38054 );
and \U$37741 ( \38056 , \22613 , \22435 );
and \U$37742 ( \38057 , \22624 , \22433 );
nor \U$37743 ( \38058 , \38056 , \38057 );
xnor \U$37744 ( \38059 , \38058 , \22445 );
xor \U$37745 ( \38060 , \38055 , \38059 );
xor \U$37746 ( \38061 , \38046 , \38060 );
xor \U$37747 ( \38062 , \38029 , \38061 );
xor \U$37748 ( \38063 , \37974 , \38062 );
xor \U$37749 ( \38064 , \37945 , \38063 );
and \U$37750 ( \38065 , \37907 , \37911 );
and \U$37751 ( \38066 , \37911 , \37916 );
and \U$37752 ( \38067 , \37907 , \37916 );
or \U$37753 ( \38068 , \38065 , \38066 , \38067 );
and \U$37754 ( \38069 , \37812 , \37856 );
and \U$37755 ( \38070 , \37856 , \37901 );
and \U$37756 ( \38071 , \37812 , \37901 );
or \U$37757 ( \38072 , \38069 , \38070 , \38071 );
xor \U$37758 ( \38073 , \38068 , \38072 );
and \U$37759 ( \38074 , \37778 , \37792 );
and \U$37760 ( \38075 , \37792 , \37807 );
and \U$37761 ( \38076 , \37778 , \37807 );
or \U$37762 ( \38077 , \38074 , \38075 , \38076 );
xor \U$37763 ( \38078 , \38073 , \38077 );
xor \U$37764 ( \38079 , \38064 , \38078 );
xor \U$37765 ( \38080 , \37931 , \38079 );
and \U$37766 ( \38081 , \37744 , \37748 );
and \U$37767 ( \38082 , \37748 , \37753 );
and \U$37768 ( \38083 , \37744 , \37753 );
or \U$37769 ( \38084 , \38081 , \38082 , \38083 );
and \U$37770 ( \38085 , \37808 , \37902 );
and \U$37771 ( \38086 , \37902 , \37917 );
and \U$37772 ( \38087 , \37808 , \37917 );
or \U$37773 ( \38088 , \38085 , \38086 , \38087 );
xor \U$37774 ( \38089 , \38084 , \38088 );
and \U$37775 ( \38090 , \37871 , \37885 );
and \U$37776 ( \38091 , \37885 , \37900 );
and \U$37777 ( \38092 , \37871 , \37900 );
or \U$37778 ( \38093 , \38090 , \38091 , \38092 );
and \U$37779 ( \38094 , \37826 , \37840 );
and \U$37780 ( \38095 , \37840 , \37855 );
and \U$37781 ( \38096 , \37826 , \37855 );
or \U$37782 ( \38097 , \38094 , \38095 , \38096 );
xor \U$37783 ( \38098 , \38093 , \38097 );
and \U$37784 ( \38099 , \22294 , \22119 );
and \U$37785 ( \38100 , \22305 , \22117 );
nor \U$37786 ( \38101 , \38099 , \38100 );
xnor \U$37787 ( \38102 , \38101 , \22129 );
and \U$37788 ( \38103 , \22318 , \22140 );
and \U$37789 ( \38104 , \22329 , \22138 );
nor \U$37790 ( \38105 , \38103 , \38104 );
xnor \U$37791 ( \38106 , \38105 , \22150 );
xor \U$37792 ( \38107 , \38102 , \38106 );
and \U$37793 ( \38108 , \22339 , \22162 );
and \U$37794 ( \38109 , \22350 , \22160 );
nor \U$37795 ( \38110 , \38108 , \38109 );
xnor \U$37796 ( \38111 , \38110 , \22172 );
xor \U$37797 ( \38112 , \38107 , \38111 );
xor \U$37798 ( \38113 , \38098 , \38112 );
xor \U$37799 ( \38114 , \38089 , \38113 );
xor \U$37800 ( \38115 , \38080 , \38114 );
xor \U$37801 ( \38116 , \37927 , \38115 );
and \U$37802 ( \38117 , \37736 , \37920 );
nor \U$37803 ( \38118 , \38116 , \38117 );
nor \U$37804 ( \38119 , \37923 , \38118 );
and \U$37805 ( \38120 , \37931 , \38079 );
and \U$37806 ( \38121 , \38079 , \38114 );
and \U$37807 ( \38122 , \37931 , \38114 );
or \U$37808 ( \38123 , \38120 , \38121 , \38122 );
and \U$37809 ( \38124 , \38068 , \38072 );
and \U$37810 ( \38125 , \38072 , \38077 );
and \U$37811 ( \38126 , \38068 , \38077 );
or \U$37812 ( \38127 , \38124 , \38125 , \38126 );
and \U$37813 ( \38128 , \37959 , \37973 );
and \U$37814 ( \38129 , \37973 , \38062 );
and \U$37815 ( \38130 , \37959 , \38062 );
or \U$37816 ( \38131 , \38128 , \38129 , \38130 );
xor \U$37817 ( \38132 , \38127 , \38131 );
and \U$37818 ( \38133 , \38035 , \38039 );
and \U$37819 ( \38134 , \38039 , \38044 );
and \U$37820 ( \38135 , \38035 , \38044 );
or \U$37821 ( \38136 , \38133 , \38134 , \38135 );
and \U$37822 ( \38137 , \22676 , \22484 );
and \U$37823 ( \38138 , \22635 , \22482 );
nor \U$37824 ( \38139 , \38137 , \38138 );
xnor \U$37825 ( \38140 , \38139 , \22494 );
and \U$37826 ( \38141 , \22696 , \22506 );
and \U$37827 ( \38142 , \22665 , \22504 );
nor \U$37828 ( \38143 , \38141 , \38142 );
xnor \U$37829 ( \38144 , \38143 , \22516 );
xor \U$37830 ( \38145 , \38140 , \38144 );
and \U$37831 ( \38146 , \22706 , \22530 );
and \U$37832 ( \38147 , \22686 , \22528 );
nor \U$37833 ( \38148 , \38146 , \38147 );
xnor \U$37834 ( \38149 , \38148 , \22540 );
xor \U$37835 ( \38150 , \38145 , \38149 );
xor \U$37836 ( \38151 , \38136 , \38150 );
and \U$37837 ( \38152 , \22603 , \22413 );
and \U$37838 ( \38153 , \22567 , \22411 );
nor \U$37839 ( \38154 , \38152 , \38153 );
xnor \U$37840 ( \38155 , \38154 , \22423 );
and \U$37841 ( \38156 , \22624 , \22435 );
and \U$37842 ( \38157 , \22592 , \22433 );
nor \U$37843 ( \38158 , \38156 , \38157 );
xnor \U$37844 ( \38159 , \38158 , \22445 );
xor \U$37845 ( \38160 , \38155 , \38159 );
and \U$37846 ( \38161 , \22646 , \22463 );
and \U$37847 ( \38162 , \22613 , \22461 );
nor \U$37848 ( \38163 , \38161 , \38162 );
xnor \U$37849 ( \38164 , \38163 , \22473 );
xor \U$37850 ( \38165 , \38160 , \38164 );
xor \U$37851 ( \38166 , \38151 , \38165 );
and \U$37852 ( \38167 , \38002 , \38006 );
and \U$37853 ( \38168 , \38006 , \38011 );
and \U$37854 ( \38169 , \38002 , \38011 );
or \U$37855 ( \38170 , \38167 , \38168 , \38169 );
and \U$37856 ( \38171 , \37988 , \37992 );
and \U$37857 ( \38172 , \37992 , \37997 );
and \U$37858 ( \38173 , \37988 , \37997 );
or \U$37859 ( \38174 , \38171 , \38172 , \38173 );
xor \U$37860 ( \38175 , \38170 , \38174 );
and \U$37861 ( \38176 , \38050 , \38054 );
and \U$37862 ( \38177 , \38054 , \38059 );
and \U$37863 ( \38178 , \38050 , \38059 );
or \U$37864 ( \38179 , \38176 , \38177 , \38178 );
xor \U$37865 ( \38180 , \38175 , \38179 );
xor \U$37866 ( \38181 , \38166 , \38180 );
and \U$37867 ( \38182 , \22540 , \37978 );
and \U$37868 ( \38183 , \37978 , \37983 );
and \U$37869 ( \38184 , \22540 , \37983 );
or \U$37870 ( \38185 , \38182 , \38183 , \38184 );
and \U$37871 ( \38186 , \38102 , \38106 );
and \U$37872 ( \38187 , \38106 , \38111 );
and \U$37873 ( \38188 , \38102 , \38111 );
or \U$37874 ( \38189 , \38186 , \38187 , \38188 );
xor \U$37875 ( \38190 , \38185 , \38189 );
and \U$37876 ( \38191 , \38017 , \38021 );
and \U$37877 ( \38192 , \38021 , \38026 );
and \U$37878 ( \38193 , \38017 , \38026 );
or \U$37879 ( \38194 , \38191 , \38192 , \38193 );
xor \U$37880 ( \38195 , \38190 , \38194 );
xor \U$37881 ( \38196 , \38181 , \38195 );
and \U$37882 ( \38197 , \37998 , \38012 );
and \U$37883 ( \38198 , \38012 , \38027 );
and \U$37884 ( \38199 , \37998 , \38027 );
or \U$37885 ( \38200 , \38197 , \38198 , \38199 );
and \U$37886 ( \38201 , \22329 , \22140 );
and \U$37887 ( \38202 , \22294 , \22138 );
nor \U$37888 ( \38203 , \38201 , \38202 );
xnor \U$37889 ( \38204 , \38203 , \22150 );
and \U$37890 ( \38205 , \22350 , \22162 );
and \U$37891 ( \38206 , \22318 , \22160 );
nor \U$37892 ( \38207 , \38205 , \38206 );
xnor \U$37893 ( \38208 , \38207 , \22172 );
xor \U$37894 ( \38209 , \38204 , \38208 );
and \U$37895 ( \38210 , \22372 , \22187 );
and \U$37896 ( \38211 , \22339 , \22185 );
nor \U$37897 ( \38212 , \38210 , \38211 );
xnor \U$37898 ( \38213 , \38212 , \22197 );
xor \U$37899 ( \38214 , \38209 , \38213 );
and \U$37900 ( \38215 , \22262 , \22076 );
and \U$37901 ( \38216 , \22224 , \22073 );
nor \U$37902 ( \38217 , \38215 , \38216 );
xnor \U$37903 ( \38218 , \38217 , \22072 );
and \U$37904 ( \38219 , \22283 , \22095 );
and \U$37905 ( \38220 , \22251 , \22093 );
nor \U$37906 ( \38221 , \38219 , \38220 );
xnor \U$37907 ( \38222 , \38221 , \22105 );
xor \U$37908 ( \38223 , \38218 , \38222 );
and \U$37909 ( \38224 , \22305 , \22119 );
and \U$37910 ( \38225 , \22272 , \22117 );
nor \U$37911 ( \38226 , \38224 , \38225 );
xnor \U$37912 ( \38227 , \38226 , \22129 );
xor \U$37913 ( \38228 , \38223 , \38227 );
xor \U$37914 ( \38229 , \38214 , \38228 );
xor \U$37915 ( \38230 , \38200 , \38229 );
and \U$37916 ( \38231 , \22535 , \22345 );
and \U$37917 ( \38232 , \22500 , \22343 );
nor \U$37918 ( \38233 , \38231 , \38232 );
xnor \U$37919 ( \38234 , \38233 , \22355 );
and \U$37920 ( \38235 , \22556 , \22367 );
and \U$37921 ( \38236 , \22524 , \22365 );
nor \U$37922 ( \38237 , \38235 , \38236 );
xnor \U$37923 ( \38238 , \38237 , \22377 );
xor \U$37924 ( \38239 , \38234 , \38238 );
and \U$37925 ( \38240 , \22578 , \22392 );
and \U$37926 ( \38241 , \22545 , \22390 );
nor \U$37927 ( \38242 , \38240 , \38241 );
xnor \U$37928 ( \38243 , \38242 , \22402 );
xor \U$37929 ( \38244 , \38239 , \38243 );
and \U$37930 ( \38245 , \22468 , \22278 );
and \U$37931 ( \38246 , \22429 , \22276 );
nor \U$37932 ( \38247 , \38245 , \38246 );
xnor \U$37933 ( \38248 , \38247 , \22288 );
and \U$37934 ( \38249 , \22489 , \22300 );
and \U$37935 ( \38250 , \22457 , \22298 );
nor \U$37936 ( \38251 , \38249 , \38250 );
xnor \U$37937 ( \38252 , \38251 , \22310 );
xor \U$37938 ( \38253 , \38248 , \38252 );
and \U$37939 ( \38254 , \22511 , \22324 );
and \U$37940 ( \38255 , \22478 , \22322 );
nor \U$37941 ( \38256 , \38254 , \38255 );
xnor \U$37942 ( \38257 , \38256 , \22334 );
xor \U$37943 ( \38258 , \38253 , \38257 );
xor \U$37944 ( \38259 , \38244 , \38258 );
and \U$37945 ( \38260 , \22397 , \22208 );
and \U$37946 ( \38261 , \22361 , \22206 );
nor \U$37947 ( \38262 , \38260 , \38261 );
xnor \U$37948 ( \38263 , \38262 , \22218 );
and \U$37949 ( \38264 , \22418 , \22230 );
and \U$37950 ( \38265 , \22386 , \22228 );
nor \U$37951 ( \38266 , \38264 , \38265 );
xnor \U$37952 ( \38267 , \38266 , \22240 );
xor \U$37953 ( \38268 , \38263 , \38267 );
and \U$37954 ( \38269 , \22440 , \22257 );
and \U$37955 ( \38270 , \22407 , \22255 );
nor \U$37956 ( \38271 , \38269 , \38270 );
xnor \U$37957 ( \38272 , \38271 , \22267 );
xor \U$37958 ( \38273 , \38268 , \38272 );
xor \U$37959 ( \38274 , \38259 , \38273 );
xor \U$37960 ( \38275 , \38230 , \38274 );
xor \U$37961 ( \38276 , \38196 , \38275 );
and \U$37962 ( \38277 , \37963 , \37967 );
and \U$37963 ( \38278 , \37967 , \37972 );
and \U$37964 ( \38279 , \37963 , \37972 );
or \U$37965 ( \38280 , \38277 , \38278 , \38279 );
and \U$37966 ( \38281 , \37949 , \37953 );
and \U$37967 ( \38282 , \37953 , \37958 );
and \U$37968 ( \38283 , \37949 , \37958 );
or \U$37969 ( \38284 , \38281 , \38282 , \38283 );
xor \U$37970 ( \38285 , \38280 , \38284 );
and \U$37971 ( \38286 , \38031 , \38045 );
and \U$37972 ( \38287 , \38045 , \38060 );
and \U$37973 ( \38288 , \38031 , \38060 );
or \U$37974 ( \38289 , \38286 , \38287 , \38288 );
xor \U$37975 ( \38290 , \38285 , \38289 );
xor \U$37976 ( \38291 , \38276 , \38290 );
xor \U$37977 ( \38292 , \38132 , \38291 );
xor \U$37978 ( \38293 , \38123 , \38292 );
and \U$37979 ( \38294 , \38084 , \38088 );
and \U$37980 ( \38295 , \38088 , \38113 );
and \U$37981 ( \38296 , \38084 , \38113 );
or \U$37982 ( \38297 , \38294 , \38295 , \38296 );
and \U$37983 ( \38298 , \37945 , \38063 );
and \U$37984 ( \38299 , \38063 , \38078 );
and \U$37985 ( \38300 , \37945 , \38078 );
or \U$37986 ( \38301 , \38298 , \38299 , \38300 );
xor \U$37987 ( \38302 , \38297 , \38301 );
and \U$37988 ( \38303 , \37935 , \37939 );
and \U$37989 ( \38304 , \37939 , \37944 );
and \U$37990 ( \38305 , \37935 , \37944 );
or \U$37991 ( \38306 , \38303 , \38304 , \38305 );
and \U$37992 ( \38307 , \38093 , \38097 );
and \U$37993 ( \38308 , \38097 , \38112 );
and \U$37994 ( \38309 , \38093 , \38112 );
or \U$37995 ( \38310 , \38307 , \38308 , \38309 );
xor \U$37996 ( \38311 , \38306 , \38310 );
and \U$37997 ( \38312 , \37984 , \38028 );
and \U$37998 ( \38313 , \38028 , \38061 );
and \U$37999 ( \38314 , \37984 , \38061 );
or \U$38000 ( \38315 , \38312 , \38313 , \38314 );
xor \U$38001 ( \38316 , \38311 , \38315 );
xor \U$38002 ( \38317 , \38302 , \38316 );
xor \U$38003 ( \38318 , \38293 , \38317 );
and \U$38004 ( \38319 , \37927 , \38115 );
nor \U$38005 ( \38320 , \38318 , \38319 );
and \U$38006 ( \38321 , \38297 , \38301 );
and \U$38007 ( \38322 , \38301 , \38316 );
and \U$38008 ( \38323 , \38297 , \38316 );
or \U$38009 ( \38324 , \38321 , \38322 , \38323 );
and \U$38010 ( \38325 , \38127 , \38131 );
and \U$38011 ( \38326 , \38131 , \38291 );
and \U$38012 ( \38327 , \38127 , \38291 );
or \U$38013 ( \38328 , \38325 , \38326 , \38327 );
and \U$38014 ( \38329 , \38218 , \38222 );
and \U$38015 ( \38330 , \38222 , \38227 );
and \U$38016 ( \38331 , \38218 , \38227 );
or \U$38017 ( \38332 , \38329 , \38330 , \38331 );
and \U$38018 ( \38333 , \38204 , \38208 );
and \U$38019 ( \38334 , \38208 , \38213 );
and \U$38020 ( \38335 , \38204 , \38213 );
or \U$38021 ( \38336 , \38333 , \38334 , \38335 );
xor \U$38022 ( \38337 , \38332 , \38336 );
and \U$38023 ( \38338 , \38263 , \38267 );
and \U$38024 ( \38339 , \38267 , \38272 );
and \U$38025 ( \38340 , \38263 , \38272 );
or \U$38026 ( \38341 , \38338 , \38339 , \38340 );
xor \U$38027 ( \38342 , \38337 , \38341 );
and \U$38028 ( \38343 , \22545 , \22392 );
and \U$38029 ( \38344 , \22556 , \22390 );
nor \U$38030 ( \38345 , \38343 , \38344 );
xnor \U$38031 ( \38346 , \38345 , \22402 );
and \U$38032 ( \38347 , \22567 , \22413 );
and \U$38033 ( \38348 , \22578 , \22411 );
nor \U$38034 ( \38349 , \38347 , \38348 );
xnor \U$38035 ( \38350 , \38349 , \22423 );
xor \U$38036 ( \38351 , \38346 , \38350 );
and \U$38037 ( \38352 , \22592 , \22435 );
and \U$38038 ( \38353 , \22603 , \22433 );
nor \U$38039 ( \38354 , \38352 , \38353 );
xnor \U$38040 ( \38355 , \38354 , \22445 );
xor \U$38041 ( \38356 , \38351 , \38355 );
and \U$38042 ( \38357 , \22478 , \22324 );
and \U$38043 ( \38358 , \22489 , \22322 );
nor \U$38044 ( \38359 , \38357 , \38358 );
xnor \U$38045 ( \38360 , \38359 , \22334 );
and \U$38046 ( \38361 , \22500 , \22345 );
and \U$38047 ( \38362 , \22511 , \22343 );
nor \U$38048 ( \38363 , \38361 , \38362 );
xnor \U$38049 ( \38364 , \38363 , \22355 );
xor \U$38050 ( \38365 , \38360 , \38364 );
and \U$38051 ( \38366 , \22524 , \22367 );
and \U$38052 ( \38367 , \22535 , \22365 );
nor \U$38053 ( \38368 , \38366 , \38367 );
xnor \U$38054 ( \38369 , \38368 , \22377 );
xor \U$38055 ( \38370 , \38365 , \38369 );
xor \U$38056 ( \38371 , \38356 , \38370 );
and \U$38057 ( \38372 , \22407 , \22257 );
and \U$38058 ( \38373 , \22418 , \22255 );
nor \U$38059 ( \38374 , \38372 , \38373 );
xnor \U$38060 ( \38375 , \38374 , \22267 );
and \U$38061 ( \38376 , \22429 , \22278 );
and \U$38062 ( \38377 , \22440 , \22276 );
nor \U$38063 ( \38378 , \38376 , \38377 );
xnor \U$38064 ( \38379 , \38378 , \22288 );
xor \U$38065 ( \38380 , \38375 , \38379 );
and \U$38066 ( \38381 , \22457 , \22300 );
and \U$38067 ( \38382 , \22468 , \22298 );
nor \U$38068 ( \38383 , \38381 , \38382 );
xnor \U$38069 ( \38384 , \38383 , \22310 );
xor \U$38070 ( \38385 , \38380 , \38384 );
xor \U$38071 ( \38386 , \38371 , \38385 );
and \U$38072 ( \38387 , \38140 , \38144 );
and \U$38073 ( \38388 , \38144 , \38149 );
and \U$38074 ( \38389 , \38140 , \38149 );
or \U$38075 ( \38390 , \38387 , \38388 , \38389 );
and \U$38076 ( \38391 , \22686 , \22530 );
and \U$38077 ( \38392 , \22696 , \22528 );
nor \U$38078 ( \38393 , \38391 , \38392 );
xnor \U$38079 ( \38394 , \38393 , \22540 );
nand \U$38080 ( \38395 , \22706 , \22549 );
xnor \U$38081 ( \38396 , \38395 , \22561 );
xor \U$38082 ( \38397 , \38394 , \38396 );
xor \U$38083 ( \38398 , \38390 , \38397 );
and \U$38084 ( \38399 , \22613 , \22463 );
and \U$38085 ( \38400 , \22624 , \22461 );
nor \U$38086 ( \38401 , \38399 , \38400 );
xnor \U$38087 ( \38402 , \38401 , \22473 );
and \U$38088 ( \38403 , \22635 , \22484 );
and \U$38089 ( \38404 , \22646 , \22482 );
nor \U$38090 ( \38405 , \38403 , \38404 );
xnor \U$38091 ( \38406 , \38405 , \22494 );
xor \U$38092 ( \38407 , \38402 , \38406 );
and \U$38093 ( \38408 , \22665 , \22506 );
and \U$38094 ( \38409 , \22676 , \22504 );
nor \U$38095 ( \38410 , \38408 , \38409 );
xnor \U$38096 ( \38411 , \38410 , \22516 );
xor \U$38097 ( \38412 , \38407 , \38411 );
xor \U$38098 ( \38413 , \38398 , \38412 );
xor \U$38099 ( \38414 , \38386 , \38413 );
and \U$38100 ( \38415 , \38248 , \38252 );
and \U$38101 ( \38416 , \38252 , \38257 );
and \U$38102 ( \38417 , \38248 , \38257 );
or \U$38103 ( \38418 , \38415 , \38416 , \38417 );
and \U$38104 ( \38419 , \38234 , \38238 );
and \U$38105 ( \38420 , \38238 , \38243 );
and \U$38106 ( \38421 , \38234 , \38243 );
or \U$38107 ( \38422 , \38419 , \38420 , \38421 );
xor \U$38108 ( \38423 , \38418 , \38422 );
and \U$38109 ( \38424 , \38155 , \38159 );
and \U$38110 ( \38425 , \38159 , \38164 );
and \U$38111 ( \38426 , \38155 , \38164 );
or \U$38112 ( \38427 , \38424 , \38425 , \38426 );
xor \U$38113 ( \38428 , \38423 , \38427 );
xor \U$38114 ( \38429 , \38414 , \38428 );
xor \U$38115 ( \38430 , \38342 , \38429 );
and \U$38116 ( \38431 , \38244 , \38258 );
and \U$38117 ( \38432 , \38258 , \38273 );
and \U$38118 ( \38433 , \38244 , \38273 );
or \U$38119 ( \38434 , \38431 , \38432 , \38433 );
and \U$38120 ( \38435 , \38214 , \38228 );
xor \U$38121 ( \38436 , \38434 , \38435 );
and \U$38122 ( \38437 , \22339 , \22187 );
and \U$38123 ( \38438 , \22350 , \22185 );
nor \U$38124 ( \38439 , \38437 , \38438 );
xnor \U$38125 ( \38440 , \38439 , \22197 );
and \U$38126 ( \38441 , \22361 , \22208 );
and \U$38127 ( \38442 , \22372 , \22206 );
nor \U$38128 ( \38443 , \38441 , \38442 );
xnor \U$38129 ( \38444 , \38443 , \22218 );
xor \U$38130 ( \38445 , \38440 , \38444 );
and \U$38131 ( \38446 , \22386 , \22230 );
and \U$38132 ( \38447 , \22397 , \22228 );
nor \U$38133 ( \38448 , \38446 , \38447 );
xnor \U$38134 ( \38449 , \38448 , \22240 );
xor \U$38135 ( \38450 , \38445 , \38449 );
and \U$38136 ( \38451 , \22272 , \22119 );
and \U$38137 ( \38452 , \22283 , \22117 );
nor \U$38138 ( \38453 , \38451 , \38452 );
xnor \U$38139 ( \38454 , \38453 , \22129 );
and \U$38140 ( \38455 , \22294 , \22140 );
and \U$38141 ( \38456 , \22305 , \22138 );
nor \U$38142 ( \38457 , \38455 , \38456 );
xnor \U$38143 ( \38458 , \38457 , \22150 );
xor \U$38144 ( \38459 , \38454 , \38458 );
and \U$38145 ( \38460 , \22318 , \22162 );
and \U$38146 ( \38461 , \22329 , \22160 );
nor \U$38147 ( \38462 , \38460 , \38461 );
xnor \U$38148 ( \38463 , \38462 , \22172 );
xor \U$38149 ( \38464 , \38459 , \38463 );
xor \U$38150 ( \38465 , \38450 , \38464 );
and \U$38151 ( \38466 , \22224 , \22076 );
and \U$38152 ( \38467 , \22235 , \22073 );
nor \U$38153 ( \38468 , \38466 , \38467 );
xnor \U$38154 ( \38469 , \38468 , \22072 );
xor \U$38155 ( \38470 , \22561 , \38469 );
and \U$38156 ( \38471 , \22251 , \22095 );
and \U$38157 ( \38472 , \22262 , \22093 );
nor \U$38158 ( \38473 , \38471 , \38472 );
xnor \U$38159 ( \38474 , \38473 , \22105 );
xor \U$38160 ( \38475 , \38470 , \38474 );
xor \U$38161 ( \38476 , \38465 , \38475 );
xor \U$38162 ( \38477 , \38436 , \38476 );
xor \U$38163 ( \38478 , \38430 , \38477 );
and \U$38164 ( \38479 , \38280 , \38284 );
and \U$38165 ( \38480 , \38284 , \38289 );
and \U$38166 ( \38481 , \38280 , \38289 );
or \U$38167 ( \38482 , \38479 , \38480 , \38481 );
and \U$38168 ( \38483 , \38200 , \38229 );
and \U$38169 ( \38484 , \38229 , \38274 );
and \U$38170 ( \38485 , \38200 , \38274 );
or \U$38171 ( \38486 , \38483 , \38484 , \38485 );
xor \U$38172 ( \38487 , \38482 , \38486 );
and \U$38173 ( \38488 , \38166 , \38180 );
and \U$38174 ( \38489 , \38180 , \38195 );
and \U$38175 ( \38490 , \38166 , \38195 );
or \U$38176 ( \38491 , \38488 , \38489 , \38490 );
xor \U$38177 ( \38492 , \38487 , \38491 );
xor \U$38178 ( \38493 , \38478 , \38492 );
xor \U$38179 ( \38494 , \38328 , \38493 );
and \U$38180 ( \38495 , \38306 , \38310 );
and \U$38181 ( \38496 , \38310 , \38315 );
and \U$38182 ( \38497 , \38306 , \38315 );
or \U$38183 ( \38498 , \38495 , \38496 , \38497 );
and \U$38184 ( \38499 , \38196 , \38275 );
and \U$38185 ( \38500 , \38275 , \38290 );
and \U$38186 ( \38501 , \38196 , \38290 );
or \U$38187 ( \38502 , \38499 , \38500 , \38501 );
xor \U$38188 ( \38503 , \38498 , \38502 );
and \U$38189 ( \38504 , \38185 , \38189 );
and \U$38190 ( \38505 , \38189 , \38194 );
and \U$38191 ( \38506 , \38185 , \38194 );
or \U$38192 ( \38507 , \38504 , \38505 , \38506 );
and \U$38193 ( \38508 , \38170 , \38174 );
and \U$38194 ( \38509 , \38174 , \38179 );
and \U$38195 ( \38510 , \38170 , \38179 );
or \U$38196 ( \38511 , \38508 , \38509 , \38510 );
xor \U$38197 ( \38512 , \38507 , \38511 );
and \U$38198 ( \38513 , \38136 , \38150 );
and \U$38199 ( \38514 , \38150 , \38165 );
and \U$38200 ( \38515 , \38136 , \38165 );
or \U$38201 ( \38516 , \38513 , \38514 , \38515 );
xor \U$38202 ( \38517 , \38512 , \38516 );
xor \U$38203 ( \38518 , \38503 , \38517 );
xor \U$38204 ( \38519 , \38494 , \38518 );
xor \U$38205 ( \38520 , \38324 , \38519 );
and \U$38206 ( \38521 , \38123 , \38292 );
and \U$38207 ( \38522 , \38292 , \38317 );
and \U$38208 ( \38523 , \38123 , \38317 );
or \U$38209 ( \38524 , \38521 , \38522 , \38523 );
nor \U$38210 ( \38525 , \38520 , \38524 );
nor \U$38211 ( \38526 , \38320 , \38525 );
nand \U$38212 ( \38527 , \38119 , \38526 );
and \U$38213 ( \38528 , \38328 , \38493 );
and \U$38214 ( \38529 , \38493 , \38518 );
and \U$38215 ( \38530 , \38328 , \38518 );
or \U$38216 ( \38531 , \38528 , \38529 , \38530 );
and \U$38217 ( \38532 , \38482 , \38486 );
and \U$38218 ( \38533 , \38486 , \38491 );
and \U$38219 ( \38534 , \38482 , \38491 );
or \U$38220 ( \38535 , \38532 , \38533 , \38534 );
and \U$38221 ( \38536 , \38342 , \38429 );
and \U$38222 ( \38537 , \38429 , \38477 );
and \U$38223 ( \38538 , \38342 , \38477 );
or \U$38224 ( \38539 , \38536 , \38537 , \38538 );
xor \U$38225 ( \38540 , \38535 , \38539 );
and \U$38226 ( \38541 , \38356 , \38370 );
and \U$38227 ( \38542 , \38370 , \38385 );
and \U$38228 ( \38543 , \38356 , \38385 );
or \U$38229 ( \38544 , \38541 , \38542 , \38543 );
and \U$38230 ( \38545 , \38450 , \38464 );
and \U$38231 ( \38546 , \38464 , \38475 );
and \U$38232 ( \38547 , \38450 , \38475 );
or \U$38233 ( \38548 , \38545 , \38546 , \38547 );
xor \U$38234 ( \38549 , \38544 , \38548 );
and \U$38235 ( \38550 , \22235 , \22076 );
and \U$38236 ( \38551 , \22202 , \22073 );
nor \U$38237 ( \38552 , \38550 , \38551 );
xnor \U$38238 ( \38553 , \38552 , \22072 );
and \U$38239 ( \38554 , \22262 , \22095 );
and \U$38240 ( \38555 , \22224 , \22093 );
nor \U$38241 ( \38556 , \38554 , \38555 );
xnor \U$38242 ( \38557 , \38556 , \22105 );
xor \U$38243 ( \38558 , \38553 , \38557 );
and \U$38244 ( \38559 , \22283 , \22119 );
and \U$38245 ( \38560 , \22251 , \22117 );
nor \U$38246 ( \38561 , \38559 , \38560 );
xnor \U$38247 ( \38562 , \38561 , \22129 );
xor \U$38248 ( \38563 , \38558 , \38562 );
xor \U$38249 ( \38564 , \38549 , \38563 );
xor \U$38250 ( \38565 , \38540 , \38564 );
xor \U$38251 ( \38566 , \38531 , \38565 );
and \U$38252 ( \38567 , \38498 , \38502 );
and \U$38253 ( \38568 , \38502 , \38517 );
and \U$38254 ( \38569 , \38498 , \38517 );
or \U$38255 ( \38570 , \38567 , \38568 , \38569 );
and \U$38256 ( \38571 , \38478 , \38492 );
xor \U$38257 ( \38572 , \38570 , \38571 );
and \U$38258 ( \38573 , \38332 , \38336 );
and \U$38259 ( \38574 , \38336 , \38341 );
and \U$38260 ( \38575 , \38332 , \38341 );
or \U$38261 ( \38576 , \38573 , \38574 , \38575 );
and \U$38262 ( \38577 , \38418 , \38422 );
and \U$38263 ( \38578 , \38422 , \38427 );
and \U$38264 ( \38579 , \38418 , \38427 );
or \U$38265 ( \38580 , \38577 , \38578 , \38579 );
xor \U$38266 ( \38581 , \38576 , \38580 );
and \U$38267 ( \38582 , \38390 , \38397 );
and \U$38268 ( \38583 , \38397 , \38412 );
and \U$38269 ( \38584 , \38390 , \38412 );
or \U$38270 ( \38585 , \38582 , \38583 , \38584 );
xor \U$38271 ( \38586 , \38581 , \38585 );
and \U$38272 ( \38587 , \38375 , \38379 );
and \U$38273 ( \38588 , \38379 , \38384 );
and \U$38274 ( \38589 , \38375 , \38384 );
or \U$38275 ( \38590 , \38587 , \38588 , \38589 );
and \U$38276 ( \38591 , \38360 , \38364 );
and \U$38277 ( \38592 , \38364 , \38369 );
and \U$38278 ( \38593 , \38360 , \38369 );
or \U$38279 ( \38594 , \38591 , \38592 , \38593 );
xor \U$38280 ( \38595 , \38590 , \38594 );
and \U$38281 ( \38596 , \38346 , \38350 );
and \U$38282 ( \38597 , \38350 , \38355 );
and \U$38283 ( \38598 , \38346 , \38355 );
or \U$38284 ( \38599 , \38596 , \38597 , \38598 );
xor \U$38285 ( \38600 , \38595 , \38599 );
and \U$38286 ( \38601 , \22561 , \38469 );
and \U$38287 ( \38602 , \38469 , \38474 );
and \U$38288 ( \38603 , \22561 , \38474 );
or \U$38289 ( \38604 , \38601 , \38602 , \38603 );
and \U$38290 ( \38605 , \38454 , \38458 );
and \U$38291 ( \38606 , \38458 , \38463 );
and \U$38292 ( \38607 , \38454 , \38463 );
or \U$38293 ( \38608 , \38605 , \38606 , \38607 );
xor \U$38294 ( \38609 , \38604 , \38608 );
and \U$38295 ( \38610 , \38440 , \38444 );
and \U$38296 ( \38611 , \38444 , \38449 );
and \U$38297 ( \38612 , \38440 , \38449 );
or \U$38298 ( \38613 , \38610 , \38611 , \38612 );
xor \U$38299 ( \38614 , \38609 , \38613 );
xor \U$38300 ( \38615 , \38600 , \38614 );
and \U$38301 ( \38616 , \22440 , \22278 );
and \U$38302 ( \38617 , \22407 , \22276 );
nor \U$38303 ( \38618 , \38616 , \38617 );
xnor \U$38304 ( \38619 , \38618 , \22288 );
and \U$38305 ( \38620 , \22468 , \22300 );
and \U$38306 ( \38621 , \22429 , \22298 );
nor \U$38307 ( \38622 , \38620 , \38621 );
xnor \U$38308 ( \38623 , \38622 , \22310 );
xor \U$38309 ( \38624 , \38619 , \38623 );
and \U$38310 ( \38625 , \22489 , \22324 );
and \U$38311 ( \38626 , \22457 , \22322 );
nor \U$38312 ( \38627 , \38625 , \38626 );
xnor \U$38313 ( \38628 , \38627 , \22334 );
xor \U$38314 ( \38629 , \38624 , \38628 );
and \U$38315 ( \38630 , \22372 , \22208 );
and \U$38316 ( \38631 , \22339 , \22206 );
nor \U$38317 ( \38632 , \38630 , \38631 );
xnor \U$38318 ( \38633 , \38632 , \22218 );
and \U$38319 ( \38634 , \22397 , \22230 );
and \U$38320 ( \38635 , \22361 , \22228 );
nor \U$38321 ( \38636 , \38634 , \38635 );
xnor \U$38322 ( \38637 , \38636 , \22240 );
xor \U$38323 ( \38638 , \38633 , \38637 );
and \U$38324 ( \38639 , \22418 , \22257 );
and \U$38325 ( \38640 , \22386 , \22255 );
nor \U$38326 ( \38641 , \38639 , \38640 );
xnor \U$38327 ( \38642 , \38641 , \22267 );
xor \U$38328 ( \38643 , \38638 , \38642 );
xor \U$38329 ( \38644 , \38629 , \38643 );
and \U$38330 ( \38645 , \22305 , \22140 );
and \U$38331 ( \38646 , \22272 , \22138 );
nor \U$38332 ( \38647 , \38645 , \38646 );
xnor \U$38333 ( \38648 , \38647 , \22150 );
and \U$38334 ( \38649 , \22329 , \22162 );
and \U$38335 ( \38650 , \22294 , \22160 );
nor \U$38336 ( \38651 , \38649 , \38650 );
xnor \U$38337 ( \38652 , \38651 , \22172 );
xor \U$38338 ( \38653 , \38648 , \38652 );
and \U$38339 ( \38654 , \22350 , \22187 );
and \U$38340 ( \38655 , \22318 , \22185 );
nor \U$38341 ( \38656 , \38654 , \38655 );
xnor \U$38342 ( \38657 , \38656 , \22197 );
xor \U$38343 ( \38658 , \38653 , \38657 );
xor \U$38344 ( \38659 , \38644 , \38658 );
and \U$38345 ( \38660 , \22646 , \22484 );
and \U$38346 ( \38661 , \22613 , \22482 );
nor \U$38347 ( \38662 , \38660 , \38661 );
xnor \U$38348 ( \38663 , \38662 , \22494 );
and \U$38349 ( \38664 , \22676 , \22506 );
and \U$38350 ( \38665 , \22635 , \22504 );
nor \U$38351 ( \38666 , \38664 , \38665 );
xnor \U$38352 ( \38667 , \38666 , \22516 );
xor \U$38353 ( \38668 , \38663 , \38667 );
and \U$38354 ( \38669 , \22696 , \22530 );
and \U$38355 ( \38670 , \22665 , \22528 );
nor \U$38356 ( \38671 , \38669 , \38670 );
xnor \U$38357 ( \38672 , \38671 , \22540 );
xor \U$38358 ( \38673 , \38668 , \38672 );
and \U$38359 ( \38674 , \22578 , \22413 );
and \U$38360 ( \38675 , \22545 , \22411 );
nor \U$38361 ( \38676 , \38674 , \38675 );
xnor \U$38362 ( \38677 , \38676 , \22423 );
and \U$38363 ( \38678 , \22603 , \22435 );
and \U$38364 ( \38679 , \22567 , \22433 );
nor \U$38365 ( \38680 , \38678 , \38679 );
xnor \U$38366 ( \38681 , \38680 , \22445 );
xor \U$38367 ( \38682 , \38677 , \38681 );
and \U$38368 ( \38683 , \22624 , \22463 );
and \U$38369 ( \38684 , \22592 , \22461 );
nor \U$38370 ( \38685 , \38683 , \38684 );
xnor \U$38371 ( \38686 , \38685 , \22473 );
xor \U$38372 ( \38687 , \38682 , \38686 );
xor \U$38373 ( \38688 , \38673 , \38687 );
and \U$38374 ( \38689 , \22511 , \22345 );
and \U$38375 ( \38690 , \22478 , \22343 );
nor \U$38376 ( \38691 , \38689 , \38690 );
xnor \U$38377 ( \38692 , \38691 , \22355 );
and \U$38378 ( \38693 , \22535 , \22367 );
and \U$38379 ( \38694 , \22500 , \22365 );
nor \U$38380 ( \38695 , \38693 , \38694 );
xnor \U$38381 ( \38696 , \38695 , \22377 );
xor \U$38382 ( \38697 , \38692 , \38696 );
and \U$38383 ( \38698 , \22556 , \22392 );
and \U$38384 ( \38699 , \22524 , \22390 );
nor \U$38385 ( \38700 , \38698 , \38699 );
xnor \U$38386 ( \38701 , \38700 , \22402 );
xor \U$38387 ( \38702 , \38697 , \38701 );
xor \U$38388 ( \38703 , \38688 , \38702 );
xor \U$38389 ( \38704 , \38659 , \38703 );
and \U$38390 ( \38705 , \38402 , \38406 );
and \U$38391 ( \38706 , \38406 , \38411 );
and \U$38392 ( \38707 , \38402 , \38411 );
or \U$38393 ( \38708 , \38705 , \38706 , \38707 );
and \U$38394 ( \38709 , \38394 , \38396 );
xor \U$38395 ( \38710 , \38708 , \38709 );
and \U$38396 ( \38711 , \22706 , \22551 );
and \U$38397 ( \38712 , \22686 , \22549 );
nor \U$38398 ( \38713 , \38711 , \38712 );
xnor \U$38399 ( \38714 , \38713 , \22561 );
xor \U$38400 ( \38715 , \38710 , \38714 );
xor \U$38401 ( \38716 , \38704 , \38715 );
xor \U$38402 ( \38717 , \38615 , \38716 );
xor \U$38403 ( \38718 , \38586 , \38717 );
and \U$38404 ( \38719 , \38507 , \38511 );
and \U$38405 ( \38720 , \38511 , \38516 );
and \U$38406 ( \38721 , \38507 , \38516 );
or \U$38407 ( \38722 , \38719 , \38720 , \38721 );
and \U$38408 ( \38723 , \38434 , \38435 );
and \U$38409 ( \38724 , \38435 , \38476 );
and \U$38410 ( \38725 , \38434 , \38476 );
or \U$38411 ( \38726 , \38723 , \38724 , \38725 );
xor \U$38412 ( \38727 , \38722 , \38726 );
and \U$38413 ( \38728 , \38386 , \38413 );
and \U$38414 ( \38729 , \38413 , \38428 );
and \U$38415 ( \38730 , \38386 , \38428 );
or \U$38416 ( \38731 , \38728 , \38729 , \38730 );
xor \U$38417 ( \38732 , \38727 , \38731 );
xor \U$38418 ( \38733 , \38718 , \38732 );
xor \U$38419 ( \38734 , \38572 , \38733 );
xor \U$38420 ( \38735 , \38566 , \38734 );
and \U$38421 ( \38736 , \38324 , \38519 );
nor \U$38422 ( \38737 , \38735 , \38736 );
and \U$38423 ( \38738 , \38570 , \38571 );
and \U$38424 ( \38739 , \38571 , \38733 );
and \U$38425 ( \38740 , \38570 , \38733 );
or \U$38426 ( \38741 , \38738 , \38739 , \38740 );
and \U$38427 ( \38742 , \38576 , \38580 );
and \U$38428 ( \38743 , \38580 , \38585 );
and \U$38429 ( \38744 , \38576 , \38585 );
or \U$38430 ( \38745 , \38742 , \38743 , \38744 );
and \U$38431 ( \38746 , \38544 , \38548 );
and \U$38432 ( \38747 , \38548 , \38563 );
and \U$38433 ( \38748 , \38544 , \38563 );
or \U$38434 ( \38749 , \38746 , \38747 , \38748 );
xor \U$38435 ( \38750 , \38745 , \38749 );
and \U$38436 ( \38751 , \38659 , \38703 );
and \U$38437 ( \38752 , \38703 , \38715 );
and \U$38438 ( \38753 , \38659 , \38715 );
or \U$38439 ( \38754 , \38751 , \38752 , \38753 );
xor \U$38440 ( \38755 , \38750 , \38754 );
and \U$38441 ( \38756 , \38722 , \38726 );
and \U$38442 ( \38757 , \38726 , \38731 );
and \U$38443 ( \38758 , \38722 , \38731 );
or \U$38444 ( \38759 , \38756 , \38757 , \38758 );
and \U$38445 ( \38760 , \38600 , \38614 );
and \U$38446 ( \38761 , \38614 , \38716 );
and \U$38447 ( \38762 , \38600 , \38716 );
or \U$38448 ( \38763 , \38760 , \38761 , \38762 );
xor \U$38449 ( \38764 , \38759 , \38763 );
and \U$38450 ( \38765 , \38604 , \38608 );
and \U$38451 ( \38766 , \38608 , \38613 );
and \U$38452 ( \38767 , \38604 , \38613 );
or \U$38453 ( \38768 , \38765 , \38766 , \38767 );
and \U$38454 ( \38769 , \38590 , \38594 );
and \U$38455 ( \38770 , \38594 , \38599 );
and \U$38456 ( \38771 , \38590 , \38599 );
or \U$38457 ( \38772 , \38769 , \38770 , \38771 );
xor \U$38458 ( \38773 , \38768 , \38772 );
and \U$38459 ( \38774 , \38708 , \38709 );
and \U$38460 ( \38775 , \38709 , \38714 );
and \U$38461 ( \38776 , \38708 , \38714 );
or \U$38462 ( \38777 , \38774 , \38775 , \38776 );
xor \U$38463 ( \38778 , \38773 , \38777 );
xor \U$38464 ( \38779 , \38764 , \38778 );
xor \U$38465 ( \38780 , \38755 , \38779 );
xor \U$38466 ( \38781 , \38741 , \38780 );
and \U$38467 ( \38782 , \38535 , \38539 );
and \U$38468 ( \38783 , \38539 , \38564 );
and \U$38469 ( \38784 , \38535 , \38564 );
or \U$38470 ( \38785 , \38782 , \38783 , \38784 );
and \U$38471 ( \38786 , \38586 , \38717 );
and \U$38472 ( \38787 , \38717 , \38732 );
and \U$38473 ( \38788 , \38586 , \38732 );
or \U$38474 ( \38789 , \38786 , \38787 , \38788 );
xor \U$38475 ( \38790 , \38785 , \38789 );
and \U$38476 ( \38791 , \38553 , \38557 );
and \U$38477 ( \38792 , \38557 , \38562 );
and \U$38478 ( \38793 , \38553 , \38562 );
or \U$38479 ( \38794 , \38791 , \38792 , \38793 );
and \U$38480 ( \38795 , \38648 , \38652 );
and \U$38481 ( \38796 , \38652 , \38657 );
and \U$38482 ( \38797 , \38648 , \38657 );
or \U$38483 ( \38798 , \38795 , \38796 , \38797 );
xor \U$38484 ( \38799 , \38794 , \38798 );
and \U$38485 ( \38800 , \38633 , \38637 );
and \U$38486 ( \38801 , \38637 , \38642 );
and \U$38487 ( \38802 , \38633 , \38642 );
or \U$38488 ( \38803 , \38800 , \38801 , \38802 );
xor \U$38489 ( \38804 , \38799 , \38803 );
and \U$38490 ( \38805 , \22524 , \22392 );
and \U$38491 ( \38806 , \22535 , \22390 );
nor \U$38492 ( \38807 , \38805 , \38806 );
xnor \U$38493 ( \38808 , \38807 , \22402 );
and \U$38494 ( \38809 , \22545 , \22413 );
and \U$38495 ( \38810 , \22556 , \22411 );
nor \U$38496 ( \38811 , \38809 , \38810 );
xnor \U$38497 ( \38812 , \38811 , \22423 );
xor \U$38498 ( \38813 , \38808 , \38812 );
and \U$38499 ( \38814 , \22567 , \22435 );
and \U$38500 ( \38815 , \22578 , \22433 );
nor \U$38501 ( \38816 , \38814 , \38815 );
xnor \U$38502 ( \38817 , \38816 , \22445 );
xor \U$38503 ( \38818 , \38813 , \38817 );
and \U$38504 ( \38819 , \22457 , \22324 );
and \U$38505 ( \38820 , \22468 , \22322 );
nor \U$38506 ( \38821 , \38819 , \38820 );
xnor \U$38507 ( \38822 , \38821 , \22334 );
and \U$38508 ( \38823 , \22478 , \22345 );
and \U$38509 ( \38824 , \22489 , \22343 );
nor \U$38510 ( \38825 , \38823 , \38824 );
xnor \U$38511 ( \38826 , \38825 , \22355 );
xor \U$38512 ( \38827 , \38822 , \38826 );
and \U$38513 ( \38828 , \22500 , \22367 );
and \U$38514 ( \38829 , \22511 , \22365 );
nor \U$38515 ( \38830 , \38828 , \38829 );
xnor \U$38516 ( \38831 , \38830 , \22377 );
xor \U$38517 ( \38832 , \38827 , \38831 );
xor \U$38518 ( \38833 , \38818 , \38832 );
and \U$38519 ( \38834 , \22386 , \22257 );
and \U$38520 ( \38835 , \22397 , \22255 );
nor \U$38521 ( \38836 , \38834 , \38835 );
xnor \U$38522 ( \38837 , \38836 , \22267 );
and \U$38523 ( \38838 , \22407 , \22278 );
and \U$38524 ( \38839 , \22418 , \22276 );
nor \U$38525 ( \38840 , \38838 , \38839 );
xnor \U$38526 ( \38841 , \38840 , \22288 );
xor \U$38527 ( \38842 , \38837 , \38841 );
and \U$38528 ( \38843 , \22429 , \22300 );
and \U$38529 ( \38844 , \22440 , \22298 );
nor \U$38530 ( \38845 , \38843 , \38844 );
xnor \U$38531 ( \38846 , \38845 , \22310 );
xor \U$38532 ( \38847 , \38842 , \38846 );
xor \U$38533 ( \38848 , \38833 , \38847 );
and \U$38534 ( \38849 , \38663 , \38667 );
and \U$38535 ( \38850 , \38667 , \38672 );
and \U$38536 ( \38851 , \38663 , \38672 );
or \U$38537 ( \38852 , \38849 , \38850 , \38851 );
and \U$38538 ( \38853 , \22665 , \22530 );
and \U$38539 ( \38854 , \22676 , \22528 );
nor \U$38540 ( \38855 , \38853 , \38854 );
xnor \U$38541 ( \38856 , \38855 , \22540 );
and \U$38542 ( \38857 , \22686 , \22551 );
and \U$38543 ( \38858 , \22696 , \22549 );
nor \U$38544 ( \38859 , \38857 , \38858 );
xnor \U$38545 ( \38860 , \38859 , \22561 );
xor \U$38546 ( \38861 , \38856 , \38860 );
nand \U$38547 ( \38862 , \22706 , \22571 );
xnor \U$38548 ( \38863 , \38862 , \22583 );
xor \U$38549 ( \38864 , \38861 , \38863 );
xor \U$38550 ( \38865 , \38852 , \38864 );
and \U$38551 ( \38866 , \22592 , \22463 );
and \U$38552 ( \38867 , \22603 , \22461 );
nor \U$38553 ( \38868 , \38866 , \38867 );
xnor \U$38554 ( \38869 , \38868 , \22473 );
and \U$38555 ( \38870 , \22613 , \22484 );
and \U$38556 ( \38871 , \22624 , \22482 );
nor \U$38557 ( \38872 , \38870 , \38871 );
xnor \U$38558 ( \38873 , \38872 , \22494 );
xor \U$38559 ( \38874 , \38869 , \38873 );
and \U$38560 ( \38875 , \22635 , \22506 );
and \U$38561 ( \38876 , \22646 , \22504 );
nor \U$38562 ( \38877 , \38875 , \38876 );
xnor \U$38563 ( \38878 , \38877 , \22516 );
xor \U$38564 ( \38879 , \38874 , \38878 );
xor \U$38565 ( \38880 , \38865 , \38879 );
xor \U$38566 ( \38881 , \38848 , \38880 );
and \U$38567 ( \38882 , \38619 , \38623 );
and \U$38568 ( \38883 , \38623 , \38628 );
and \U$38569 ( \38884 , \38619 , \38628 );
or \U$38570 ( \38885 , \38882 , \38883 , \38884 );
and \U$38571 ( \38886 , \38692 , \38696 );
and \U$38572 ( \38887 , \38696 , \38701 );
and \U$38573 ( \38888 , \38692 , \38701 );
or \U$38574 ( \38889 , \38886 , \38887 , \38888 );
xor \U$38575 ( \38890 , \38885 , \38889 );
and \U$38576 ( \38891 , \38677 , \38681 );
and \U$38577 ( \38892 , \38681 , \38686 );
and \U$38578 ( \38893 , \38677 , \38686 );
or \U$38579 ( \38894 , \38891 , \38892 , \38893 );
xor \U$38580 ( \38895 , \38890 , \38894 );
xor \U$38581 ( \38896 , \38881 , \38895 );
xor \U$38582 ( \38897 , \38804 , \38896 );
and \U$38583 ( \38898 , \38673 , \38687 );
and \U$38584 ( \38899 , \38687 , \38702 );
and \U$38585 ( \38900 , \38673 , \38702 );
or \U$38586 ( \38901 , \38898 , \38899 , \38900 );
and \U$38587 ( \38902 , \38629 , \38643 );
and \U$38588 ( \38903 , \38643 , \38658 );
and \U$38589 ( \38904 , \38629 , \38658 );
or \U$38590 ( \38905 , \38902 , \38903 , \38904 );
xor \U$38591 ( \38906 , \38901 , \38905 );
and \U$38592 ( \38907 , \22318 , \22187 );
and \U$38593 ( \38908 , \22329 , \22185 );
nor \U$38594 ( \38909 , \38907 , \38908 );
xnor \U$38595 ( \38910 , \38909 , \22197 );
and \U$38596 ( \38911 , \22339 , \22208 );
and \U$38597 ( \38912 , \22350 , \22206 );
nor \U$38598 ( \38913 , \38911 , \38912 );
xnor \U$38599 ( \38914 , \38913 , \22218 );
xor \U$38600 ( \38915 , \38910 , \38914 );
and \U$38601 ( \38916 , \22361 , \22230 );
and \U$38602 ( \38917 , \22372 , \22228 );
nor \U$38603 ( \38918 , \38916 , \38917 );
xnor \U$38604 ( \38919 , \38918 , \22240 );
xor \U$38605 ( \38920 , \38915 , \38919 );
and \U$38606 ( \38921 , \22251 , \22119 );
and \U$38607 ( \38922 , \22262 , \22117 );
nor \U$38608 ( \38923 , \38921 , \38922 );
xnor \U$38609 ( \38924 , \38923 , \22129 );
and \U$38610 ( \38925 , \22272 , \22140 );
and \U$38611 ( \38926 , \22283 , \22138 );
nor \U$38612 ( \38927 , \38925 , \38926 );
xnor \U$38613 ( \38928 , \38927 , \22150 );
xor \U$38614 ( \38929 , \38924 , \38928 );
and \U$38615 ( \38930 , \22294 , \22162 );
and \U$38616 ( \38931 , \22305 , \22160 );
nor \U$38617 ( \38932 , \38930 , \38931 );
xnor \U$38618 ( \38933 , \38932 , \22172 );
xor \U$38619 ( \38934 , \38929 , \38933 );
xor \U$38620 ( \38935 , \38920 , \38934 );
and \U$38621 ( \38936 , \22202 , \22076 );
and \U$38622 ( \38937 , \22213 , \22073 );
nor \U$38623 ( \38938 , \38936 , \38937 );
xnor \U$38624 ( \38939 , \38938 , \22072 );
xor \U$38625 ( \38940 , \22583 , \38939 );
and \U$38626 ( \38941 , \22224 , \22095 );
and \U$38627 ( \38942 , \22235 , \22093 );
nor \U$38628 ( \38943 , \38941 , \38942 );
xnor \U$38629 ( \38944 , \38943 , \22105 );
xor \U$38630 ( \38945 , \38940 , \38944 );
xor \U$38631 ( \38946 , \38935 , \38945 );
xor \U$38632 ( \38947 , \38906 , \38946 );
xor \U$38633 ( \38948 , \38897 , \38947 );
xor \U$38634 ( \38949 , \38790 , \38948 );
xor \U$38635 ( \38950 , \38781 , \38949 );
and \U$38636 ( \38951 , \38531 , \38565 );
and \U$38637 ( \38952 , \38565 , \38734 );
and \U$38638 ( \38953 , \38531 , \38734 );
or \U$38639 ( \38954 , \38951 , \38952 , \38953 );
nor \U$38640 ( \38955 , \38950 , \38954 );
nor \U$38641 ( \38956 , \38737 , \38955 );
and \U$38642 ( \38957 , \38785 , \38789 );
and \U$38643 ( \38958 , \38789 , \38948 );
and \U$38644 ( \38959 , \38785 , \38948 );
or \U$38645 ( \38960 , \38957 , \38958 , \38959 );
and \U$38646 ( \38961 , \38755 , \38779 );
xor \U$38647 ( \38962 , \38960 , \38961 );
and \U$38648 ( \38963 , \38759 , \38763 );
and \U$38649 ( \38964 , \38763 , \38778 );
and \U$38650 ( \38965 , \38759 , \38778 );
or \U$38651 ( \38966 , \38963 , \38964 , \38965 );
and \U$38652 ( \38967 , \38869 , \38873 );
and \U$38653 ( \38968 , \38873 , \38878 );
and \U$38654 ( \38969 , \38869 , \38878 );
or \U$38655 ( \38970 , \38967 , \38968 , \38969 );
and \U$38656 ( \38971 , \38856 , \38860 );
and \U$38657 ( \38972 , \38860 , \38863 );
and \U$38658 ( \38973 , \38856 , \38863 );
or \U$38659 ( \38974 , \38971 , \38972 , \38973 );
xor \U$38660 ( \38975 , \38970 , \38974 );
and \U$38661 ( \38976 , \22696 , \22551 );
and \U$38662 ( \38977 , \22665 , \22549 );
nor \U$38663 ( \38978 , \38976 , \38977 );
xnor \U$38664 ( \38979 , \38978 , \22561 );
xor \U$38665 ( \38980 , \38975 , \38979 );
and \U$38666 ( \38981 , \38837 , \38841 );
and \U$38667 ( \38982 , \38841 , \38846 );
and \U$38668 ( \38983 , \38837 , \38846 );
or \U$38669 ( \38984 , \38981 , \38982 , \38983 );
and \U$38670 ( \38985 , \38822 , \38826 );
and \U$38671 ( \38986 , \38826 , \38831 );
and \U$38672 ( \38987 , \38822 , \38831 );
or \U$38673 ( \38988 , \38985 , \38986 , \38987 );
xor \U$38674 ( \38989 , \38984 , \38988 );
and \U$38675 ( \38990 , \38808 , \38812 );
and \U$38676 ( \38991 , \38812 , \38817 );
and \U$38677 ( \38992 , \38808 , \38817 );
or \U$38678 ( \38993 , \38990 , \38991 , \38992 );
xor \U$38679 ( \38994 , \38989 , \38993 );
xor \U$38680 ( \38995 , \38980 , \38994 );
and \U$38681 ( \38996 , \22583 , \38939 );
and \U$38682 ( \38997 , \38939 , \38944 );
and \U$38683 ( \38998 , \22583 , \38944 );
or \U$38684 ( \38999 , \38996 , \38997 , \38998 );
and \U$38685 ( \39000 , \38924 , \38928 );
and \U$38686 ( \39001 , \38928 , \38933 );
and \U$38687 ( \39002 , \38924 , \38933 );
or \U$38688 ( \39003 , \39000 , \39001 , \39002 );
xor \U$38689 ( \39004 , \38999 , \39003 );
and \U$38690 ( \39005 , \38910 , \38914 );
and \U$38691 ( \39006 , \38914 , \38919 );
and \U$38692 ( \39007 , \38910 , \38919 );
or \U$38693 ( \39008 , \39005 , \39006 , \39007 );
xor \U$38694 ( \39009 , \39004 , \39008 );
xor \U$38695 ( \39010 , \38995 , \39009 );
and \U$38696 ( \39011 , \22213 , \22076 );
and \U$38697 ( \39012 , \22181 , \22073 );
nor \U$38698 ( \39013 , \39011 , \39012 );
xnor \U$38699 ( \39014 , \39013 , \22072 );
and \U$38700 ( \39015 , \22235 , \22095 );
and \U$38701 ( \39016 , \22202 , \22093 );
nor \U$38702 ( \39017 , \39015 , \39016 );
xnor \U$38703 ( \39018 , \39017 , \22105 );
xor \U$38704 ( \39019 , \39014 , \39018 );
and \U$38705 ( \39020 , \22262 , \22119 );
and \U$38706 ( \39021 , \22224 , \22117 );
nor \U$38707 ( \39022 , \39020 , \39021 );
xnor \U$38708 ( \39023 , \39022 , \22129 );
xor \U$38709 ( \39024 , \39019 , \39023 );
and \U$38710 ( \39025 , \22489 , \22345 );
and \U$38711 ( \39026 , \22457 , \22343 );
nor \U$38712 ( \39027 , \39025 , \39026 );
xnor \U$38713 ( \39028 , \39027 , \22355 );
and \U$38714 ( \39029 , \22511 , \22367 );
and \U$38715 ( \39030 , \22478 , \22365 );
nor \U$38716 ( \39031 , \39029 , \39030 );
xnor \U$38717 ( \39032 , \39031 , \22377 );
xor \U$38718 ( \39033 , \39028 , \39032 );
and \U$38719 ( \39034 , \22535 , \22392 );
and \U$38720 ( \39035 , \22500 , \22390 );
nor \U$38721 ( \39036 , \39034 , \39035 );
xnor \U$38722 ( \39037 , \39036 , \22402 );
xor \U$38723 ( \39038 , \39033 , \39037 );
and \U$38724 ( \39039 , \22418 , \22278 );
and \U$38725 ( \39040 , \22386 , \22276 );
nor \U$38726 ( \39041 , \39039 , \39040 );
xnor \U$38727 ( \39042 , \39041 , \22288 );
and \U$38728 ( \39043 , \22440 , \22300 );
and \U$38729 ( \39044 , \22407 , \22298 );
nor \U$38730 ( \39045 , \39043 , \39044 );
xnor \U$38731 ( \39046 , \39045 , \22310 );
xor \U$38732 ( \39047 , \39042 , \39046 );
and \U$38733 ( \39048 , \22468 , \22324 );
and \U$38734 ( \39049 , \22429 , \22322 );
nor \U$38735 ( \39050 , \39048 , \39049 );
xnor \U$38736 ( \39051 , \39050 , \22334 );
xor \U$38737 ( \39052 , \39047 , \39051 );
xor \U$38738 ( \39053 , \39038 , \39052 );
and \U$38739 ( \39054 , \22350 , \22208 );
and \U$38740 ( \39055 , \22318 , \22206 );
nor \U$38741 ( \39056 , \39054 , \39055 );
xnor \U$38742 ( \39057 , \39056 , \22218 );
and \U$38743 ( \39058 , \22372 , \22230 );
and \U$38744 ( \39059 , \22339 , \22228 );
nor \U$38745 ( \39060 , \39058 , \39059 );
xnor \U$38746 ( \39061 , \39060 , \22240 );
xor \U$38747 ( \39062 , \39057 , \39061 );
and \U$38748 ( \39063 , \22397 , \22257 );
and \U$38749 ( \39064 , \22361 , \22255 );
nor \U$38750 ( \39065 , \39063 , \39064 );
xnor \U$38751 ( \39066 , \39065 , \22267 );
xor \U$38752 ( \39067 , \39062 , \39066 );
xor \U$38753 ( \39068 , \39053 , \39067 );
xor \U$38754 ( \39069 , \39024 , \39068 );
and \U$38755 ( \39070 , \22706 , \22573 );
and \U$38756 ( \39071 , \22686 , \22571 );
nor \U$38757 ( \39072 , \39070 , \39071 );
xnor \U$38758 ( \39073 , \39072 , \22583 );
and \U$38759 ( \39074 , \22624 , \22484 );
and \U$38760 ( \39075 , \22592 , \22482 );
nor \U$38761 ( \39076 , \39074 , \39075 );
xnor \U$38762 ( \39077 , \39076 , \22494 );
and \U$38763 ( \39078 , \22646 , \22506 );
and \U$38764 ( \39079 , \22613 , \22504 );
nor \U$38765 ( \39080 , \39078 , \39079 );
xnor \U$38766 ( \39081 , \39080 , \22516 );
xor \U$38767 ( \39082 , \39077 , \39081 );
and \U$38768 ( \39083 , \22676 , \22530 );
and \U$38769 ( \39084 , \22635 , \22528 );
nor \U$38770 ( \39085 , \39083 , \39084 );
xnor \U$38771 ( \39086 , \39085 , \22540 );
xor \U$38772 ( \39087 , \39082 , \39086 );
xor \U$38773 ( \39088 , \39073 , \39087 );
and \U$38774 ( \39089 , \22556 , \22413 );
and \U$38775 ( \39090 , \22524 , \22411 );
nor \U$38776 ( \39091 , \39089 , \39090 );
xnor \U$38777 ( \39092 , \39091 , \22423 );
and \U$38778 ( \39093 , \22578 , \22435 );
and \U$38779 ( \39094 , \22545 , \22433 );
nor \U$38780 ( \39095 , \39093 , \39094 );
xnor \U$38781 ( \39096 , \39095 , \22445 );
xor \U$38782 ( \39097 , \39092 , \39096 );
and \U$38783 ( \39098 , \22603 , \22463 );
and \U$38784 ( \39099 , \22567 , \22461 );
nor \U$38785 ( \39100 , \39098 , \39099 );
xnor \U$38786 ( \39101 , \39100 , \22473 );
xor \U$38787 ( \39102 , \39097 , \39101 );
xor \U$38788 ( \39103 , \39088 , \39102 );
xor \U$38789 ( \39104 , \39069 , \39103 );
xor \U$38790 ( \39105 , \39010 , \39104 );
and \U$38791 ( \39106 , \38818 , \38832 );
and \U$38792 ( \39107 , \38832 , \38847 );
and \U$38793 ( \39108 , \38818 , \38847 );
or \U$38794 ( \39109 , \39106 , \39107 , \39108 );
and \U$38795 ( \39110 , \38920 , \38934 );
and \U$38796 ( \39111 , \38934 , \38945 );
and \U$38797 ( \39112 , \38920 , \38945 );
or \U$38798 ( \39113 , \39110 , \39111 , \39112 );
xor \U$38799 ( \39114 , \39109 , \39113 );
and \U$38800 ( \39115 , \22283 , \22140 );
and \U$38801 ( \39116 , \22251 , \22138 );
nor \U$38802 ( \39117 , \39115 , \39116 );
xnor \U$38803 ( \39118 , \39117 , \22150 );
and \U$38804 ( \39119 , \22305 , \22162 );
and \U$38805 ( \39120 , \22272 , \22160 );
nor \U$38806 ( \39121 , \39119 , \39120 );
xnor \U$38807 ( \39122 , \39121 , \22172 );
xor \U$38808 ( \39123 , \39118 , \39122 );
and \U$38809 ( \39124 , \22329 , \22187 );
and \U$38810 ( \39125 , \22294 , \22185 );
nor \U$38811 ( \39126 , \39124 , \39125 );
xnor \U$38812 ( \39127 , \39126 , \22197 );
xor \U$38813 ( \39128 , \39123 , \39127 );
xor \U$38814 ( \39129 , \39114 , \39128 );
xor \U$38815 ( \39130 , \39105 , \39129 );
and \U$38816 ( \39131 , \38768 , \38772 );
and \U$38817 ( \39132 , \38772 , \38777 );
and \U$38818 ( \39133 , \38768 , \38777 );
or \U$38819 ( \39134 , \39131 , \39132 , \39133 );
and \U$38820 ( \39135 , \38901 , \38905 );
and \U$38821 ( \39136 , \38905 , \38946 );
and \U$38822 ( \39137 , \38901 , \38946 );
or \U$38823 ( \39138 , \39135 , \39136 , \39137 );
xor \U$38824 ( \39139 , \39134 , \39138 );
and \U$38825 ( \39140 , \38848 , \38880 );
and \U$38826 ( \39141 , \38880 , \38895 );
and \U$38827 ( \39142 , \38848 , \38895 );
or \U$38828 ( \39143 , \39140 , \39141 , \39142 );
xor \U$38829 ( \39144 , \39139 , \39143 );
xor \U$38830 ( \39145 , \39130 , \39144 );
xor \U$38831 ( \39146 , \38966 , \39145 );
and \U$38832 ( \39147 , \38745 , \38749 );
and \U$38833 ( \39148 , \38749 , \38754 );
and \U$38834 ( \39149 , \38745 , \38754 );
or \U$38835 ( \39150 , \39147 , \39148 , \39149 );
and \U$38836 ( \39151 , \38804 , \38896 );
and \U$38837 ( \39152 , \38896 , \38947 );
and \U$38838 ( \39153 , \38804 , \38947 );
or \U$38839 ( \39154 , \39151 , \39152 , \39153 );
xor \U$38840 ( \39155 , \39150 , \39154 );
and \U$38841 ( \39156 , \38794 , \38798 );
and \U$38842 ( \39157 , \38798 , \38803 );
and \U$38843 ( \39158 , \38794 , \38803 );
or \U$38844 ( \39159 , \39156 , \39157 , \39158 );
and \U$38845 ( \39160 , \38885 , \38889 );
and \U$38846 ( \39161 , \38889 , \38894 );
and \U$38847 ( \39162 , \38885 , \38894 );
or \U$38848 ( \39163 , \39160 , \39161 , \39162 );
xor \U$38849 ( \39164 , \39159 , \39163 );
and \U$38850 ( \39165 , \38852 , \38864 );
and \U$38851 ( \39166 , \38864 , \38879 );
and \U$38852 ( \39167 , \38852 , \38879 );
or \U$38853 ( \39168 , \39165 , \39166 , \39167 );
xor \U$38854 ( \39169 , \39164 , \39168 );
xor \U$38855 ( \39170 , \39155 , \39169 );
xor \U$38856 ( \39171 , \39146 , \39170 );
xor \U$38857 ( \39172 , \38962 , \39171 );
and \U$38858 ( \39173 , \38741 , \38780 );
and \U$38859 ( \39174 , \38780 , \38949 );
and \U$38860 ( \39175 , \38741 , \38949 );
or \U$38861 ( \39176 , \39173 , \39174 , \39175 );
nor \U$38862 ( \39177 , \39172 , \39176 );
and \U$38863 ( \39178 , \38966 , \39145 );
and \U$38864 ( \39179 , \39145 , \39170 );
and \U$38865 ( \39180 , \38966 , \39170 );
or \U$38866 ( \39181 , \39178 , \39179 , \39180 );
and \U$38867 ( \39182 , \39159 , \39163 );
and \U$38868 ( \39183 , \39163 , \39168 );
and \U$38869 ( \39184 , \39159 , \39168 );
or \U$38870 ( \39185 , \39182 , \39183 , \39184 );
and \U$38871 ( \39186 , \39109 , \39113 );
and \U$38872 ( \39187 , \39113 , \39128 );
and \U$38873 ( \39188 , \39109 , \39128 );
or \U$38874 ( \39189 , \39186 , \39187 , \39188 );
xor \U$38875 ( \39190 , \39185 , \39189 );
and \U$38876 ( \39191 , \39024 , \39068 );
and \U$38877 ( \39192 , \39068 , \39103 );
and \U$38878 ( \39193 , \39024 , \39103 );
or \U$38879 ( \39194 , \39191 , \39192 , \39193 );
xor \U$38880 ( \39195 , \39190 , \39194 );
and \U$38881 ( \39196 , \39134 , \39138 );
and \U$38882 ( \39197 , \39138 , \39143 );
and \U$38883 ( \39198 , \39134 , \39143 );
or \U$38884 ( \39199 , \39196 , \39197 , \39198 );
and \U$38885 ( \39200 , \39010 , \39104 );
and \U$38886 ( \39201 , \39104 , \39129 );
and \U$38887 ( \39202 , \39010 , \39129 );
or \U$38888 ( \39203 , \39200 , \39201 , \39202 );
xor \U$38889 ( \39204 , \39199 , \39203 );
and \U$38890 ( \39205 , \22361 , \22257 );
and \U$38891 ( \39206 , \22372 , \22255 );
nor \U$38892 ( \39207 , \39205 , \39206 );
xnor \U$38893 ( \39208 , \39207 , \22267 );
and \U$38894 ( \39209 , \22386 , \22278 );
and \U$38895 ( \39210 , \22397 , \22276 );
nor \U$38896 ( \39211 , \39209 , \39210 );
xnor \U$38897 ( \39212 , \39211 , \22288 );
xor \U$38898 ( \39213 , \39208 , \39212 );
and \U$38899 ( \39214 , \22407 , \22300 );
and \U$38900 ( \39215 , \22418 , \22298 );
nor \U$38901 ( \39216 , \39214 , \39215 );
xnor \U$38902 ( \39217 , \39216 , \22310 );
xor \U$38903 ( \39218 , \39213 , \39217 );
and \U$38904 ( \39219 , \22294 , \22187 );
and \U$38905 ( \39220 , \22305 , \22185 );
nor \U$38906 ( \39221 , \39219 , \39220 );
xnor \U$38907 ( \39222 , \39221 , \22197 );
and \U$38908 ( \39223 , \22318 , \22208 );
and \U$38909 ( \39224 , \22329 , \22206 );
nor \U$38910 ( \39225 , \39223 , \39224 );
xnor \U$38911 ( \39226 , \39225 , \22218 );
xor \U$38912 ( \39227 , \39222 , \39226 );
and \U$38913 ( \39228 , \22339 , \22230 );
and \U$38914 ( \39229 , \22350 , \22228 );
nor \U$38915 ( \39230 , \39228 , \39229 );
xnor \U$38916 ( \39231 , \39230 , \22240 );
xor \U$38917 ( \39232 , \39227 , \39231 );
xor \U$38918 ( \39233 , \39218 , \39232 );
and \U$38919 ( \39234 , \22224 , \22119 );
and \U$38920 ( \39235 , \22235 , \22117 );
nor \U$38921 ( \39236 , \39234 , \39235 );
xnor \U$38922 ( \39237 , \39236 , \22129 );
and \U$38923 ( \39238 , \22251 , \22140 );
and \U$38924 ( \39239 , \22262 , \22138 );
nor \U$38925 ( \39240 , \39238 , \39239 );
xnor \U$38926 ( \39241 , \39240 , \22150 );
xor \U$38927 ( \39242 , \39237 , \39241 );
and \U$38928 ( \39243 , \22272 , \22162 );
and \U$38929 ( \39244 , \22283 , \22160 );
nor \U$38930 ( \39245 , \39243 , \39244 );
xnor \U$38931 ( \39246 , \39245 , \22172 );
xor \U$38932 ( \39247 , \39242 , \39246 );
xor \U$38933 ( \39248 , \39233 , \39247 );
and \U$38934 ( \39249 , \22567 , \22463 );
and \U$38935 ( \39250 , \22578 , \22461 );
nor \U$38936 ( \39251 , \39249 , \39250 );
xnor \U$38937 ( \39252 , \39251 , \22473 );
and \U$38938 ( \39253 , \22592 , \22484 );
and \U$38939 ( \39254 , \22603 , \22482 );
nor \U$38940 ( \39255 , \39253 , \39254 );
xnor \U$38941 ( \39256 , \39255 , \22494 );
xor \U$38942 ( \39257 , \39252 , \39256 );
and \U$38943 ( \39258 , \22613 , \22506 );
and \U$38944 ( \39259 , \22624 , \22504 );
nor \U$38945 ( \39260 , \39258 , \39259 );
xnor \U$38946 ( \39261 , \39260 , \22516 );
xor \U$38947 ( \39262 , \39257 , \39261 );
and \U$38948 ( \39263 , \22500 , \22392 );
and \U$38949 ( \39264 , \22511 , \22390 );
nor \U$38950 ( \39265 , \39263 , \39264 );
xnor \U$38951 ( \39266 , \39265 , \22402 );
and \U$38952 ( \39267 , \22524 , \22413 );
and \U$38953 ( \39268 , \22535 , \22411 );
nor \U$38954 ( \39269 , \39267 , \39268 );
xnor \U$38955 ( \39270 , \39269 , \22423 );
xor \U$38956 ( \39271 , \39266 , \39270 );
and \U$38957 ( \39272 , \22545 , \22435 );
and \U$38958 ( \39273 , \22556 , \22433 );
nor \U$38959 ( \39274 , \39272 , \39273 );
xnor \U$38960 ( \39275 , \39274 , \22445 );
xor \U$38961 ( \39276 , \39271 , \39275 );
xor \U$38962 ( \39277 , \39262 , \39276 );
and \U$38963 ( \39278 , \22429 , \22324 );
and \U$38964 ( \39279 , \22440 , \22322 );
nor \U$38965 ( \39280 , \39278 , \39279 );
xnor \U$38966 ( \39281 , \39280 , \22334 );
and \U$38967 ( \39282 , \22457 , \22345 );
and \U$38968 ( \39283 , \22468 , \22343 );
nor \U$38969 ( \39284 , \39282 , \39283 );
xnor \U$38970 ( \39285 , \39284 , \22355 );
xor \U$38971 ( \39286 , \39281 , \39285 );
and \U$38972 ( \39287 , \22478 , \22367 );
and \U$38973 ( \39288 , \22489 , \22365 );
nor \U$38974 ( \39289 , \39287 , \39288 );
xnor \U$38975 ( \39290 , \39289 , \22377 );
xor \U$38976 ( \39291 , \39286 , \39290 );
xor \U$38977 ( \39292 , \39277 , \39291 );
xor \U$38978 ( \39293 , \39248 , \39292 );
and \U$38979 ( \39294 , \39077 , \39081 );
and \U$38980 ( \39295 , \39081 , \39086 );
and \U$38981 ( \39296 , \39077 , \39086 );
or \U$38982 ( \39297 , \39294 , \39295 , \39296 );
nand \U$38983 ( \39298 , \22706 , \22596 );
xnor \U$38984 ( \39299 , \39298 , \22608 );
xor \U$38985 ( \39300 , \39297 , \39299 );
and \U$38986 ( \39301 , \22635 , \22530 );
and \U$38987 ( \39302 , \22646 , \22528 );
nor \U$38988 ( \39303 , \39301 , \39302 );
xnor \U$38989 ( \39304 , \39303 , \22540 );
and \U$38990 ( \39305 , \22665 , \22551 );
and \U$38991 ( \39306 , \22676 , \22549 );
nor \U$38992 ( \39307 , \39305 , \39306 );
xnor \U$38993 ( \39308 , \39307 , \22561 );
xor \U$38994 ( \39309 , \39304 , \39308 );
and \U$38995 ( \39310 , \22686 , \22573 );
and \U$38996 ( \39311 , \22696 , \22571 );
nor \U$38997 ( \39312 , \39310 , \39311 );
xnor \U$38998 ( \39313 , \39312 , \22583 );
xor \U$38999 ( \39314 , \39309 , \39313 );
xor \U$39000 ( \39315 , \39300 , \39314 );
xor \U$39001 ( \39316 , \39293 , \39315 );
and \U$39002 ( \39317 , \39073 , \39087 );
and \U$39003 ( \39318 , \39087 , \39102 );
and \U$39004 ( \39319 , \39073 , \39102 );
or \U$39005 ( \39320 , \39317 , \39318 , \39319 );
and \U$39006 ( \39321 , \39038 , \39052 );
and \U$39007 ( \39322 , \39052 , \39067 );
and \U$39008 ( \39323 , \39038 , \39067 );
or \U$39009 ( \39324 , \39321 , \39322 , \39323 );
xor \U$39010 ( \39325 , \39320 , \39324 );
and \U$39011 ( \39326 , \22181 , \22076 );
and \U$39012 ( \39327 , \22192 , \22073 );
nor \U$39013 ( \39328 , \39326 , \39327 );
xnor \U$39014 ( \39329 , \39328 , \22072 );
xor \U$39015 ( \39330 , \22608 , \39329 );
and \U$39016 ( \39331 , \22202 , \22095 );
and \U$39017 ( \39332 , \22213 , \22093 );
nor \U$39018 ( \39333 , \39331 , \39332 );
xnor \U$39019 ( \39334 , \39333 , \22105 );
xor \U$39020 ( \39335 , \39330 , \39334 );
xor \U$39021 ( \39336 , \39325 , \39335 );
xor \U$39022 ( \39337 , \39316 , \39336 );
and \U$39023 ( \39338 , \38999 , \39003 );
and \U$39024 ( \39339 , \39003 , \39008 );
and \U$39025 ( \39340 , \38999 , \39008 );
or \U$39026 ( \39341 , \39338 , \39339 , \39340 );
and \U$39027 ( \39342 , \38984 , \38988 );
and \U$39028 ( \39343 , \38988 , \38993 );
and \U$39029 ( \39344 , \38984 , \38993 );
or \U$39030 ( \39345 , \39342 , \39343 , \39344 );
xor \U$39031 ( \39346 , \39341 , \39345 );
and \U$39032 ( \39347 , \38970 , \38974 );
and \U$39033 ( \39348 , \38974 , \38979 );
and \U$39034 ( \39349 , \38970 , \38979 );
or \U$39035 ( \39350 , \39347 , \39348 , \39349 );
xor \U$39036 ( \39351 , \39346 , \39350 );
xor \U$39037 ( \39352 , \39337 , \39351 );
xor \U$39038 ( \39353 , \39204 , \39352 );
xor \U$39039 ( \39354 , \39195 , \39353 );
xor \U$39040 ( \39355 , \39181 , \39354 );
and \U$39041 ( \39356 , \39150 , \39154 );
and \U$39042 ( \39357 , \39154 , \39169 );
and \U$39043 ( \39358 , \39150 , \39169 );
or \U$39044 ( \39359 , \39356 , \39357 , \39358 );
and \U$39045 ( \39360 , \39130 , \39144 );
xor \U$39046 ( \39361 , \39359 , \39360 );
and \U$39047 ( \39362 , \38980 , \38994 );
and \U$39048 ( \39363 , \38994 , \39009 );
and \U$39049 ( \39364 , \38980 , \39009 );
or \U$39050 ( \39365 , \39362 , \39363 , \39364 );
and \U$39051 ( \39366 , \39042 , \39046 );
and \U$39052 ( \39367 , \39046 , \39051 );
and \U$39053 ( \39368 , \39042 , \39051 );
or \U$39054 ( \39369 , \39366 , \39367 , \39368 );
and \U$39055 ( \39370 , \39028 , \39032 );
and \U$39056 ( \39371 , \39032 , \39037 );
and \U$39057 ( \39372 , \39028 , \39037 );
or \U$39058 ( \39373 , \39370 , \39371 , \39372 );
xor \U$39059 ( \39374 , \39369 , \39373 );
and \U$39060 ( \39375 , \39092 , \39096 );
and \U$39061 ( \39376 , \39096 , \39101 );
and \U$39062 ( \39377 , \39092 , \39101 );
or \U$39063 ( \39378 , \39375 , \39376 , \39377 );
xor \U$39064 ( \39379 , \39374 , \39378 );
xor \U$39065 ( \39380 , \39365 , \39379 );
and \U$39066 ( \39381 , \39014 , \39018 );
and \U$39067 ( \39382 , \39018 , \39023 );
and \U$39068 ( \39383 , \39014 , \39023 );
or \U$39069 ( \39384 , \39381 , \39382 , \39383 );
and \U$39070 ( \39385 , \39118 , \39122 );
and \U$39071 ( \39386 , \39122 , \39127 );
and \U$39072 ( \39387 , \39118 , \39127 );
or \U$39073 ( \39388 , \39385 , \39386 , \39387 );
xor \U$39074 ( \39389 , \39384 , \39388 );
and \U$39075 ( \39390 , \39057 , \39061 );
and \U$39076 ( \39391 , \39061 , \39066 );
and \U$39077 ( \39392 , \39057 , \39066 );
or \U$39078 ( \39393 , \39390 , \39391 , \39392 );
xor \U$39079 ( \39394 , \39389 , \39393 );
xor \U$39080 ( \39395 , \39380 , \39394 );
xor \U$39081 ( \39396 , \39361 , \39395 );
xor \U$39082 ( \39397 , \39355 , \39396 );
and \U$39083 ( \39398 , \38960 , \38961 );
and \U$39084 ( \39399 , \38961 , \39171 );
and \U$39085 ( \39400 , \38960 , \39171 );
or \U$39086 ( \39401 , \39398 , \39399 , \39400 );
nor \U$39087 ( \39402 , \39397 , \39401 );
nor \U$39088 ( \39403 , \39177 , \39402 );
nand \U$39089 ( \39404 , \38956 , \39403 );
nor \U$39090 ( \39405 , \38527 , \39404 );
nand \U$39091 ( \39406 , \37732 , \39405 );
and \U$39092 ( \39407 , \39359 , \39360 );
and \U$39093 ( \39408 , \39360 , \39395 );
and \U$39094 ( \39409 , \39359 , \39395 );
or \U$39095 ( \39410 , \39407 , \39408 , \39409 );
and \U$39096 ( \39411 , \39195 , \39353 );
xor \U$39097 ( \39412 , \39410 , \39411 );
and \U$39098 ( \39413 , \39199 , \39203 );
and \U$39099 ( \39414 , \39203 , \39352 );
and \U$39100 ( \39415 , \39199 , \39352 );
or \U$39101 ( \39416 , \39413 , \39414 , \39415 );
and \U$39102 ( \39417 , \39262 , \39276 );
and \U$39103 ( \39418 , \39276 , \39291 );
and \U$39104 ( \39419 , \39262 , \39291 );
or \U$39105 ( \39420 , \39417 , \39418 , \39419 );
and \U$39106 ( \39421 , \39218 , \39232 );
and \U$39107 ( \39422 , \39232 , \39247 );
and \U$39108 ( \39423 , \39218 , \39247 );
or \U$39109 ( \39424 , \39421 , \39422 , \39423 );
xor \U$39110 ( \39425 , \39420 , \39424 );
and \U$39111 ( \39426 , \22192 , \22076 );
and \U$39112 ( \39427 , \22156 , \22073 );
nor \U$39113 ( \39428 , \39426 , \39427 );
xnor \U$39114 ( \39429 , \39428 , \22072 );
and \U$39115 ( \39430 , \22213 , \22095 );
and \U$39116 ( \39431 , \22181 , \22093 );
nor \U$39117 ( \39432 , \39430 , \39431 );
xnor \U$39118 ( \39433 , \39432 , \22105 );
xor \U$39119 ( \39434 , \39429 , \39433 );
and \U$39120 ( \39435 , \22235 , \22119 );
and \U$39121 ( \39436 , \22202 , \22117 );
nor \U$39122 ( \39437 , \39435 , \39436 );
xnor \U$39123 ( \39438 , \39437 , \22129 );
xor \U$39124 ( \39439 , \39434 , \39438 );
xor \U$39125 ( \39440 , \39425 , \39439 );
and \U$39126 ( \39441 , \39384 , \39388 );
and \U$39127 ( \39442 , \39388 , \39393 );
and \U$39128 ( \39443 , \39384 , \39393 );
or \U$39129 ( \39444 , \39441 , \39442 , \39443 );
and \U$39130 ( \39445 , \39369 , \39373 );
and \U$39131 ( \39446 , \39373 , \39378 );
and \U$39132 ( \39447 , \39369 , \39378 );
or \U$39133 ( \39448 , \39445 , \39446 , \39447 );
xor \U$39134 ( \39449 , \39444 , \39448 );
and \U$39135 ( \39450 , \39297 , \39299 );
and \U$39136 ( \39451 , \39299 , \39314 );
and \U$39137 ( \39452 , \39297 , \39314 );
or \U$39138 ( \39453 , \39450 , \39451 , \39452 );
xor \U$39139 ( \39454 , \39449 , \39453 );
xor \U$39140 ( \39455 , \39440 , \39454 );
and \U$39141 ( \39456 , \39208 , \39212 );
and \U$39142 ( \39457 , \39212 , \39217 );
and \U$39143 ( \39458 , \39208 , \39217 );
or \U$39144 ( \39459 , \39456 , \39457 , \39458 );
and \U$39145 ( \39460 , \39281 , \39285 );
and \U$39146 ( \39461 , \39285 , \39290 );
and \U$39147 ( \39462 , \39281 , \39290 );
or \U$39148 ( \39463 , \39460 , \39461 , \39462 );
xor \U$39149 ( \39464 , \39459 , \39463 );
and \U$39150 ( \39465 , \39266 , \39270 );
and \U$39151 ( \39466 , \39270 , \39275 );
and \U$39152 ( \39467 , \39266 , \39275 );
or \U$39153 ( \39468 , \39465 , \39466 , \39467 );
xor \U$39154 ( \39469 , \39464 , \39468 );
and \U$39155 ( \39470 , \22608 , \39329 );
and \U$39156 ( \39471 , \39329 , \39334 );
and \U$39157 ( \39472 , \22608 , \39334 );
or \U$39158 ( \39473 , \39470 , \39471 , \39472 );
and \U$39159 ( \39474 , \39237 , \39241 );
and \U$39160 ( \39475 , \39241 , \39246 );
and \U$39161 ( \39476 , \39237 , \39246 );
or \U$39162 ( \39477 , \39474 , \39475 , \39476 );
xor \U$39163 ( \39478 , \39473 , \39477 );
and \U$39164 ( \39479 , \39222 , \39226 );
and \U$39165 ( \39480 , \39226 , \39231 );
and \U$39166 ( \39481 , \39222 , \39231 );
or \U$39167 ( \39482 , \39479 , \39480 , \39481 );
xor \U$39168 ( \39483 , \39478 , \39482 );
xor \U$39169 ( \39484 , \39469 , \39483 );
and \U$39170 ( \39485 , \22397 , \22278 );
and \U$39171 ( \39486 , \22361 , \22276 );
nor \U$39172 ( \39487 , \39485 , \39486 );
xnor \U$39173 ( \39488 , \39487 , \22288 );
and \U$39174 ( \39489 , \22418 , \22300 );
and \U$39175 ( \39490 , \22386 , \22298 );
nor \U$39176 ( \39491 , \39489 , \39490 );
xnor \U$39177 ( \39492 , \39491 , \22310 );
xor \U$39178 ( \39493 , \39488 , \39492 );
and \U$39179 ( \39494 , \22440 , \22324 );
and \U$39180 ( \39495 , \22407 , \22322 );
nor \U$39181 ( \39496 , \39494 , \39495 );
xnor \U$39182 ( \39497 , \39496 , \22334 );
xor \U$39183 ( \39498 , \39493 , \39497 );
and \U$39184 ( \39499 , \22329 , \22208 );
and \U$39185 ( \39500 , \22294 , \22206 );
nor \U$39186 ( \39501 , \39499 , \39500 );
xnor \U$39187 ( \39502 , \39501 , \22218 );
and \U$39188 ( \39503 , \22350 , \22230 );
and \U$39189 ( \39504 , \22318 , \22228 );
nor \U$39190 ( \39505 , \39503 , \39504 );
xnor \U$39191 ( \39506 , \39505 , \22240 );
xor \U$39192 ( \39507 , \39502 , \39506 );
and \U$39193 ( \39508 , \22372 , \22257 );
and \U$39194 ( \39509 , \22339 , \22255 );
nor \U$39195 ( \39510 , \39508 , \39509 );
xnor \U$39196 ( \39511 , \39510 , \22267 );
xor \U$39197 ( \39512 , \39507 , \39511 );
xor \U$39198 ( \39513 , \39498 , \39512 );
and \U$39199 ( \39514 , \22262 , \22140 );
and \U$39200 ( \39515 , \22224 , \22138 );
nor \U$39201 ( \39516 , \39514 , \39515 );
xnor \U$39202 ( \39517 , \39516 , \22150 );
and \U$39203 ( \39518 , \22283 , \22162 );
and \U$39204 ( \39519 , \22251 , \22160 );
nor \U$39205 ( \39520 , \39518 , \39519 );
xnor \U$39206 ( \39521 , \39520 , \22172 );
xor \U$39207 ( \39522 , \39517 , \39521 );
and \U$39208 ( \39523 , \22305 , \22187 );
and \U$39209 ( \39524 , \22272 , \22185 );
nor \U$39210 ( \39525 , \39523 , \39524 );
xnor \U$39211 ( \39526 , \39525 , \22197 );
xor \U$39212 ( \39527 , \39522 , \39526 );
xor \U$39213 ( \39528 , \39513 , \39527 );
and \U$39214 ( \39529 , \22603 , \22484 );
and \U$39215 ( \39530 , \22567 , \22482 );
nor \U$39216 ( \39531 , \39529 , \39530 );
xnor \U$39217 ( \39532 , \39531 , \22494 );
and \U$39218 ( \39533 , \22624 , \22506 );
and \U$39219 ( \39534 , \22592 , \22504 );
nor \U$39220 ( \39535 , \39533 , \39534 );
xnor \U$39221 ( \39536 , \39535 , \22516 );
xor \U$39222 ( \39537 , \39532 , \39536 );
and \U$39223 ( \39538 , \22646 , \22530 );
and \U$39224 ( \39539 , \22613 , \22528 );
nor \U$39225 ( \39540 , \39538 , \39539 );
xnor \U$39226 ( \39541 , \39540 , \22540 );
xor \U$39227 ( \39542 , \39537 , \39541 );
and \U$39228 ( \39543 , \22535 , \22413 );
and \U$39229 ( \39544 , \22500 , \22411 );
nor \U$39230 ( \39545 , \39543 , \39544 );
xnor \U$39231 ( \39546 , \39545 , \22423 );
and \U$39232 ( \39547 , \22556 , \22435 );
and \U$39233 ( \39548 , \22524 , \22433 );
nor \U$39234 ( \39549 , \39547 , \39548 );
xnor \U$39235 ( \39550 , \39549 , \22445 );
xor \U$39236 ( \39551 , \39546 , \39550 );
and \U$39237 ( \39552 , \22578 , \22463 );
and \U$39238 ( \39553 , \22545 , \22461 );
nor \U$39239 ( \39554 , \39552 , \39553 );
xnor \U$39240 ( \39555 , \39554 , \22473 );
xor \U$39241 ( \39556 , \39551 , \39555 );
xor \U$39242 ( \39557 , \39542 , \39556 );
and \U$39243 ( \39558 , \22468 , \22345 );
and \U$39244 ( \39559 , \22429 , \22343 );
nor \U$39245 ( \39560 , \39558 , \39559 );
xnor \U$39246 ( \39561 , \39560 , \22355 );
and \U$39247 ( \39562 , \22489 , \22367 );
and \U$39248 ( \39563 , \22457 , \22365 );
nor \U$39249 ( \39564 , \39562 , \39563 );
xnor \U$39250 ( \39565 , \39564 , \22377 );
xor \U$39251 ( \39566 , \39561 , \39565 );
and \U$39252 ( \39567 , \22511 , \22392 );
and \U$39253 ( \39568 , \22478 , \22390 );
nor \U$39254 ( \39569 , \39567 , \39568 );
xnor \U$39255 ( \39570 , \39569 , \22402 );
xor \U$39256 ( \39571 , \39566 , \39570 );
xor \U$39257 ( \39572 , \39557 , \39571 );
xor \U$39258 ( \39573 , \39528 , \39572 );
and \U$39259 ( \39574 , \39252 , \39256 );
and \U$39260 ( \39575 , \39256 , \39261 );
and \U$39261 ( \39576 , \39252 , \39261 );
or \U$39262 ( \39577 , \39574 , \39575 , \39576 );
and \U$39263 ( \39578 , \39304 , \39308 );
and \U$39264 ( \39579 , \39308 , \39313 );
and \U$39265 ( \39580 , \39304 , \39313 );
or \U$39266 ( \39581 , \39578 , \39579 , \39580 );
xor \U$39267 ( \39582 , \39577 , \39581 );
and \U$39268 ( \39583 , \22676 , \22551 );
and \U$39269 ( \39584 , \22635 , \22549 );
nor \U$39270 ( \39585 , \39583 , \39584 );
xnor \U$39271 ( \39586 , \39585 , \22561 );
and \U$39272 ( \39587 , \22696 , \22573 );
and \U$39273 ( \39588 , \22665 , \22571 );
nor \U$39274 ( \39589 , \39587 , \39588 );
xnor \U$39275 ( \39590 , \39589 , \22583 );
xor \U$39276 ( \39591 , \39586 , \39590 );
and \U$39277 ( \39592 , \22706 , \22598 );
and \U$39278 ( \39593 , \22686 , \22596 );
nor \U$39279 ( \39594 , \39592 , \39593 );
xnor \U$39280 ( \39595 , \39594 , \22608 );
xor \U$39281 ( \39596 , \39591 , \39595 );
xor \U$39282 ( \39597 , \39582 , \39596 );
xor \U$39283 ( \39598 , \39573 , \39597 );
xor \U$39284 ( \39599 , \39484 , \39598 );
xor \U$39285 ( \39600 , \39455 , \39599 );
and \U$39286 ( \39601 , \39341 , \39345 );
and \U$39287 ( \39602 , \39345 , \39350 );
and \U$39288 ( \39603 , \39341 , \39350 );
or \U$39289 ( \39604 , \39601 , \39602 , \39603 );
and \U$39290 ( \39605 , \39320 , \39324 );
and \U$39291 ( \39606 , \39324 , \39335 );
and \U$39292 ( \39607 , \39320 , \39335 );
or \U$39293 ( \39608 , \39605 , \39606 , \39607 );
xor \U$39294 ( \39609 , \39604 , \39608 );
and \U$39295 ( \39610 , \39248 , \39292 );
and \U$39296 ( \39611 , \39292 , \39315 );
and \U$39297 ( \39612 , \39248 , \39315 );
or \U$39298 ( \39613 , \39610 , \39611 , \39612 );
xor \U$39299 ( \39614 , \39609 , \39613 );
xor \U$39300 ( \39615 , \39600 , \39614 );
xor \U$39301 ( \39616 , \39416 , \39615 );
and \U$39302 ( \39617 , \39185 , \39189 );
and \U$39303 ( \39618 , \39189 , \39194 );
and \U$39304 ( \39619 , \39185 , \39194 );
or \U$39305 ( \39620 , \39617 , \39618 , \39619 );
and \U$39306 ( \39621 , \39365 , \39379 );
and \U$39307 ( \39622 , \39379 , \39394 );
and \U$39308 ( \39623 , \39365 , \39394 );
or \U$39309 ( \39624 , \39621 , \39622 , \39623 );
xor \U$39310 ( \39625 , \39620 , \39624 );
and \U$39311 ( \39626 , \39316 , \39336 );
and \U$39312 ( \39627 , \39336 , \39351 );
and \U$39313 ( \39628 , \39316 , \39351 );
or \U$39314 ( \39629 , \39626 , \39627 , \39628 );
xor \U$39315 ( \39630 , \39625 , \39629 );
xor \U$39316 ( \39631 , \39616 , \39630 );
xor \U$39317 ( \39632 , \39412 , \39631 );
and \U$39318 ( \39633 , \39181 , \39354 );
and \U$39319 ( \39634 , \39354 , \39396 );
and \U$39320 ( \39635 , \39181 , \39396 );
or \U$39321 ( \39636 , \39633 , \39634 , \39635 );
nor \U$39322 ( \39637 , \39632 , \39636 );
and \U$39323 ( \39638 , \39416 , \39615 );
and \U$39324 ( \39639 , \39615 , \39630 );
and \U$39325 ( \39640 , \39416 , \39630 );
or \U$39326 ( \39641 , \39638 , \39639 , \39640 );
and \U$39327 ( \39642 , \39604 , \39608 );
and \U$39328 ( \39643 , \39608 , \39613 );
and \U$39329 ( \39644 , \39604 , \39613 );
or \U$39330 ( \39645 , \39642 , \39643 , \39644 );
and \U$39331 ( \39646 , \39469 , \39483 );
and \U$39332 ( \39647 , \39483 , \39598 );
and \U$39333 ( \39648 , \39469 , \39598 );
or \U$39334 ( \39649 , \39646 , \39647 , \39648 );
xor \U$39335 ( \39650 , \39645 , \39649 );
and \U$39336 ( \39651 , \39440 , \39454 );
xor \U$39337 ( \39652 , \39650 , \39651 );
xor \U$39338 ( \39653 , \39641 , \39652 );
and \U$39339 ( \39654 , \39620 , \39624 );
and \U$39340 ( \39655 , \39624 , \39629 );
and \U$39341 ( \39656 , \39620 , \39629 );
or \U$39342 ( \39657 , \39654 , \39655 , \39656 );
and \U$39343 ( \39658 , \39455 , \39599 );
and \U$39344 ( \39659 , \39599 , \39614 );
and \U$39345 ( \39660 , \39455 , \39614 );
or \U$39346 ( \39661 , \39658 , \39659 , \39660 );
xor \U$39347 ( \39662 , \39657 , \39661 );
and \U$39348 ( \39663 , \39542 , \39556 );
and \U$39349 ( \39664 , \39556 , \39571 );
and \U$39350 ( \39665 , \39542 , \39571 );
or \U$39351 ( \39666 , \39663 , \39664 , \39665 );
and \U$39352 ( \39667 , \39498 , \39512 );
and \U$39353 ( \39668 , \39512 , \39527 );
and \U$39354 ( \39669 , \39498 , \39527 );
or \U$39355 ( \39670 , \39667 , \39668 , \39669 );
xor \U$39356 ( \39671 , \39666 , \39670 );
and \U$39357 ( \39672 , \22272 , \22187 );
and \U$39358 ( \39673 , \22283 , \22185 );
nor \U$39359 ( \39674 , \39672 , \39673 );
xnor \U$39360 ( \39675 , \39674 , \22197 );
and \U$39361 ( \39676 , \22294 , \22208 );
and \U$39362 ( \39677 , \22305 , \22206 );
nor \U$39363 ( \39678 , \39676 , \39677 );
xnor \U$39364 ( \39679 , \39678 , \22218 );
xor \U$39365 ( \39680 , \39675 , \39679 );
and \U$39366 ( \39681 , \22318 , \22230 );
and \U$39367 ( \39682 , \22329 , \22228 );
nor \U$39368 ( \39683 , \39681 , \39682 );
xnor \U$39369 ( \39684 , \39683 , \22240 );
xor \U$39370 ( \39685 , \39680 , \39684 );
and \U$39371 ( \39686 , \22202 , \22119 );
and \U$39372 ( \39687 , \22213 , \22117 );
nor \U$39373 ( \39688 , \39686 , \39687 );
xnor \U$39374 ( \39689 , \39688 , \22129 );
and \U$39375 ( \39690 , \22224 , \22140 );
and \U$39376 ( \39691 , \22235 , \22138 );
nor \U$39377 ( \39692 , \39690 , \39691 );
xnor \U$39378 ( \39693 , \39692 , \22150 );
xor \U$39379 ( \39694 , \39689 , \39693 );
and \U$39380 ( \39695 , \22251 , \22162 );
and \U$39381 ( \39696 , \22262 , \22160 );
nor \U$39382 ( \39697 , \39695 , \39696 );
xnor \U$39383 ( \39698 , \39697 , \22172 );
xor \U$39384 ( \39699 , \39694 , \39698 );
xor \U$39385 ( \39700 , \39685 , \39699 );
and \U$39386 ( \39701 , \22156 , \22076 );
and \U$39387 ( \39702 , \22167 , \22073 );
nor \U$39388 ( \39703 , \39701 , \39702 );
xnor \U$39389 ( \39704 , \39703 , \22072 );
xor \U$39390 ( \39705 , \22629 , \39704 );
and \U$39391 ( \39706 , \22181 , \22095 );
and \U$39392 ( \39707 , \22192 , \22093 );
nor \U$39393 ( \39708 , \39706 , \39707 );
xnor \U$39394 ( \39709 , \39708 , \22105 );
xor \U$39395 ( \39710 , \39705 , \39709 );
xor \U$39396 ( \39711 , \39700 , \39710 );
xor \U$39397 ( \39712 , \39671 , \39711 );
and \U$39398 ( \39713 , \39473 , \39477 );
and \U$39399 ( \39714 , \39477 , \39482 );
and \U$39400 ( \39715 , \39473 , \39482 );
or \U$39401 ( \39716 , \39713 , \39714 , \39715 );
and \U$39402 ( \39717 , \39459 , \39463 );
and \U$39403 ( \39718 , \39463 , \39468 );
and \U$39404 ( \39719 , \39459 , \39468 );
or \U$39405 ( \39720 , \39717 , \39718 , \39719 );
xor \U$39406 ( \39721 , \39716 , \39720 );
and \U$39407 ( \39722 , \39577 , \39581 );
and \U$39408 ( \39723 , \39581 , \39596 );
and \U$39409 ( \39724 , \39577 , \39596 );
or \U$39410 ( \39725 , \39722 , \39723 , \39724 );
xor \U$39411 ( \39726 , \39721 , \39725 );
xor \U$39412 ( \39727 , \39712 , \39726 );
and \U$39413 ( \39728 , \39488 , \39492 );
and \U$39414 ( \39729 , \39492 , \39497 );
and \U$39415 ( \39730 , \39488 , \39497 );
or \U$39416 ( \39731 , \39728 , \39729 , \39730 );
and \U$39417 ( \39732 , \39561 , \39565 );
and \U$39418 ( \39733 , \39565 , \39570 );
and \U$39419 ( \39734 , \39561 , \39570 );
or \U$39420 ( \39735 , \39732 , \39733 , \39734 );
xor \U$39421 ( \39736 , \39731 , \39735 );
and \U$39422 ( \39737 , \39546 , \39550 );
and \U$39423 ( \39738 , \39550 , \39555 );
and \U$39424 ( \39739 , \39546 , \39555 );
or \U$39425 ( \39740 , \39737 , \39738 , \39739 );
xor \U$39426 ( \39741 , \39736 , \39740 );
and \U$39427 ( \39742 , \39429 , \39433 );
and \U$39428 ( \39743 , \39433 , \39438 );
and \U$39429 ( \39744 , \39429 , \39438 );
or \U$39430 ( \39745 , \39742 , \39743 , \39744 );
and \U$39431 ( \39746 , \39517 , \39521 );
and \U$39432 ( \39747 , \39521 , \39526 );
and \U$39433 ( \39748 , \39517 , \39526 );
or \U$39434 ( \39749 , \39746 , \39747 , \39748 );
xor \U$39435 ( \39750 , \39745 , \39749 );
and \U$39436 ( \39751 , \39502 , \39506 );
and \U$39437 ( \39752 , \39506 , \39511 );
and \U$39438 ( \39753 , \39502 , \39511 );
or \U$39439 ( \39754 , \39751 , \39752 , \39753 );
xor \U$39440 ( \39755 , \39750 , \39754 );
xor \U$39441 ( \39756 , \39741 , \39755 );
and \U$39442 ( \39757 , \22478 , \22392 );
and \U$39443 ( \39758 , \22489 , \22390 );
nor \U$39444 ( \39759 , \39757 , \39758 );
xnor \U$39445 ( \39760 , \39759 , \22402 );
and \U$39446 ( \39761 , \22500 , \22413 );
and \U$39447 ( \39762 , \22511 , \22411 );
nor \U$39448 ( \39763 , \39761 , \39762 );
xnor \U$39449 ( \39764 , \39763 , \22423 );
xor \U$39450 ( \39765 , \39760 , \39764 );
and \U$39451 ( \39766 , \22524 , \22435 );
and \U$39452 ( \39767 , \22535 , \22433 );
nor \U$39453 ( \39768 , \39766 , \39767 );
xnor \U$39454 ( \39769 , \39768 , \22445 );
xor \U$39455 ( \39770 , \39765 , \39769 );
and \U$39456 ( \39771 , \22407 , \22324 );
and \U$39457 ( \39772 , \22418 , \22322 );
nor \U$39458 ( \39773 , \39771 , \39772 );
xnor \U$39459 ( \39774 , \39773 , \22334 );
and \U$39460 ( \39775 , \22429 , \22345 );
and \U$39461 ( \39776 , \22440 , \22343 );
nor \U$39462 ( \39777 , \39775 , \39776 );
xnor \U$39463 ( \39778 , \39777 , \22355 );
xor \U$39464 ( \39779 , \39774 , \39778 );
and \U$39465 ( \39780 , \22457 , \22367 );
and \U$39466 ( \39781 , \22468 , \22365 );
nor \U$39467 ( \39782 , \39780 , \39781 );
xnor \U$39468 ( \39783 , \39782 , \22377 );
xor \U$39469 ( \39784 , \39779 , \39783 );
xor \U$39470 ( \39785 , \39770 , \39784 );
and \U$39471 ( \39786 , \22339 , \22257 );
and \U$39472 ( \39787 , \22350 , \22255 );
nor \U$39473 ( \39788 , \39786 , \39787 );
xnor \U$39474 ( \39789 , \39788 , \22267 );
and \U$39475 ( \39790 , \22361 , \22278 );
and \U$39476 ( \39791 , \22372 , \22276 );
nor \U$39477 ( \39792 , \39790 , \39791 );
xnor \U$39478 ( \39793 , \39792 , \22288 );
xor \U$39479 ( \39794 , \39789 , \39793 );
and \U$39480 ( \39795 , \22386 , \22300 );
and \U$39481 ( \39796 , \22397 , \22298 );
nor \U$39482 ( \39797 , \39795 , \39796 );
xnor \U$39483 ( \39798 , \39797 , \22310 );
xor \U$39484 ( \39799 , \39794 , \39798 );
xor \U$39485 ( \39800 , \39785 , \39799 );
nand \U$39486 ( \39801 , \22706 , \22617 );
xnor \U$39487 ( \39802 , \39801 , \22629 );
and \U$39488 ( \39803 , \22613 , \22530 );
and \U$39489 ( \39804 , \22624 , \22528 );
nor \U$39490 ( \39805 , \39803 , \39804 );
xnor \U$39491 ( \39806 , \39805 , \22540 );
and \U$39492 ( \39807 , \22635 , \22551 );
and \U$39493 ( \39808 , \22646 , \22549 );
nor \U$39494 ( \39809 , \39807 , \39808 );
xnor \U$39495 ( \39810 , \39809 , \22561 );
xor \U$39496 ( \39811 , \39806 , \39810 );
and \U$39497 ( \39812 , \22665 , \22573 );
and \U$39498 ( \39813 , \22676 , \22571 );
nor \U$39499 ( \39814 , \39812 , \39813 );
xnor \U$39500 ( \39815 , \39814 , \22583 );
xor \U$39501 ( \39816 , \39811 , \39815 );
xor \U$39502 ( \39817 , \39802 , \39816 );
and \U$39503 ( \39818 , \22545 , \22463 );
and \U$39504 ( \39819 , \22556 , \22461 );
nor \U$39505 ( \39820 , \39818 , \39819 );
xnor \U$39506 ( \39821 , \39820 , \22473 );
and \U$39507 ( \39822 , \22567 , \22484 );
and \U$39508 ( \39823 , \22578 , \22482 );
nor \U$39509 ( \39824 , \39822 , \39823 );
xnor \U$39510 ( \39825 , \39824 , \22494 );
xor \U$39511 ( \39826 , \39821 , \39825 );
and \U$39512 ( \39827 , \22592 , \22506 );
and \U$39513 ( \39828 , \22603 , \22504 );
nor \U$39514 ( \39829 , \39827 , \39828 );
xnor \U$39515 ( \39830 , \39829 , \22516 );
xor \U$39516 ( \39831 , \39826 , \39830 );
xor \U$39517 ( \39832 , \39817 , \39831 );
xor \U$39518 ( \39833 , \39800 , \39832 );
and \U$39519 ( \39834 , \39532 , \39536 );
and \U$39520 ( \39835 , \39536 , \39541 );
and \U$39521 ( \39836 , \39532 , \39541 );
or \U$39522 ( \39837 , \39834 , \39835 , \39836 );
and \U$39523 ( \39838 , \39586 , \39590 );
and \U$39524 ( \39839 , \39590 , \39595 );
and \U$39525 ( \39840 , \39586 , \39595 );
or \U$39526 ( \39841 , \39838 , \39839 , \39840 );
xor \U$39527 ( \39842 , \39837 , \39841 );
and \U$39528 ( \39843 , \22686 , \22598 );
and \U$39529 ( \39844 , \22696 , \22596 );
nor \U$39530 ( \39845 , \39843 , \39844 );
xnor \U$39531 ( \39846 , \39845 , \22608 );
xor \U$39532 ( \39847 , \39842 , \39846 );
xor \U$39533 ( \39848 , \39833 , \39847 );
xor \U$39534 ( \39849 , \39756 , \39848 );
xor \U$39535 ( \39850 , \39727 , \39849 );
and \U$39536 ( \39851 , \39444 , \39448 );
and \U$39537 ( \39852 , \39448 , \39453 );
and \U$39538 ( \39853 , \39444 , \39453 );
or \U$39539 ( \39854 , \39851 , \39852 , \39853 );
and \U$39540 ( \39855 , \39420 , \39424 );
and \U$39541 ( \39856 , \39424 , \39439 );
and \U$39542 ( \39857 , \39420 , \39439 );
or \U$39543 ( \39858 , \39855 , \39856 , \39857 );
xor \U$39544 ( \39859 , \39854 , \39858 );
and \U$39545 ( \39860 , \39528 , \39572 );
and \U$39546 ( \39861 , \39572 , \39597 );
and \U$39547 ( \39862 , \39528 , \39597 );
or \U$39548 ( \39863 , \39860 , \39861 , \39862 );
xor \U$39549 ( \39864 , \39859 , \39863 );
xor \U$39550 ( \39865 , \39850 , \39864 );
xor \U$39551 ( \39866 , \39662 , \39865 );
xor \U$39552 ( \39867 , \39653 , \39866 );
and \U$39553 ( \39868 , \39410 , \39411 );
and \U$39554 ( \39869 , \39411 , \39631 );
and \U$39555 ( \39870 , \39410 , \39631 );
or \U$39556 ( \39871 , \39868 , \39869 , \39870 );
nor \U$39557 ( \39872 , \39867 , \39871 );
nor \U$39558 ( \39873 , \39637 , \39872 );
and \U$39559 ( \39874 , \39657 , \39661 );
and \U$39560 ( \39875 , \39661 , \39865 );
and \U$39561 ( \39876 , \39657 , \39865 );
or \U$39562 ( \39877 , \39874 , \39875 , \39876 );
and \U$39563 ( \39878 , \39854 , \39858 );
and \U$39564 ( \39879 , \39858 , \39863 );
and \U$39565 ( \39880 , \39854 , \39863 );
or \U$39566 ( \39881 , \39878 , \39879 , \39880 );
and \U$39567 ( \39882 , \39741 , \39755 );
and \U$39568 ( \39883 , \39755 , \39848 );
and \U$39569 ( \39884 , \39741 , \39848 );
or \U$39570 ( \39885 , \39882 , \39883 , \39884 );
xor \U$39571 ( \39886 , \39881 , \39885 );
and \U$39572 ( \39887 , \39712 , \39726 );
xor \U$39573 ( \39888 , \39886 , \39887 );
xor \U$39574 ( \39889 , \39877 , \39888 );
and \U$39575 ( \39890 , \39645 , \39649 );
and \U$39576 ( \39891 , \39649 , \39651 );
and \U$39577 ( \39892 , \39645 , \39651 );
or \U$39578 ( \39893 , \39890 , \39891 , \39892 );
and \U$39579 ( \39894 , \39727 , \39849 );
and \U$39580 ( \39895 , \39849 , \39864 );
and \U$39581 ( \39896 , \39727 , \39864 );
or \U$39582 ( \39897 , \39894 , \39895 , \39896 );
xor \U$39583 ( \39898 , \39893 , \39897 );
and \U$39584 ( \39899 , \39745 , \39749 );
and \U$39585 ( \39900 , \39749 , \39754 );
and \U$39586 ( \39901 , \39745 , \39754 );
or \U$39587 ( \39902 , \39899 , \39900 , \39901 );
and \U$39588 ( \39903 , \39731 , \39735 );
and \U$39589 ( \39904 , \39735 , \39740 );
and \U$39590 ( \39905 , \39731 , \39740 );
or \U$39591 ( \39906 , \39903 , \39904 , \39905 );
xor \U$39592 ( \39907 , \39902 , \39906 );
and \U$39593 ( \39908 , \39837 , \39841 );
and \U$39594 ( \39909 , \39841 , \39846 );
and \U$39595 ( \39910 , \39837 , \39846 );
or \U$39596 ( \39911 , \39908 , \39909 , \39910 );
xor \U$39597 ( \39912 , \39907 , \39911 );
and \U$39598 ( \39913 , \39821 , \39825 );
and \U$39599 ( \39914 , \39825 , \39830 );
and \U$39600 ( \39915 , \39821 , \39830 );
or \U$39601 ( \39916 , \39913 , \39914 , \39915 );
and \U$39602 ( \39917 , \39806 , \39810 );
and \U$39603 ( \39918 , \39810 , \39815 );
and \U$39604 ( \39919 , \39806 , \39815 );
or \U$39605 ( \39920 , \39917 , \39918 , \39919 );
xor \U$39606 ( \39921 , \39916 , \39920 );
and \U$39607 ( \39922 , \22706 , \22619 );
and \U$39608 ( \39923 , \22686 , \22617 );
nor \U$39609 ( \39924 , \39922 , \39923 );
xnor \U$39610 ( \39925 , \39924 , \22629 );
xor \U$39611 ( \39926 , \39921 , \39925 );
and \U$39612 ( \39927 , \39789 , \39793 );
and \U$39613 ( \39928 , \39793 , \39798 );
and \U$39614 ( \39929 , \39789 , \39798 );
or \U$39615 ( \39930 , \39927 , \39928 , \39929 );
and \U$39616 ( \39931 , \39774 , \39778 );
and \U$39617 ( \39932 , \39778 , \39783 );
and \U$39618 ( \39933 , \39774 , \39783 );
or \U$39619 ( \39934 , \39931 , \39932 , \39933 );
xor \U$39620 ( \39935 , \39930 , \39934 );
and \U$39621 ( \39936 , \39760 , \39764 );
and \U$39622 ( \39937 , \39764 , \39769 );
and \U$39623 ( \39938 , \39760 , \39769 );
or \U$39624 ( \39939 , \39936 , \39937 , \39938 );
xor \U$39625 ( \39940 , \39935 , \39939 );
xor \U$39626 ( \39941 , \39926 , \39940 );
and \U$39627 ( \39942 , \22629 , \39704 );
and \U$39628 ( \39943 , \39704 , \39709 );
and \U$39629 ( \39944 , \22629 , \39709 );
or \U$39630 ( \39945 , \39942 , \39943 , \39944 );
and \U$39631 ( \39946 , \39689 , \39693 );
and \U$39632 ( \39947 , \39693 , \39698 );
and \U$39633 ( \39948 , \39689 , \39698 );
or \U$39634 ( \39949 , \39946 , \39947 , \39948 );
xor \U$39635 ( \39950 , \39945 , \39949 );
and \U$39636 ( \39951 , \39675 , \39679 );
and \U$39637 ( \39952 , \39679 , \39684 );
and \U$39638 ( \39953 , \39675 , \39684 );
or \U$39639 ( \39954 , \39951 , \39952 , \39953 );
xor \U$39640 ( \39955 , \39950 , \39954 );
xor \U$39641 ( \39956 , \39941 , \39955 );
and \U$39642 ( \39957 , \22235 , \22140 );
and \U$39643 ( \39958 , \22202 , \22138 );
nor \U$39644 ( \39959 , \39957 , \39958 );
xnor \U$39645 ( \39960 , \39959 , \22150 );
and \U$39646 ( \39961 , \22262 , \22162 );
and \U$39647 ( \39962 , \22224 , \22160 );
nor \U$39648 ( \39963 , \39961 , \39962 );
xnor \U$39649 ( \39964 , \39963 , \22172 );
xor \U$39650 ( \39965 , \39960 , \39964 );
and \U$39651 ( \39966 , \22283 , \22187 );
and \U$39652 ( \39967 , \22251 , \22185 );
nor \U$39653 ( \39968 , \39966 , \39967 );
xnor \U$39654 ( \39969 , \39968 , \22197 );
xor \U$39655 ( \39970 , \39965 , \39969 );
and \U$39656 ( \39971 , \22167 , \22076 );
and \U$39657 ( \39972 , \22134 , \22073 );
nor \U$39658 ( \39973 , \39971 , \39972 );
xnor \U$39659 ( \39974 , \39973 , \22072 );
and \U$39660 ( \39975 , \22192 , \22095 );
and \U$39661 ( \39976 , \22156 , \22093 );
nor \U$39662 ( \39977 , \39975 , \39976 );
xnor \U$39663 ( \39978 , \39977 , \22105 );
xor \U$39664 ( \39979 , \39974 , \39978 );
and \U$39665 ( \39980 , \22213 , \22119 );
and \U$39666 ( \39981 , \22181 , \22117 );
nor \U$39667 ( \39982 , \39980 , \39981 );
xnor \U$39668 ( \39983 , \39982 , \22129 );
xor \U$39669 ( \39984 , \39979 , \39983 );
xor \U$39670 ( \39985 , \39970 , \39984 );
and \U$39671 ( \39986 , \22440 , \22345 );
and \U$39672 ( \39987 , \22407 , \22343 );
nor \U$39673 ( \39988 , \39986 , \39987 );
xnor \U$39674 ( \39989 , \39988 , \22355 );
and \U$39675 ( \39990 , \22468 , \22367 );
and \U$39676 ( \39991 , \22429 , \22365 );
nor \U$39677 ( \39992 , \39990 , \39991 );
xnor \U$39678 ( \39993 , \39992 , \22377 );
xor \U$39679 ( \39994 , \39989 , \39993 );
and \U$39680 ( \39995 , \22489 , \22392 );
and \U$39681 ( \39996 , \22457 , \22390 );
nor \U$39682 ( \39997 , \39995 , \39996 );
xnor \U$39683 ( \39998 , \39997 , \22402 );
xor \U$39684 ( \39999 , \39994 , \39998 );
and \U$39685 ( \40000 , \22372 , \22278 );
and \U$39686 ( \40001 , \22339 , \22276 );
nor \U$39687 ( \40002 , \40000 , \40001 );
xnor \U$39688 ( \40003 , \40002 , \22288 );
and \U$39689 ( \40004 , \22397 , \22300 );
and \U$39690 ( \40005 , \22361 , \22298 );
nor \U$39691 ( \40006 , \40004 , \40005 );
xnor \U$39692 ( \40007 , \40006 , \22310 );
xor \U$39693 ( \40008 , \40003 , \40007 );
and \U$39694 ( \40009 , \22418 , \22324 );
and \U$39695 ( \40010 , \22386 , \22322 );
nor \U$39696 ( \40011 , \40009 , \40010 );
xnor \U$39697 ( \40012 , \40011 , \22334 );
xor \U$39698 ( \40013 , \40008 , \40012 );
xor \U$39699 ( \40014 , \39999 , \40013 );
and \U$39700 ( \40015 , \22305 , \22208 );
and \U$39701 ( \40016 , \22272 , \22206 );
nor \U$39702 ( \40017 , \40015 , \40016 );
xnor \U$39703 ( \40018 , \40017 , \22218 );
and \U$39704 ( \40019 , \22329 , \22230 );
and \U$39705 ( \40020 , \22294 , \22228 );
nor \U$39706 ( \40021 , \40019 , \40020 );
xnor \U$39707 ( \40022 , \40021 , \22240 );
xor \U$39708 ( \40023 , \40018 , \40022 );
and \U$39709 ( \40024 , \22350 , \22257 );
and \U$39710 ( \40025 , \22318 , \22255 );
nor \U$39711 ( \40026 , \40024 , \40025 );
xnor \U$39712 ( \40027 , \40026 , \22267 );
xor \U$39713 ( \40028 , \40023 , \40027 );
xor \U$39714 ( \40029 , \40014 , \40028 );
xor \U$39715 ( \40030 , \39985 , \40029 );
and \U$39716 ( \40031 , \22646 , \22551 );
and \U$39717 ( \40032 , \22613 , \22549 );
nor \U$39718 ( \40033 , \40031 , \40032 );
xnor \U$39719 ( \40034 , \40033 , \22561 );
and \U$39720 ( \40035 , \22676 , \22573 );
and \U$39721 ( \40036 , \22635 , \22571 );
nor \U$39722 ( \40037 , \40035 , \40036 );
xnor \U$39723 ( \40038 , \40037 , \22583 );
xor \U$39724 ( \40039 , \40034 , \40038 );
and \U$39725 ( \40040 , \22696 , \22598 );
and \U$39726 ( \40041 , \22665 , \22596 );
nor \U$39727 ( \40042 , \40040 , \40041 );
xnor \U$39728 ( \40043 , \40042 , \22608 );
xor \U$39729 ( \40044 , \40039 , \40043 );
and \U$39730 ( \40045 , \22578 , \22484 );
and \U$39731 ( \40046 , \22545 , \22482 );
nor \U$39732 ( \40047 , \40045 , \40046 );
xnor \U$39733 ( \40048 , \40047 , \22494 );
and \U$39734 ( \40049 , \22603 , \22506 );
and \U$39735 ( \40050 , \22567 , \22504 );
nor \U$39736 ( \40051 , \40049 , \40050 );
xnor \U$39737 ( \40052 , \40051 , \22516 );
xor \U$39738 ( \40053 , \40048 , \40052 );
and \U$39739 ( \40054 , \22624 , \22530 );
and \U$39740 ( \40055 , \22592 , \22528 );
nor \U$39741 ( \40056 , \40054 , \40055 );
xnor \U$39742 ( \40057 , \40056 , \22540 );
xor \U$39743 ( \40058 , \40053 , \40057 );
xor \U$39744 ( \40059 , \40044 , \40058 );
and \U$39745 ( \40060 , \22511 , \22413 );
and \U$39746 ( \40061 , \22478 , \22411 );
nor \U$39747 ( \40062 , \40060 , \40061 );
xnor \U$39748 ( \40063 , \40062 , \22423 );
and \U$39749 ( \40064 , \22535 , \22435 );
and \U$39750 ( \40065 , \22500 , \22433 );
nor \U$39751 ( \40066 , \40064 , \40065 );
xnor \U$39752 ( \40067 , \40066 , \22445 );
xor \U$39753 ( \40068 , \40063 , \40067 );
and \U$39754 ( \40069 , \22556 , \22463 );
and \U$39755 ( \40070 , \22524 , \22461 );
nor \U$39756 ( \40071 , \40069 , \40070 );
xnor \U$39757 ( \40072 , \40071 , \22473 );
xor \U$39758 ( \40073 , \40068 , \40072 );
xor \U$39759 ( \40074 , \40059 , \40073 );
xor \U$39760 ( \40075 , \40030 , \40074 );
xor \U$39761 ( \40076 , \39956 , \40075 );
and \U$39762 ( \40077 , \39802 , \39816 );
and \U$39763 ( \40078 , \39816 , \39831 );
and \U$39764 ( \40079 , \39802 , \39831 );
or \U$39765 ( \40080 , \40077 , \40078 , \40079 );
and \U$39766 ( \40081 , \39770 , \39784 );
and \U$39767 ( \40082 , \39784 , \39799 );
and \U$39768 ( \40083 , \39770 , \39799 );
or \U$39769 ( \40084 , \40081 , \40082 , \40083 );
xor \U$39770 ( \40085 , \40080 , \40084 );
and \U$39771 ( \40086 , \39685 , \39699 );
and \U$39772 ( \40087 , \39699 , \39710 );
and \U$39773 ( \40088 , \39685 , \39710 );
or \U$39774 ( \40089 , \40086 , \40087 , \40088 );
xor \U$39775 ( \40090 , \40085 , \40089 );
xor \U$39776 ( \40091 , \40076 , \40090 );
xor \U$39777 ( \40092 , \39912 , \40091 );
and \U$39778 ( \40093 , \39716 , \39720 );
and \U$39779 ( \40094 , \39720 , \39725 );
and \U$39780 ( \40095 , \39716 , \39725 );
or \U$39781 ( \40096 , \40093 , \40094 , \40095 );
and \U$39782 ( \40097 , \39666 , \39670 );
and \U$39783 ( \40098 , \39670 , \39711 );
and \U$39784 ( \40099 , \39666 , \39711 );
or \U$39785 ( \40100 , \40097 , \40098 , \40099 );
xor \U$39786 ( \40101 , \40096 , \40100 );
and \U$39787 ( \40102 , \39800 , \39832 );
and \U$39788 ( \40103 , \39832 , \39847 );
and \U$39789 ( \40104 , \39800 , \39847 );
or \U$39790 ( \40105 , \40102 , \40103 , \40104 );
xor \U$39791 ( \40106 , \40101 , \40105 );
xor \U$39792 ( \40107 , \40092 , \40106 );
xor \U$39793 ( \40108 , \39898 , \40107 );
xor \U$39794 ( \40109 , \39889 , \40108 );
and \U$39795 ( \40110 , \39641 , \39652 );
and \U$39796 ( \40111 , \39652 , \39866 );
and \U$39797 ( \40112 , \39641 , \39866 );
or \U$39798 ( \40113 , \40110 , \40111 , \40112 );
nor \U$39799 ( \40114 , \40109 , \40113 );
and \U$39800 ( \40115 , \39893 , \39897 );
and \U$39801 ( \40116 , \39897 , \40107 );
and \U$39802 ( \40117 , \39893 , \40107 );
or \U$39803 ( \40118 , \40115 , \40116 , \40117 );
and \U$39804 ( \40119 , \40096 , \40100 );
and \U$39805 ( \40120 , \40100 , \40105 );
and \U$39806 ( \40121 , \40096 , \40105 );
or \U$39807 ( \40122 , \40119 , \40120 , \40121 );
and \U$39808 ( \40123 , \39956 , \40075 );
and \U$39809 ( \40124 , \40075 , \40090 );
and \U$39810 ( \40125 , \39956 , \40090 );
or \U$39811 ( \40126 , \40123 , \40124 , \40125 );
xor \U$39812 ( \40127 , \40122 , \40126 );
and \U$39813 ( \40128 , \40044 , \40058 );
and \U$39814 ( \40129 , \40058 , \40073 );
and \U$39815 ( \40130 , \40044 , \40073 );
or \U$39816 ( \40131 , \40128 , \40129 , \40130 );
and \U$39817 ( \40132 , \39999 , \40013 );
and \U$39818 ( \40133 , \40013 , \40028 );
and \U$39819 ( \40134 , \39999 , \40028 );
or \U$39820 ( \40135 , \40132 , \40133 , \40134 );
xor \U$39821 ( \40136 , \40131 , \40135 );
and \U$39822 ( \40137 , \39970 , \39984 );
xor \U$39823 ( \40138 , \40136 , \40137 );
xor \U$39824 ( \40139 , \40127 , \40138 );
xor \U$39825 ( \40140 , \40118 , \40139 );
and \U$39826 ( \40141 , \39881 , \39885 );
and \U$39827 ( \40142 , \39885 , \39887 );
and \U$39828 ( \40143 , \39881 , \39887 );
or \U$39829 ( \40144 , \40141 , \40142 , \40143 );
and \U$39830 ( \40145 , \39912 , \40091 );
and \U$39831 ( \40146 , \40091 , \40106 );
and \U$39832 ( \40147 , \39912 , \40106 );
or \U$39833 ( \40148 , \40145 , \40146 , \40147 );
xor \U$39834 ( \40149 , \40144 , \40148 );
and \U$39835 ( \40150 , \39945 , \39949 );
and \U$39836 ( \40151 , \39949 , \39954 );
and \U$39837 ( \40152 , \39945 , \39954 );
or \U$39838 ( \40153 , \40150 , \40151 , \40152 );
and \U$39839 ( \40154 , \39930 , \39934 );
and \U$39840 ( \40155 , \39934 , \39939 );
and \U$39841 ( \40156 , \39930 , \39939 );
or \U$39842 ( \40157 , \40154 , \40155 , \40156 );
xor \U$39843 ( \40158 , \40153 , \40157 );
and \U$39844 ( \40159 , \39916 , \39920 );
and \U$39845 ( \40160 , \39920 , \39925 );
and \U$39846 ( \40161 , \39916 , \39925 );
or \U$39847 ( \40162 , \40159 , \40160 , \40161 );
xor \U$39848 ( \40163 , \40158 , \40162 );
and \U$39849 ( \40164 , \39926 , \39940 );
and \U$39850 ( \40165 , \39940 , \39955 );
and \U$39851 ( \40166 , \39926 , \39955 );
or \U$39852 ( \40167 , \40164 , \40165 , \40166 );
and \U$39853 ( \40168 , \40048 , \40052 );
and \U$39854 ( \40169 , \40052 , \40057 );
and \U$39855 ( \40170 , \40048 , \40057 );
or \U$39856 ( \40171 , \40168 , \40169 , \40170 );
and \U$39857 ( \40172 , \40034 , \40038 );
and \U$39858 ( \40173 , \40038 , \40043 );
and \U$39859 ( \40174 , \40034 , \40043 );
or \U$39860 ( \40175 , \40172 , \40173 , \40174 );
xor \U$39861 ( \40176 , \40171 , \40175 );
and \U$39862 ( \40177 , \22665 , \22598 );
and \U$39863 ( \40178 , \22676 , \22596 );
nor \U$39864 ( \40179 , \40177 , \40178 );
xnor \U$39865 ( \40180 , \40179 , \22608 );
and \U$39866 ( \40181 , \22686 , \22619 );
and \U$39867 ( \40182 , \22696 , \22617 );
nor \U$39868 ( \40183 , \40181 , \40182 );
xnor \U$39869 ( \40184 , \40183 , \22629 );
xor \U$39870 ( \40185 , \40180 , \40184 );
nand \U$39871 ( \40186 , \22706 , \22639 );
xnor \U$39872 ( \40187 , \40186 , \22651 );
xor \U$39873 ( \40188 , \40185 , \40187 );
xor \U$39874 ( \40189 , \40176 , \40188 );
and \U$39875 ( \40190 , \40003 , \40007 );
and \U$39876 ( \40191 , \40007 , \40012 );
and \U$39877 ( \40192 , \40003 , \40012 );
or \U$39878 ( \40193 , \40190 , \40191 , \40192 );
and \U$39879 ( \40194 , \39989 , \39993 );
and \U$39880 ( \40195 , \39993 , \39998 );
and \U$39881 ( \40196 , \39989 , \39998 );
or \U$39882 ( \40197 , \40194 , \40195 , \40196 );
xor \U$39883 ( \40198 , \40193 , \40197 );
and \U$39884 ( \40199 , \40063 , \40067 );
and \U$39885 ( \40200 , \40067 , \40072 );
and \U$39886 ( \40201 , \40063 , \40072 );
or \U$39887 ( \40202 , \40199 , \40200 , \40201 );
xor \U$39888 ( \40203 , \40198 , \40202 );
xor \U$39889 ( \40204 , \40189 , \40203 );
and \U$39890 ( \40205 , \39974 , \39978 );
and \U$39891 ( \40206 , \39978 , \39983 );
and \U$39892 ( \40207 , \39974 , \39983 );
or \U$39893 ( \40208 , \40205 , \40206 , \40207 );
and \U$39894 ( \40209 , \39960 , \39964 );
and \U$39895 ( \40210 , \39964 , \39969 );
and \U$39896 ( \40211 , \39960 , \39969 );
or \U$39897 ( \40212 , \40209 , \40210 , \40211 );
xor \U$39898 ( \40213 , \40208 , \40212 );
and \U$39899 ( \40214 , \40018 , \40022 );
and \U$39900 ( \40215 , \40022 , \40027 );
and \U$39901 ( \40216 , \40018 , \40027 );
or \U$39902 ( \40217 , \40214 , \40215 , \40216 );
xor \U$39903 ( \40218 , \40213 , \40217 );
xor \U$39904 ( \40219 , \40204 , \40218 );
xor \U$39905 ( \40220 , \40167 , \40219 );
and \U$39906 ( \40221 , \22181 , \22119 );
and \U$39907 ( \40222 , \22192 , \22117 );
nor \U$39908 ( \40223 , \40221 , \40222 );
xnor \U$39909 ( \40224 , \40223 , \22129 );
and \U$39910 ( \40225 , \22202 , \22140 );
and \U$39911 ( \40226 , \22213 , \22138 );
nor \U$39912 ( \40227 , \40225 , \40226 );
xnor \U$39913 ( \40228 , \40227 , \22150 );
xor \U$39914 ( \40229 , \40224 , \40228 );
and \U$39915 ( \40230 , \22224 , \22162 );
and \U$39916 ( \40231 , \22235 , \22160 );
nor \U$39917 ( \40232 , \40230 , \40231 );
xnor \U$39918 ( \40233 , \40232 , \22172 );
xor \U$39919 ( \40234 , \40229 , \40233 );
and \U$39920 ( \40235 , \22134 , \22076 );
and \U$39921 ( \40236 , \22145 , \22073 );
nor \U$39922 ( \40237 , \40235 , \40236 );
xnor \U$39923 ( \40238 , \40237 , \22072 );
xor \U$39924 ( \40239 , \22651 , \40238 );
and \U$39925 ( \40240 , \22156 , \22095 );
and \U$39926 ( \40241 , \22167 , \22093 );
nor \U$39927 ( \40242 , \40240 , \40241 );
xnor \U$39928 ( \40243 , \40242 , \22105 );
xor \U$39929 ( \40244 , \40239 , \40243 );
xor \U$39930 ( \40245 , \40234 , \40244 );
and \U$39931 ( \40246 , \22386 , \22324 );
and \U$39932 ( \40247 , \22397 , \22322 );
nor \U$39933 ( \40248 , \40246 , \40247 );
xnor \U$39934 ( \40249 , \40248 , \22334 );
and \U$39935 ( \40250 , \22407 , \22345 );
and \U$39936 ( \40251 , \22418 , \22343 );
nor \U$39937 ( \40252 , \40250 , \40251 );
xnor \U$39938 ( \40253 , \40252 , \22355 );
xor \U$39939 ( \40254 , \40249 , \40253 );
and \U$39940 ( \40255 , \22429 , \22367 );
and \U$39941 ( \40256 , \22440 , \22365 );
nor \U$39942 ( \40257 , \40255 , \40256 );
xnor \U$39943 ( \40258 , \40257 , \22377 );
xor \U$39944 ( \40259 , \40254 , \40258 );
and \U$39945 ( \40260 , \22318 , \22257 );
and \U$39946 ( \40261 , \22329 , \22255 );
nor \U$39947 ( \40262 , \40260 , \40261 );
xnor \U$39948 ( \40263 , \40262 , \22267 );
and \U$39949 ( \40264 , \22339 , \22278 );
and \U$39950 ( \40265 , \22350 , \22276 );
nor \U$39951 ( \40266 , \40264 , \40265 );
xnor \U$39952 ( \40267 , \40266 , \22288 );
xor \U$39953 ( \40268 , \40263 , \40267 );
and \U$39954 ( \40269 , \22361 , \22300 );
and \U$39955 ( \40270 , \22372 , \22298 );
nor \U$39956 ( \40271 , \40269 , \40270 );
xnor \U$39957 ( \40272 , \40271 , \22310 );
xor \U$39958 ( \40273 , \40268 , \40272 );
xor \U$39959 ( \40274 , \40259 , \40273 );
and \U$39960 ( \40275 , \22251 , \22187 );
and \U$39961 ( \40276 , \22262 , \22185 );
nor \U$39962 ( \40277 , \40275 , \40276 );
xnor \U$39963 ( \40278 , \40277 , \22197 );
and \U$39964 ( \40279 , \22272 , \22208 );
and \U$39965 ( \40280 , \22283 , \22206 );
nor \U$39966 ( \40281 , \40279 , \40280 );
xnor \U$39967 ( \40282 , \40281 , \22218 );
xor \U$39968 ( \40283 , \40278 , \40282 );
and \U$39969 ( \40284 , \22294 , \22230 );
and \U$39970 ( \40285 , \22305 , \22228 );
nor \U$39971 ( \40286 , \40284 , \40285 );
xnor \U$39972 ( \40287 , \40286 , \22240 );
xor \U$39973 ( \40288 , \40283 , \40287 );
xor \U$39974 ( \40289 , \40274 , \40288 );
xor \U$39975 ( \40290 , \40245 , \40289 );
and \U$39976 ( \40291 , \22592 , \22530 );
and \U$39977 ( \40292 , \22603 , \22528 );
nor \U$39978 ( \40293 , \40291 , \40292 );
xnor \U$39979 ( \40294 , \40293 , \22540 );
and \U$39980 ( \40295 , \22613 , \22551 );
and \U$39981 ( \40296 , \22624 , \22549 );
nor \U$39982 ( \40297 , \40295 , \40296 );
xnor \U$39983 ( \40298 , \40297 , \22561 );
xor \U$39984 ( \40299 , \40294 , \40298 );
and \U$39985 ( \40300 , \22635 , \22573 );
and \U$39986 ( \40301 , \22646 , \22571 );
nor \U$39987 ( \40302 , \40300 , \40301 );
xnor \U$39988 ( \40303 , \40302 , \22583 );
xor \U$39989 ( \40304 , \40299 , \40303 );
and \U$39990 ( \40305 , \22524 , \22463 );
and \U$39991 ( \40306 , \22535 , \22461 );
nor \U$39992 ( \40307 , \40305 , \40306 );
xnor \U$39993 ( \40308 , \40307 , \22473 );
and \U$39994 ( \40309 , \22545 , \22484 );
and \U$39995 ( \40310 , \22556 , \22482 );
nor \U$39996 ( \40311 , \40309 , \40310 );
xnor \U$39997 ( \40312 , \40311 , \22494 );
xor \U$39998 ( \40313 , \40308 , \40312 );
and \U$39999 ( \40314 , \22567 , \22506 );
and \U$40000 ( \40315 , \22578 , \22504 );
nor \U$40001 ( \40316 , \40314 , \40315 );
xnor \U$40002 ( \40317 , \40316 , \22516 );
xor \U$40003 ( \40318 , \40313 , \40317 );
xor \U$40004 ( \40319 , \40304 , \40318 );
and \U$40005 ( \40320 , \22457 , \22392 );
and \U$40006 ( \40321 , \22468 , \22390 );
nor \U$40007 ( \40322 , \40320 , \40321 );
xnor \U$40008 ( \40323 , \40322 , \22402 );
and \U$40009 ( \40324 , \22478 , \22413 );
and \U$40010 ( \40325 , \22489 , \22411 );
nor \U$40011 ( \40326 , \40324 , \40325 );
xnor \U$40012 ( \40327 , \40326 , \22423 );
xor \U$40013 ( \40328 , \40323 , \40327 );
and \U$40014 ( \40329 , \22500 , \22435 );
and \U$40015 ( \40330 , \22511 , \22433 );
nor \U$40016 ( \40331 , \40329 , \40330 );
xnor \U$40017 ( \40332 , \40331 , \22445 );
xor \U$40018 ( \40333 , \40328 , \40332 );
xor \U$40019 ( \40334 , \40319 , \40333 );
xor \U$40020 ( \40335 , \40290 , \40334 );
xor \U$40021 ( \40336 , \40220 , \40335 );
xor \U$40022 ( \40337 , \40163 , \40336 );
and \U$40023 ( \40338 , \39902 , \39906 );
and \U$40024 ( \40339 , \39906 , \39911 );
and \U$40025 ( \40340 , \39902 , \39911 );
or \U$40026 ( \40341 , \40338 , \40339 , \40340 );
and \U$40027 ( \40342 , \40080 , \40084 );
and \U$40028 ( \40343 , \40084 , \40089 );
and \U$40029 ( \40344 , \40080 , \40089 );
or \U$40030 ( \40345 , \40342 , \40343 , \40344 );
xor \U$40031 ( \40346 , \40341 , \40345 );
and \U$40032 ( \40347 , \39985 , \40029 );
and \U$40033 ( \40348 , \40029 , \40074 );
and \U$40034 ( \40349 , \39985 , \40074 );
or \U$40035 ( \40350 , \40347 , \40348 , \40349 );
xor \U$40036 ( \40351 , \40346 , \40350 );
xor \U$40037 ( \40352 , \40337 , \40351 );
xor \U$40038 ( \40353 , \40149 , \40352 );
xor \U$40039 ( \40354 , \40140 , \40353 );
and \U$40040 ( \40355 , \39877 , \39888 );
and \U$40041 ( \40356 , \39888 , \40108 );
and \U$40042 ( \40357 , \39877 , \40108 );
or \U$40043 ( \40358 , \40355 , \40356 , \40357 );
nor \U$40044 ( \40359 , \40354 , \40358 );
nor \U$40045 ( \40360 , \40114 , \40359 );
nand \U$40046 ( \40361 , \39873 , \40360 );
and \U$40047 ( \40362 , \40144 , \40148 );
and \U$40048 ( \40363 , \40148 , \40352 );
and \U$40049 ( \40364 , \40144 , \40352 );
or \U$40050 ( \40365 , \40362 , \40363 , \40364 );
and \U$40051 ( \40366 , \40341 , \40345 );
and \U$40052 ( \40367 , \40345 , \40350 );
and \U$40053 ( \40368 , \40341 , \40350 );
or \U$40054 ( \40369 , \40366 , \40367 , \40368 );
and \U$40055 ( \40370 , \40167 , \40219 );
and \U$40056 ( \40371 , \40219 , \40335 );
and \U$40057 ( \40372 , \40167 , \40335 );
or \U$40058 ( \40373 , \40370 , \40371 , \40372 );
xor \U$40059 ( \40374 , \40369 , \40373 );
and \U$40060 ( \40375 , \40304 , \40318 );
and \U$40061 ( \40376 , \40318 , \40333 );
and \U$40062 ( \40377 , \40304 , \40333 );
or \U$40063 ( \40378 , \40375 , \40376 , \40377 );
and \U$40064 ( \40379 , \40259 , \40273 );
and \U$40065 ( \40380 , \40273 , \40288 );
and \U$40066 ( \40381 , \40259 , \40288 );
or \U$40067 ( \40382 , \40379 , \40380 , \40381 );
xor \U$40068 ( \40383 , \40378 , \40382 );
and \U$40069 ( \40384 , \40234 , \40244 );
xor \U$40070 ( \40385 , \40383 , \40384 );
xor \U$40071 ( \40386 , \40374 , \40385 );
xor \U$40072 ( \40387 , \40365 , \40386 );
and \U$40073 ( \40388 , \40122 , \40126 );
and \U$40074 ( \40389 , \40126 , \40138 );
and \U$40075 ( \40390 , \40122 , \40138 );
or \U$40076 ( \40391 , \40388 , \40389 , \40390 );
and \U$40077 ( \40392 , \40163 , \40336 );
and \U$40078 ( \40393 , \40336 , \40351 );
and \U$40079 ( \40394 , \40163 , \40351 );
or \U$40080 ( \40395 , \40392 , \40393 , \40394 );
xor \U$40081 ( \40396 , \40391 , \40395 );
and \U$40082 ( \40397 , \40208 , \40212 );
and \U$40083 ( \40398 , \40212 , \40217 );
and \U$40084 ( \40399 , \40208 , \40217 );
or \U$40085 ( \40400 , \40397 , \40398 , \40399 );
and \U$40086 ( \40401 , \40193 , \40197 );
and \U$40087 ( \40402 , \40197 , \40202 );
and \U$40088 ( \40403 , \40193 , \40202 );
or \U$40089 ( \40404 , \40401 , \40402 , \40403 );
xor \U$40090 ( \40405 , \40400 , \40404 );
and \U$40091 ( \40406 , \40171 , \40175 );
and \U$40092 ( \40407 , \40175 , \40188 );
and \U$40093 ( \40408 , \40171 , \40188 );
or \U$40094 ( \40409 , \40406 , \40407 , \40408 );
xor \U$40095 ( \40410 , \40405 , \40409 );
and \U$40096 ( \40411 , \40189 , \40203 );
and \U$40097 ( \40412 , \40203 , \40218 );
and \U$40098 ( \40413 , \40189 , \40218 );
or \U$40099 ( \40414 , \40411 , \40412 , \40413 );
and \U$40100 ( \40415 , \40308 , \40312 );
and \U$40101 ( \40416 , \40312 , \40317 );
and \U$40102 ( \40417 , \40308 , \40317 );
or \U$40103 ( \40418 , \40415 , \40416 , \40417 );
and \U$40104 ( \40419 , \40294 , \40298 );
and \U$40105 ( \40420 , \40298 , \40303 );
and \U$40106 ( \40421 , \40294 , \40303 );
or \U$40107 ( \40422 , \40419 , \40420 , \40421 );
xor \U$40108 ( \40423 , \40418 , \40422 );
and \U$40109 ( \40424 , \40180 , \40184 );
and \U$40110 ( \40425 , \40184 , \40187 );
and \U$40111 ( \40426 , \40180 , \40187 );
or \U$40112 ( \40427 , \40424 , \40425 , \40426 );
xor \U$40113 ( \40428 , \40423 , \40427 );
and \U$40114 ( \40429 , \40263 , \40267 );
and \U$40115 ( \40430 , \40267 , \40272 );
and \U$40116 ( \40431 , \40263 , \40272 );
or \U$40117 ( \40432 , \40429 , \40430 , \40431 );
and \U$40118 ( \40433 , \40249 , \40253 );
and \U$40119 ( \40434 , \40253 , \40258 );
and \U$40120 ( \40435 , \40249 , \40258 );
or \U$40121 ( \40436 , \40433 , \40434 , \40435 );
xor \U$40122 ( \40437 , \40432 , \40436 );
and \U$40123 ( \40438 , \40323 , \40327 );
and \U$40124 ( \40439 , \40327 , \40332 );
and \U$40125 ( \40440 , \40323 , \40332 );
or \U$40126 ( \40441 , \40438 , \40439 , \40440 );
xor \U$40127 ( \40442 , \40437 , \40441 );
xor \U$40128 ( \40443 , \40428 , \40442 );
and \U$40129 ( \40444 , \22651 , \40238 );
and \U$40130 ( \40445 , \40238 , \40243 );
and \U$40131 ( \40446 , \22651 , \40243 );
or \U$40132 ( \40447 , \40444 , \40445 , \40446 );
and \U$40133 ( \40448 , \40224 , \40228 );
and \U$40134 ( \40449 , \40228 , \40233 );
and \U$40135 ( \40450 , \40224 , \40233 );
or \U$40136 ( \40451 , \40448 , \40449 , \40450 );
xor \U$40137 ( \40452 , \40447 , \40451 );
and \U$40138 ( \40453 , \40278 , \40282 );
and \U$40139 ( \40454 , \40282 , \40287 );
and \U$40140 ( \40455 , \40278 , \40287 );
or \U$40141 ( \40456 , \40453 , \40454 , \40455 );
xor \U$40142 ( \40457 , \40452 , \40456 );
xor \U$40143 ( \40458 , \40443 , \40457 );
xor \U$40144 ( \40459 , \40414 , \40458 );
and \U$40145 ( \40460 , \22283 , \22208 );
and \U$40146 ( \40461 , \22251 , \22206 );
nor \U$40147 ( \40462 , \40460 , \40461 );
xnor \U$40148 ( \40463 , \40462 , \22218 );
and \U$40149 ( \40464 , \22305 , \22230 );
and \U$40150 ( \40465 , \22272 , \22228 );
nor \U$40151 ( \40466 , \40464 , \40465 );
xnor \U$40152 ( \40467 , \40466 , \22240 );
xor \U$40153 ( \40468 , \40463 , \40467 );
and \U$40154 ( \40469 , \22329 , \22257 );
and \U$40155 ( \40470 , \22294 , \22255 );
nor \U$40156 ( \40471 , \40469 , \40470 );
xnor \U$40157 ( \40472 , \40471 , \22267 );
xor \U$40158 ( \40473 , \40468 , \40472 );
and \U$40159 ( \40474 , \22213 , \22140 );
and \U$40160 ( \40475 , \22181 , \22138 );
nor \U$40161 ( \40476 , \40474 , \40475 );
xnor \U$40162 ( \40477 , \40476 , \22150 );
and \U$40163 ( \40478 , \22235 , \22162 );
and \U$40164 ( \40479 , \22202 , \22160 );
nor \U$40165 ( \40480 , \40478 , \40479 );
xnor \U$40166 ( \40481 , \40480 , \22172 );
xor \U$40167 ( \40482 , \40477 , \40481 );
and \U$40168 ( \40483 , \22262 , \22187 );
and \U$40169 ( \40484 , \22224 , \22185 );
nor \U$40170 ( \40485 , \40483 , \40484 );
xnor \U$40171 ( \40486 , \40485 , \22197 );
xor \U$40172 ( \40487 , \40482 , \40486 );
xor \U$40173 ( \40488 , \40473 , \40487 );
and \U$40174 ( \40489 , \22145 , \22076 );
and \U$40175 ( \40490 , \22113 , \22073 );
nor \U$40176 ( \40491 , \40489 , \40490 );
xnor \U$40177 ( \40492 , \40491 , \22072 );
and \U$40178 ( \40493 , \22167 , \22095 );
and \U$40179 ( \40494 , \22134 , \22093 );
nor \U$40180 ( \40495 , \40493 , \40494 );
xnor \U$40181 ( \40496 , \40495 , \22105 );
xor \U$40182 ( \40497 , \40492 , \40496 );
and \U$40183 ( \40498 , \22192 , \22119 );
and \U$40184 ( \40499 , \22156 , \22117 );
nor \U$40185 ( \40500 , \40498 , \40499 );
xnor \U$40186 ( \40501 , \40500 , \22129 );
xor \U$40187 ( \40502 , \40497 , \40501 );
xor \U$40188 ( \40503 , \40488 , \40502 );
and \U$40189 ( \40504 , \22489 , \22413 );
and \U$40190 ( \40505 , \22457 , \22411 );
nor \U$40191 ( \40506 , \40504 , \40505 );
xnor \U$40192 ( \40507 , \40506 , \22423 );
and \U$40193 ( \40508 , \22511 , \22435 );
and \U$40194 ( \40509 , \22478 , \22433 );
nor \U$40195 ( \40510 , \40508 , \40509 );
xnor \U$40196 ( \40511 , \40510 , \22445 );
xor \U$40197 ( \40512 , \40507 , \40511 );
and \U$40198 ( \40513 , \22535 , \22463 );
and \U$40199 ( \40514 , \22500 , \22461 );
nor \U$40200 ( \40515 , \40513 , \40514 );
xnor \U$40201 ( \40516 , \40515 , \22473 );
xor \U$40202 ( \40517 , \40512 , \40516 );
and \U$40203 ( \40518 , \22418 , \22345 );
and \U$40204 ( \40519 , \22386 , \22343 );
nor \U$40205 ( \40520 , \40518 , \40519 );
xnor \U$40206 ( \40521 , \40520 , \22355 );
and \U$40207 ( \40522 , \22440 , \22367 );
and \U$40208 ( \40523 , \22407 , \22365 );
nor \U$40209 ( \40524 , \40522 , \40523 );
xnor \U$40210 ( \40525 , \40524 , \22377 );
xor \U$40211 ( \40526 , \40521 , \40525 );
and \U$40212 ( \40527 , \22468 , \22392 );
and \U$40213 ( \40528 , \22429 , \22390 );
nor \U$40214 ( \40529 , \40527 , \40528 );
xnor \U$40215 ( \40530 , \40529 , \22402 );
xor \U$40216 ( \40531 , \40526 , \40530 );
xor \U$40217 ( \40532 , \40517 , \40531 );
and \U$40218 ( \40533 , \22350 , \22278 );
and \U$40219 ( \40534 , \22318 , \22276 );
nor \U$40220 ( \40535 , \40533 , \40534 );
xnor \U$40221 ( \40536 , \40535 , \22288 );
and \U$40222 ( \40537 , \22372 , \22300 );
and \U$40223 ( \40538 , \22339 , \22298 );
nor \U$40224 ( \40539 , \40537 , \40538 );
xnor \U$40225 ( \40540 , \40539 , \22310 );
xor \U$40226 ( \40541 , \40536 , \40540 );
and \U$40227 ( \40542 , \22397 , \22324 );
and \U$40228 ( \40543 , \22361 , \22322 );
nor \U$40229 ( \40544 , \40542 , \40543 );
xnor \U$40230 ( \40545 , \40544 , \22334 );
xor \U$40231 ( \40546 , \40541 , \40545 );
xor \U$40232 ( \40547 , \40532 , \40546 );
xor \U$40233 ( \40548 , \40503 , \40547 );
and \U$40234 ( \40549 , \22696 , \22619 );
and \U$40235 ( \40550 , \22665 , \22617 );
nor \U$40236 ( \40551 , \40549 , \40550 );
xnor \U$40237 ( \40552 , \40551 , \22629 );
and \U$40238 ( \40553 , \22706 , \22641 );
and \U$40239 ( \40554 , \22686 , \22639 );
nor \U$40240 ( \40555 , \40553 , \40554 );
xnor \U$40241 ( \40556 , \40555 , \22651 );
xor \U$40242 ( \40557 , \40552 , \40556 );
and \U$40243 ( \40558 , \22624 , \22551 );
and \U$40244 ( \40559 , \22592 , \22549 );
nor \U$40245 ( \40560 , \40558 , \40559 );
xnor \U$40246 ( \40561 , \40560 , \22561 );
and \U$40247 ( \40562 , \22646 , \22573 );
and \U$40248 ( \40563 , \22613 , \22571 );
nor \U$40249 ( \40564 , \40562 , \40563 );
xnor \U$40250 ( \40565 , \40564 , \22583 );
xor \U$40251 ( \40566 , \40561 , \40565 );
and \U$40252 ( \40567 , \22676 , \22598 );
and \U$40253 ( \40568 , \22635 , \22596 );
nor \U$40254 ( \40569 , \40567 , \40568 );
xnor \U$40255 ( \40570 , \40569 , \22608 );
xor \U$40256 ( \40571 , \40566 , \40570 );
xor \U$40257 ( \40572 , \40557 , \40571 );
and \U$40258 ( \40573 , \22556 , \22484 );
and \U$40259 ( \40574 , \22524 , \22482 );
nor \U$40260 ( \40575 , \40573 , \40574 );
xnor \U$40261 ( \40576 , \40575 , \22494 );
and \U$40262 ( \40577 , \22578 , \22506 );
and \U$40263 ( \40578 , \22545 , \22504 );
nor \U$40264 ( \40579 , \40577 , \40578 );
xnor \U$40265 ( \40580 , \40579 , \22516 );
xor \U$40266 ( \40581 , \40576 , \40580 );
and \U$40267 ( \40582 , \22603 , \22530 );
and \U$40268 ( \40583 , \22567 , \22528 );
nor \U$40269 ( \40584 , \40582 , \40583 );
xnor \U$40270 ( \40585 , \40584 , \22540 );
xor \U$40271 ( \40586 , \40581 , \40585 );
xor \U$40272 ( \40587 , \40572 , \40586 );
xor \U$40273 ( \40588 , \40548 , \40587 );
xor \U$40274 ( \40589 , \40459 , \40588 );
xor \U$40275 ( \40590 , \40410 , \40589 );
and \U$40276 ( \40591 , \40153 , \40157 );
and \U$40277 ( \40592 , \40157 , \40162 );
and \U$40278 ( \40593 , \40153 , \40162 );
or \U$40279 ( \40594 , \40591 , \40592 , \40593 );
and \U$40280 ( \40595 , \40131 , \40135 );
and \U$40281 ( \40596 , \40135 , \40137 );
and \U$40282 ( \40597 , \40131 , \40137 );
or \U$40283 ( \40598 , \40595 , \40596 , \40597 );
xor \U$40284 ( \40599 , \40594 , \40598 );
and \U$40285 ( \40600 , \40245 , \40289 );
and \U$40286 ( \40601 , \40289 , \40334 );
and \U$40287 ( \40602 , \40245 , \40334 );
or \U$40288 ( \40603 , \40600 , \40601 , \40602 );
xor \U$40289 ( \40604 , \40599 , \40603 );
xor \U$40290 ( \40605 , \40590 , \40604 );
xor \U$40291 ( \40606 , \40396 , \40605 );
xor \U$40292 ( \40607 , \40387 , \40606 );
and \U$40293 ( \40608 , \40118 , \40139 );
and \U$40294 ( \40609 , \40139 , \40353 );
and \U$40295 ( \40610 , \40118 , \40353 );
or \U$40296 ( \40611 , \40608 , \40609 , \40610 );
nor \U$40297 ( \40612 , \40607 , \40611 );
and \U$40298 ( \40613 , \40391 , \40395 );
and \U$40299 ( \40614 , \40395 , \40605 );
and \U$40300 ( \40615 , \40391 , \40605 );
or \U$40301 ( \40616 , \40613 , \40614 , \40615 );
and \U$40302 ( \40617 , \40400 , \40404 );
and \U$40303 ( \40618 , \40404 , \40409 );
and \U$40304 ( \40619 , \40400 , \40409 );
or \U$40305 ( \40620 , \40617 , \40618 , \40619 );
and \U$40306 ( \40621 , \40378 , \40382 );
and \U$40307 ( \40622 , \40382 , \40384 );
and \U$40308 ( \40623 , \40378 , \40384 );
or \U$40309 ( \40624 , \40621 , \40622 , \40623 );
xor \U$40310 ( \40625 , \40620 , \40624 );
and \U$40311 ( \40626 , \40503 , \40547 );
and \U$40312 ( \40627 , \40547 , \40587 );
and \U$40313 ( \40628 , \40503 , \40587 );
or \U$40314 ( \40629 , \40626 , \40627 , \40628 );
xor \U$40315 ( \40630 , \40625 , \40629 );
and \U$40316 ( \40631 , \40594 , \40598 );
and \U$40317 ( \40632 , \40598 , \40603 );
and \U$40318 ( \40633 , \40594 , \40603 );
or \U$40319 ( \40634 , \40631 , \40632 , \40633 );
and \U$40320 ( \40635 , \40414 , \40458 );
and \U$40321 ( \40636 , \40458 , \40588 );
and \U$40322 ( \40637 , \40414 , \40588 );
or \U$40323 ( \40638 , \40635 , \40636 , \40637 );
xor \U$40324 ( \40639 , \40634 , \40638 );
and \U$40325 ( \40640 , \22113 , \22076 );
and \U$40326 ( \40641 , \22124 , \22073 );
nor \U$40327 ( \40642 , \40640 , \40641 );
xnor \U$40328 ( \40643 , \40642 , \22072 );
xor \U$40329 ( \40644 , \22681 , \40643 );
and \U$40330 ( \40645 , \22134 , \22095 );
and \U$40331 ( \40646 , \22145 , \22093 );
nor \U$40332 ( \40647 , \40645 , \40646 );
xnor \U$40333 ( \40648 , \40647 , \22105 );
xor \U$40334 ( \40649 , \40644 , \40648 );
and \U$40335 ( \40650 , \22294 , \22257 );
and \U$40336 ( \40651 , \22305 , \22255 );
nor \U$40337 ( \40652 , \40650 , \40651 );
xnor \U$40338 ( \40653 , \40652 , \22267 );
and \U$40339 ( \40654 , \22318 , \22278 );
and \U$40340 ( \40655 , \22329 , \22276 );
nor \U$40341 ( \40656 , \40654 , \40655 );
xnor \U$40342 ( \40657 , \40656 , \22288 );
xor \U$40343 ( \40658 , \40653 , \40657 );
and \U$40344 ( \40659 , \22339 , \22300 );
and \U$40345 ( \40660 , \22350 , \22298 );
nor \U$40346 ( \40661 , \40659 , \40660 );
xnor \U$40347 ( \40662 , \40661 , \22310 );
xor \U$40348 ( \40663 , \40658 , \40662 );
and \U$40349 ( \40664 , \22224 , \22187 );
and \U$40350 ( \40665 , \22235 , \22185 );
nor \U$40351 ( \40666 , \40664 , \40665 );
xnor \U$40352 ( \40667 , \40666 , \22197 );
and \U$40353 ( \40668 , \22251 , \22208 );
and \U$40354 ( \40669 , \22262 , \22206 );
nor \U$40355 ( \40670 , \40668 , \40669 );
xnor \U$40356 ( \40671 , \40670 , \22218 );
xor \U$40357 ( \40672 , \40667 , \40671 );
and \U$40358 ( \40673 , \22272 , \22230 );
and \U$40359 ( \40674 , \22283 , \22228 );
nor \U$40360 ( \40675 , \40673 , \40674 );
xnor \U$40361 ( \40676 , \40675 , \22240 );
xor \U$40362 ( \40677 , \40672 , \40676 );
xor \U$40363 ( \40678 , \40663 , \40677 );
and \U$40364 ( \40679 , \22156 , \22119 );
and \U$40365 ( \40680 , \22167 , \22117 );
nor \U$40366 ( \40681 , \40679 , \40680 );
xnor \U$40367 ( \40682 , \40681 , \22129 );
and \U$40368 ( \40683 , \22181 , \22140 );
and \U$40369 ( \40684 , \22192 , \22138 );
nor \U$40370 ( \40685 , \40683 , \40684 );
xnor \U$40371 ( \40686 , \40685 , \22150 );
xor \U$40372 ( \40687 , \40682 , \40686 );
and \U$40373 ( \40688 , \22202 , \22162 );
and \U$40374 ( \40689 , \22213 , \22160 );
nor \U$40375 ( \40690 , \40688 , \40689 );
xnor \U$40376 ( \40691 , \40690 , \22172 );
xor \U$40377 ( \40692 , \40687 , \40691 );
xor \U$40378 ( \40693 , \40678 , \40692 );
xor \U$40379 ( \40694 , \40649 , \40693 );
and \U$40380 ( \40695 , \22500 , \22463 );
and \U$40381 ( \40696 , \22511 , \22461 );
nor \U$40382 ( \40697 , \40695 , \40696 );
xnor \U$40383 ( \40698 , \40697 , \22473 );
and \U$40384 ( \40699 , \22524 , \22484 );
and \U$40385 ( \40700 , \22535 , \22482 );
nor \U$40386 ( \40701 , \40699 , \40700 );
xnor \U$40387 ( \40702 , \40701 , \22494 );
xor \U$40388 ( \40703 , \40698 , \40702 );
and \U$40389 ( \40704 , \22545 , \22506 );
and \U$40390 ( \40705 , \22556 , \22504 );
nor \U$40391 ( \40706 , \40704 , \40705 );
xnor \U$40392 ( \40707 , \40706 , \22516 );
xor \U$40393 ( \40708 , \40703 , \40707 );
and \U$40394 ( \40709 , \22429 , \22392 );
and \U$40395 ( \40710 , \22440 , \22390 );
nor \U$40396 ( \40711 , \40709 , \40710 );
xnor \U$40397 ( \40712 , \40711 , \22402 );
and \U$40398 ( \40713 , \22457 , \22413 );
and \U$40399 ( \40714 , \22468 , \22411 );
nor \U$40400 ( \40715 , \40713 , \40714 );
xnor \U$40401 ( \40716 , \40715 , \22423 );
xor \U$40402 ( \40717 , \40712 , \40716 );
and \U$40403 ( \40718 , \22478 , \22435 );
and \U$40404 ( \40719 , \22489 , \22433 );
nor \U$40405 ( \40720 , \40718 , \40719 );
xnor \U$40406 ( \40721 , \40720 , \22445 );
xor \U$40407 ( \40722 , \40717 , \40721 );
xor \U$40408 ( \40723 , \40708 , \40722 );
and \U$40409 ( \40724 , \22361 , \22324 );
and \U$40410 ( \40725 , \22372 , \22322 );
nor \U$40411 ( \40726 , \40724 , \40725 );
xnor \U$40412 ( \40727 , \40726 , \22334 );
and \U$40413 ( \40728 , \22386 , \22345 );
and \U$40414 ( \40729 , \22397 , \22343 );
nor \U$40415 ( \40730 , \40728 , \40729 );
xnor \U$40416 ( \40731 , \40730 , \22355 );
xor \U$40417 ( \40732 , \40727 , \40731 );
and \U$40418 ( \40733 , \22407 , \22367 );
and \U$40419 ( \40734 , \22418 , \22365 );
nor \U$40420 ( \40735 , \40733 , \40734 );
xnor \U$40421 ( \40736 , \40735 , \22377 );
xor \U$40422 ( \40737 , \40732 , \40736 );
xor \U$40423 ( \40738 , \40723 , \40737 );
xor \U$40424 ( \40739 , \40694 , \40738 );
and \U$40425 ( \40740 , \40557 , \40571 );
and \U$40426 ( \40741 , \40571 , \40586 );
and \U$40427 ( \40742 , \40557 , \40586 );
or \U$40428 ( \40743 , \40740 , \40741 , \40742 );
and \U$40429 ( \40744 , \40517 , \40531 );
and \U$40430 ( \40745 , \40531 , \40546 );
and \U$40431 ( \40746 , \40517 , \40546 );
or \U$40432 ( \40747 , \40744 , \40745 , \40746 );
xor \U$40433 ( \40748 , \40743 , \40747 );
and \U$40434 ( \40749 , \40473 , \40487 );
and \U$40435 ( \40750 , \40487 , \40502 );
and \U$40436 ( \40751 , \40473 , \40502 );
or \U$40437 ( \40752 , \40749 , \40750 , \40751 );
xor \U$40438 ( \40753 , \40748 , \40752 );
xor \U$40439 ( \40754 , \40739 , \40753 );
and \U$40440 ( \40755 , \40447 , \40451 );
and \U$40441 ( \40756 , \40451 , \40456 );
and \U$40442 ( \40757 , \40447 , \40456 );
or \U$40443 ( \40758 , \40755 , \40756 , \40757 );
and \U$40444 ( \40759 , \40432 , \40436 );
and \U$40445 ( \40760 , \40436 , \40441 );
and \U$40446 ( \40761 , \40432 , \40441 );
or \U$40447 ( \40762 , \40759 , \40760 , \40761 );
xor \U$40448 ( \40763 , \40758 , \40762 );
and \U$40449 ( \40764 , \40418 , \40422 );
and \U$40450 ( \40765 , \40422 , \40427 );
and \U$40451 ( \40766 , \40418 , \40427 );
or \U$40452 ( \40767 , \40764 , \40765 , \40766 );
xor \U$40453 ( \40768 , \40763 , \40767 );
xor \U$40454 ( \40769 , \40754 , \40768 );
xor \U$40455 ( \40770 , \40639 , \40769 );
xor \U$40456 ( \40771 , \40630 , \40770 );
xor \U$40457 ( \40772 , \40616 , \40771 );
and \U$40458 ( \40773 , \40369 , \40373 );
and \U$40459 ( \40774 , \40373 , \40385 );
and \U$40460 ( \40775 , \40369 , \40385 );
or \U$40461 ( \40776 , \40773 , \40774 , \40775 );
and \U$40462 ( \40777 , \40410 , \40589 );
and \U$40463 ( \40778 , \40589 , \40604 );
and \U$40464 ( \40779 , \40410 , \40604 );
or \U$40465 ( \40780 , \40777 , \40778 , \40779 );
xor \U$40466 ( \40781 , \40776 , \40780 );
and \U$40467 ( \40782 , \40428 , \40442 );
and \U$40468 ( \40783 , \40442 , \40457 );
and \U$40469 ( \40784 , \40428 , \40457 );
or \U$40470 ( \40785 , \40782 , \40783 , \40784 );
and \U$40471 ( \40786 , \40492 , \40496 );
and \U$40472 ( \40787 , \40496 , \40501 );
and \U$40473 ( \40788 , \40492 , \40501 );
or \U$40474 ( \40789 , \40786 , \40787 , \40788 );
and \U$40475 ( \40790 , \40477 , \40481 );
and \U$40476 ( \40791 , \40481 , \40486 );
and \U$40477 ( \40792 , \40477 , \40486 );
or \U$40478 ( \40793 , \40790 , \40791 , \40792 );
xor \U$40479 ( \40794 , \40789 , \40793 );
and \U$40480 ( \40795 , \40463 , \40467 );
and \U$40481 ( \40796 , \40467 , \40472 );
and \U$40482 ( \40797 , \40463 , \40472 );
or \U$40483 ( \40798 , \40795 , \40796 , \40797 );
xor \U$40484 ( \40799 , \40794 , \40798 );
xor \U$40485 ( \40800 , \40785 , \40799 );
nand \U$40486 ( \40801 , \22706 , \22669 );
xnor \U$40487 ( \40802 , \40801 , \22681 );
and \U$40488 ( \40803 , \22635 , \22598 );
and \U$40489 ( \40804 , \22646 , \22596 );
nor \U$40490 ( \40805 , \40803 , \40804 );
xnor \U$40491 ( \40806 , \40805 , \22608 );
and \U$40492 ( \40807 , \22665 , \22619 );
and \U$40493 ( \40808 , \22676 , \22617 );
nor \U$40494 ( \40809 , \40807 , \40808 );
xnor \U$40495 ( \40810 , \40809 , \22629 );
xor \U$40496 ( \40811 , \40806 , \40810 );
and \U$40497 ( \40812 , \22686 , \22641 );
and \U$40498 ( \40813 , \22696 , \22639 );
nor \U$40499 ( \40814 , \40812 , \40813 );
xnor \U$40500 ( \40815 , \40814 , \22651 );
xor \U$40501 ( \40816 , \40811 , \40815 );
xor \U$40502 ( \40817 , \40802 , \40816 );
and \U$40503 ( \40818 , \22567 , \22530 );
and \U$40504 ( \40819 , \22578 , \22528 );
nor \U$40505 ( \40820 , \40818 , \40819 );
xnor \U$40506 ( \40821 , \40820 , \22540 );
and \U$40507 ( \40822 , \22592 , \22551 );
and \U$40508 ( \40823 , \22603 , \22549 );
nor \U$40509 ( \40824 , \40822 , \40823 );
xnor \U$40510 ( \40825 , \40824 , \22561 );
xor \U$40511 ( \40826 , \40821 , \40825 );
and \U$40512 ( \40827 , \22613 , \22573 );
and \U$40513 ( \40828 , \22624 , \22571 );
nor \U$40514 ( \40829 , \40827 , \40828 );
xnor \U$40515 ( \40830 , \40829 , \22583 );
xor \U$40516 ( \40831 , \40826 , \40830 );
xor \U$40517 ( \40832 , \40817 , \40831 );
and \U$40518 ( \40833 , \40576 , \40580 );
and \U$40519 ( \40834 , \40580 , \40585 );
and \U$40520 ( \40835 , \40576 , \40585 );
or \U$40521 ( \40836 , \40833 , \40834 , \40835 );
and \U$40522 ( \40837 , \40561 , \40565 );
and \U$40523 ( \40838 , \40565 , \40570 );
and \U$40524 ( \40839 , \40561 , \40570 );
or \U$40525 ( \40840 , \40837 , \40838 , \40839 );
xor \U$40526 ( \40841 , \40836 , \40840 );
and \U$40527 ( \40842 , \40552 , \40556 );
xor \U$40528 ( \40843 , \40841 , \40842 );
xor \U$40529 ( \40844 , \40832 , \40843 );
and \U$40530 ( \40845 , \40536 , \40540 );
and \U$40531 ( \40846 , \40540 , \40545 );
and \U$40532 ( \40847 , \40536 , \40545 );
or \U$40533 ( \40848 , \40845 , \40846 , \40847 );
and \U$40534 ( \40849 , \40521 , \40525 );
and \U$40535 ( \40850 , \40525 , \40530 );
and \U$40536 ( \40851 , \40521 , \40530 );
or \U$40537 ( \40852 , \40849 , \40850 , \40851 );
xor \U$40538 ( \40853 , \40848 , \40852 );
and \U$40539 ( \40854 , \40507 , \40511 );
and \U$40540 ( \40855 , \40511 , \40516 );
and \U$40541 ( \40856 , \40507 , \40516 );
or \U$40542 ( \40857 , \40854 , \40855 , \40856 );
xor \U$40543 ( \40858 , \40853 , \40857 );
xor \U$40544 ( \40859 , \40844 , \40858 );
xor \U$40545 ( \40860 , \40800 , \40859 );
xor \U$40546 ( \40861 , \40781 , \40860 );
xor \U$40547 ( \40862 , \40772 , \40861 );
and \U$40548 ( \40863 , \40365 , \40386 );
and \U$40549 ( \40864 , \40386 , \40606 );
and \U$40550 ( \40865 , \40365 , \40606 );
or \U$40551 ( \40866 , \40863 , \40864 , \40865 );
nor \U$40552 ( \40867 , \40862 , \40866 );
nor \U$40553 ( \40868 , \40612 , \40867 );
and \U$40554 ( \40869 , \40776 , \40780 );
and \U$40555 ( \40870 , \40780 , \40860 );
and \U$40556 ( \40871 , \40776 , \40860 );
or \U$40557 ( \40872 , \40869 , \40870 , \40871 );
and \U$40558 ( \40873 , \40630 , \40770 );
xor \U$40559 ( \40874 , \40872 , \40873 );
and \U$40560 ( \40875 , \40634 , \40638 );
and \U$40561 ( \40876 , \40638 , \40769 );
and \U$40562 ( \40877 , \40634 , \40769 );
or \U$40563 ( \40878 , \40875 , \40876 , \40877 );
and \U$40564 ( \40879 , \40802 , \40816 );
and \U$40565 ( \40880 , \40816 , \40831 );
and \U$40566 ( \40881 , \40802 , \40831 );
or \U$40567 ( \40882 , \40879 , \40880 , \40881 );
and \U$40568 ( \40883 , \40708 , \40722 );
and \U$40569 ( \40884 , \40722 , \40737 );
and \U$40570 ( \40885 , \40708 , \40737 );
or \U$40571 ( \40886 , \40883 , \40884 , \40885 );
xor \U$40572 ( \40887 , \40882 , \40886 );
and \U$40573 ( \40888 , \40663 , \40677 );
and \U$40574 ( \40889 , \40677 , \40692 );
and \U$40575 ( \40890 , \40663 , \40692 );
or \U$40576 ( \40891 , \40888 , \40889 , \40890 );
xor \U$40577 ( \40892 , \40887 , \40891 );
and \U$40578 ( \40893 , \40789 , \40793 );
and \U$40579 ( \40894 , \40793 , \40798 );
and \U$40580 ( \40895 , \40789 , \40798 );
or \U$40581 ( \40896 , \40893 , \40894 , \40895 );
and \U$40582 ( \40897 , \40848 , \40852 );
and \U$40583 ( \40898 , \40852 , \40857 );
and \U$40584 ( \40899 , \40848 , \40857 );
or \U$40585 ( \40900 , \40897 , \40898 , \40899 );
xor \U$40586 ( \40901 , \40896 , \40900 );
and \U$40587 ( \40902 , \40836 , \40840 );
and \U$40588 ( \40903 , \40840 , \40842 );
and \U$40589 ( \40904 , \40836 , \40842 );
or \U$40590 ( \40905 , \40902 , \40903 , \40904 );
xor \U$40591 ( \40906 , \40901 , \40905 );
xor \U$40592 ( \40907 , \40892 , \40906 );
and \U$40593 ( \40908 , \40832 , \40843 );
and \U$40594 ( \40909 , \40843 , \40858 );
and \U$40595 ( \40910 , \40832 , \40858 );
or \U$40596 ( \40911 , \40908 , \40909 , \40910 );
and \U$40597 ( \40912 , \40698 , \40702 );
and \U$40598 ( \40913 , \40702 , \40707 );
and \U$40599 ( \40914 , \40698 , \40707 );
or \U$40600 ( \40915 , \40912 , \40913 , \40914 );
and \U$40601 ( \40916 , \40821 , \40825 );
and \U$40602 ( \40917 , \40825 , \40830 );
and \U$40603 ( \40918 , \40821 , \40830 );
or \U$40604 ( \40919 , \40916 , \40917 , \40918 );
xor \U$40605 ( \40920 , \40915 , \40919 );
and \U$40606 ( \40921 , \40806 , \40810 );
and \U$40607 ( \40922 , \40810 , \40815 );
and \U$40608 ( \40923 , \40806 , \40815 );
or \U$40609 ( \40924 , \40921 , \40922 , \40923 );
xor \U$40610 ( \40925 , \40920 , \40924 );
and \U$40611 ( \40926 , \40653 , \40657 );
and \U$40612 ( \40927 , \40657 , \40662 );
and \U$40613 ( \40928 , \40653 , \40662 );
or \U$40614 ( \40929 , \40926 , \40927 , \40928 );
and \U$40615 ( \40930 , \40727 , \40731 );
and \U$40616 ( \40931 , \40731 , \40736 );
and \U$40617 ( \40932 , \40727 , \40736 );
or \U$40618 ( \40933 , \40930 , \40931 , \40932 );
xor \U$40619 ( \40934 , \40929 , \40933 );
and \U$40620 ( \40935 , \40712 , \40716 );
and \U$40621 ( \40936 , \40716 , \40721 );
and \U$40622 ( \40937 , \40712 , \40721 );
or \U$40623 ( \40938 , \40935 , \40936 , \40937 );
xor \U$40624 ( \40939 , \40934 , \40938 );
xor \U$40625 ( \40940 , \40925 , \40939 );
and \U$40626 ( \40941 , \22681 , \40643 );
and \U$40627 ( \40942 , \40643 , \40648 );
and \U$40628 ( \40943 , \22681 , \40648 );
or \U$40629 ( \40944 , \40941 , \40942 , \40943 );
and \U$40630 ( \40945 , \40682 , \40686 );
and \U$40631 ( \40946 , \40686 , \40691 );
and \U$40632 ( \40947 , \40682 , \40691 );
or \U$40633 ( \40948 , \40945 , \40946 , \40947 );
xor \U$40634 ( \40949 , \40944 , \40948 );
and \U$40635 ( \40950 , \40667 , \40671 );
and \U$40636 ( \40951 , \40671 , \40676 );
and \U$40637 ( \40952 , \40667 , \40676 );
or \U$40638 ( \40953 , \40950 , \40951 , \40952 );
xor \U$40639 ( \40954 , \40949 , \40953 );
xor \U$40640 ( \40955 , \40940 , \40954 );
xor \U$40641 ( \40956 , \40911 , \40955 );
and \U$40642 ( \40957 , \22262 , \22208 );
and \U$40643 ( \40958 , \22224 , \22206 );
nor \U$40644 ( \40959 , \40957 , \40958 );
xnor \U$40645 ( \40960 , \40959 , \22218 );
and \U$40646 ( \40961 , \22283 , \22230 );
and \U$40647 ( \40962 , \22251 , \22228 );
nor \U$40648 ( \40963 , \40961 , \40962 );
xnor \U$40649 ( \40964 , \40963 , \22240 );
xor \U$40650 ( \40965 , \40960 , \40964 );
and \U$40651 ( \40966 , \22305 , \22257 );
and \U$40652 ( \40967 , \22272 , \22255 );
nor \U$40653 ( \40968 , \40966 , \40967 );
xnor \U$40654 ( \40969 , \40968 , \22267 );
xor \U$40655 ( \40970 , \40965 , \40969 );
and \U$40656 ( \40971 , \22192 , \22140 );
and \U$40657 ( \40972 , \22156 , \22138 );
nor \U$40658 ( \40973 , \40971 , \40972 );
xnor \U$40659 ( \40974 , \40973 , \22150 );
and \U$40660 ( \40975 , \22213 , \22162 );
and \U$40661 ( \40976 , \22181 , \22160 );
nor \U$40662 ( \40977 , \40975 , \40976 );
xnor \U$40663 ( \40978 , \40977 , \22172 );
xor \U$40664 ( \40979 , \40974 , \40978 );
and \U$40665 ( \40980 , \22235 , \22187 );
and \U$40666 ( \40981 , \22202 , \22185 );
nor \U$40667 ( \40982 , \40980 , \40981 );
xnor \U$40668 ( \40983 , \40982 , \22197 );
xor \U$40669 ( \40984 , \40979 , \40983 );
xor \U$40670 ( \40985 , \40970 , \40984 );
and \U$40671 ( \40986 , \22124 , \22076 );
and \U$40672 ( \40987 , \22089 , \22073 );
nor \U$40673 ( \40988 , \40986 , \40987 );
xnor \U$40674 ( \40989 , \40988 , \22072 );
and \U$40675 ( \40990 , \22145 , \22095 );
and \U$40676 ( \40991 , \22113 , \22093 );
nor \U$40677 ( \40992 , \40990 , \40991 );
xnor \U$40678 ( \40993 , \40992 , \22105 );
xor \U$40679 ( \40994 , \40989 , \40993 );
and \U$40680 ( \40995 , \22167 , \22119 );
and \U$40681 ( \40996 , \22134 , \22117 );
nor \U$40682 ( \40997 , \40995 , \40996 );
xnor \U$40683 ( \40998 , \40997 , \22129 );
xor \U$40684 ( \40999 , \40994 , \40998 );
xor \U$40685 ( \41000 , \40985 , \40999 );
and \U$40686 ( \41001 , \22468 , \22413 );
and \U$40687 ( \41002 , \22429 , \22411 );
nor \U$40688 ( \41003 , \41001 , \41002 );
xnor \U$40689 ( \41004 , \41003 , \22423 );
and \U$40690 ( \41005 , \22489 , \22435 );
and \U$40691 ( \41006 , \22457 , \22433 );
nor \U$40692 ( \41007 , \41005 , \41006 );
xnor \U$40693 ( \41008 , \41007 , \22445 );
xor \U$40694 ( \41009 , \41004 , \41008 );
and \U$40695 ( \41010 , \22511 , \22463 );
and \U$40696 ( \41011 , \22478 , \22461 );
nor \U$40697 ( \41012 , \41010 , \41011 );
xnor \U$40698 ( \41013 , \41012 , \22473 );
xor \U$40699 ( \41014 , \41009 , \41013 );
and \U$40700 ( \41015 , \22397 , \22345 );
and \U$40701 ( \41016 , \22361 , \22343 );
nor \U$40702 ( \41017 , \41015 , \41016 );
xnor \U$40703 ( \41018 , \41017 , \22355 );
and \U$40704 ( \41019 , \22418 , \22367 );
and \U$40705 ( \41020 , \22386 , \22365 );
nor \U$40706 ( \41021 , \41019 , \41020 );
xnor \U$40707 ( \41022 , \41021 , \22377 );
xor \U$40708 ( \41023 , \41018 , \41022 );
and \U$40709 ( \41024 , \22440 , \22392 );
and \U$40710 ( \41025 , \22407 , \22390 );
nor \U$40711 ( \41026 , \41024 , \41025 );
xnor \U$40712 ( \41027 , \41026 , \22402 );
xor \U$40713 ( \41028 , \41023 , \41027 );
xor \U$40714 ( \41029 , \41014 , \41028 );
and \U$40715 ( \41030 , \22329 , \22278 );
and \U$40716 ( \41031 , \22294 , \22276 );
nor \U$40717 ( \41032 , \41030 , \41031 );
xnor \U$40718 ( \41033 , \41032 , \22288 );
and \U$40719 ( \41034 , \22350 , \22300 );
and \U$40720 ( \41035 , \22318 , \22298 );
nor \U$40721 ( \41036 , \41034 , \41035 );
xnor \U$40722 ( \41037 , \41036 , \22310 );
xor \U$40723 ( \41038 , \41033 , \41037 );
and \U$40724 ( \41039 , \22372 , \22324 );
and \U$40725 ( \41040 , \22339 , \22322 );
nor \U$40726 ( \41041 , \41039 , \41040 );
xnor \U$40727 ( \41042 , \41041 , \22334 );
xor \U$40728 ( \41043 , \41038 , \41042 );
xor \U$40729 ( \41044 , \41029 , \41043 );
xor \U$40730 ( \41045 , \41000 , \41044 );
and \U$40731 ( \41046 , \22676 , \22619 );
and \U$40732 ( \41047 , \22635 , \22617 );
nor \U$40733 ( \41048 , \41046 , \41047 );
xnor \U$40734 ( \41049 , \41048 , \22629 );
and \U$40735 ( \41050 , \22696 , \22641 );
and \U$40736 ( \41051 , \22665 , \22639 );
nor \U$40737 ( \41052 , \41050 , \41051 );
xnor \U$40738 ( \41053 , \41052 , \22651 );
xor \U$40739 ( \41054 , \41049 , \41053 );
and \U$40740 ( \41055 , \22706 , \22671 );
and \U$40741 ( \41056 , \22686 , \22669 );
nor \U$40742 ( \41057 , \41055 , \41056 );
xnor \U$40743 ( \41058 , \41057 , \22681 );
xor \U$40744 ( \41059 , \41054 , \41058 );
and \U$40745 ( \41060 , \22603 , \22551 );
and \U$40746 ( \41061 , \22567 , \22549 );
nor \U$40747 ( \41062 , \41060 , \41061 );
xnor \U$40748 ( \41063 , \41062 , \22561 );
and \U$40749 ( \41064 , \22624 , \22573 );
and \U$40750 ( \41065 , \22592 , \22571 );
nor \U$40751 ( \41066 , \41064 , \41065 );
xnor \U$40752 ( \41067 , \41066 , \22583 );
xor \U$40753 ( \41068 , \41063 , \41067 );
and \U$40754 ( \41069 , \22646 , \22598 );
and \U$40755 ( \41070 , \22613 , \22596 );
nor \U$40756 ( \41071 , \41069 , \41070 );
xnor \U$40757 ( \41072 , \41071 , \22608 );
xor \U$40758 ( \41073 , \41068 , \41072 );
xor \U$40759 ( \41074 , \41059 , \41073 );
and \U$40760 ( \41075 , \22535 , \22484 );
and \U$40761 ( \41076 , \22500 , \22482 );
nor \U$40762 ( \41077 , \41075 , \41076 );
xnor \U$40763 ( \41078 , \41077 , \22494 );
and \U$40764 ( \41079 , \22556 , \22506 );
and \U$40765 ( \41080 , \22524 , \22504 );
nor \U$40766 ( \41081 , \41079 , \41080 );
xnor \U$40767 ( \41082 , \41081 , \22516 );
xor \U$40768 ( \41083 , \41078 , \41082 );
and \U$40769 ( \41084 , \22578 , \22530 );
and \U$40770 ( \41085 , \22545 , \22528 );
nor \U$40771 ( \41086 , \41084 , \41085 );
xnor \U$40772 ( \41087 , \41086 , \22540 );
xor \U$40773 ( \41088 , \41083 , \41087 );
xor \U$40774 ( \41089 , \41074 , \41088 );
xor \U$40775 ( \41090 , \41045 , \41089 );
xor \U$40776 ( \41091 , \40956 , \41090 );
xor \U$40777 ( \41092 , \40907 , \41091 );
and \U$40778 ( \41093 , \40758 , \40762 );
and \U$40779 ( \41094 , \40762 , \40767 );
and \U$40780 ( \41095 , \40758 , \40767 );
or \U$40781 ( \41096 , \41093 , \41094 , \41095 );
and \U$40782 ( \41097 , \40743 , \40747 );
and \U$40783 ( \41098 , \40747 , \40752 );
and \U$40784 ( \41099 , \40743 , \40752 );
or \U$40785 ( \41100 , \41097 , \41098 , \41099 );
xor \U$40786 ( \41101 , \41096 , \41100 );
and \U$40787 ( \41102 , \40649 , \40693 );
and \U$40788 ( \41103 , \40693 , \40738 );
and \U$40789 ( \41104 , \40649 , \40738 );
or \U$40790 ( \41105 , \41102 , \41103 , \41104 );
xor \U$40791 ( \41106 , \41101 , \41105 );
xor \U$40792 ( \41107 , \41092 , \41106 );
xor \U$40793 ( \41108 , \40878 , \41107 );
and \U$40794 ( \41109 , \40620 , \40624 );
and \U$40795 ( \41110 , \40624 , \40629 );
and \U$40796 ( \41111 , \40620 , \40629 );
or \U$40797 ( \41112 , \41109 , \41110 , \41111 );
and \U$40798 ( \41113 , \40785 , \40799 );
and \U$40799 ( \41114 , \40799 , \40859 );
and \U$40800 ( \41115 , \40785 , \40859 );
or \U$40801 ( \41116 , \41113 , \41114 , \41115 );
xor \U$40802 ( \41117 , \41112 , \41116 );
and \U$40803 ( \41118 , \40739 , \40753 );
and \U$40804 ( \41119 , \40753 , \40768 );
and \U$40805 ( \41120 , \40739 , \40768 );
or \U$40806 ( \41121 , \41118 , \41119 , \41120 );
xor \U$40807 ( \41122 , \41117 , \41121 );
xor \U$40808 ( \41123 , \41108 , \41122 );
xor \U$40809 ( \41124 , \40874 , \41123 );
and \U$40810 ( \41125 , \40616 , \40771 );
and \U$40811 ( \41126 , \40771 , \40861 );
and \U$40812 ( \41127 , \40616 , \40861 );
or \U$40813 ( \41128 , \41125 , \41126 , \41127 );
nor \U$40814 ( \41129 , \41124 , \41128 );
and \U$40815 ( \41130 , \40878 , \41107 );
and \U$40816 ( \41131 , \41107 , \41122 );
and \U$40817 ( \41132 , \40878 , \41122 );
or \U$40818 ( \41133 , \41130 , \41131 , \41132 );
and \U$40819 ( \41134 , \41096 , \41100 );
and \U$40820 ( \41135 , \41100 , \41105 );
and \U$40821 ( \41136 , \41096 , \41105 );
or \U$40822 ( \41137 , \41134 , \41135 , \41136 );
and \U$40823 ( \41138 , \40911 , \40955 );
and \U$40824 ( \41139 , \40955 , \41090 );
and \U$40825 ( \41140 , \40911 , \41090 );
or \U$40826 ( \41141 , \41138 , \41139 , \41140 );
xor \U$40827 ( \41142 , \41137 , \41141 );
and \U$40828 ( \41143 , \40892 , \40906 );
xor \U$40829 ( \41144 , \41142 , \41143 );
xor \U$40830 ( \41145 , \41133 , \41144 );
and \U$40831 ( \41146 , \41112 , \41116 );
and \U$40832 ( \41147 , \41116 , \41121 );
and \U$40833 ( \41148 , \41112 , \41121 );
or \U$40834 ( \41149 , \41146 , \41147 , \41148 );
and \U$40835 ( \41150 , \40907 , \41091 );
and \U$40836 ( \41151 , \41091 , \41106 );
and \U$40837 ( \41152 , \40907 , \41106 );
or \U$40838 ( \41153 , \41150 , \41151 , \41152 );
xor \U$40839 ( \41154 , \41149 , \41153 );
and \U$40840 ( \41155 , \22134 , \22119 );
and \U$40841 ( \41156 , \22145 , \22117 );
nor \U$40842 ( \41157 , \41155 , \41156 );
xnor \U$40843 ( \41158 , \41157 , \22129 );
and \U$40844 ( \41159 , \22156 , \22140 );
and \U$40845 ( \41160 , \22167 , \22138 );
nor \U$40846 ( \41161 , \41159 , \41160 );
xnor \U$40847 ( \41162 , \41161 , \22150 );
xor \U$40848 ( \41163 , \41158 , \41162 );
and \U$40849 ( \41164 , \22181 , \22162 );
and \U$40850 ( \41165 , \22192 , \22160 );
nor \U$40851 ( \41166 , \41164 , \41165 );
xnor \U$40852 ( \41167 , \41166 , \22172 );
xor \U$40853 ( \41168 , \41163 , \41167 );
and \U$40854 ( \41169 , \22089 , \22076 );
and \U$40855 ( \41170 , \22100 , \22073 );
nor \U$40856 ( \41171 , \41169 , \41170 );
xnor \U$40857 ( \41172 , \41171 , \22072 );
xor \U$40858 ( \41173 , \22701 , \41172 );
and \U$40859 ( \41174 , \22113 , \22095 );
and \U$40860 ( \41175 , \22124 , \22093 );
nor \U$40861 ( \41176 , \41174 , \41175 );
xnor \U$40862 ( \41177 , \41176 , \22105 );
xor \U$40863 ( \41178 , \41173 , \41177 );
xor \U$40864 ( \41179 , \41168 , \41178 );
and \U$40865 ( \41180 , \22339 , \22324 );
and \U$40866 ( \41181 , \22350 , \22322 );
nor \U$40867 ( \41182 , \41180 , \41181 );
xnor \U$40868 ( \41183 , \41182 , \22334 );
and \U$40869 ( \41184 , \22361 , \22345 );
and \U$40870 ( \41185 , \22372 , \22343 );
nor \U$40871 ( \41186 , \41184 , \41185 );
xnor \U$40872 ( \41187 , \41186 , \22355 );
xor \U$40873 ( \41188 , \41183 , \41187 );
and \U$40874 ( \41189 , \22386 , \22367 );
and \U$40875 ( \41190 , \22397 , \22365 );
nor \U$40876 ( \41191 , \41189 , \41190 );
xnor \U$40877 ( \41192 , \41191 , \22377 );
xor \U$40878 ( \41193 , \41188 , \41192 );
and \U$40879 ( \41194 , \22272 , \22257 );
and \U$40880 ( \41195 , \22283 , \22255 );
nor \U$40881 ( \41196 , \41194 , \41195 );
xnor \U$40882 ( \41197 , \41196 , \22267 );
and \U$40883 ( \41198 , \22294 , \22278 );
and \U$40884 ( \41199 , \22305 , \22276 );
nor \U$40885 ( \41200 , \41198 , \41199 );
xnor \U$40886 ( \41201 , \41200 , \22288 );
xor \U$40887 ( \41202 , \41197 , \41201 );
and \U$40888 ( \41203 , \22318 , \22300 );
and \U$40889 ( \41204 , \22329 , \22298 );
nor \U$40890 ( \41205 , \41203 , \41204 );
xnor \U$40891 ( \41206 , \41205 , \22310 );
xor \U$40892 ( \41207 , \41202 , \41206 );
xor \U$40893 ( \41208 , \41193 , \41207 );
and \U$40894 ( \41209 , \22202 , \22187 );
and \U$40895 ( \41210 , \22213 , \22185 );
nor \U$40896 ( \41211 , \41209 , \41210 );
xnor \U$40897 ( \41212 , \41211 , \22197 );
and \U$40898 ( \41213 , \22224 , \22208 );
and \U$40899 ( \41214 , \22235 , \22206 );
nor \U$40900 ( \41215 , \41213 , \41214 );
xnor \U$40901 ( \41216 , \41215 , \22218 );
xor \U$40902 ( \41217 , \41212 , \41216 );
and \U$40903 ( \41218 , \22251 , \22230 );
and \U$40904 ( \41219 , \22262 , \22228 );
nor \U$40905 ( \41220 , \41218 , \41219 );
xnor \U$40906 ( \41221 , \41220 , \22240 );
xor \U$40907 ( \41222 , \41217 , \41221 );
xor \U$40908 ( \41223 , \41208 , \41222 );
xor \U$40909 ( \41224 , \41179 , \41223 );
and \U$40910 ( \41225 , \41059 , \41073 );
and \U$40911 ( \41226 , \41073 , \41088 );
and \U$40912 ( \41227 , \41059 , \41088 );
or \U$40913 ( \41228 , \41225 , \41226 , \41227 );
and \U$40914 ( \41229 , \41014 , \41028 );
and \U$40915 ( \41230 , \41028 , \41043 );
and \U$40916 ( \41231 , \41014 , \41043 );
or \U$40917 ( \41232 , \41229 , \41230 , \41231 );
xor \U$40918 ( \41233 , \41228 , \41232 );
and \U$40919 ( \41234 , \40970 , \40984 );
and \U$40920 ( \41235 , \40984 , \40999 );
and \U$40921 ( \41236 , \40970 , \40999 );
or \U$40922 ( \41237 , \41234 , \41235 , \41236 );
xor \U$40923 ( \41238 , \41233 , \41237 );
xor \U$40924 ( \41239 , \41224 , \41238 );
and \U$40925 ( \41240 , \40944 , \40948 );
and \U$40926 ( \41241 , \40948 , \40953 );
and \U$40927 ( \41242 , \40944 , \40953 );
or \U$40928 ( \41243 , \41240 , \41241 , \41242 );
and \U$40929 ( \41244 , \40929 , \40933 );
and \U$40930 ( \41245 , \40933 , \40938 );
and \U$40931 ( \41246 , \40929 , \40938 );
or \U$40932 ( \41247 , \41244 , \41245 , \41246 );
xor \U$40933 ( \41248 , \41243 , \41247 );
and \U$40934 ( \41249 , \40915 , \40919 );
and \U$40935 ( \41250 , \40919 , \40924 );
and \U$40936 ( \41251 , \40915 , \40924 );
or \U$40937 ( \41252 , \41249 , \41250 , \41251 );
xor \U$40938 ( \41253 , \41248 , \41252 );
xor \U$40939 ( \41254 , \41239 , \41253 );
and \U$40940 ( \41255 , \40925 , \40939 );
and \U$40941 ( \41256 , \40939 , \40954 );
and \U$40942 ( \41257 , \40925 , \40954 );
or \U$40943 ( \41258 , \41255 , \41256 , \41257 );
and \U$40944 ( \41259 , \41033 , \41037 );
and \U$40945 ( \41260 , \41037 , \41042 );
and \U$40946 ( \41261 , \41033 , \41042 );
or \U$40947 ( \41262 , \41259 , \41260 , \41261 );
and \U$40948 ( \41263 , \41018 , \41022 );
and \U$40949 ( \41264 , \41022 , \41027 );
and \U$40950 ( \41265 , \41018 , \41027 );
or \U$40951 ( \41266 , \41263 , \41264 , \41265 );
xor \U$40952 ( \41267 , \41262 , \41266 );
and \U$40953 ( \41268 , \41004 , \41008 );
and \U$40954 ( \41269 , \41008 , \41013 );
and \U$40955 ( \41270 , \41004 , \41013 );
or \U$40956 ( \41271 , \41268 , \41269 , \41270 );
xor \U$40957 ( \41272 , \41267 , \41271 );
and \U$40958 ( \41273 , \40989 , \40993 );
and \U$40959 ( \41274 , \40993 , \40998 );
and \U$40960 ( \41275 , \40989 , \40998 );
or \U$40961 ( \41276 , \41273 , \41274 , \41275 );
and \U$40962 ( \41277 , \40974 , \40978 );
and \U$40963 ( \41278 , \40978 , \40983 );
and \U$40964 ( \41279 , \40974 , \40983 );
or \U$40965 ( \41280 , \41277 , \41278 , \41279 );
xor \U$40966 ( \41281 , \41276 , \41280 );
and \U$40967 ( \41282 , \40960 , \40964 );
and \U$40968 ( \41283 , \40964 , \40969 );
and \U$40969 ( \41284 , \40960 , \40969 );
or \U$40970 ( \41285 , \41282 , \41283 , \41284 );
xor \U$40971 ( \41286 , \41281 , \41285 );
xor \U$40972 ( \41287 , \41272 , \41286 );
xor \U$40973 ( \41288 , \41258 , \41287 );
and \U$40974 ( \41289 , \22545 , \22530 );
and \U$40975 ( \41290 , \22556 , \22528 );
nor \U$40976 ( \41291 , \41289 , \41290 );
xnor \U$40977 ( \41292 , \41291 , \22540 );
and \U$40978 ( \41293 , \22567 , \22551 );
and \U$40979 ( \41294 , \22578 , \22549 );
nor \U$40980 ( \41295 , \41293 , \41294 );
xnor \U$40981 ( \41296 , \41295 , \22561 );
xor \U$40982 ( \41297 , \41292 , \41296 );
and \U$40983 ( \41298 , \22592 , \22573 );
and \U$40984 ( \41299 , \22603 , \22571 );
nor \U$40985 ( \41300 , \41298 , \41299 );
xnor \U$40986 ( \41301 , \41300 , \22583 );
xor \U$40987 ( \41302 , \41297 , \41301 );
and \U$40988 ( \41303 , \22478 , \22463 );
and \U$40989 ( \41304 , \22489 , \22461 );
nor \U$40990 ( \41305 , \41303 , \41304 );
xnor \U$40991 ( \41306 , \41305 , \22473 );
and \U$40992 ( \41307 , \22500 , \22484 );
and \U$40993 ( \41308 , \22511 , \22482 );
nor \U$40994 ( \41309 , \41307 , \41308 );
xnor \U$40995 ( \41310 , \41309 , \22494 );
xor \U$40996 ( \41311 , \41306 , \41310 );
and \U$40997 ( \41312 , \22524 , \22506 );
and \U$40998 ( \41313 , \22535 , \22504 );
nor \U$40999 ( \41314 , \41312 , \41313 );
xnor \U$41000 ( \41315 , \41314 , \22516 );
xor \U$41001 ( \41316 , \41311 , \41315 );
xor \U$41002 ( \41317 , \41302 , \41316 );
and \U$41003 ( \41318 , \22407 , \22392 );
and \U$41004 ( \41319 , \22418 , \22390 );
nor \U$41005 ( \41320 , \41318 , \41319 );
xnor \U$41006 ( \41321 , \41320 , \22402 );
and \U$41007 ( \41322 , \22429 , \22413 );
and \U$41008 ( \41323 , \22440 , \22411 );
nor \U$41009 ( \41324 , \41322 , \41323 );
xnor \U$41010 ( \41325 , \41324 , \22423 );
xor \U$41011 ( \41326 , \41321 , \41325 );
and \U$41012 ( \41327 , \22457 , \22435 );
and \U$41013 ( \41328 , \22468 , \22433 );
nor \U$41014 ( \41329 , \41327 , \41328 );
xnor \U$41015 ( \41330 , \41329 , \22445 );
xor \U$41016 ( \41331 , \41326 , \41330 );
xor \U$41017 ( \41332 , \41317 , \41331 );
and \U$41018 ( \41333 , \22686 , \22671 );
and \U$41019 ( \41334 , \22696 , \22669 );
nor \U$41020 ( \41335 , \41333 , \41334 );
xnor \U$41021 ( \41336 , \41335 , \22681 );
nand \U$41022 ( \41337 , \22706 , \22689 );
xnor \U$41023 ( \41338 , \41337 , \22701 );
xor \U$41024 ( \41339 , \41336 , \41338 );
and \U$41025 ( \41340 , \22613 , \22598 );
and \U$41026 ( \41341 , \22624 , \22596 );
nor \U$41027 ( \41342 , \41340 , \41341 );
xnor \U$41028 ( \41343 , \41342 , \22608 );
and \U$41029 ( \41344 , \22635 , \22619 );
and \U$41030 ( \41345 , \22646 , \22617 );
nor \U$41031 ( \41346 , \41344 , \41345 );
xnor \U$41032 ( \41347 , \41346 , \22629 );
xor \U$41033 ( \41348 , \41343 , \41347 );
and \U$41034 ( \41349 , \22665 , \22641 );
and \U$41035 ( \41350 , \22676 , \22639 );
nor \U$41036 ( \41351 , \41349 , \41350 );
xnor \U$41037 ( \41352 , \41351 , \22651 );
xor \U$41038 ( \41353 , \41348 , \41352 );
xor \U$41039 ( \41354 , \41339 , \41353 );
xor \U$41040 ( \41355 , \41332 , \41354 );
and \U$41041 ( \41356 , \41078 , \41082 );
and \U$41042 ( \41357 , \41082 , \41087 );
and \U$41043 ( \41358 , \41078 , \41087 );
or \U$41044 ( \41359 , \41356 , \41357 , \41358 );
and \U$41045 ( \41360 , \41063 , \41067 );
and \U$41046 ( \41361 , \41067 , \41072 );
and \U$41047 ( \41362 , \41063 , \41072 );
or \U$41048 ( \41363 , \41360 , \41361 , \41362 );
xor \U$41049 ( \41364 , \41359 , \41363 );
and \U$41050 ( \41365 , \41049 , \41053 );
and \U$41051 ( \41366 , \41053 , \41058 );
and \U$41052 ( \41367 , \41049 , \41058 );
or \U$41053 ( \41368 , \41365 , \41366 , \41367 );
xor \U$41054 ( \41369 , \41364 , \41368 );
xor \U$41055 ( \41370 , \41355 , \41369 );
xor \U$41056 ( \41371 , \41288 , \41370 );
xor \U$41057 ( \41372 , \41254 , \41371 );
and \U$41058 ( \41373 , \40896 , \40900 );
and \U$41059 ( \41374 , \40900 , \40905 );
and \U$41060 ( \41375 , \40896 , \40905 );
or \U$41061 ( \41376 , \41373 , \41374 , \41375 );
and \U$41062 ( \41377 , \40882 , \40886 );
and \U$41063 ( \41378 , \40886 , \40891 );
and \U$41064 ( \41379 , \40882 , \40891 );
or \U$41065 ( \41380 , \41377 , \41378 , \41379 );
xor \U$41066 ( \41381 , \41376 , \41380 );
and \U$41067 ( \41382 , \41000 , \41044 );
and \U$41068 ( \41383 , \41044 , \41089 );
and \U$41069 ( \41384 , \41000 , \41089 );
or \U$41070 ( \41385 , \41382 , \41383 , \41384 );
xor \U$41071 ( \41386 , \41381 , \41385 );
xor \U$41072 ( \41387 , \41372 , \41386 );
xor \U$41073 ( \41388 , \41154 , \41387 );
xor \U$41074 ( \41389 , \41145 , \41388 );
and \U$41075 ( \41390 , \40872 , \40873 );
and \U$41076 ( \41391 , \40873 , \41123 );
and \U$41077 ( \41392 , \40872 , \41123 );
or \U$41078 ( \41393 , \41390 , \41391 , \41392 );
nor \U$41079 ( \41394 , \41389 , \41393 );
nor \U$41080 ( \41395 , \41129 , \41394 );
nand \U$41081 ( \41396 , \40868 , \41395 );
nor \U$41082 ( \41397 , \40361 , \41396 );
and \U$41083 ( \41398 , \41149 , \41153 );
and \U$41084 ( \41399 , \41153 , \41387 );
and \U$41085 ( \41400 , \41149 , \41387 );
or \U$41086 ( \41401 , \41398 , \41399 , \41400 );
and \U$41087 ( \41402 , \41276 , \41280 );
and \U$41088 ( \41403 , \41280 , \41285 );
and \U$41089 ( \41404 , \41276 , \41285 );
or \U$41090 ( \41405 , \41402 , \41403 , \41404 );
and \U$41091 ( \41406 , \41262 , \41266 );
and \U$41092 ( \41407 , \41266 , \41271 );
and \U$41093 ( \41408 , \41262 , \41271 );
or \U$41094 ( \41409 , \41406 , \41407 , \41408 );
xor \U$41095 ( \41410 , \41405 , \41409 );
and \U$41096 ( \41411 , \41359 , \41363 );
and \U$41097 ( \41412 , \41363 , \41368 );
and \U$41098 ( \41413 , \41359 , \41368 );
or \U$41099 ( \41414 , \41411 , \41412 , \41413 );
xor \U$41100 ( \41415 , \41410 , \41414 );
and \U$41101 ( \41416 , \22706 , \22691 );
and \U$41102 ( \41417 , \22686 , \22689 );
nor \U$41103 ( \41418 , \41416 , \41417 );
xnor \U$41104 ( \41419 , \41418 , \22701 );
xor \U$41105 ( \41420 , \24598 , \24602 );
xor \U$41106 ( \41421 , \41420 , \24607 );
xor \U$41107 ( \41422 , \41419 , \41421 );
xor \U$41108 ( \41423 , \24581 , \24585 );
xor \U$41109 ( \41424 , \41423 , \24590 );
xor \U$41110 ( \41425 , \41422 , \41424 );
and \U$41111 ( \41426 , \41306 , \41310 );
and \U$41112 ( \41427 , \41310 , \41315 );
and \U$41113 ( \41428 , \41306 , \41315 );
or \U$41114 ( \41429 , \41426 , \41427 , \41428 );
and \U$41115 ( \41430 , \41292 , \41296 );
and \U$41116 ( \41431 , \41296 , \41301 );
and \U$41117 ( \41432 , \41292 , \41301 );
or \U$41118 ( \41433 , \41430 , \41431 , \41432 );
xor \U$41119 ( \41434 , \41429 , \41433 );
and \U$41120 ( \41435 , \41343 , \41347 );
and \U$41121 ( \41436 , \41347 , \41352 );
and \U$41122 ( \41437 , \41343 , \41352 );
or \U$41123 ( \41438 , \41435 , \41436 , \41437 );
xor \U$41124 ( \41439 , \41434 , \41438 );
xor \U$41125 ( \41440 , \41425 , \41439 );
and \U$41126 ( \41441 , \41197 , \41201 );
and \U$41127 ( \41442 , \41201 , \41206 );
and \U$41128 ( \41443 , \41197 , \41206 );
or \U$41129 ( \41444 , \41441 , \41442 , \41443 );
and \U$41130 ( \41445 , \41183 , \41187 );
and \U$41131 ( \41446 , \41187 , \41192 );
and \U$41132 ( \41447 , \41183 , \41192 );
or \U$41133 ( \41448 , \41445 , \41446 , \41447 );
xor \U$41134 ( \41449 , \41444 , \41448 );
and \U$41135 ( \41450 , \41321 , \41325 );
and \U$41136 ( \41451 , \41325 , \41330 );
and \U$41137 ( \41452 , \41321 , \41330 );
or \U$41138 ( \41453 , \41450 , \41451 , \41452 );
xor \U$41139 ( \41454 , \41449 , \41453 );
xor \U$41140 ( \41455 , \41440 , \41454 );
xor \U$41141 ( \41456 , \24460 , \24464 );
xor \U$41142 ( \41457 , \41456 , \24469 );
xor \U$41143 ( \41458 , \24512 , \24516 );
xor \U$41144 ( \41459 , \41458 , \24521 );
xor \U$41145 ( \41460 , \24493 , \24497 );
xor \U$41146 ( \41461 , \41460 , \24502 );
xor \U$41147 ( \41462 , \41459 , \41461 );
xor \U$41148 ( \41463 , \24476 , \24480 );
xor \U$41149 ( \41464 , \41463 , \24485 );
xor \U$41150 ( \41465 , \41462 , \41464 );
xor \U$41151 ( \41466 , \41457 , \41465 );
xor \U$41152 ( \41467 , \24565 , \24569 );
xor \U$41153 ( \41468 , \41467 , \24574 );
xor \U$41154 ( \41469 , \24545 , \24549 );
xor \U$41155 ( \41470 , \41469 , \24554 );
xor \U$41156 ( \41471 , \41468 , \41470 );
xor \U$41157 ( \41472 , \24528 , \24532 );
xor \U$41158 ( \41473 , \41472 , \24537 );
xor \U$41159 ( \41474 , \41471 , \41473 );
xor \U$41160 ( \41475 , \41466 , \41474 );
xor \U$41161 ( \41476 , \41455 , \41475 );
and \U$41162 ( \41477 , \41336 , \41338 );
and \U$41163 ( \41478 , \41338 , \41353 );
and \U$41164 ( \41479 , \41336 , \41353 );
or \U$41165 ( \41480 , \41477 , \41478 , \41479 );
and \U$41166 ( \41481 , \41302 , \41316 );
and \U$41167 ( \41482 , \41316 , \41331 );
and \U$41168 ( \41483 , \41302 , \41331 );
or \U$41169 ( \41484 , \41481 , \41482 , \41483 );
xor \U$41170 ( \41485 , \41480 , \41484 );
and \U$41171 ( \41486 , \41193 , \41207 );
and \U$41172 ( \41487 , \41207 , \41222 );
and \U$41173 ( \41488 , \41193 , \41222 );
or \U$41174 ( \41489 , \41486 , \41487 , \41488 );
xor \U$41175 ( \41490 , \41485 , \41489 );
xor \U$41176 ( \41491 , \41476 , \41490 );
xor \U$41177 ( \41492 , \41415 , \41491 );
and \U$41178 ( \41493 , \41332 , \41354 );
and \U$41179 ( \41494 , \41354 , \41369 );
and \U$41180 ( \41495 , \41332 , \41369 );
or \U$41181 ( \41496 , \41493 , \41494 , \41495 );
and \U$41182 ( \41497 , \41272 , \41286 );
xor \U$41183 ( \41498 , \41496 , \41497 );
and \U$41184 ( \41499 , \22701 , \41172 );
and \U$41185 ( \41500 , \41172 , \41177 );
and \U$41186 ( \41501 , \22701 , \41177 );
or \U$41187 ( \41502 , \41499 , \41500 , \41501 );
and \U$41188 ( \41503 , \41158 , \41162 );
and \U$41189 ( \41504 , \41162 , \41167 );
and \U$41190 ( \41505 , \41158 , \41167 );
or \U$41191 ( \41506 , \41503 , \41504 , \41505 );
xor \U$41192 ( \41507 , \41502 , \41506 );
and \U$41193 ( \41508 , \41212 , \41216 );
and \U$41194 ( \41509 , \41216 , \41221 );
and \U$41195 ( \41510 , \41212 , \41221 );
or \U$41196 ( \41511 , \41508 , \41509 , \41510 );
xor \U$41197 ( \41512 , \41507 , \41511 );
xor \U$41198 ( \41513 , \41498 , \41512 );
xor \U$41199 ( \41514 , \41492 , \41513 );
and \U$41200 ( \41515 , \41376 , \41380 );
and \U$41201 ( \41516 , \41380 , \41385 );
and \U$41202 ( \41517 , \41376 , \41385 );
or \U$41203 ( \41518 , \41515 , \41516 , \41517 );
and \U$41204 ( \41519 , \41258 , \41287 );
and \U$41205 ( \41520 , \41287 , \41370 );
and \U$41206 ( \41521 , \41258 , \41370 );
or \U$41207 ( \41522 , \41519 , \41520 , \41521 );
xor \U$41208 ( \41523 , \41518 , \41522 );
and \U$41209 ( \41524 , \41224 , \41238 );
and \U$41210 ( \41525 , \41238 , \41253 );
and \U$41211 ( \41526 , \41224 , \41253 );
or \U$41212 ( \41527 , \41524 , \41525 , \41526 );
xor \U$41213 ( \41528 , \41523 , \41527 );
xor \U$41214 ( \41529 , \41514 , \41528 );
xor \U$41215 ( \41530 , \41401 , \41529 );
and \U$41216 ( \41531 , \41137 , \41141 );
and \U$41217 ( \41532 , \41141 , \41143 );
and \U$41218 ( \41533 , \41137 , \41143 );
or \U$41219 ( \41534 , \41531 , \41532 , \41533 );
and \U$41220 ( \41535 , \41254 , \41371 );
and \U$41221 ( \41536 , \41371 , \41386 );
and \U$41222 ( \41537 , \41254 , \41386 );
or \U$41223 ( \41538 , \41535 , \41536 , \41537 );
xor \U$41224 ( \41539 , \41534 , \41538 );
and \U$41225 ( \41540 , \41243 , \41247 );
and \U$41226 ( \41541 , \41247 , \41252 );
and \U$41227 ( \41542 , \41243 , \41252 );
or \U$41228 ( \41543 , \41540 , \41541 , \41542 );
and \U$41229 ( \41544 , \41228 , \41232 );
and \U$41230 ( \41545 , \41232 , \41237 );
and \U$41231 ( \41546 , \41228 , \41237 );
or \U$41232 ( \41547 , \41544 , \41545 , \41546 );
xor \U$41233 ( \41548 , \41543 , \41547 );
and \U$41234 ( \41549 , \41168 , \41178 );
and \U$41235 ( \41550 , \41178 , \41223 );
and \U$41236 ( \41551 , \41168 , \41223 );
or \U$41237 ( \41552 , \41549 , \41550 , \41551 );
xor \U$41238 ( \41553 , \41548 , \41552 );
xor \U$41239 ( \41554 , \41539 , \41553 );
xor \U$41240 ( \41555 , \41530 , \41554 );
and \U$41241 ( \41556 , \41133 , \41144 );
and \U$41242 ( \41557 , \41144 , \41388 );
and \U$41243 ( \41558 , \41133 , \41388 );
or \U$41244 ( \41559 , \41556 , \41557 , \41558 );
nor \U$41245 ( \41560 , \41555 , \41559 );
and \U$41246 ( \41561 , \41518 , \41522 );
and \U$41247 ( \41562 , \41522 , \41527 );
and \U$41248 ( \41563 , \41518 , \41527 );
or \U$41249 ( \41564 , \41561 , \41562 , \41563 );
and \U$41250 ( \41565 , \41415 , \41491 );
and \U$41251 ( \41566 , \41491 , \41513 );
and \U$41252 ( \41567 , \41415 , \41513 );
or \U$41253 ( \41568 , \41565 , \41566 , \41567 );
xor \U$41254 ( \41569 , \41564 , \41568 );
xor \U$41255 ( \41570 , \22067 , \22084 );
xor \U$41256 ( \41571 , \41570 , \22106 );
xor \U$41257 ( \41572 , \24639 , \24641 );
xor \U$41258 ( \41573 , \41572 , \24644 );
xor \U$41259 ( \41574 , \41571 , \41573 );
xor \U$41260 ( \41575 , \24628 , \24630 );
xor \U$41261 ( \41576 , \41575 , \24633 );
xor \U$41262 ( \41577 , \41574 , \41576 );
and \U$41263 ( \41578 , \41419 , \41421 );
and \U$41264 ( \41579 , \41421 , \41424 );
and \U$41265 ( \41580 , \41419 , \41424 );
or \U$41266 ( \41581 , \41578 , \41579 , \41580 );
and \U$41267 ( \41582 , \41468 , \41470 );
and \U$41268 ( \41583 , \41470 , \41473 );
and \U$41269 ( \41584 , \41468 , \41473 );
or \U$41270 ( \41585 , \41582 , \41583 , \41584 );
xor \U$41271 ( \41586 , \41581 , \41585 );
and \U$41272 ( \41587 , \41459 , \41461 );
and \U$41273 ( \41588 , \41461 , \41464 );
and \U$41274 ( \41589 , \41459 , \41464 );
or \U$41275 ( \41590 , \41587 , \41588 , \41589 );
xor \U$41276 ( \41591 , \41586 , \41590 );
xor \U$41277 ( \41592 , \41577 , \41591 );
and \U$41278 ( \41593 , \41502 , \41506 );
and \U$41279 ( \41594 , \41506 , \41511 );
and \U$41280 ( \41595 , \41502 , \41511 );
or \U$41281 ( \41596 , \41593 , \41594 , \41595 );
and \U$41282 ( \41597 , \41444 , \41448 );
and \U$41283 ( \41598 , \41448 , \41453 );
and \U$41284 ( \41599 , \41444 , \41453 );
or \U$41285 ( \41600 , \41597 , \41598 , \41599 );
xor \U$41286 ( \41601 , \41596 , \41600 );
and \U$41287 ( \41602 , \41429 , \41433 );
and \U$41288 ( \41603 , \41433 , \41438 );
and \U$41289 ( \41604 , \41429 , \41438 );
or \U$41290 ( \41605 , \41602 , \41603 , \41604 );
xor \U$41291 ( \41606 , \41601 , \41605 );
xor \U$41292 ( \41607 , \41592 , \41606 );
and \U$41293 ( \41608 , \41425 , \41439 );
and \U$41294 ( \41609 , \41439 , \41454 );
and \U$41295 ( \41610 , \41425 , \41454 );
or \U$41296 ( \41611 , \41608 , \41609 , \41610 );
xor \U$41297 ( \41612 , \24472 , \24488 );
xor \U$41298 ( \41613 , \41612 , \24505 );
xor \U$41299 ( \41614 , \41611 , \41613 );
xor \U$41300 ( \41615 , \24618 , \24620 );
xor \U$41301 ( \41616 , \41615 , \24623 );
xor \U$41302 ( \41617 , \24577 , \24593 );
xor \U$41303 ( \41618 , \41617 , \24610 );
xor \U$41304 ( \41619 , \41616 , \41618 );
xor \U$41305 ( \41620 , \24524 , \24540 );
xor \U$41306 ( \41621 , \41620 , \24557 );
xor \U$41307 ( \41622 , \41619 , \41621 );
xor \U$41308 ( \41623 , \41614 , \41622 );
xor \U$41309 ( \41624 , \41607 , \41623 );
and \U$41310 ( \41625 , \41405 , \41409 );
and \U$41311 ( \41626 , \41409 , \41414 );
and \U$41312 ( \41627 , \41405 , \41414 );
or \U$41313 ( \41628 , \41625 , \41626 , \41627 );
and \U$41314 ( \41629 , \41480 , \41484 );
and \U$41315 ( \41630 , \41484 , \41489 );
and \U$41316 ( \41631 , \41480 , \41489 );
or \U$41317 ( \41632 , \41629 , \41630 , \41631 );
xor \U$41318 ( \41633 , \41628 , \41632 );
and \U$41319 ( \41634 , \41457 , \41465 );
and \U$41320 ( \41635 , \41465 , \41474 );
and \U$41321 ( \41636 , \41457 , \41474 );
or \U$41322 ( \41637 , \41634 , \41635 , \41636 );
xor \U$41323 ( \41638 , \41633 , \41637 );
xor \U$41324 ( \41639 , \41624 , \41638 );
xor \U$41325 ( \41640 , \41569 , \41639 );
and \U$41326 ( \41641 , \41534 , \41538 );
and \U$41327 ( \41642 , \41538 , \41553 );
and \U$41328 ( \41643 , \41534 , \41553 );
or \U$41329 ( \41644 , \41641 , \41642 , \41643 );
and \U$41330 ( \41645 , \41514 , \41528 );
xor \U$41331 ( \41646 , \41644 , \41645 );
and \U$41332 ( \41647 , \41543 , \41547 );
and \U$41333 ( \41648 , \41547 , \41552 );
and \U$41334 ( \41649 , \41543 , \41552 );
or \U$41335 ( \41650 , \41647 , \41648 , \41649 );
and \U$41336 ( \41651 , \41496 , \41497 );
and \U$41337 ( \41652 , \41497 , \41512 );
and \U$41338 ( \41653 , \41496 , \41512 );
or \U$41339 ( \41654 , \41651 , \41652 , \41653 );
xor \U$41340 ( \41655 , \41650 , \41654 );
and \U$41341 ( \41656 , \41455 , \41475 );
and \U$41342 ( \41657 , \41475 , \41490 );
and \U$41343 ( \41658 , \41455 , \41490 );
or \U$41344 ( \41659 , \41656 , \41657 , \41658 );
xor \U$41345 ( \41660 , \41655 , \41659 );
xor \U$41346 ( \41661 , \41646 , \41660 );
xor \U$41347 ( \41662 , \41640 , \41661 );
and \U$41348 ( \41663 , \41401 , \41529 );
and \U$41349 ( \41664 , \41529 , \41554 );
and \U$41350 ( \41665 , \41401 , \41554 );
or \U$41351 ( \41666 , \41663 , \41664 , \41665 );
nor \U$41352 ( \41667 , \41662 , \41666 );
nor \U$41353 ( \41668 , \41560 , \41667 );
and \U$41354 ( \41669 , \41644 , \41645 );
and \U$41355 ( \41670 , \41645 , \41660 );
and \U$41356 ( \41671 , \41644 , \41660 );
or \U$41357 ( \41672 , \41669 , \41670 , \41671 );
and \U$41358 ( \41673 , \41564 , \41568 );
and \U$41359 ( \41674 , \41568 , \41639 );
and \U$41360 ( \41675 , \41564 , \41639 );
or \U$41361 ( \41676 , \41673 , \41674 , \41675 );
and \U$41362 ( \41677 , \41628 , \41632 );
and \U$41363 ( \41678 , \41632 , \41637 );
and \U$41364 ( \41679 , \41628 , \41637 );
or \U$41365 ( \41680 , \41677 , \41678 , \41679 );
and \U$41366 ( \41681 , \41611 , \41613 );
and \U$41367 ( \41682 , \41613 , \41622 );
and \U$41368 ( \41683 , \41611 , \41622 );
or \U$41369 ( \41684 , \41681 , \41682 , \41683 );
xor \U$41370 ( \41685 , \41680 , \41684 );
and \U$41371 ( \41686 , \41577 , \41591 );
and \U$41372 ( \41687 , \41591 , \41606 );
and \U$41373 ( \41688 , \41577 , \41606 );
or \U$41374 ( \41689 , \41686 , \41687 , \41688 );
xor \U$41375 ( \41690 , \41685 , \41689 );
xor \U$41376 ( \41691 , \41676 , \41690 );
and \U$41377 ( \41692 , \41650 , \41654 );
and \U$41378 ( \41693 , \41654 , \41659 );
and \U$41379 ( \41694 , \41650 , \41659 );
or \U$41380 ( \41695 , \41692 , \41693 , \41694 );
and \U$41381 ( \41696 , \41607 , \41623 );
and \U$41382 ( \41697 , \41623 , \41638 );
and \U$41383 ( \41698 , \41607 , \41638 );
or \U$41384 ( \41699 , \41696 , \41697 , \41698 );
xor \U$41385 ( \41700 , \41695 , \41699 );
xor \U$41386 ( \41701 , \24653 , \24655 );
xor \U$41387 ( \41702 , \41701 , \24658 );
xor \U$41388 ( \41703 , \24626 , \24636 );
xor \U$41389 ( \41704 , \41703 , \24647 );
xor \U$41390 ( \41705 , \41702 , \41704 );
xor \U$41391 ( \41706 , \24508 , \24560 );
xor \U$41392 ( \41707 , \41706 , \24613 );
xor \U$41393 ( \41708 , \41705 , \41707 );
and \U$41394 ( \41709 , \41616 , \41618 );
and \U$41395 ( \41710 , \41618 , \41621 );
and \U$41396 ( \41711 , \41616 , \41621 );
or \U$41397 ( \41712 , \41709 , \41710 , \41711 );
xor \U$41398 ( \41713 , \22109 , \22176 );
xor \U$41399 ( \41714 , \41713 , \22244 );
xor \U$41400 ( \41715 , \41712 , \41714 );
xor \U$41401 ( \41716 , \24666 , \24668 );
xor \U$41402 ( \41717 , \41716 , \24671 );
xor \U$41403 ( \41718 , \41715 , \41717 );
xor \U$41404 ( \41719 , \41708 , \41718 );
and \U$41405 ( \41720 , \41596 , \41600 );
and \U$41406 ( \41721 , \41600 , \41605 );
and \U$41407 ( \41722 , \41596 , \41605 );
or \U$41408 ( \41723 , \41720 , \41721 , \41722 );
and \U$41409 ( \41724 , \41581 , \41585 );
and \U$41410 ( \41725 , \41585 , \41590 );
and \U$41411 ( \41726 , \41581 , \41590 );
or \U$41412 ( \41727 , \41724 , \41725 , \41726 );
xor \U$41413 ( \41728 , \41723 , \41727 );
and \U$41414 ( \41729 , \41571 , \41573 );
and \U$41415 ( \41730 , \41573 , \41576 );
and \U$41416 ( \41731 , \41571 , \41576 );
or \U$41417 ( \41732 , \41729 , \41730 , \41731 );
xor \U$41418 ( \41733 , \41728 , \41732 );
xor \U$41419 ( \41734 , \41719 , \41733 );
xor \U$41420 ( \41735 , \41700 , \41734 );
xor \U$41421 ( \41736 , \41691 , \41735 );
xor \U$41422 ( \41737 , \41672 , \41736 );
and \U$41423 ( \41738 , \41640 , \41661 );
nor \U$41424 ( \41739 , \41737 , \41738 );
and \U$41425 ( \41740 , \41676 , \41690 );
and \U$41426 ( \41741 , \41690 , \41735 );
and \U$41427 ( \41742 , \41676 , \41735 );
or \U$41428 ( \41743 , \41740 , \41741 , \41742 );
and \U$41429 ( \41744 , \41695 , \41699 );
and \U$41430 ( \41745 , \41699 , \41734 );
and \U$41431 ( \41746 , \41695 , \41734 );
or \U$41432 ( \41747 , \41744 , \41745 , \41746 );
and \U$41433 ( \41748 , \41723 , \41727 );
and \U$41434 ( \41749 , \41727 , \41732 );
and \U$41435 ( \41750 , \41723 , \41732 );
or \U$41436 ( \41751 , \41748 , \41749 , \41750 );
and \U$41437 ( \41752 , \41712 , \41714 );
and \U$41438 ( \41753 , \41714 , \41717 );
and \U$41439 ( \41754 , \41712 , \41717 );
or \U$41440 ( \41755 , \41752 , \41753 , \41754 );
xor \U$41441 ( \41756 , \41751 , \41755 );
and \U$41442 ( \41757 , \41702 , \41704 );
and \U$41443 ( \41758 , \41704 , \41707 );
and \U$41444 ( \41759 , \41702 , \41707 );
or \U$41445 ( \41760 , \41757 , \41758 , \41759 );
xor \U$41446 ( \41761 , \41756 , \41760 );
xor \U$41447 ( \41762 , \41747 , \41761 );
and \U$41448 ( \41763 , \41680 , \41684 );
and \U$41449 ( \41764 , \41684 , \41689 );
and \U$41450 ( \41765 , \41680 , \41689 );
or \U$41451 ( \41766 , \41763 , \41764 , \41765 );
and \U$41452 ( \41767 , \41708 , \41718 );
and \U$41453 ( \41768 , \41718 , \41733 );
and \U$41454 ( \41769 , \41708 , \41733 );
or \U$41455 ( \41770 , \41767 , \41768 , \41769 );
xor \U$41456 ( \41771 , \41766 , \41770 );
xor \U$41457 ( \41772 , \24685 , \24687 );
xor \U$41458 ( \41773 , \41772 , \24690 );
xor \U$41459 ( \41774 , \24674 , \24676 );
xor \U$41460 ( \41775 , \41774 , \24679 );
xor \U$41461 ( \41776 , \41773 , \41775 );
xor \U$41462 ( \41777 , \24616 , \24650 );
xor \U$41463 ( \41778 , \41777 , \24661 );
xor \U$41464 ( \41779 , \41776 , \41778 );
xor \U$41465 ( \41780 , \41771 , \41779 );
xor \U$41466 ( \41781 , \41762 , \41780 );
xor \U$41467 ( \41782 , \41743 , \41781 );
and \U$41468 ( \41783 , \41672 , \41736 );
nor \U$41469 ( \41784 , \41782 , \41783 );
nor \U$41470 ( \41785 , \41739 , \41784 );
nand \U$41471 ( \41786 , \41668 , \41785 );
and \U$41472 ( \41787 , \41747 , \41761 );
and \U$41473 ( \41788 , \41761 , \41780 );
and \U$41474 ( \41789 , \41747 , \41780 );
or \U$41475 ( \41790 , \41787 , \41788 , \41789 );
and \U$41476 ( \41791 , \41766 , \41770 );
and \U$41477 ( \41792 , \41770 , \41779 );
and \U$41478 ( \41793 , \41766 , \41779 );
or \U$41479 ( \41794 , \41791 , \41792 , \41793 );
xor \U$41480 ( \41795 , \22661 , \22823 );
xor \U$41481 ( \41796 , \41795 , \22906 );
xor \U$41482 ( \41797 , \24698 , \24700 );
xor \U$41483 ( \41798 , \41797 , \24703 );
xor \U$41484 ( \41799 , \41796 , \41798 );
xor \U$41485 ( \41800 , \24664 , \24682 );
xor \U$41486 ( \41801 , \41800 , \24693 );
xor \U$41487 ( \41802 , \41799 , \41801 );
xor \U$41488 ( \41803 , \41794 , \41802 );
and \U$41489 ( \41804 , \41751 , \41755 );
and \U$41490 ( \41805 , \41755 , \41760 );
and \U$41491 ( \41806 , \41751 , \41760 );
or \U$41492 ( \41807 , \41804 , \41805 , \41806 );
and \U$41493 ( \41808 , \41773 , \41775 );
and \U$41494 ( \41809 , \41775 , \41778 );
and \U$41495 ( \41810 , \41773 , \41778 );
or \U$41496 ( \41811 , \41808 , \41809 , \41810 );
xor \U$41497 ( \41812 , \41807 , \41811 );
xor \U$41498 ( \41813 , \23034 , \23080 );
xor \U$41499 ( \41814 , \41813 , \23095 );
xor \U$41500 ( \41815 , \41812 , \41814 );
xor \U$41501 ( \41816 , \41803 , \41815 );
xor \U$41502 ( \41817 , \41790 , \41816 );
and \U$41503 ( \41818 , \41743 , \41781 );
nor \U$41504 ( \41819 , \41817 , \41818 );
and \U$41505 ( \41820 , \41794 , \41802 );
and \U$41506 ( \41821 , \41802 , \41815 );
and \U$41507 ( \41822 , \41794 , \41815 );
or \U$41508 ( \41823 , \41820 , \41821 , \41822 );
xor \U$41509 ( \41824 , \24696 , \24706 );
xor \U$41510 ( \41825 , \41824 , \24709 );
xor \U$41511 ( \41826 , \41823 , \41825 );
and \U$41512 ( \41827 , \41807 , \41811 );
and \U$41513 ( \41828 , \41811 , \41814 );
and \U$41514 ( \41829 , \41807 , \41814 );
or \U$41515 ( \41830 , \41827 , \41828 , \41829 );
and \U$41516 ( \41831 , \41796 , \41798 );
and \U$41517 ( \41832 , \41798 , \41801 );
and \U$41518 ( \41833 , \41796 , \41801 );
or \U$41519 ( \41834 , \41831 , \41832 , \41833 );
xor \U$41520 ( \41835 , \41830 , \41834 );
xor \U$41521 ( \41836 , \22909 , \23098 );
xor \U$41522 ( \41837 , \41836 , \23292 );
xor \U$41523 ( \41838 , \41835 , \41837 );
xor \U$41524 ( \41839 , \41826 , \41838 );
and \U$41525 ( \41840 , \41790 , \41816 );
nor \U$41526 ( \41841 , \41839 , \41840 );
nor \U$41527 ( \41842 , \41819 , \41841 );
and \U$41528 ( \41843 , \41830 , \41834 );
and \U$41529 ( \41844 , \41834 , \41837 );
and \U$41530 ( \41845 , \41830 , \41837 );
or \U$41531 ( \41846 , \41843 , \41844 , \41845 );
xor \U$41532 ( \41847 , \24712 , \24714 );
xor \U$41533 ( \41848 , \41847 , \24717 );
xor \U$41534 ( \41849 , \41846 , \41848 );
and \U$41535 ( \41850 , \41823 , \41825 );
and \U$41536 ( \41851 , \41825 , \41838 );
and \U$41537 ( \41852 , \41823 , \41838 );
or \U$41538 ( \41853 , \41850 , \41851 , \41852 );
nor \U$41539 ( \41854 , \41849 , \41853 );
xor \U$41540 ( \41855 , \24720 , \24722 );
and \U$41541 ( \41856 , \41846 , \41848 );
nor \U$41542 ( \41857 , \41855 , \41856 );
nor \U$41543 ( \41858 , \41854 , \41857 );
nand \U$41544 ( \41859 , \41842 , \41858 );
nor \U$41545 ( \41860 , \41786 , \41859 );
nand \U$41546 ( \41861 , \41397 , \41860 );
nor \U$41547 ( \41862 , \39406 , \41861 );
and \U$41548 ( \41863 , \22567 , \22076 );
and \U$41549 ( \41864 , \22578 , \22073 );
nor \U$41550 ( \41865 , \41863 , \41864 );
xnor \U$41551 ( \41866 , \41865 , \22072 );
and \U$41552 ( \41867 , \22218 , \41866 );
and \U$41553 ( \41868 , \22592 , \22095 );
and \U$41554 ( \41869 , \22603 , \22093 );
nor \U$41555 ( \41870 , \41868 , \41869 );
xnor \U$41556 ( \41871 , \41870 , \22105 );
and \U$41557 ( \41872 , \41866 , \41871 );
and \U$41558 ( \41873 , \22218 , \41871 );
or \U$41559 ( \41874 , \41867 , \41872 , \41873 );
and \U$41560 ( \41875 , \22613 , \22119 );
and \U$41561 ( \41876 , \22624 , \22117 );
nor \U$41562 ( \41877 , \41875 , \41876 );
xnor \U$41563 ( \41878 , \41877 , \22129 );
and \U$41564 ( \41879 , \22635 , \22140 );
and \U$41565 ( \41880 , \22646 , \22138 );
nor \U$41566 ( \41881 , \41879 , \41880 );
xnor \U$41567 ( \41882 , \41881 , \22150 );
and \U$41568 ( \41883 , \41878 , \41882 );
and \U$41569 ( \41884 , \22665 , \22162 );
and \U$41570 ( \41885 , \22676 , \22160 );
nor \U$41571 ( \41886 , \41884 , \41885 );
xnor \U$41572 ( \41887 , \41886 , \22172 );
and \U$41573 ( \41888 , \41882 , \41887 );
and \U$41574 ( \41889 , \41878 , \41887 );
or \U$41575 ( \41890 , \41883 , \41888 , \41889 );
and \U$41576 ( \41891 , \41874 , \41890 );
and \U$41577 ( \41892 , \22706 , \22208 );
and \U$41578 ( \41893 , \22686 , \22206 );
nor \U$41579 ( \41894 , \41892 , \41893 );
xnor \U$41580 ( \41895 , \41894 , \22218 );
and \U$41581 ( \41896 , \41890 , \41895 );
and \U$41582 ( \41897 , \41874 , \41895 );
or \U$41583 ( \41898 , \41891 , \41896 , \41897 );
and \U$41584 ( \41899 , \22592 , \22119 );
and \U$41585 ( \41900 , \22603 , \22117 );
nor \U$41586 ( \41901 , \41899 , \41900 );
xnor \U$41587 ( \41902 , \41901 , \22129 );
and \U$41588 ( \41903 , \22613 , \22140 );
and \U$41589 ( \41904 , \22624 , \22138 );
nor \U$41590 ( \41905 , \41903 , \41904 );
xnor \U$41591 ( \41906 , \41905 , \22150 );
xor \U$41592 ( \41907 , \41902 , \41906 );
and \U$41593 ( \41908 , \22635 , \22162 );
and \U$41594 ( \41909 , \22646 , \22160 );
nor \U$41595 ( \41910 , \41908 , \41909 );
xnor \U$41596 ( \41911 , \41910 , \22172 );
xor \U$41597 ( \41912 , \41907 , \41911 );
and \U$41598 ( \41913 , \22545 , \22076 );
and \U$41599 ( \41914 , \22556 , \22073 );
nor \U$41600 ( \41915 , \41913 , \41914 );
xnor \U$41601 ( \41916 , \41915 , \22072 );
xor \U$41602 ( \41917 , \22240 , \41916 );
and \U$41603 ( \41918 , \22567 , \22095 );
and \U$41604 ( \41919 , \22578 , \22093 );
nor \U$41605 ( \41920 , \41918 , \41919 );
xnor \U$41606 ( \41921 , \41920 , \22105 );
xor \U$41607 ( \41922 , \41917 , \41921 );
xor \U$41608 ( \41923 , \41912 , \41922 );
and \U$41609 ( \41924 , \41898 , \41923 );
and \U$41610 ( \41925 , \22578 , \22076 );
and \U$41611 ( \41926 , \22545 , \22073 );
nor \U$41612 ( \41927 , \41925 , \41926 );
xnor \U$41613 ( \41928 , \41927 , \22072 );
and \U$41614 ( \41929 , \22603 , \22095 );
and \U$41615 ( \41930 , \22567 , \22093 );
nor \U$41616 ( \41931 , \41929 , \41930 );
xnor \U$41617 ( \41932 , \41931 , \22105 );
and \U$41618 ( \41933 , \41928 , \41932 );
and \U$41619 ( \41934 , \22624 , \22119 );
and \U$41620 ( \41935 , \22592 , \22117 );
nor \U$41621 ( \41936 , \41934 , \41935 );
xnor \U$41622 ( \41937 , \41936 , \22129 );
and \U$41623 ( \41938 , \41932 , \41937 );
and \U$41624 ( \41939 , \41928 , \41937 );
or \U$41625 ( \41940 , \41933 , \41938 , \41939 );
and \U$41626 ( \41941 , \22646 , \22140 );
and \U$41627 ( \41942 , \22613 , \22138 );
nor \U$41628 ( \41943 , \41941 , \41942 );
xnor \U$41629 ( \41944 , \41943 , \22150 );
and \U$41630 ( \41945 , \22676 , \22162 );
and \U$41631 ( \41946 , \22635 , \22160 );
nor \U$41632 ( \41947 , \41945 , \41946 );
xnor \U$41633 ( \41948 , \41947 , \22172 );
and \U$41634 ( \41949 , \41944 , \41948 );
and \U$41635 ( \41950 , \22696 , \22187 );
and \U$41636 ( \41951 , \22665 , \22185 );
nor \U$41637 ( \41952 , \41950 , \41951 );
xnor \U$41638 ( \41953 , \41952 , \22197 );
and \U$41639 ( \41954 , \41948 , \41953 );
and \U$41640 ( \41955 , \41944 , \41953 );
or \U$41641 ( \41956 , \41949 , \41954 , \41955 );
xor \U$41642 ( \41957 , \41940 , \41956 );
and \U$41643 ( \41958 , \22665 , \22187 );
and \U$41644 ( \41959 , \22676 , \22185 );
nor \U$41645 ( \41960 , \41958 , \41959 );
xnor \U$41646 ( \41961 , \41960 , \22197 );
and \U$41647 ( \41962 , \22686 , \22208 );
and \U$41648 ( \41963 , \22696 , \22206 );
nor \U$41649 ( \41964 , \41962 , \41963 );
xnor \U$41650 ( \41965 , \41964 , \22218 );
xor \U$41651 ( \41966 , \41961 , \41965 );
nand \U$41652 ( \41967 , \22706 , \22228 );
xnor \U$41653 ( \41968 , \41967 , \22240 );
xor \U$41654 ( \41969 , \41966 , \41968 );
xor \U$41655 ( \41970 , \41957 , \41969 );
and \U$41656 ( \41971 , \41923 , \41970 );
and \U$41657 ( \41972 , \41898 , \41970 );
or \U$41658 ( \41973 , \41924 , \41971 , \41972 );
and \U$41659 ( \41974 , \22240 , \41916 );
and \U$41660 ( \41975 , \41916 , \41921 );
and \U$41661 ( \41976 , \22240 , \41921 );
or \U$41662 ( \41977 , \41974 , \41975 , \41976 );
and \U$41663 ( \41978 , \41902 , \41906 );
and \U$41664 ( \41979 , \41906 , \41911 );
and \U$41665 ( \41980 , \41902 , \41911 );
or \U$41666 ( \41981 , \41978 , \41979 , \41980 );
xor \U$41667 ( \41982 , \41977 , \41981 );
and \U$41668 ( \41983 , \41961 , \41965 );
and \U$41669 ( \41984 , \41965 , \41968 );
and \U$41670 ( \41985 , \41961 , \41968 );
or \U$41671 ( \41986 , \41983 , \41984 , \41985 );
xor \U$41672 ( \41987 , \41982 , \41986 );
xor \U$41673 ( \41988 , \41973 , \41987 );
and \U$41674 ( \41989 , \41940 , \41956 );
and \U$41675 ( \41990 , \41956 , \41969 );
and \U$41676 ( \41991 , \41940 , \41969 );
or \U$41677 ( \41992 , \41989 , \41990 , \41991 );
and \U$41678 ( \41993 , \41912 , \41922 );
xor \U$41679 ( \41994 , \41992 , \41993 );
and \U$41680 ( \41995 , \22696 , \22208 );
and \U$41681 ( \41996 , \22665 , \22206 );
nor \U$41682 ( \41997 , \41995 , \41996 );
xnor \U$41683 ( \41998 , \41997 , \22218 );
and \U$41684 ( \41999 , \22706 , \22230 );
and \U$41685 ( \42000 , \22686 , \22228 );
nor \U$41686 ( \42001 , \41999 , \42000 );
xnor \U$41687 ( \42002 , \42001 , \22240 );
xor \U$41688 ( \42003 , \41998 , \42002 );
and \U$41689 ( \42004 , \22624 , \22140 );
and \U$41690 ( \42005 , \22592 , \22138 );
nor \U$41691 ( \42006 , \42004 , \42005 );
xnor \U$41692 ( \42007 , \42006 , \22150 );
and \U$41693 ( \42008 , \22646 , \22162 );
and \U$41694 ( \42009 , \22613 , \22160 );
nor \U$41695 ( \42010 , \42008 , \42009 );
xnor \U$41696 ( \42011 , \42010 , \22172 );
xor \U$41697 ( \42012 , \42007 , \42011 );
and \U$41698 ( \42013 , \22676 , \22187 );
and \U$41699 ( \42014 , \22635 , \22185 );
nor \U$41700 ( \42015 , \42013 , \42014 );
xnor \U$41701 ( \42016 , \42015 , \22197 );
xor \U$41702 ( \42017 , \42012 , \42016 );
xor \U$41703 ( \42018 , \42003 , \42017 );
and \U$41704 ( \42019 , \22556 , \22076 );
and \U$41705 ( \42020 , \22524 , \22073 );
nor \U$41706 ( \42021 , \42019 , \42020 );
xnor \U$41707 ( \42022 , \42021 , \22072 );
and \U$41708 ( \42023 , \22578 , \22095 );
and \U$41709 ( \42024 , \22545 , \22093 );
nor \U$41710 ( \42025 , \42023 , \42024 );
xnor \U$41711 ( \42026 , \42025 , \22105 );
xor \U$41712 ( \42027 , \42022 , \42026 );
and \U$41713 ( \42028 , \22603 , \22119 );
and \U$41714 ( \42029 , \22567 , \22117 );
nor \U$41715 ( \42030 , \42028 , \42029 );
xnor \U$41716 ( \42031 , \42030 , \22129 );
xor \U$41717 ( \42032 , \42027 , \42031 );
xor \U$41718 ( \42033 , \42018 , \42032 );
xor \U$41719 ( \42034 , \41994 , \42033 );
xor \U$41720 ( \42035 , \41988 , \42034 );
and \U$41721 ( \42036 , \22603 , \22076 );
and \U$41722 ( \42037 , \22567 , \22073 );
nor \U$41723 ( \42038 , \42036 , \42037 );
xnor \U$41724 ( \42039 , \42038 , \22072 );
and \U$41725 ( \42040 , \22624 , \22095 );
and \U$41726 ( \42041 , \22592 , \22093 );
nor \U$41727 ( \42042 , \42040 , \42041 );
xnor \U$41728 ( \42043 , \42042 , \22105 );
and \U$41729 ( \42044 , \42039 , \42043 );
and \U$41730 ( \42045 , \22646 , \22119 );
and \U$41731 ( \42046 , \22613 , \22117 );
nor \U$41732 ( \42047 , \42045 , \42046 );
xnor \U$41733 ( \42048 , \42047 , \22129 );
and \U$41734 ( \42049 , \42043 , \42048 );
and \U$41735 ( \42050 , \42039 , \42048 );
or \U$41736 ( \42051 , \42044 , \42049 , \42050 );
and \U$41737 ( \42052 , \22676 , \22140 );
and \U$41738 ( \42053 , \22635 , \22138 );
nor \U$41739 ( \42054 , \42052 , \42053 );
xnor \U$41740 ( \42055 , \42054 , \22150 );
and \U$41741 ( \42056 , \22696 , \22162 );
and \U$41742 ( \42057 , \22665 , \22160 );
nor \U$41743 ( \42058 , \42056 , \42057 );
xnor \U$41744 ( \42059 , \42058 , \22172 );
and \U$41745 ( \42060 , \42055 , \42059 );
and \U$41746 ( \42061 , \22706 , \22187 );
and \U$41747 ( \42062 , \22686 , \22185 );
nor \U$41748 ( \42063 , \42061 , \42062 );
xnor \U$41749 ( \42064 , \42063 , \22197 );
and \U$41750 ( \42065 , \42059 , \42064 );
and \U$41751 ( \42066 , \42055 , \42064 );
or \U$41752 ( \42067 , \42060 , \42065 , \42066 );
and \U$41753 ( \42068 , \42051 , \42067 );
and \U$41754 ( \42069 , \22686 , \22187 );
and \U$41755 ( \42070 , \22696 , \22185 );
nor \U$41756 ( \42071 , \42069 , \42070 );
xnor \U$41757 ( \42072 , \42071 , \22197 );
and \U$41758 ( \42073 , \42067 , \42072 );
and \U$41759 ( \42074 , \42051 , \42072 );
or \U$41760 ( \42075 , \42068 , \42073 , \42074 );
nand \U$41761 ( \42076 , \22706 , \22206 );
xnor \U$41762 ( \42077 , \42076 , \22218 );
xor \U$41763 ( \42078 , \41878 , \41882 );
xor \U$41764 ( \42079 , \42078 , \41887 );
and \U$41765 ( \42080 , \42077 , \42079 );
xor \U$41766 ( \42081 , \22218 , \41866 );
xor \U$41767 ( \42082 , \42081 , \41871 );
and \U$41768 ( \42083 , \42079 , \42082 );
and \U$41769 ( \42084 , \42077 , \42082 );
or \U$41770 ( \42085 , \42080 , \42083 , \42084 );
and \U$41771 ( \42086 , \42075 , \42085 );
xor \U$41772 ( \42087 , \41944 , \41948 );
xor \U$41773 ( \42088 , \42087 , \41953 );
and \U$41774 ( \42089 , \42085 , \42088 );
and \U$41775 ( \42090 , \42075 , \42088 );
or \U$41776 ( \42091 , \42086 , \42089 , \42090 );
xor \U$41777 ( \42092 , \41928 , \41932 );
xor \U$41778 ( \42093 , \42092 , \41937 );
xor \U$41779 ( \42094 , \41874 , \41890 );
xor \U$41780 ( \42095 , \42094 , \41895 );
and \U$41781 ( \42096 , \42093 , \42095 );
and \U$41782 ( \42097 , \42091 , \42096 );
xor \U$41783 ( \42098 , \41898 , \41923 );
xor \U$41784 ( \42099 , \42098 , \41970 );
and \U$41785 ( \42100 , \42096 , \42099 );
and \U$41786 ( \42101 , \42091 , \42099 );
or \U$41787 ( \42102 , \42097 , \42100 , \42101 );
nor \U$41788 ( \42103 , \42035 , \42102 );
and \U$41789 ( \42104 , \41992 , \41993 );
and \U$41790 ( \42105 , \41993 , \42033 );
and \U$41791 ( \42106 , \41992 , \42033 );
or \U$41792 ( \42107 , \42104 , \42105 , \42106 );
nand \U$41793 ( \42108 , \22706 , \22255 );
xnor \U$41794 ( \42109 , \42108 , \22267 );
and \U$41795 ( \42110 , \22635 , \22187 );
and \U$41796 ( \42111 , \22646 , \22185 );
nor \U$41797 ( \42112 , \42110 , \42111 );
xnor \U$41798 ( \42113 , \42112 , \22197 );
and \U$41799 ( \42114 , \22665 , \22208 );
and \U$41800 ( \42115 , \22676 , \22206 );
nor \U$41801 ( \42116 , \42114 , \42115 );
xnor \U$41802 ( \42117 , \42116 , \22218 );
xor \U$41803 ( \42118 , \42113 , \42117 );
and \U$41804 ( \42119 , \22686 , \22230 );
and \U$41805 ( \42120 , \22696 , \22228 );
nor \U$41806 ( \42121 , \42119 , \42120 );
xnor \U$41807 ( \42122 , \42121 , \22240 );
xor \U$41808 ( \42123 , \42118 , \42122 );
xor \U$41809 ( \42124 , \42109 , \42123 );
and \U$41810 ( \42125 , \22567 , \22119 );
and \U$41811 ( \42126 , \22578 , \22117 );
nor \U$41812 ( \42127 , \42125 , \42126 );
xnor \U$41813 ( \42128 , \42127 , \22129 );
and \U$41814 ( \42129 , \22592 , \22140 );
and \U$41815 ( \42130 , \22603 , \22138 );
nor \U$41816 ( \42131 , \42129 , \42130 );
xnor \U$41817 ( \42132 , \42131 , \22150 );
xor \U$41818 ( \42133 , \42128 , \42132 );
and \U$41819 ( \42134 , \22613 , \22162 );
and \U$41820 ( \42135 , \22624 , \22160 );
nor \U$41821 ( \42136 , \42134 , \42135 );
xnor \U$41822 ( \42137 , \42136 , \22172 );
xor \U$41823 ( \42138 , \42133 , \42137 );
xor \U$41824 ( \42139 , \42124 , \42138 );
and \U$41825 ( \42140 , \42022 , \42026 );
and \U$41826 ( \42141 , \42026 , \42031 );
and \U$41827 ( \42142 , \42022 , \42031 );
or \U$41828 ( \42143 , \42140 , \42141 , \42142 );
and \U$41829 ( \42144 , \42007 , \42011 );
and \U$41830 ( \42145 , \42011 , \42016 );
and \U$41831 ( \42146 , \42007 , \42016 );
or \U$41832 ( \42147 , \42144 , \42145 , \42146 );
xor \U$41833 ( \42148 , \42143 , \42147 );
and \U$41834 ( \42149 , \41998 , \42002 );
xor \U$41835 ( \42150 , \42148 , \42149 );
xor \U$41836 ( \42151 , \42139 , \42150 );
xor \U$41837 ( \42152 , \42107 , \42151 );
and \U$41838 ( \42153 , \41977 , \41981 );
and \U$41839 ( \42154 , \41981 , \41986 );
and \U$41840 ( \42155 , \41977 , \41986 );
or \U$41841 ( \42156 , \42153 , \42154 , \42155 );
and \U$41842 ( \42157 , \42003 , \42017 );
and \U$41843 ( \42158 , \42017 , \42032 );
and \U$41844 ( \42159 , \42003 , \42032 );
or \U$41845 ( \42160 , \42157 , \42158 , \42159 );
xor \U$41846 ( \42161 , \42156 , \42160 );
and \U$41847 ( \42162 , \22524 , \22076 );
and \U$41848 ( \42163 , \22535 , \22073 );
nor \U$41849 ( \42164 , \42162 , \42163 );
xnor \U$41850 ( \42165 , \42164 , \22072 );
xor \U$41851 ( \42166 , \22267 , \42165 );
and \U$41852 ( \42167 , \22545 , \22095 );
and \U$41853 ( \42168 , \22556 , \22093 );
nor \U$41854 ( \42169 , \42167 , \42168 );
xnor \U$41855 ( \42170 , \42169 , \22105 );
xor \U$41856 ( \42171 , \42166 , \42170 );
xor \U$41857 ( \42172 , \42161 , \42171 );
xor \U$41858 ( \42173 , \42152 , \42172 );
and \U$41859 ( \42174 , \41973 , \41987 );
and \U$41860 ( \42175 , \41987 , \42034 );
and \U$41861 ( \42176 , \41973 , \42034 );
or \U$41862 ( \42177 , \42174 , \42175 , \42176 );
nor \U$41863 ( \42178 , \42173 , \42177 );
nor \U$41864 ( \42179 , \42103 , \42178 );
and \U$41865 ( \42180 , \42143 , \42147 );
and \U$41866 ( \42181 , \42147 , \42149 );
and \U$41867 ( \42182 , \42143 , \42149 );
or \U$41868 ( \42183 , \42180 , \42181 , \42182 );
and \U$41869 ( \42184 , \42109 , \42123 );
and \U$41870 ( \42185 , \42123 , \42138 );
and \U$41871 ( \42186 , \42109 , \42138 );
or \U$41872 ( \42187 , \42184 , \42185 , \42186 );
xor \U$41873 ( \42188 , \42183 , \42187 );
and \U$41874 ( \42189 , \22676 , \22208 );
and \U$41875 ( \42190 , \22635 , \22206 );
nor \U$41876 ( \42191 , \42189 , \42190 );
xnor \U$41877 ( \42192 , \42191 , \22218 );
and \U$41878 ( \42193 , \22696 , \22230 );
and \U$41879 ( \42194 , \22665 , \22228 );
nor \U$41880 ( \42195 , \42193 , \42194 );
xnor \U$41881 ( \42196 , \42195 , \22240 );
xor \U$41882 ( \42197 , \42192 , \42196 );
and \U$41883 ( \42198 , \22706 , \22257 );
and \U$41884 ( \42199 , \22686 , \22255 );
nor \U$41885 ( \42200 , \42198 , \42199 );
xnor \U$41886 ( \42201 , \42200 , \22267 );
xor \U$41887 ( \42202 , \42197 , \42201 );
and \U$41888 ( \42203 , \22603 , \22140 );
and \U$41889 ( \42204 , \22567 , \22138 );
nor \U$41890 ( \42205 , \42203 , \42204 );
xnor \U$41891 ( \42206 , \42205 , \22150 );
and \U$41892 ( \42207 , \22624 , \22162 );
and \U$41893 ( \42208 , \22592 , \22160 );
nor \U$41894 ( \42209 , \42207 , \42208 );
xnor \U$41895 ( \42210 , \42209 , \22172 );
xor \U$41896 ( \42211 , \42206 , \42210 );
and \U$41897 ( \42212 , \22646 , \22187 );
and \U$41898 ( \42213 , \22613 , \22185 );
nor \U$41899 ( \42214 , \42212 , \42213 );
xnor \U$41900 ( \42215 , \42214 , \22197 );
xor \U$41901 ( \42216 , \42211 , \42215 );
xor \U$41902 ( \42217 , \42202 , \42216 );
and \U$41903 ( \42218 , \22535 , \22076 );
and \U$41904 ( \42219 , \22500 , \22073 );
nor \U$41905 ( \42220 , \42218 , \42219 );
xnor \U$41906 ( \42221 , \42220 , \22072 );
and \U$41907 ( \42222 , \22556 , \22095 );
and \U$41908 ( \42223 , \22524 , \22093 );
nor \U$41909 ( \42224 , \42222 , \42223 );
xnor \U$41910 ( \42225 , \42224 , \22105 );
xor \U$41911 ( \42226 , \42221 , \42225 );
and \U$41912 ( \42227 , \22578 , \22119 );
and \U$41913 ( \42228 , \22545 , \22117 );
nor \U$41914 ( \42229 , \42227 , \42228 );
xnor \U$41915 ( \42230 , \42229 , \22129 );
xor \U$41916 ( \42231 , \42226 , \42230 );
xor \U$41917 ( \42232 , \42217 , \42231 );
xor \U$41918 ( \42233 , \42188 , \42232 );
and \U$41919 ( \42234 , \42156 , \42160 );
and \U$41920 ( \42235 , \42160 , \42171 );
and \U$41921 ( \42236 , \42156 , \42171 );
or \U$41922 ( \42237 , \42234 , \42235 , \42236 );
and \U$41923 ( \42238 , \42139 , \42150 );
xor \U$41924 ( \42239 , \42237 , \42238 );
and \U$41925 ( \42240 , \22267 , \42165 );
and \U$41926 ( \42241 , \42165 , \42170 );
and \U$41927 ( \42242 , \22267 , \42170 );
or \U$41928 ( \42243 , \42240 , \42241 , \42242 );
and \U$41929 ( \42244 , \42128 , \42132 );
and \U$41930 ( \42245 , \42132 , \42137 );
and \U$41931 ( \42246 , \42128 , \42137 );
or \U$41932 ( \42247 , \42244 , \42245 , \42246 );
xor \U$41933 ( \42248 , \42243 , \42247 );
and \U$41934 ( \42249 , \42113 , \42117 );
and \U$41935 ( \42250 , \42117 , \42122 );
and \U$41936 ( \42251 , \42113 , \42122 );
or \U$41937 ( \42252 , \42249 , \42250 , \42251 );
xor \U$41938 ( \42253 , \42248 , \42252 );
xor \U$41939 ( \42254 , \42239 , \42253 );
xor \U$41940 ( \42255 , \42233 , \42254 );
and \U$41941 ( \42256 , \42107 , \42151 );
and \U$41942 ( \42257 , \42151 , \42172 );
and \U$41943 ( \42258 , \42107 , \42172 );
or \U$41944 ( \42259 , \42256 , \42257 , \42258 );
nor \U$41945 ( \42260 , \42255 , \42259 );
and \U$41946 ( \42261 , \42237 , \42238 );
and \U$41947 ( \42262 , \42238 , \42253 );
and \U$41948 ( \42263 , \42237 , \42253 );
or \U$41949 ( \42264 , \42261 , \42262 , \42263 );
and \U$41950 ( \42265 , \42183 , \42187 );
and \U$41951 ( \42266 , \42187 , \42232 );
and \U$41952 ( \42267 , \42183 , \42232 );
or \U$41953 ( \42268 , \42265 , \42266 , \42267 );
and \U$41954 ( \42269 , \22500 , \22076 );
and \U$41955 ( \42270 , \22511 , \22073 );
nor \U$41956 ( \42271 , \42269 , \42270 );
xnor \U$41957 ( \42272 , \42271 , \22072 );
xor \U$41958 ( \42273 , \22288 , \42272 );
and \U$41959 ( \42274 , \22524 , \22095 );
and \U$41960 ( \42275 , \22535 , \22093 );
nor \U$41961 ( \42276 , \42274 , \42275 );
xnor \U$41962 ( \42277 , \42276 , \22105 );
xor \U$41963 ( \42278 , \42273 , \42277 );
and \U$41964 ( \42279 , \22686 , \22257 );
and \U$41965 ( \42280 , \22696 , \22255 );
nor \U$41966 ( \42281 , \42279 , \42280 );
xnor \U$41967 ( \42282 , \42281 , \22267 );
nand \U$41968 ( \42283 , \22706 , \22276 );
xnor \U$41969 ( \42284 , \42283 , \22288 );
xor \U$41970 ( \42285 , \42282 , \42284 );
and \U$41971 ( \42286 , \22613 , \22187 );
and \U$41972 ( \42287 , \22624 , \22185 );
nor \U$41973 ( \42288 , \42286 , \42287 );
xnor \U$41974 ( \42289 , \42288 , \22197 );
and \U$41975 ( \42290 , \22635 , \22208 );
and \U$41976 ( \42291 , \22646 , \22206 );
nor \U$41977 ( \42292 , \42290 , \42291 );
xnor \U$41978 ( \42293 , \42292 , \22218 );
xor \U$41979 ( \42294 , \42289 , \42293 );
and \U$41980 ( \42295 , \22665 , \22230 );
and \U$41981 ( \42296 , \22676 , \22228 );
nor \U$41982 ( \42297 , \42295 , \42296 );
xnor \U$41983 ( \42298 , \42297 , \22240 );
xor \U$41984 ( \42299 , \42294 , \42298 );
xor \U$41985 ( \42300 , \42285 , \42299 );
xor \U$41986 ( \42301 , \42278 , \42300 );
and \U$41987 ( \42302 , \42221 , \42225 );
and \U$41988 ( \42303 , \42225 , \42230 );
and \U$41989 ( \42304 , \42221 , \42230 );
or \U$41990 ( \42305 , \42302 , \42303 , \42304 );
and \U$41991 ( \42306 , \42206 , \42210 );
and \U$41992 ( \42307 , \42210 , \42215 );
and \U$41993 ( \42308 , \42206 , \42215 );
or \U$41994 ( \42309 , \42306 , \42307 , \42308 );
xor \U$41995 ( \42310 , \42305 , \42309 );
and \U$41996 ( \42311 , \42192 , \42196 );
and \U$41997 ( \42312 , \42196 , \42201 );
and \U$41998 ( \42313 , \42192 , \42201 );
or \U$41999 ( \42314 , \42311 , \42312 , \42313 );
xor \U$42000 ( \42315 , \42310 , \42314 );
xor \U$42001 ( \42316 , \42301 , \42315 );
xor \U$42002 ( \42317 , \42268 , \42316 );
and \U$42003 ( \42318 , \42243 , \42247 );
and \U$42004 ( \42319 , \42247 , \42252 );
and \U$42005 ( \42320 , \42243 , \42252 );
or \U$42006 ( \42321 , \42318 , \42319 , \42320 );
and \U$42007 ( \42322 , \42202 , \42216 );
and \U$42008 ( \42323 , \42216 , \42231 );
and \U$42009 ( \42324 , \42202 , \42231 );
or \U$42010 ( \42325 , \42322 , \42323 , \42324 );
xor \U$42011 ( \42326 , \42321 , \42325 );
and \U$42012 ( \42327 , \22545 , \22119 );
and \U$42013 ( \42328 , \22556 , \22117 );
nor \U$42014 ( \42329 , \42327 , \42328 );
xnor \U$42015 ( \42330 , \42329 , \22129 );
and \U$42016 ( \42331 , \22567 , \22140 );
and \U$42017 ( \42332 , \22578 , \22138 );
nor \U$42018 ( \42333 , \42331 , \42332 );
xnor \U$42019 ( \42334 , \42333 , \22150 );
xor \U$42020 ( \42335 , \42330 , \42334 );
and \U$42021 ( \42336 , \22592 , \22162 );
and \U$42022 ( \42337 , \22603 , \22160 );
nor \U$42023 ( \42338 , \42336 , \42337 );
xnor \U$42024 ( \42339 , \42338 , \22172 );
xor \U$42025 ( \42340 , \42335 , \42339 );
xor \U$42026 ( \42341 , \42326 , \42340 );
xor \U$42027 ( \42342 , \42317 , \42341 );
xor \U$42028 ( \42343 , \42264 , \42342 );
and \U$42029 ( \42344 , \42233 , \42254 );
nor \U$42030 ( \42345 , \42343 , \42344 );
nor \U$42031 ( \42346 , \42260 , \42345 );
nand \U$42032 ( \42347 , \42179 , \42346 );
and \U$42033 ( \42348 , \42268 , \42316 );
and \U$42034 ( \42349 , \42316 , \42341 );
and \U$42035 ( \42350 , \42268 , \42341 );
or \U$42036 ( \42351 , \42348 , \42349 , \42350 );
and \U$42037 ( \42352 , \22288 , \42272 );
and \U$42038 ( \42353 , \42272 , \42277 );
and \U$42039 ( \42354 , \22288 , \42277 );
or \U$42040 ( \42355 , \42352 , \42353 , \42354 );
and \U$42041 ( \42356 , \42330 , \42334 );
and \U$42042 ( \42357 , \42334 , \42339 );
and \U$42043 ( \42358 , \42330 , \42339 );
or \U$42044 ( \42359 , \42356 , \42357 , \42358 );
xor \U$42045 ( \42360 , \42355 , \42359 );
and \U$42046 ( \42361 , \42289 , \42293 );
and \U$42047 ( \42362 , \42293 , \42298 );
and \U$42048 ( \42363 , \42289 , \42298 );
or \U$42049 ( \42364 , \42361 , \42362 , \42363 );
xor \U$42050 ( \42365 , \42360 , \42364 );
and \U$42051 ( \42366 , \42305 , \42309 );
and \U$42052 ( \42367 , \42309 , \42314 );
and \U$42053 ( \42368 , \42305 , \42314 );
or \U$42054 ( \42369 , \42366 , \42367 , \42368 );
and \U$42055 ( \42370 , \42282 , \42284 );
and \U$42056 ( \42371 , \42284 , \42299 );
and \U$42057 ( \42372 , \42282 , \42299 );
or \U$42058 ( \42373 , \42370 , \42371 , \42372 );
xor \U$42059 ( \42374 , \42369 , \42373 );
and \U$42060 ( \42375 , \22511 , \22076 );
and \U$42061 ( \42376 , \22478 , \22073 );
nor \U$42062 ( \42377 , \42375 , \42376 );
xnor \U$42063 ( \42378 , \42377 , \22072 );
and \U$42064 ( \42379 , \22535 , \22095 );
and \U$42065 ( \42380 , \22500 , \22093 );
nor \U$42066 ( \42381 , \42379 , \42380 );
xnor \U$42067 ( \42382 , \42381 , \22105 );
xor \U$42068 ( \42383 , \42378 , \42382 );
and \U$42069 ( \42384 , \22556 , \22119 );
and \U$42070 ( \42385 , \22524 , \22117 );
nor \U$42071 ( \42386 , \42384 , \42385 );
xnor \U$42072 ( \42387 , \42386 , \22129 );
xor \U$42073 ( \42388 , \42383 , \42387 );
xor \U$42074 ( \42389 , \42374 , \42388 );
xor \U$42075 ( \42390 , \42365 , \42389 );
xor \U$42076 ( \42391 , \42351 , \42390 );
and \U$42077 ( \42392 , \42321 , \42325 );
and \U$42078 ( \42393 , \42325 , \42340 );
and \U$42079 ( \42394 , \42321 , \42340 );
or \U$42080 ( \42395 , \42392 , \42393 , \42394 );
and \U$42081 ( \42396 , \42278 , \42300 );
and \U$42082 ( \42397 , \42300 , \42315 );
and \U$42083 ( \42398 , \42278 , \42315 );
or \U$42084 ( \42399 , \42396 , \42397 , \42398 );
xor \U$42085 ( \42400 , \42395 , \42399 );
and \U$42086 ( \42401 , \22706 , \22278 );
and \U$42087 ( \42402 , \22686 , \22276 );
nor \U$42088 ( \42403 , \42401 , \42402 );
xnor \U$42089 ( \42404 , \42403 , \22288 );
and \U$42090 ( \42405 , \22646 , \22208 );
and \U$42091 ( \42406 , \22613 , \22206 );
nor \U$42092 ( \42407 , \42405 , \42406 );
xnor \U$42093 ( \42408 , \42407 , \22218 );
and \U$42094 ( \42409 , \22676 , \22230 );
and \U$42095 ( \42410 , \22635 , \22228 );
nor \U$42096 ( \42411 , \42409 , \42410 );
xnor \U$42097 ( \42412 , \42411 , \22240 );
xor \U$42098 ( \42413 , \42408 , \42412 );
and \U$42099 ( \42414 , \22696 , \22257 );
and \U$42100 ( \42415 , \22665 , \22255 );
nor \U$42101 ( \42416 , \42414 , \42415 );
xnor \U$42102 ( \42417 , \42416 , \22267 );
xor \U$42103 ( \42418 , \42413 , \42417 );
xor \U$42104 ( \42419 , \42404 , \42418 );
and \U$42105 ( \42420 , \22578 , \22140 );
and \U$42106 ( \42421 , \22545 , \22138 );
nor \U$42107 ( \42422 , \42420 , \42421 );
xnor \U$42108 ( \42423 , \42422 , \22150 );
and \U$42109 ( \42424 , \22603 , \22162 );
and \U$42110 ( \42425 , \22567 , \22160 );
nor \U$42111 ( \42426 , \42424 , \42425 );
xnor \U$42112 ( \42427 , \42426 , \22172 );
xor \U$42113 ( \42428 , \42423 , \42427 );
and \U$42114 ( \42429 , \22624 , \22187 );
and \U$42115 ( \42430 , \22592 , \22185 );
nor \U$42116 ( \42431 , \42429 , \42430 );
xnor \U$42117 ( \42432 , \42431 , \22197 );
xor \U$42118 ( \42433 , \42428 , \42432 );
xor \U$42119 ( \42434 , \42419 , \42433 );
xor \U$42120 ( \42435 , \42400 , \42434 );
xor \U$42121 ( \42436 , \42391 , \42435 );
and \U$42122 ( \42437 , \42264 , \42342 );
nor \U$42123 ( \42438 , \42436 , \42437 );
and \U$42124 ( \42439 , \42395 , \42399 );
and \U$42125 ( \42440 , \42399 , \42434 );
and \U$42126 ( \42441 , \42395 , \42434 );
or \U$42127 ( \42442 , \42439 , \42440 , \42441 );
and \U$42128 ( \42443 , \42365 , \42389 );
xor \U$42129 ( \42444 , \42442 , \42443 );
and \U$42130 ( \42445 , \42369 , \42373 );
and \U$42131 ( \42446 , \42373 , \42388 );
and \U$42132 ( \42447 , \42369 , \42388 );
or \U$42133 ( \42448 , \42445 , \42446 , \42447 );
and \U$42134 ( \42449 , \22665 , \22257 );
and \U$42135 ( \42450 , \22676 , \22255 );
nor \U$42136 ( \42451 , \42449 , \42450 );
xnor \U$42137 ( \42452 , \42451 , \22267 );
and \U$42138 ( \42453 , \22686 , \22278 );
and \U$42139 ( \42454 , \22696 , \22276 );
nor \U$42140 ( \42455 , \42453 , \42454 );
xnor \U$42141 ( \42456 , \42455 , \22288 );
xor \U$42142 ( \42457 , \42452 , \42456 );
nand \U$42143 ( \42458 , \22706 , \22298 );
xnor \U$42144 ( \42459 , \42458 , \22310 );
xor \U$42145 ( \42460 , \42457 , \42459 );
and \U$42146 ( \42461 , \22592 , \22187 );
and \U$42147 ( \42462 , \22603 , \22185 );
nor \U$42148 ( \42463 , \42461 , \42462 );
xnor \U$42149 ( \42464 , \42463 , \22197 );
and \U$42150 ( \42465 , \22613 , \22208 );
and \U$42151 ( \42466 , \22624 , \22206 );
nor \U$42152 ( \42467 , \42465 , \42466 );
xnor \U$42153 ( \42468 , \42467 , \22218 );
xor \U$42154 ( \42469 , \42464 , \42468 );
and \U$42155 ( \42470 , \22635 , \22230 );
and \U$42156 ( \42471 , \22646 , \22228 );
nor \U$42157 ( \42472 , \42470 , \42471 );
xnor \U$42158 ( \42473 , \42472 , \22240 );
xor \U$42159 ( \42474 , \42469 , \42473 );
xor \U$42160 ( \42475 , \42460 , \42474 );
and \U$42161 ( \42476 , \22524 , \22119 );
and \U$42162 ( \42477 , \22535 , \22117 );
nor \U$42163 ( \42478 , \42476 , \42477 );
xnor \U$42164 ( \42479 , \42478 , \22129 );
and \U$42165 ( \42480 , \22545 , \22140 );
and \U$42166 ( \42481 , \22556 , \22138 );
nor \U$42167 ( \42482 , \42480 , \42481 );
xnor \U$42168 ( \42483 , \42482 , \22150 );
xor \U$42169 ( \42484 , \42479 , \42483 );
and \U$42170 ( \42485 , \22567 , \22162 );
and \U$42171 ( \42486 , \22578 , \22160 );
nor \U$42172 ( \42487 , \42485 , \42486 );
xnor \U$42173 ( \42488 , \42487 , \22172 );
xor \U$42174 ( \42489 , \42484 , \42488 );
xor \U$42175 ( \42490 , \42475 , \42489 );
and \U$42176 ( \42491 , \42378 , \42382 );
and \U$42177 ( \42492 , \42382 , \42387 );
and \U$42178 ( \42493 , \42378 , \42387 );
or \U$42179 ( \42494 , \42491 , \42492 , \42493 );
and \U$42180 ( \42495 , \42423 , \42427 );
and \U$42181 ( \42496 , \42427 , \42432 );
and \U$42182 ( \42497 , \42423 , \42432 );
or \U$42183 ( \42498 , \42495 , \42496 , \42497 );
xor \U$42184 ( \42499 , \42494 , \42498 );
and \U$42185 ( \42500 , \42408 , \42412 );
and \U$42186 ( \42501 , \42412 , \42417 );
and \U$42187 ( \42502 , \42408 , \42417 );
or \U$42188 ( \42503 , \42500 , \42501 , \42502 );
xor \U$42189 ( \42504 , \42499 , \42503 );
xor \U$42190 ( \42505 , \42490 , \42504 );
xor \U$42191 ( \42506 , \42448 , \42505 );
and \U$42192 ( \42507 , \42355 , \42359 );
and \U$42193 ( \42508 , \42359 , \42364 );
and \U$42194 ( \42509 , \42355 , \42364 );
or \U$42195 ( \42510 , \42507 , \42508 , \42509 );
and \U$42196 ( \42511 , \42404 , \42418 );
and \U$42197 ( \42512 , \42418 , \42433 );
and \U$42198 ( \42513 , \42404 , \42433 );
or \U$42199 ( \42514 , \42511 , \42512 , \42513 );
xor \U$42200 ( \42515 , \42510 , \42514 );
and \U$42201 ( \42516 , \22478 , \22076 );
and \U$42202 ( \42517 , \22489 , \22073 );
nor \U$42203 ( \42518 , \42516 , \42517 );
xnor \U$42204 ( \42519 , \42518 , \22072 );
xor \U$42205 ( \42520 , \22310 , \42519 );
and \U$42206 ( \42521 , \22500 , \22095 );
and \U$42207 ( \42522 , \22511 , \22093 );
nor \U$42208 ( \42523 , \42521 , \42522 );
xnor \U$42209 ( \42524 , \42523 , \22105 );
xor \U$42210 ( \42525 , \42520 , \42524 );
xor \U$42211 ( \42526 , \42515 , \42525 );
xor \U$42212 ( \42527 , \42506 , \42526 );
xor \U$42213 ( \42528 , \42444 , \42527 );
and \U$42214 ( \42529 , \42351 , \42390 );
and \U$42215 ( \42530 , \42390 , \42435 );
and \U$42216 ( \42531 , \42351 , \42435 );
or \U$42217 ( \42532 , \42529 , \42530 , \42531 );
nor \U$42218 ( \42533 , \42528 , \42532 );
nor \U$42219 ( \42534 , \42438 , \42533 );
and \U$42220 ( \42535 , \42448 , \42505 );
and \U$42221 ( \42536 , \42505 , \42526 );
and \U$42222 ( \42537 , \42448 , \42526 );
or \U$42223 ( \42538 , \42535 , \42536 , \42537 );
and \U$42224 ( \42539 , \22310 , \42519 );
and \U$42225 ( \42540 , \42519 , \42524 );
and \U$42226 ( \42541 , \22310 , \42524 );
or \U$42227 ( \42542 , \42539 , \42540 , \42541 );
and \U$42228 ( \42543 , \42479 , \42483 );
and \U$42229 ( \42544 , \42483 , \42488 );
and \U$42230 ( \42545 , \42479 , \42488 );
or \U$42231 ( \42546 , \42543 , \42544 , \42545 );
xor \U$42232 ( \42547 , \42542 , \42546 );
and \U$42233 ( \42548 , \42464 , \42468 );
and \U$42234 ( \42549 , \42468 , \42473 );
and \U$42235 ( \42550 , \42464 , \42473 );
or \U$42236 ( \42551 , \42548 , \42549 , \42550 );
xor \U$42237 ( \42552 , \42547 , \42551 );
and \U$42238 ( \42553 , \42494 , \42498 );
and \U$42239 ( \42554 , \42498 , \42503 );
and \U$42240 ( \42555 , \42494 , \42503 );
or \U$42241 ( \42556 , \42553 , \42554 , \42555 );
and \U$42242 ( \42557 , \42460 , \42474 );
and \U$42243 ( \42558 , \42474 , \42489 );
and \U$42244 ( \42559 , \42460 , \42489 );
or \U$42245 ( \42560 , \42557 , \42558 , \42559 );
xor \U$42246 ( \42561 , \42556 , \42560 );
and \U$42247 ( \42562 , \22624 , \22208 );
and \U$42248 ( \42563 , \22592 , \22206 );
nor \U$42249 ( \42564 , \42562 , \42563 );
xnor \U$42250 ( \42565 , \42564 , \22218 );
and \U$42251 ( \42566 , \22646 , \22230 );
and \U$42252 ( \42567 , \22613 , \22228 );
nor \U$42253 ( \42568 , \42566 , \42567 );
xnor \U$42254 ( \42569 , \42568 , \22240 );
xor \U$42255 ( \42570 , \42565 , \42569 );
and \U$42256 ( \42571 , \22676 , \22257 );
and \U$42257 ( \42572 , \22635 , \22255 );
nor \U$42258 ( \42573 , \42571 , \42572 );
xnor \U$42259 ( \42574 , \42573 , \22267 );
xor \U$42260 ( \42575 , \42570 , \42574 );
and \U$42261 ( \42576 , \22556 , \22140 );
and \U$42262 ( \42577 , \22524 , \22138 );
nor \U$42263 ( \42578 , \42576 , \42577 );
xnor \U$42264 ( \42579 , \42578 , \22150 );
and \U$42265 ( \42580 , \22578 , \22162 );
and \U$42266 ( \42581 , \22545 , \22160 );
nor \U$42267 ( \42582 , \42580 , \42581 );
xnor \U$42268 ( \42583 , \42582 , \22172 );
xor \U$42269 ( \42584 , \42579 , \42583 );
and \U$42270 ( \42585 , \22603 , \22187 );
and \U$42271 ( \42586 , \22567 , \22185 );
nor \U$42272 ( \42587 , \42585 , \42586 );
xnor \U$42273 ( \42588 , \42587 , \22197 );
xor \U$42274 ( \42589 , \42584 , \42588 );
xor \U$42275 ( \42590 , \42575 , \42589 );
and \U$42276 ( \42591 , \22489 , \22076 );
and \U$42277 ( \42592 , \22457 , \22073 );
nor \U$42278 ( \42593 , \42591 , \42592 );
xnor \U$42279 ( \42594 , \42593 , \22072 );
and \U$42280 ( \42595 , \22511 , \22095 );
and \U$42281 ( \42596 , \22478 , \22093 );
nor \U$42282 ( \42597 , \42595 , \42596 );
xnor \U$42283 ( \42598 , \42597 , \22105 );
xor \U$42284 ( \42599 , \42594 , \42598 );
and \U$42285 ( \42600 , \22535 , \22119 );
and \U$42286 ( \42601 , \22500 , \22117 );
nor \U$42287 ( \42602 , \42600 , \42601 );
xnor \U$42288 ( \42603 , \42602 , \22129 );
xor \U$42289 ( \42604 , \42599 , \42603 );
xor \U$42290 ( \42605 , \42590 , \42604 );
xor \U$42291 ( \42606 , \42561 , \42605 );
xor \U$42292 ( \42607 , \42552 , \42606 );
xor \U$42293 ( \42608 , \42538 , \42607 );
and \U$42294 ( \42609 , \42510 , \42514 );
and \U$42295 ( \42610 , \42514 , \42525 );
and \U$42296 ( \42611 , \42510 , \42525 );
or \U$42297 ( \42612 , \42609 , \42610 , \42611 );
and \U$42298 ( \42613 , \42490 , \42504 );
xor \U$42299 ( \42614 , \42612 , \42613 );
and \U$42300 ( \42615 , \42452 , \42456 );
and \U$42301 ( \42616 , \42456 , \42459 );
and \U$42302 ( \42617 , \42452 , \42459 );
or \U$42303 ( \42618 , \42615 , \42616 , \42617 );
and \U$42304 ( \42619 , \22696 , \22278 );
and \U$42305 ( \42620 , \22665 , \22276 );
nor \U$42306 ( \42621 , \42619 , \42620 );
xnor \U$42307 ( \42622 , \42621 , \22288 );
xor \U$42308 ( \42623 , \42618 , \42622 );
and \U$42309 ( \42624 , \22706 , \22300 );
and \U$42310 ( \42625 , \22686 , \22298 );
nor \U$42311 ( \42626 , \42624 , \42625 );
xnor \U$42312 ( \42627 , \42626 , \22310 );
xor \U$42313 ( \42628 , \42623 , \42627 );
xor \U$42314 ( \42629 , \42614 , \42628 );
xor \U$42315 ( \42630 , \42608 , \42629 );
and \U$42316 ( \42631 , \42442 , \42443 );
and \U$42317 ( \42632 , \42443 , \42527 );
and \U$42318 ( \42633 , \42442 , \42527 );
or \U$42319 ( \42634 , \42631 , \42632 , \42633 );
nor \U$42320 ( \42635 , \42630 , \42634 );
and \U$42321 ( \42636 , \42612 , \42613 );
and \U$42322 ( \42637 , \42613 , \42628 );
and \U$42323 ( \42638 , \42612 , \42628 );
or \U$42324 ( \42639 , \42636 , \42637 , \42638 );
and \U$42325 ( \42640 , \42552 , \42606 );
xor \U$42326 ( \42641 , \42639 , \42640 );
and \U$42327 ( \42642 , \42556 , \42560 );
and \U$42328 ( \42643 , \42560 , \42605 );
and \U$42329 ( \42644 , \42556 , \42605 );
or \U$42330 ( \42645 , \42642 , \42643 , \42644 );
and \U$42331 ( \42646 , \22500 , \22119 );
and \U$42332 ( \42647 , \22511 , \22117 );
nor \U$42333 ( \42648 , \42646 , \42647 );
xnor \U$42334 ( \42649 , \42648 , \22129 );
and \U$42335 ( \42650 , \22524 , \22140 );
and \U$42336 ( \42651 , \22535 , \22138 );
nor \U$42337 ( \42652 , \42650 , \42651 );
xnor \U$42338 ( \42653 , \42652 , \22150 );
xor \U$42339 ( \42654 , \42649 , \42653 );
and \U$42340 ( \42655 , \22545 , \22162 );
and \U$42341 ( \42656 , \22556 , \22160 );
nor \U$42342 ( \42657 , \42655 , \42656 );
xnor \U$42343 ( \42658 , \42657 , \22172 );
xor \U$42344 ( \42659 , \42654 , \42658 );
and \U$42345 ( \42660 , \22457 , \22076 );
and \U$42346 ( \42661 , \22468 , \22073 );
nor \U$42347 ( \42662 , \42660 , \42661 );
xnor \U$42348 ( \42663 , \42662 , \22072 );
xor \U$42349 ( \42664 , \22334 , \42663 );
and \U$42350 ( \42665 , \22478 , \22095 );
and \U$42351 ( \42666 , \22489 , \22093 );
nor \U$42352 ( \42667 , \42665 , \42666 );
xnor \U$42353 ( \42668 , \42667 , \22105 );
xor \U$42354 ( \42669 , \42664 , \42668 );
xor \U$42355 ( \42670 , \42659 , \42669 );
nand \U$42356 ( \42671 , \22706 , \22322 );
xnor \U$42357 ( \42672 , \42671 , \22334 );
and \U$42358 ( \42673 , \22635 , \22257 );
and \U$42359 ( \42674 , \22646 , \22255 );
nor \U$42360 ( \42675 , \42673 , \42674 );
xnor \U$42361 ( \42676 , \42675 , \22267 );
and \U$42362 ( \42677 , \22665 , \22278 );
and \U$42363 ( \42678 , \22676 , \22276 );
nor \U$42364 ( \42679 , \42677 , \42678 );
xnor \U$42365 ( \42680 , \42679 , \22288 );
xor \U$42366 ( \42681 , \42676 , \42680 );
and \U$42367 ( \42682 , \22686 , \22300 );
and \U$42368 ( \42683 , \22696 , \22298 );
nor \U$42369 ( \42684 , \42682 , \42683 );
xnor \U$42370 ( \42685 , \42684 , \22310 );
xor \U$42371 ( \42686 , \42681 , \42685 );
xor \U$42372 ( \42687 , \42672 , \42686 );
and \U$42373 ( \42688 , \22567 , \22187 );
and \U$42374 ( \42689 , \22578 , \22185 );
nor \U$42375 ( \42690 , \42688 , \42689 );
xnor \U$42376 ( \42691 , \42690 , \22197 );
and \U$42377 ( \42692 , \22592 , \22208 );
and \U$42378 ( \42693 , \22603 , \22206 );
nor \U$42379 ( \42694 , \42692 , \42693 );
xnor \U$42380 ( \42695 , \42694 , \22218 );
xor \U$42381 ( \42696 , \42691 , \42695 );
and \U$42382 ( \42697 , \22613 , \22230 );
and \U$42383 ( \42698 , \22624 , \22228 );
nor \U$42384 ( \42699 , \42697 , \42698 );
xnor \U$42385 ( \42700 , \42699 , \22240 );
xor \U$42386 ( \42701 , \42696 , \42700 );
xor \U$42387 ( \42702 , \42687 , \42701 );
xor \U$42388 ( \42703 , \42670 , \42702 );
and \U$42389 ( \42704 , \42594 , \42598 );
and \U$42390 ( \42705 , \42598 , \42603 );
and \U$42391 ( \42706 , \42594 , \42603 );
or \U$42392 ( \42707 , \42704 , \42705 , \42706 );
and \U$42393 ( \42708 , \42579 , \42583 );
and \U$42394 ( \42709 , \42583 , \42588 );
and \U$42395 ( \42710 , \42579 , \42588 );
or \U$42396 ( \42711 , \42708 , \42709 , \42710 );
xor \U$42397 ( \42712 , \42707 , \42711 );
and \U$42398 ( \42713 , \42565 , \42569 );
and \U$42399 ( \42714 , \42569 , \42574 );
and \U$42400 ( \42715 , \42565 , \42574 );
or \U$42401 ( \42716 , \42713 , \42714 , \42715 );
xor \U$42402 ( \42717 , \42712 , \42716 );
xor \U$42403 ( \42718 , \42703 , \42717 );
xor \U$42404 ( \42719 , \42645 , \42718 );
and \U$42405 ( \42720 , \42542 , \42546 );
and \U$42406 ( \42721 , \42546 , \42551 );
and \U$42407 ( \42722 , \42542 , \42551 );
or \U$42408 ( \42723 , \42720 , \42721 , \42722 );
and \U$42409 ( \42724 , \42618 , \42622 );
and \U$42410 ( \42725 , \42622 , \42627 );
and \U$42411 ( \42726 , \42618 , \42627 );
or \U$42412 ( \42727 , \42724 , \42725 , \42726 );
xor \U$42413 ( \42728 , \42723 , \42727 );
and \U$42414 ( \42729 , \42575 , \42589 );
and \U$42415 ( \42730 , \42589 , \42604 );
and \U$42416 ( \42731 , \42575 , \42604 );
or \U$42417 ( \42732 , \42729 , \42730 , \42731 );
xor \U$42418 ( \42733 , \42728 , \42732 );
xor \U$42419 ( \42734 , \42719 , \42733 );
xor \U$42420 ( \42735 , \42641 , \42734 );
and \U$42421 ( \42736 , \42538 , \42607 );
and \U$42422 ( \42737 , \42607 , \42629 );
and \U$42423 ( \42738 , \42538 , \42629 );
or \U$42424 ( \42739 , \42736 , \42737 , \42738 );
nor \U$42425 ( \42740 , \42735 , \42739 );
nor \U$42426 ( \42741 , \42635 , \42740 );
nand \U$42427 ( \42742 , \42534 , \42741 );
nor \U$42428 ( \42743 , \42347 , \42742 );
and \U$42429 ( \42744 , \42645 , \42718 );
and \U$42430 ( \42745 , \42718 , \42733 );
and \U$42431 ( \42746 , \42645 , \42733 );
or \U$42432 ( \42747 , \42744 , \42745 , \42746 );
and \U$42433 ( \42748 , \42707 , \42711 );
and \U$42434 ( \42749 , \42711 , \42716 );
and \U$42435 ( \42750 , \42707 , \42716 );
or \U$42436 ( \42751 , \42748 , \42749 , \42750 );
and \U$42437 ( \42752 , \42672 , \42686 );
and \U$42438 ( \42753 , \42686 , \42701 );
and \U$42439 ( \42754 , \42672 , \42701 );
or \U$42440 ( \42755 , \42752 , \42753 , \42754 );
xor \U$42441 ( \42756 , \42751 , \42755 );
and \U$42442 ( \42757 , \42659 , \42669 );
xor \U$42443 ( \42758 , \42756 , \42757 );
xor \U$42444 ( \42759 , \42747 , \42758 );
and \U$42445 ( \42760 , \42723 , \42727 );
and \U$42446 ( \42761 , \42727 , \42732 );
and \U$42447 ( \42762 , \42723 , \42732 );
or \U$42448 ( \42763 , \42760 , \42761 , \42762 );
and \U$42449 ( \42764 , \42670 , \42702 );
and \U$42450 ( \42765 , \42702 , \42717 );
and \U$42451 ( \42766 , \42670 , \42717 );
or \U$42452 ( \42767 , \42764 , \42765 , \42766 );
xor \U$42453 ( \42768 , \42763 , \42767 );
and \U$42454 ( \42769 , \22535 , \22140 );
and \U$42455 ( \42770 , \22500 , \22138 );
nor \U$42456 ( \42771 , \42769 , \42770 );
xnor \U$42457 ( \42772 , \42771 , \22150 );
and \U$42458 ( \42773 , \22556 , \22162 );
and \U$42459 ( \42774 , \22524 , \22160 );
nor \U$42460 ( \42775 , \42773 , \42774 );
xnor \U$42461 ( \42776 , \42775 , \22172 );
xor \U$42462 ( \42777 , \42772 , \42776 );
and \U$42463 ( \42778 , \22578 , \22187 );
and \U$42464 ( \42779 , \22545 , \22185 );
nor \U$42465 ( \42780 , \42778 , \42779 );
xnor \U$42466 ( \42781 , \42780 , \22197 );
xor \U$42467 ( \42782 , \42777 , \42781 );
and \U$42468 ( \42783 , \22468 , \22076 );
and \U$42469 ( \42784 , \22429 , \22073 );
nor \U$42470 ( \42785 , \42783 , \42784 );
xnor \U$42471 ( \42786 , \42785 , \22072 );
and \U$42472 ( \42787 , \22489 , \22095 );
and \U$42473 ( \42788 , \22457 , \22093 );
nor \U$42474 ( \42789 , \42787 , \42788 );
xnor \U$42475 ( \42790 , \42789 , \22105 );
xor \U$42476 ( \42791 , \42786 , \42790 );
and \U$42477 ( \42792 , \22511 , \22119 );
and \U$42478 ( \42793 , \22478 , \22117 );
nor \U$42479 ( \42794 , \42792 , \42793 );
xnor \U$42480 ( \42795 , \42794 , \22129 );
xor \U$42481 ( \42796 , \42791 , \42795 );
xor \U$42482 ( \42797 , \42782 , \42796 );
and \U$42483 ( \42798 , \42676 , \42680 );
and \U$42484 ( \42799 , \42680 , \42685 );
and \U$42485 ( \42800 , \42676 , \42685 );
or \U$42486 ( \42801 , \42798 , \42799 , \42800 );
and \U$42487 ( \42802 , \22676 , \22278 );
and \U$42488 ( \42803 , \22635 , \22276 );
nor \U$42489 ( \42804 , \42802 , \42803 );
xnor \U$42490 ( \42805 , \42804 , \22288 );
and \U$42491 ( \42806 , \22696 , \22300 );
and \U$42492 ( \42807 , \22665 , \22298 );
nor \U$42493 ( \42808 , \42806 , \42807 );
xnor \U$42494 ( \42809 , \42808 , \22310 );
xor \U$42495 ( \42810 , \42805 , \42809 );
and \U$42496 ( \42811 , \22706 , \22324 );
and \U$42497 ( \42812 , \22686 , \22322 );
nor \U$42498 ( \42813 , \42811 , \42812 );
xnor \U$42499 ( \42814 , \42813 , \22334 );
xor \U$42500 ( \42815 , \42810 , \42814 );
xor \U$42501 ( \42816 , \42801 , \42815 );
and \U$42502 ( \42817 , \22603 , \22208 );
and \U$42503 ( \42818 , \22567 , \22206 );
nor \U$42504 ( \42819 , \42817 , \42818 );
xnor \U$42505 ( \42820 , \42819 , \22218 );
and \U$42506 ( \42821 , \22624 , \22230 );
and \U$42507 ( \42822 , \22592 , \22228 );
nor \U$42508 ( \42823 , \42821 , \42822 );
xnor \U$42509 ( \42824 , \42823 , \22240 );
xor \U$42510 ( \42825 , \42820 , \42824 );
and \U$42511 ( \42826 , \22646 , \22257 );
and \U$42512 ( \42827 , \22613 , \22255 );
nor \U$42513 ( \42828 , \42826 , \42827 );
xnor \U$42514 ( \42829 , \42828 , \22267 );
xor \U$42515 ( \42830 , \42825 , \42829 );
xor \U$42516 ( \42831 , \42816 , \42830 );
xor \U$42517 ( \42832 , \42797 , \42831 );
and \U$42518 ( \42833 , \22334 , \42663 );
and \U$42519 ( \42834 , \42663 , \42668 );
and \U$42520 ( \42835 , \22334 , \42668 );
or \U$42521 ( \42836 , \42833 , \42834 , \42835 );
and \U$42522 ( \42837 , \42649 , \42653 );
and \U$42523 ( \42838 , \42653 , \42658 );
and \U$42524 ( \42839 , \42649 , \42658 );
or \U$42525 ( \42840 , \42837 , \42838 , \42839 );
xor \U$42526 ( \42841 , \42836 , \42840 );
and \U$42527 ( \42842 , \42691 , \42695 );
and \U$42528 ( \42843 , \42695 , \42700 );
and \U$42529 ( \42844 , \42691 , \42700 );
or \U$42530 ( \42845 , \42842 , \42843 , \42844 );
xor \U$42531 ( \42846 , \42841 , \42845 );
xor \U$42532 ( \42847 , \42832 , \42846 );
xor \U$42533 ( \42848 , \42768 , \42847 );
xor \U$42534 ( \42849 , \42759 , \42848 );
and \U$42535 ( \42850 , \42639 , \42640 );
and \U$42536 ( \42851 , \42640 , \42734 );
and \U$42537 ( \42852 , \42639 , \42734 );
or \U$42538 ( \42853 , \42850 , \42851 , \42852 );
nor \U$42539 ( \42854 , \42849 , \42853 );
and \U$42540 ( \42855 , \42763 , \42767 );
and \U$42541 ( \42856 , \42767 , \42847 );
and \U$42542 ( \42857 , \42763 , \42847 );
or \U$42543 ( \42858 , \42855 , \42856 , \42857 );
and \U$42544 ( \42859 , \42836 , \42840 );
and \U$42545 ( \42860 , \42840 , \42845 );
and \U$42546 ( \42861 , \42836 , \42845 );
or \U$42547 ( \42862 , \42859 , \42860 , \42861 );
and \U$42548 ( \42863 , \42801 , \42815 );
and \U$42549 ( \42864 , \42815 , \42830 );
and \U$42550 ( \42865 , \42801 , \42830 );
or \U$42551 ( \42866 , \42863 , \42864 , \42865 );
xor \U$42552 ( \42867 , \42862 , \42866 );
and \U$42553 ( \42868 , \42782 , \42796 );
xor \U$42554 ( \42869 , \42867 , \42868 );
xor \U$42555 ( \42870 , \42858 , \42869 );
and \U$42556 ( \42871 , \42751 , \42755 );
and \U$42557 ( \42872 , \42755 , \42757 );
and \U$42558 ( \42873 , \42751 , \42757 );
or \U$42559 ( \42874 , \42871 , \42872 , \42873 );
and \U$42560 ( \42875 , \42797 , \42831 );
and \U$42561 ( \42876 , \42831 , \42846 );
and \U$42562 ( \42877 , \42797 , \42846 );
or \U$42563 ( \42878 , \42875 , \42876 , \42877 );
xor \U$42564 ( \42879 , \42874 , \42878 );
and \U$42565 ( \42880 , \22545 , \22187 );
and \U$42566 ( \42881 , \22556 , \22185 );
nor \U$42567 ( \42882 , \42880 , \42881 );
xnor \U$42568 ( \42883 , \42882 , \22197 );
and \U$42569 ( \42884 , \22567 , \22208 );
and \U$42570 ( \42885 , \22578 , \22206 );
nor \U$42571 ( \42886 , \42884 , \42885 );
xnor \U$42572 ( \42887 , \42886 , \22218 );
xor \U$42573 ( \42888 , \42883 , \42887 );
and \U$42574 ( \42889 , \22592 , \22230 );
and \U$42575 ( \42890 , \22603 , \22228 );
nor \U$42576 ( \42891 , \42889 , \42890 );
xnor \U$42577 ( \42892 , \42891 , \22240 );
xor \U$42578 ( \42893 , \42888 , \42892 );
and \U$42579 ( \42894 , \22478 , \22119 );
and \U$42580 ( \42895 , \22489 , \22117 );
nor \U$42581 ( \42896 , \42894 , \42895 );
xnor \U$42582 ( \42897 , \42896 , \22129 );
and \U$42583 ( \42898 , \22500 , \22140 );
and \U$42584 ( \42899 , \22511 , \22138 );
nor \U$42585 ( \42900 , \42898 , \42899 );
xnor \U$42586 ( \42901 , \42900 , \22150 );
xor \U$42587 ( \42902 , \42897 , \42901 );
and \U$42588 ( \42903 , \22524 , \22162 );
and \U$42589 ( \42904 , \22535 , \22160 );
nor \U$42590 ( \42905 , \42903 , \42904 );
xnor \U$42591 ( \42906 , \42905 , \22172 );
xor \U$42592 ( \42907 , \42902 , \42906 );
xor \U$42593 ( \42908 , \42893 , \42907 );
and \U$42594 ( \42909 , \22429 , \22076 );
and \U$42595 ( \42910 , \22440 , \22073 );
nor \U$42596 ( \42911 , \42909 , \42910 );
xnor \U$42597 ( \42912 , \42911 , \22072 );
xor \U$42598 ( \42913 , \22355 , \42912 );
and \U$42599 ( \42914 , \22457 , \22095 );
and \U$42600 ( \42915 , \22468 , \22093 );
nor \U$42601 ( \42916 , \42914 , \42915 );
xnor \U$42602 ( \42917 , \42916 , \22105 );
xor \U$42603 ( \42918 , \42913 , \42917 );
xor \U$42604 ( \42919 , \42908 , \42918 );
and \U$42605 ( \42920 , \42805 , \42809 );
and \U$42606 ( \42921 , \42809 , \42814 );
and \U$42607 ( \42922 , \42805 , \42814 );
or \U$42608 ( \42923 , \42920 , \42921 , \42922 );
and \U$42609 ( \42924 , \22686 , \22324 );
and \U$42610 ( \42925 , \22696 , \22322 );
nor \U$42611 ( \42926 , \42924 , \42925 );
xnor \U$42612 ( \42927 , \42926 , \22334 );
nand \U$42613 ( \42928 , \22706 , \22343 );
xnor \U$42614 ( \42929 , \42928 , \22355 );
xor \U$42615 ( \42930 , \42927 , \42929 );
xor \U$42616 ( \42931 , \42923 , \42930 );
and \U$42617 ( \42932 , \22613 , \22257 );
and \U$42618 ( \42933 , \22624 , \22255 );
nor \U$42619 ( \42934 , \42932 , \42933 );
xnor \U$42620 ( \42935 , \42934 , \22267 );
and \U$42621 ( \42936 , \22635 , \22278 );
and \U$42622 ( \42937 , \22646 , \22276 );
nor \U$42623 ( \42938 , \42936 , \42937 );
xnor \U$42624 ( \42939 , \42938 , \22288 );
xor \U$42625 ( \42940 , \42935 , \42939 );
and \U$42626 ( \42941 , \22665 , \22300 );
and \U$42627 ( \42942 , \22676 , \22298 );
nor \U$42628 ( \42943 , \42941 , \42942 );
xnor \U$42629 ( \42944 , \42943 , \22310 );
xor \U$42630 ( \42945 , \42940 , \42944 );
xor \U$42631 ( \42946 , \42931 , \42945 );
xor \U$42632 ( \42947 , \42919 , \42946 );
and \U$42633 ( \42948 , \42786 , \42790 );
and \U$42634 ( \42949 , \42790 , \42795 );
and \U$42635 ( \42950 , \42786 , \42795 );
or \U$42636 ( \42951 , \42948 , \42949 , \42950 );
and \U$42637 ( \42952 , \42772 , \42776 );
and \U$42638 ( \42953 , \42776 , \42781 );
and \U$42639 ( \42954 , \42772 , \42781 );
or \U$42640 ( \42955 , \42952 , \42953 , \42954 );
xor \U$42641 ( \42956 , \42951 , \42955 );
and \U$42642 ( \42957 , \42820 , \42824 );
and \U$42643 ( \42958 , \42824 , \42829 );
and \U$42644 ( \42959 , \42820 , \42829 );
or \U$42645 ( \42960 , \42957 , \42958 , \42959 );
xor \U$42646 ( \42961 , \42956 , \42960 );
xor \U$42647 ( \42962 , \42947 , \42961 );
xor \U$42648 ( \42963 , \42879 , \42962 );
xor \U$42649 ( \42964 , \42870 , \42963 );
and \U$42650 ( \42965 , \42747 , \42758 );
and \U$42651 ( \42966 , \42758 , \42848 );
and \U$42652 ( \42967 , \42747 , \42848 );
or \U$42653 ( \42968 , \42965 , \42966 , \42967 );
nor \U$42654 ( \42969 , \42964 , \42968 );
nor \U$42655 ( \42970 , \42854 , \42969 );
and \U$42656 ( \42971 , \42874 , \42878 );
and \U$42657 ( \42972 , \42878 , \42962 );
and \U$42658 ( \42973 , \42874 , \42962 );
or \U$42659 ( \42974 , \42971 , \42972 , \42973 );
xor \U$42660 ( \42975 , \36415 , \36419 );
xor \U$42661 ( \42976 , \42975 , \36424 );
xor \U$42662 ( \42977 , \36467 , \36471 );
xor \U$42663 ( \42978 , \42977 , \36476 );
xor \U$42664 ( \42979 , \36448 , \36452 );
xor \U$42665 ( \42980 , \42979 , \36457 );
xor \U$42666 ( \42981 , \42978 , \42980 );
xor \U$42667 ( \42982 , \36431 , \36435 );
xor \U$42668 ( \42983 , \42982 , \36440 );
xor \U$42669 ( \42984 , \42981 , \42983 );
xor \U$42670 ( \42985 , \42976 , \42984 );
and \U$42671 ( \42986 , \42935 , \42939 );
and \U$42672 ( \42987 , \42939 , \42944 );
and \U$42673 ( \42988 , \42935 , \42944 );
or \U$42674 ( \42989 , \42986 , \42987 , \42988 );
and \U$42675 ( \42990 , \42927 , \42929 );
xor \U$42676 ( \42991 , \42989 , \42990 );
and \U$42677 ( \42992 , \22706 , \22345 );
and \U$42678 ( \42993 , \22686 , \22343 );
nor \U$42679 ( \42994 , \42992 , \42993 );
xnor \U$42680 ( \42995 , \42994 , \22355 );
xor \U$42681 ( \42996 , \42991 , \42995 );
xor \U$42682 ( \42997 , \42985 , \42996 );
and \U$42683 ( \42998 , \42951 , \42955 );
and \U$42684 ( \42999 , \42955 , \42960 );
and \U$42685 ( \43000 , \42951 , \42960 );
or \U$42686 ( \43001 , \42998 , \42999 , \43000 );
and \U$42687 ( \43002 , \42923 , \42930 );
and \U$42688 ( \43003 , \42930 , \42945 );
and \U$42689 ( \43004 , \42923 , \42945 );
or \U$42690 ( \43005 , \43002 , \43003 , \43004 );
xor \U$42691 ( \43006 , \43001 , \43005 );
and \U$42692 ( \43007 , \42893 , \42907 );
and \U$42693 ( \43008 , \42907 , \42918 );
and \U$42694 ( \43009 , \42893 , \42918 );
or \U$42695 ( \43010 , \43007 , \43008 , \43009 );
xor \U$42696 ( \43011 , \43006 , \43010 );
xor \U$42697 ( \43012 , \42997 , \43011 );
xor \U$42698 ( \43013 , \42974 , \43012 );
and \U$42699 ( \43014 , \42862 , \42866 );
and \U$42700 ( \43015 , \42866 , \42868 );
and \U$42701 ( \43016 , \42862 , \42868 );
or \U$42702 ( \43017 , \43014 , \43015 , \43016 );
and \U$42703 ( \43018 , \42919 , \42946 );
and \U$42704 ( \43019 , \42946 , \42961 );
and \U$42705 ( \43020 , \42919 , \42961 );
or \U$42706 ( \43021 , \43018 , \43019 , \43020 );
xor \U$42707 ( \43022 , \43017 , \43021 );
and \U$42708 ( \43023 , \22355 , \42912 );
and \U$42709 ( \43024 , \42912 , \42917 );
and \U$42710 ( \43025 , \22355 , \42917 );
or \U$42711 ( \43026 , \43023 , \43024 , \43025 );
and \U$42712 ( \43027 , \42897 , \42901 );
and \U$42713 ( \43028 , \42901 , \42906 );
and \U$42714 ( \43029 , \42897 , \42906 );
or \U$42715 ( \43030 , \43027 , \43028 , \43029 );
xor \U$42716 ( \43031 , \43026 , \43030 );
and \U$42717 ( \43032 , \42883 , \42887 );
and \U$42718 ( \43033 , \42887 , \42892 );
and \U$42719 ( \43034 , \42883 , \42892 );
or \U$42720 ( \43035 , \43032 , \43033 , \43034 );
xor \U$42721 ( \43036 , \43031 , \43035 );
xor \U$42722 ( \43037 , \43022 , \43036 );
xor \U$42723 ( \43038 , \43013 , \43037 );
and \U$42724 ( \43039 , \42858 , \42869 );
and \U$42725 ( \43040 , \42869 , \42963 );
and \U$42726 ( \43041 , \42858 , \42963 );
or \U$42727 ( \43042 , \43039 , \43040 , \43041 );
nor \U$42728 ( \43043 , \43038 , \43042 );
and \U$42729 ( \43044 , \43001 , \43005 );
and \U$42730 ( \43045 , \43005 , \43010 );
and \U$42731 ( \43046 , \43001 , \43010 );
or \U$42732 ( \43047 , \43044 , \43045 , \43046 );
and \U$42733 ( \43048 , \42976 , \42984 );
and \U$42734 ( \43049 , \42984 , \42996 );
and \U$42735 ( \43050 , \42976 , \42996 );
or \U$42736 ( \43051 , \43048 , \43049 , \43050 );
xor \U$42737 ( \43052 , \43047 , \43051 );
xor \U$42738 ( \43053 , \36490 , \36492 );
xor \U$42739 ( \43054 , \43053 , \36495 );
xor \U$42740 ( \43055 , \36479 , \36481 );
xor \U$42741 ( \43056 , \43055 , \36484 );
xor \U$42742 ( \43057 , \43054 , \43056 );
xor \U$42743 ( \43058 , \36427 , \36443 );
xor \U$42744 ( \43059 , \43058 , \36460 );
xor \U$42745 ( \43060 , \43057 , \43059 );
xor \U$42746 ( \43061 , \43052 , \43060 );
and \U$42747 ( \43062 , \43017 , \43021 );
and \U$42748 ( \43063 , \43021 , \43036 );
and \U$42749 ( \43064 , \43017 , \43036 );
or \U$42750 ( \43065 , \43062 , \43063 , \43064 );
and \U$42751 ( \43066 , \42997 , \43011 );
xor \U$42752 ( \43067 , \43065 , \43066 );
and \U$42753 ( \43068 , \43026 , \43030 );
and \U$42754 ( \43069 , \43030 , \43035 );
and \U$42755 ( \43070 , \43026 , \43035 );
or \U$42756 ( \43071 , \43068 , \43069 , \43070 );
and \U$42757 ( \43072 , \42989 , \42990 );
and \U$42758 ( \43073 , \42990 , \42995 );
and \U$42759 ( \43074 , \42989 , \42995 );
or \U$42760 ( \43075 , \43072 , \43073 , \43074 );
xor \U$42761 ( \43076 , \43071 , \43075 );
and \U$42762 ( \43077 , \42978 , \42980 );
and \U$42763 ( \43078 , \42980 , \42983 );
and \U$42764 ( \43079 , \42978 , \42983 );
or \U$42765 ( \43080 , \43077 , \43078 , \43079 );
xor \U$42766 ( \43081 , \43076 , \43080 );
xor \U$42767 ( \43082 , \43067 , \43081 );
xor \U$42768 ( \43083 , \43061 , \43082 );
and \U$42769 ( \43084 , \42974 , \43012 );
and \U$42770 ( \43085 , \43012 , \43037 );
and \U$42771 ( \43086 , \42974 , \43037 );
or \U$42772 ( \43087 , \43084 , \43085 , \43086 );
nor \U$42773 ( \43088 , \43083 , \43087 );
nor \U$42774 ( \43089 , \43043 , \43088 );
nand \U$42775 ( \43090 , \42970 , \43089 );
and \U$42776 ( \43091 , \43065 , \43066 );
and \U$42777 ( \43092 , \43066 , \43081 );
and \U$42778 ( \43093 , \43065 , \43081 );
or \U$42779 ( \43094 , \43091 , \43092 , \43093 );
and \U$42780 ( \43095 , \43047 , \43051 );
and \U$42781 ( \43096 , \43051 , \43060 );
and \U$42782 ( \43097 , \43047 , \43060 );
or \U$42783 ( \43098 , \43095 , \43096 , \43097 );
xor \U$42784 ( \43099 , \35792 , \35808 );
xor \U$42785 ( \43100 , \43099 , \35825 );
xor \U$42786 ( \43101 , \36503 , \36505 );
xor \U$42787 ( \43102 , \43101 , \36508 );
xor \U$42788 ( \43103 , \43100 , \43102 );
xor \U$42789 ( \43104 , \36463 , \36487 );
xor \U$42790 ( \43105 , \43104 , \36498 );
xor \U$42791 ( \43106 , \43103 , \43105 );
xor \U$42792 ( \43107 , \43098 , \43106 );
and \U$42793 ( \43108 , \43071 , \43075 );
and \U$42794 ( \43109 , \43075 , \43080 );
and \U$42795 ( \43110 , \43071 , \43080 );
or \U$42796 ( \43111 , \43108 , \43109 , \43110 );
and \U$42797 ( \43112 , \43054 , \43056 );
and \U$42798 ( \43113 , \43056 , \43059 );
and \U$42799 ( \43114 , \43054 , \43059 );
or \U$42800 ( \43115 , \43112 , \43113 , \43114 );
xor \U$42801 ( \43116 , \43111 , \43115 );
xor \U$42802 ( \43117 , \35844 , \35858 );
xor \U$42803 ( \43118 , \43117 , \35863 );
xor \U$42804 ( \43119 , \43116 , \43118 );
xor \U$42805 ( \43120 , \43107 , \43119 );
xor \U$42806 ( \43121 , \43094 , \43120 );
and \U$42807 ( \43122 , \43061 , \43082 );
nor \U$42808 ( \43123 , \43121 , \43122 );
and \U$42809 ( \43124 , \43098 , \43106 );
and \U$42810 ( \43125 , \43106 , \43119 );
and \U$42811 ( \43126 , \43098 , \43119 );
or \U$42812 ( \43127 , \43124 , \43125 , \43126 );
xor \U$42813 ( \43128 , \35828 , \35866 );
xor \U$42814 ( \43129 , \43128 , \35903 );
xor \U$42815 ( \43130 , \36501 , \36511 );
xor \U$42816 ( \43131 , \43130 , \36514 );
xor \U$42817 ( \43132 , \43129 , \43131 );
xor \U$42818 ( \43133 , \43127 , \43132 );
and \U$42819 ( \43134 , \43111 , \43115 );
and \U$42820 ( \43135 , \43115 , \43118 );
and \U$42821 ( \43136 , \43111 , \43118 );
or \U$42822 ( \43137 , \43134 , \43135 , \43136 );
and \U$42823 ( \43138 , \43100 , \43102 );
and \U$42824 ( \43139 , \43102 , \43105 );
and \U$42825 ( \43140 , \43100 , \43105 );
or \U$42826 ( \43141 , \43138 , \43139 , \43140 );
xor \U$42827 ( \43142 , \43137 , \43141 );
xor \U$42828 ( \43143 , \35916 , \35960 );
xor \U$42829 ( \43144 , \43143 , \35983 );
xor \U$42830 ( \43145 , \43142 , \43144 );
xor \U$42831 ( \43146 , \43133 , \43145 );
and \U$42832 ( \43147 , \43094 , \43120 );
nor \U$42833 ( \43148 , \43146 , \43147 );
nor \U$42834 ( \43149 , \43123 , \43148 );
and \U$42835 ( \43150 , \43137 , \43141 );
and \U$42836 ( \43151 , \43141 , \43144 );
and \U$42837 ( \43152 , \43137 , \43144 );
or \U$42838 ( \43153 , \43150 , \43151 , \43152 );
and \U$42839 ( \43154 , \43129 , \43131 );
xor \U$42840 ( \43155 , \43153 , \43154 );
xor \U$42841 ( \43156 , \36517 , \36518 );
xor \U$42842 ( \43157 , \43156 , \36521 );
xor \U$42843 ( \43158 , \43155 , \43157 );
and \U$42844 ( \43159 , \43127 , \43132 );
and \U$42845 ( \43160 , \43132 , \43145 );
and \U$42846 ( \43161 , \43127 , \43145 );
or \U$42847 ( \43162 , \43159 , \43160 , \43161 );
nor \U$42848 ( \43163 , \43158 , \43162 );
xor \U$42849 ( \43164 , \36524 , \36525 );
xor \U$42850 ( \43165 , \43164 , \36528 );
and \U$42851 ( \43166 , \43153 , \43154 );
and \U$42852 ( \43167 , \43154 , \43157 );
and \U$42853 ( \43168 , \43153 , \43157 );
or \U$42854 ( \43169 , \43166 , \43167 , \43168 );
nor \U$42855 ( \43170 , \43165 , \43169 );
nor \U$42856 ( \43171 , \43163 , \43170 );
nand \U$42857 ( \43172 , \43149 , \43171 );
nor \U$42858 ( \43173 , \43090 , \43172 );
nand \U$42859 ( \43174 , \42743 , \43173 );
and \U$42860 ( \43175 , \22646 , \22076 );
and \U$42861 ( \43176 , \22613 , \22073 );
nor \U$42862 ( \43177 , \43175 , \43176 );
xnor \U$42863 ( \43178 , \43177 , \22072 );
and \U$42864 ( \43179 , \22676 , \22095 );
and \U$42865 ( \43180 , \22635 , \22093 );
nor \U$42866 ( \43181 , \43179 , \43180 );
xnor \U$42867 ( \43182 , \43181 , \22105 );
xor \U$42868 ( \43183 , \43178 , \43182 );
and \U$42869 ( \43184 , \22696 , \22119 );
and \U$42870 ( \43185 , \22665 , \22117 );
nor \U$42871 ( \43186 , \43184 , \43185 );
xnor \U$42872 ( \43187 , \43186 , \22129 );
xor \U$42873 ( \43188 , \43183 , \43187 );
and \U$42874 ( \43189 , \22635 , \22076 );
and \U$42875 ( \43190 , \22646 , \22073 );
nor \U$42876 ( \43191 , \43189 , \43190 );
xnor \U$42877 ( \43192 , \43191 , \22072 );
and \U$42878 ( \43193 , \22150 , \43192 );
and \U$42879 ( \43194 , \22665 , \22095 );
and \U$42880 ( \43195 , \22676 , \22093 );
nor \U$42881 ( \43196 , \43194 , \43195 );
xnor \U$42882 ( \43197 , \43196 , \22105 );
and \U$42883 ( \43198 , \43192 , \43197 );
and \U$42884 ( \43199 , \22150 , \43197 );
or \U$42885 ( \43200 , \43193 , \43198 , \43199 );
and \U$42886 ( \43201 , \22686 , \22119 );
and \U$42887 ( \43202 , \22696 , \22117 );
nor \U$42888 ( \43203 , \43201 , \43202 );
xnor \U$42889 ( \43204 , \43203 , \22129 );
nand \U$42890 ( \43205 , \22706 , \22138 );
xnor \U$42891 ( \43206 , \43205 , \22150 );
and \U$42892 ( \43207 , \43204 , \43206 );
xor \U$42893 ( \43208 , \43200 , \43207 );
and \U$42894 ( \43209 , \22706 , \22140 );
and \U$42895 ( \43210 , \22686 , \22138 );
nor \U$42896 ( \43211 , \43209 , \43210 );
xnor \U$42897 ( \43212 , \43211 , \22150 );
xor \U$42898 ( \43213 , \43208 , \43212 );
xor \U$42899 ( \43214 , \43188 , \43213 );
and \U$42900 ( \43215 , \22676 , \22076 );
and \U$42901 ( \43216 , \22635 , \22073 );
nor \U$42902 ( \43217 , \43215 , \43216 );
xnor \U$42903 ( \43218 , \43217 , \22072 );
and \U$42904 ( \43219 , \22696 , \22095 );
and \U$42905 ( \43220 , \22665 , \22093 );
nor \U$42906 ( \43221 , \43219 , \43220 );
xnor \U$42907 ( \43222 , \43221 , \22105 );
and \U$42908 ( \43223 , \43218 , \43222 );
and \U$42909 ( \43224 , \22706 , \22119 );
and \U$42910 ( \43225 , \22686 , \22117 );
nor \U$42911 ( \43226 , \43224 , \43225 );
xnor \U$42912 ( \43227 , \43226 , \22129 );
and \U$42913 ( \43228 , \43222 , \43227 );
and \U$42914 ( \43229 , \43218 , \43227 );
or \U$42915 ( \43230 , \43223 , \43228 , \43229 );
xor \U$42916 ( \43231 , \43204 , \43206 );
and \U$42917 ( \43232 , \43230 , \43231 );
xor \U$42918 ( \43233 , \22150 , \43192 );
xor \U$42919 ( \43234 , \43233 , \43197 );
and \U$42920 ( \43235 , \43231 , \43234 );
and \U$42921 ( \43236 , \43230 , \43234 );
or \U$42922 ( \43237 , \43232 , \43235 , \43236 );
nor \U$42923 ( \43238 , \43214 , \43237 );
and \U$42924 ( \43239 , \43200 , \43207 );
and \U$42925 ( \43240 , \43207 , \43212 );
and \U$42926 ( \43241 , \43200 , \43212 );
or \U$42927 ( \43242 , \43239 , \43240 , \43241 );
and \U$42928 ( \43243 , \43178 , \43182 );
and \U$42929 ( \43244 , \43182 , \43187 );
and \U$42930 ( \43245 , \43178 , \43187 );
or \U$42931 ( \43246 , \43243 , \43244 , \43245 );
and \U$42932 ( \43247 , \22665 , \22119 );
and \U$42933 ( \43248 , \22676 , \22117 );
nor \U$42934 ( \43249 , \43247 , \43248 );
xnor \U$42935 ( \43250 , \43249 , \22129 );
and \U$42936 ( \43251 , \22686 , \22140 );
and \U$42937 ( \43252 , \22696 , \22138 );
nor \U$42938 ( \43253 , \43251 , \43252 );
xnor \U$42939 ( \43254 , \43253 , \22150 );
xor \U$42940 ( \43255 , \43250 , \43254 );
nand \U$42941 ( \43256 , \22706 , \22160 );
xnor \U$42942 ( \43257 , \43256 , \22172 );
xor \U$42943 ( \43258 , \43255 , \43257 );
xor \U$42944 ( \43259 , \43246 , \43258 );
and \U$42945 ( \43260 , \22613 , \22076 );
and \U$42946 ( \43261 , \22624 , \22073 );
nor \U$42947 ( \43262 , \43260 , \43261 );
xnor \U$42948 ( \43263 , \43262 , \22072 );
xor \U$42949 ( \43264 , \22172 , \43263 );
and \U$42950 ( \43265 , \22635 , \22095 );
and \U$42951 ( \43266 , \22646 , \22093 );
nor \U$42952 ( \43267 , \43265 , \43266 );
xnor \U$42953 ( \43268 , \43267 , \22105 );
xor \U$42954 ( \43269 , \43264 , \43268 );
xor \U$42955 ( \43270 , \43259 , \43269 );
xor \U$42956 ( \43271 , \43242 , \43270 );
and \U$42957 ( \43272 , \43188 , \43213 );
nor \U$42958 ( \43273 , \43271 , \43272 );
nor \U$42959 ( \43274 , \43238 , \43273 );
and \U$42960 ( \43275 , \43246 , \43258 );
and \U$42961 ( \43276 , \43258 , \43269 );
and \U$42962 ( \43277 , \43246 , \43269 );
or \U$42963 ( \43278 , \43275 , \43276 , \43277 );
and \U$42964 ( \43279 , \22706 , \22162 );
and \U$42965 ( \43280 , \22686 , \22160 );
nor \U$42966 ( \43281 , \43279 , \43280 );
xnor \U$42967 ( \43282 , \43281 , \22172 );
and \U$42968 ( \43283 , \22624 , \22076 );
and \U$42969 ( \43284 , \22592 , \22073 );
nor \U$42970 ( \43285 , \43283 , \43284 );
xnor \U$42971 ( \43286 , \43285 , \22072 );
and \U$42972 ( \43287 , \22646 , \22095 );
and \U$42973 ( \43288 , \22613 , \22093 );
nor \U$42974 ( \43289 , \43287 , \43288 );
xnor \U$42975 ( \43290 , \43289 , \22105 );
xor \U$42976 ( \43291 , \43286 , \43290 );
and \U$42977 ( \43292 , \22676 , \22119 );
and \U$42978 ( \43293 , \22635 , \22117 );
nor \U$42979 ( \43294 , \43292 , \43293 );
xnor \U$42980 ( \43295 , \43294 , \22129 );
xor \U$42981 ( \43296 , \43291 , \43295 );
xor \U$42982 ( \43297 , \43282 , \43296 );
xor \U$42983 ( \43298 , \43278 , \43297 );
and \U$42984 ( \43299 , \22172 , \43263 );
and \U$42985 ( \43300 , \43263 , \43268 );
and \U$42986 ( \43301 , \22172 , \43268 );
or \U$42987 ( \43302 , \43299 , \43300 , \43301 );
and \U$42988 ( \43303 , \43250 , \43254 );
and \U$42989 ( \43304 , \43254 , \43257 );
and \U$42990 ( \43305 , \43250 , \43257 );
or \U$42991 ( \43306 , \43303 , \43304 , \43305 );
xor \U$42992 ( \43307 , \43302 , \43306 );
and \U$42993 ( \43308 , \22696 , \22140 );
and \U$42994 ( \43309 , \22665 , \22138 );
nor \U$42995 ( \43310 , \43308 , \43309 );
xnor \U$42996 ( \43311 , \43310 , \22150 );
xor \U$42997 ( \43312 , \43307 , \43311 );
xor \U$42998 ( \43313 , \43298 , \43312 );
and \U$42999 ( \43314 , \43242 , \43270 );
nor \U$43000 ( \43315 , \43313 , \43314 );
and \U$43001 ( \43316 , \43286 , \43290 );
and \U$43002 ( \43317 , \43290 , \43295 );
and \U$43003 ( \43318 , \43286 , \43295 );
or \U$43004 ( \43319 , \43316 , \43317 , \43318 );
nand \U$43005 ( \43320 , \22706 , \22185 );
xnor \U$43006 ( \43321 , \43320 , \22197 );
xor \U$43007 ( \43322 , \43319 , \43321 );
and \U$43008 ( \43323 , \22635 , \22119 );
and \U$43009 ( \43324 , \22646 , \22117 );
nor \U$43010 ( \43325 , \43323 , \43324 );
xnor \U$43011 ( \43326 , \43325 , \22129 );
and \U$43012 ( \43327 , \22665 , \22140 );
and \U$43013 ( \43328 , \22676 , \22138 );
nor \U$43014 ( \43329 , \43327 , \43328 );
xnor \U$43015 ( \43330 , \43329 , \22150 );
xor \U$43016 ( \43331 , \43326 , \43330 );
and \U$43017 ( \43332 , \22686 , \22162 );
and \U$43018 ( \43333 , \22696 , \22160 );
nor \U$43019 ( \43334 , \43332 , \43333 );
xnor \U$43020 ( \43335 , \43334 , \22172 );
xor \U$43021 ( \43336 , \43331 , \43335 );
xor \U$43022 ( \43337 , \43322 , \43336 );
and \U$43023 ( \43338 , \43302 , \43306 );
and \U$43024 ( \43339 , \43306 , \43311 );
and \U$43025 ( \43340 , \43302 , \43311 );
or \U$43026 ( \43341 , \43338 , \43339 , \43340 );
and \U$43027 ( \43342 , \43282 , \43296 );
xor \U$43028 ( \43343 , \43341 , \43342 );
and \U$43029 ( \43344 , \22592 , \22076 );
and \U$43030 ( \43345 , \22603 , \22073 );
nor \U$43031 ( \43346 , \43344 , \43345 );
xnor \U$43032 ( \43347 , \43346 , \22072 );
xor \U$43033 ( \43348 , \22197 , \43347 );
and \U$43034 ( \43349 , \22613 , \22095 );
and \U$43035 ( \43350 , \22624 , \22093 );
nor \U$43036 ( \43351 , \43349 , \43350 );
xnor \U$43037 ( \43352 , \43351 , \22105 );
xor \U$43038 ( \43353 , \43348 , \43352 );
xor \U$43039 ( \43354 , \43343 , \43353 );
xor \U$43040 ( \43355 , \43337 , \43354 );
and \U$43041 ( \43356 , \43278 , \43297 );
and \U$43042 ( \43357 , \43297 , \43312 );
and \U$43043 ( \43358 , \43278 , \43312 );
or \U$43044 ( \43359 , \43356 , \43357 , \43358 );
nor \U$43045 ( \43360 , \43355 , \43359 );
nor \U$43046 ( \43361 , \43315 , \43360 );
nand \U$43047 ( \43362 , \43274 , \43361 );
and \U$43048 ( \43363 , \43341 , \43342 );
and \U$43049 ( \43364 , \43342 , \43353 );
and \U$43050 ( \43365 , \43341 , \43353 );
or \U$43051 ( \43366 , \43363 , \43364 , \43365 );
and \U$43052 ( \43367 , \43319 , \43321 );
and \U$43053 ( \43368 , \43321 , \43336 );
and \U$43054 ( \43369 , \43319 , \43336 );
or \U$43055 ( \43370 , \43367 , \43368 , \43369 );
xor \U$43056 ( \43371 , \42039 , \42043 );
xor \U$43057 ( \43372 , \43371 , \42048 );
xor \U$43058 ( \43373 , \43370 , \43372 );
and \U$43059 ( \43374 , \22197 , \43347 );
and \U$43060 ( \43375 , \43347 , \43352 );
and \U$43061 ( \43376 , \22197 , \43352 );
or \U$43062 ( \43377 , \43374 , \43375 , \43376 );
and \U$43063 ( \43378 , \43326 , \43330 );
and \U$43064 ( \43379 , \43330 , \43335 );
and \U$43065 ( \43380 , \43326 , \43335 );
or \U$43066 ( \43381 , \43378 , \43379 , \43380 );
xor \U$43067 ( \43382 , \43377 , \43381 );
xor \U$43068 ( \43383 , \42055 , \42059 );
xor \U$43069 ( \43384 , \43383 , \42064 );
xor \U$43070 ( \43385 , \43382 , \43384 );
xor \U$43071 ( \43386 , \43373 , \43385 );
xor \U$43072 ( \43387 , \43366 , \43386 );
and \U$43073 ( \43388 , \43337 , \43354 );
nor \U$43074 ( \43389 , \43387 , \43388 );
and \U$43075 ( \43390 , \43370 , \43372 );
and \U$43076 ( \43391 , \43372 , \43385 );
and \U$43077 ( \43392 , \43370 , \43385 );
or \U$43078 ( \43393 , \43390 , \43391 , \43392 );
and \U$43079 ( \43394 , \43377 , \43381 );
and \U$43080 ( \43395 , \43381 , \43384 );
and \U$43081 ( \43396 , \43377 , \43384 );
or \U$43082 ( \43397 , \43394 , \43395 , \43396 );
xor \U$43083 ( \43398 , \42077 , \42079 );
xor \U$43084 ( \43399 , \43398 , \42082 );
xor \U$43085 ( \43400 , \43397 , \43399 );
xor \U$43086 ( \43401 , \42051 , \42067 );
xor \U$43087 ( \43402 , \43401 , \42072 );
xor \U$43088 ( \43403 , \43400 , \43402 );
xor \U$43089 ( \43404 , \43393 , \43403 );
and \U$43090 ( \43405 , \43366 , \43386 );
nor \U$43091 ( \43406 , \43404 , \43405 );
nor \U$43092 ( \43407 , \43389 , \43406 );
and \U$43093 ( \43408 , \43397 , \43399 );
and \U$43094 ( \43409 , \43399 , \43402 );
and \U$43095 ( \43410 , \43397 , \43402 );
or \U$43096 ( \43411 , \43408 , \43409 , \43410 );
xor \U$43097 ( \43412 , \42093 , \42095 );
xor \U$43098 ( \43413 , \43411 , \43412 );
xor \U$43099 ( \43414 , \42075 , \42085 );
xor \U$43100 ( \43415 , \43414 , \42088 );
xor \U$43101 ( \43416 , \43413 , \43415 );
and \U$43102 ( \43417 , \43393 , \43403 );
nor \U$43103 ( \43418 , \43416 , \43417 );
xor \U$43104 ( \43419 , \42091 , \42096 );
xor \U$43105 ( \43420 , \43419 , \42099 );
and \U$43106 ( \43421 , \43411 , \43412 );
and \U$43107 ( \43422 , \43412 , \43415 );
and \U$43108 ( \43423 , \43411 , \43415 );
or \U$43109 ( \43424 , \43421 , \43422 , \43423 );
nor \U$43110 ( \43425 , \43420 , \43424 );
nor \U$43111 ( \43426 , \43418 , \43425 );
nand \U$43112 ( \43427 , \43407 , \43426 );
nor \U$43113 ( \43428 , \43362 , \43427 );
and \U$43114 ( \43429 , \22696 , \22076 );
and \U$43115 ( \43430 , \22665 , \22073 );
nor \U$43116 ( \43431 , \43429 , \43430 );
xnor \U$43117 ( \43432 , \43431 , \22072 );
and \U$43118 ( \43433 , \22706 , \22095 );
and \U$43119 ( \43434 , \22686 , \22093 );
nor \U$43120 ( \43435 , \43433 , \43434 );
xnor \U$43121 ( \43436 , \43435 , \22105 );
xor \U$43122 ( \43437 , \43432 , \43436 );
and \U$43123 ( \43438 , \22686 , \22076 );
and \U$43124 ( \43439 , \22696 , \22073 );
nor \U$43125 ( \43440 , \43438 , \43439 );
xnor \U$43126 ( \43441 , \43440 , \22072 );
and \U$43127 ( \43442 , \43441 , \22105 );
nor \U$43128 ( \43443 , \43437 , \43442 );
nand \U$43129 ( \43444 , \22706 , \22117 );
xnor \U$43130 ( \43445 , \43444 , \22129 );
and \U$43131 ( \43446 , \22665 , \22076 );
and \U$43132 ( \43447 , \22676 , \22073 );
nor \U$43133 ( \43448 , \43446 , \43447 );
xnor \U$43134 ( \43449 , \43448 , \22072 );
xor \U$43135 ( \43450 , \22129 , \43449 );
and \U$43136 ( \43451 , \22686 , \22095 );
and \U$43137 ( \43452 , \22696 , \22093 );
nor \U$43138 ( \43453 , \43451 , \43452 );
xnor \U$43139 ( \43454 , \43453 , \22105 );
xor \U$43140 ( \43455 , \43450 , \43454 );
xor \U$43141 ( \43456 , \43445 , \43455 );
and \U$43142 ( \43457 , \43432 , \43436 );
nor \U$43143 ( \43458 , \43456 , \43457 );
nor \U$43144 ( \43459 , \43443 , \43458 );
and \U$43145 ( \43460 , \22129 , \43449 );
and \U$43146 ( \43461 , \43449 , \43454 );
and \U$43147 ( \43462 , \22129 , \43454 );
or \U$43148 ( \43463 , \43460 , \43461 , \43462 );
xor \U$43149 ( \43464 , \43218 , \43222 );
xor \U$43150 ( \43465 , \43464 , \43227 );
xor \U$43151 ( \43466 , \43463 , \43465 );
and \U$43152 ( \43467 , \43445 , \43455 );
nor \U$43153 ( \43468 , \43466 , \43467 );
xor \U$43154 ( \43469 , \43230 , \43231 );
xor \U$43155 ( \43470 , \43469 , \43234 );
and \U$43156 ( \43471 , \43463 , \43465 );
nor \U$43157 ( \43472 , \43470 , \43471 );
nor \U$43158 ( \43473 , \43468 , \43472 );
nand \U$43159 ( \43474 , \43459 , \43473 );
xor \U$43160 ( \43475 , \43441 , \22105 );
nand \U$43161 ( \43476 , \22706 , \22093 );
xnor \U$43162 ( \43477 , \43476 , \22105 );
nor \U$43163 ( \43478 , \43475 , \43477 );
and \U$43164 ( \43479 , \22706 , \22076 );
and \U$43165 ( \43480 , \22686 , \22073 );
nor \U$43166 ( \43481 , \43479 , \43480 );
xnor \U$43167 ( \43482 , \43481 , \22072 );
nand \U$43168 ( \43483 , \22706 , \22073 );
xnor \U$43169 ( \43484 , \43483 , \22072 );
and \U$43170 ( \43485 , \43484 , \22072 );
nand \U$43171 ( \43486 , \43482 , \43485 );
or \U$43172 ( \43487 , \43478 , \43486 );
nand \U$43173 ( \43488 , \43475 , \43477 );
nand \U$43174 ( \43489 , \43487 , \43488 );
not \U$43175 ( \43490 , \43489 );
or \U$43176 ( \43491 , \43474 , \43490 );
nand \U$43177 ( \43492 , \43437 , \43442 );
or \U$43178 ( \43493 , \43458 , \43492 );
nand \U$43179 ( \43494 , \43456 , \43457 );
nand \U$43180 ( \43495 , \43493 , \43494 );
and \U$43181 ( \43496 , \43473 , \43495 );
nand \U$43182 ( \43497 , \43466 , \43467 );
or \U$43183 ( \43498 , \43472 , \43497 );
nand \U$43184 ( \43499 , \43470 , \43471 );
nand \U$43185 ( \43500 , \43498 , \43499 );
nor \U$43186 ( \43501 , \43496 , \43500 );
nand \U$43187 ( \43502 , \43491 , \43501 );
and \U$43188 ( \43503 , \43428 , \43502 );
nand \U$43189 ( \43504 , \43214 , \43237 );
or \U$43190 ( \43505 , \43273 , \43504 );
nand \U$43191 ( \43506 , \43271 , \43272 );
nand \U$43192 ( \43507 , \43505 , \43506 );
and \U$43193 ( \43508 , \43361 , \43507 );
nand \U$43194 ( \43509 , \43313 , \43314 );
or \U$43195 ( \43510 , \43360 , \43509 );
nand \U$43196 ( \43511 , \43355 , \43359 );
nand \U$43197 ( \43512 , \43510 , \43511 );
nor \U$43198 ( \43513 , \43508 , \43512 );
or \U$43199 ( \43514 , \43427 , \43513 );
nand \U$43200 ( \43515 , \43387 , \43388 );
or \U$43201 ( \43516 , \43406 , \43515 );
nand \U$43202 ( \43517 , \43404 , \43405 );
nand \U$43203 ( \43518 , \43516 , \43517 );
and \U$43204 ( \43519 , \43426 , \43518 );
nand \U$43205 ( \43520 , \43416 , \43417 );
or \U$43206 ( \43521 , \43425 , \43520 );
nand \U$43207 ( \43522 , \43420 , \43424 );
nand \U$43208 ( \43523 , \43521 , \43522 );
nor \U$43209 ( \43524 , \43519 , \43523 );
nand \U$43210 ( \43525 , \43514 , \43524 );
nor \U$43211 ( \43526 , \43503 , \43525 );
or \U$43212 ( \43527 , \43174 , \43526 );
nand \U$43213 ( \43528 , \42035 , \42102 );
or \U$43214 ( \43529 , \42178 , \43528 );
nand \U$43215 ( \43530 , \42173 , \42177 );
nand \U$43216 ( \43531 , \43529 , \43530 );
and \U$43217 ( \43532 , \42346 , \43531 );
nand \U$43218 ( \43533 , \42255 , \42259 );
or \U$43219 ( \43534 , \42345 , \43533 );
nand \U$43220 ( \43535 , \42343 , \42344 );
nand \U$43221 ( \43536 , \43534 , \43535 );
nor \U$43222 ( \43537 , \43532 , \43536 );
or \U$43223 ( \43538 , \42742 , \43537 );
nand \U$43224 ( \43539 , \42436 , \42437 );
or \U$43225 ( \43540 , \42533 , \43539 );
nand \U$43226 ( \43541 , \42528 , \42532 );
nand \U$43227 ( \43542 , \43540 , \43541 );
and \U$43228 ( \43543 , \42741 , \43542 );
nand \U$43229 ( \43544 , \42630 , \42634 );
or \U$43230 ( \43545 , \42740 , \43544 );
nand \U$43231 ( \43546 , \42735 , \42739 );
nand \U$43232 ( \43547 , \43545 , \43546 );
nor \U$43233 ( \43548 , \43543 , \43547 );
nand \U$43234 ( \43549 , \43538 , \43548 );
and \U$43235 ( \43550 , \43173 , \43549 );
nand \U$43236 ( \43551 , \42849 , \42853 );
or \U$43237 ( \43552 , \42969 , \43551 );
nand \U$43238 ( \43553 , \42964 , \42968 );
nand \U$43239 ( \43554 , \43552 , \43553 );
and \U$43240 ( \43555 , \43089 , \43554 );
nand \U$43241 ( \43556 , \43038 , \43042 );
or \U$43242 ( \43557 , \43088 , \43556 );
nand \U$43243 ( \43558 , \43083 , \43087 );
nand \U$43244 ( \43559 , \43557 , \43558 );
nor \U$43245 ( \43560 , \43555 , \43559 );
or \U$43246 ( \43561 , \43172 , \43560 );
nand \U$43247 ( \43562 , \43121 , \43122 );
or \U$43248 ( \43563 , \43148 , \43562 );
nand \U$43249 ( \43564 , \43146 , \43147 );
nand \U$43250 ( \43565 , \43563 , \43564 );
and \U$43251 ( \43566 , \43171 , \43565 );
nand \U$43252 ( \43567 , \43158 , \43162 );
or \U$43253 ( \43568 , \43170 , \43567 );
nand \U$43254 ( \43569 , \43165 , \43169 );
nand \U$43255 ( \43570 , \43568 , \43569 );
nor \U$43256 ( \43571 , \43566 , \43570 );
nand \U$43257 ( \43572 , \43561 , \43571 );
nor \U$43258 ( \43573 , \43550 , \43572 );
nand \U$43259 ( \43574 , \43527 , \43573 );
and \U$43260 ( \43575 , \41862 , \43574 );
nand \U$43261 ( \43576 , \36411 , \36531 );
or \U$43262 ( \43577 , \36687 , \43576 );
nand \U$43263 ( \43578 , \36682 , \36686 );
nand \U$43264 ( \43579 , \43577 , \43578 );
and \U$43265 ( \43580 , \37015 , \43579 );
nand \U$43266 ( \43581 , \36844 , \36848 );
or \U$43267 ( \43582 , \37014 , \43581 );
nand \U$43268 ( \43583 , \37009 , \37013 );
nand \U$43269 ( \43584 , \43582 , \43583 );
nor \U$43270 ( \43585 , \43580 , \43584 );
or \U$43271 ( \43586 , \37731 , \43585 );
nand \U$43272 ( \43587 , \37182 , \37186 );
or \U$43273 ( \43588 , \37362 , \43587 );
nand \U$43274 ( \43589 , \37357 , \37361 );
nand \U$43275 ( \43590 , \43588 , \43589 );
and \U$43276 ( \43591 , \37730 , \43590 );
nand \U$43277 ( \43592 , \37539 , \37543 );
or \U$43278 ( \43593 , \37729 , \43592 );
nand \U$43279 ( \43594 , \37724 , \37728 );
nand \U$43280 ( \43595 , \43593 , \43594 );
nor \U$43281 ( \43596 , \43591 , \43595 );
nand \U$43282 ( \43597 , \43586 , \43596 );
and \U$43283 ( \43598 , \39405 , \43597 );
nand \U$43284 ( \43599 , \37921 , \37922 );
or \U$43285 ( \43600 , \38118 , \43599 );
nand \U$43286 ( \43601 , \38116 , \38117 );
nand \U$43287 ( \43602 , \43600 , \43601 );
and \U$43288 ( \43603 , \38526 , \43602 );
nand \U$43289 ( \43604 , \38318 , \38319 );
or \U$43290 ( \43605 , \38525 , \43604 );
nand \U$43291 ( \43606 , \38520 , \38524 );
nand \U$43292 ( \43607 , \43605 , \43606 );
nor \U$43293 ( \43608 , \43603 , \43607 );
or \U$43294 ( \43609 , \39404 , \43608 );
nand \U$43295 ( \43610 , \38735 , \38736 );
or \U$43296 ( \43611 , \38955 , \43610 );
nand \U$43297 ( \43612 , \38950 , \38954 );
nand \U$43298 ( \43613 , \43611 , \43612 );
and \U$43299 ( \43614 , \39403 , \43613 );
nand \U$43300 ( \43615 , \39172 , \39176 );
or \U$43301 ( \43616 , \39402 , \43615 );
nand \U$43302 ( \43617 , \39397 , \39401 );
nand \U$43303 ( \43618 , \43616 , \43617 );
nor \U$43304 ( \43619 , \43614 , \43618 );
nand \U$43305 ( \43620 , \43609 , \43619 );
nor \U$43306 ( \43621 , \43598 , \43620 );
or \U$43307 ( \43622 , \41861 , \43621 );
nand \U$43308 ( \43623 , \39632 , \39636 );
or \U$43309 ( \43624 , \39872 , \43623 );
nand \U$43310 ( \43625 , \39867 , \39871 );
nand \U$43311 ( \43626 , \43624 , \43625 );
and \U$43312 ( \43627 , \40360 , \43626 );
nand \U$43313 ( \43628 , \40109 , \40113 );
or \U$43314 ( \43629 , \40359 , \43628 );
nand \U$43315 ( \43630 , \40354 , \40358 );
nand \U$43316 ( \43631 , \43629 , \43630 );
nor \U$43317 ( \43632 , \43627 , \43631 );
or \U$43318 ( \43633 , \41396 , \43632 );
nand \U$43319 ( \43634 , \40607 , \40611 );
or \U$43320 ( \43635 , \40867 , \43634 );
nand \U$43321 ( \43636 , \40862 , \40866 );
nand \U$43322 ( \43637 , \43635 , \43636 );
and \U$43323 ( \43638 , \41395 , \43637 );
nand \U$43324 ( \43639 , \41124 , \41128 );
or \U$43325 ( \43640 , \41394 , \43639 );
nand \U$43326 ( \43641 , \41389 , \41393 );
nand \U$43327 ( \43642 , \43640 , \43641 );
nor \U$43328 ( \43643 , \43638 , \43642 );
nand \U$43329 ( \43644 , \43633 , \43643 );
and \U$43330 ( \43645 , \41860 , \43644 );
nand \U$43331 ( \43646 , \41555 , \41559 );
or \U$43332 ( \43647 , \41667 , \43646 );
nand \U$43333 ( \43648 , \41662 , \41666 );
nand \U$43334 ( \43649 , \43647 , \43648 );
and \U$43335 ( \43650 , \41785 , \43649 );
nand \U$43336 ( \43651 , \41737 , \41738 );
or \U$43337 ( \43652 , \41784 , \43651 );
nand \U$43338 ( \43653 , \41782 , \41783 );
nand \U$43339 ( \43654 , \43652 , \43653 );
nor \U$43340 ( \43655 , \43650 , \43654 );
or \U$43341 ( \43656 , \41859 , \43655 );
nand \U$43342 ( \43657 , \41817 , \41818 );
or \U$43343 ( \43658 , \41841 , \43657 );
nand \U$43344 ( \43659 , \41839 , \41840 );
nand \U$43345 ( \43660 , \43658 , \43659 );
and \U$43346 ( \43661 , \41858 , \43660 );
nand \U$43347 ( \43662 , \41849 , \41853 );
or \U$43348 ( \43663 , \41857 , \43662 );
nand \U$43349 ( \43664 , \41855 , \41856 );
nand \U$43350 ( \43665 , \43663 , \43664 );
nor \U$43351 ( \43666 , \43661 , \43665 );
nand \U$43352 ( \43667 , \43656 , \43666 );
nor \U$43353 ( \43668 , \43645 , \43667 );
nand \U$43354 ( \43669 , \43622 , \43668 );
nor \U$43355 ( \43670 , \43575 , \43669 );
or \U$43356 ( \43671 , \35780 , \43670 );
nand \U$43357 ( \43672 , \24456 , \24723 );
or \U$43358 ( \43673 , \25038 , \43672 );
nand \U$43359 ( \43674 , \25033 , \25037 );
nand \U$43360 ( \43675 , \43673 , \43674 );
and \U$43361 ( \43676 , \25669 , \43675 );
nand \U$43362 ( \43677 , \25351 , \25352 );
or \U$43363 ( \43678 , \25668 , \43677 );
nand \U$43364 ( \43679 , \25663 , \25667 );
nand \U$43365 ( \43680 , \43678 , \43679 );
nor \U$43366 ( \43681 , \43676 , \43680 );
or \U$43367 ( \43682 , \26900 , \43681 );
nand \U$43368 ( \43683 , \25976 , \25980 );
or \U$43369 ( \43684 , \26291 , \43683 );
nand \U$43370 ( \43685 , \26286 , \26290 );
nand \U$43371 ( \43686 , \43684 , \43685 );
and \U$43372 ( \43687 , \26899 , \43686 );
nand \U$43373 ( \43688 , \26592 , \26596 );
or \U$43374 ( \43689 , \26898 , \43688 );
nand \U$43375 ( \43690 , \26893 , \26897 );
nand \U$43376 ( \43691 , \43689 , \43690 );
nor \U$43377 ( \43692 , \43687 , \43691 );
nand \U$43378 ( \43693 , \43682 , \43692 );
and \U$43379 ( \43694 , \29123 , \43693 );
nand \U$43380 ( \43695 , \27193 , \27197 );
or \U$43381 ( \43696 , \27488 , \43695 );
nand \U$43382 ( \43697 , \27483 , \27487 );
nand \U$43383 ( \43698 , \43696 , \43697 );
and \U$43384 ( \43699 , \28052 , \43698 );
nand \U$43385 ( \43700 , \27769 , \27773 );
or \U$43386 ( \43701 , \28051 , \43700 );
nand \U$43387 ( \43702 , \28049 , \28050 );
nand \U$43388 ( \43703 , \43701 , \43702 );
nor \U$43389 ( \43704 , \43699 , \43703 );
or \U$43390 ( \43705 , \29122 , \43704 );
nand \U$43391 ( \43706 , \28323 , \28327 );
or \U$43392 ( \43707 , \28595 , \43706 );
nand \U$43393 ( \43708 , \28593 , \28594 );
nand \U$43394 ( \43709 , \43707 , \43708 );
and \U$43395 ( \43710 , \29121 , \43709 );
nand \U$43396 ( \43711 , \28858 , \28859 );
or \U$43397 ( \43712 , \29120 , \43711 );
nand \U$43398 ( \43713 , \29115 , \29119 );
nand \U$43399 ( \43714 , \43712 , \43713 );
nor \U$43400 ( \43715 , \43710 , \43714 );
nand \U$43401 ( \43716 , \43705 , \43715 );
nor \U$43402 ( \43717 , \43694 , \43716 );
or \U$43403 ( \43718 , \32641 , \43717 );
nand \U$43404 ( \43719 , \29376 , \29377 );
or \U$43405 ( \43720 , \29627 , \43719 );
nand \U$43406 ( \43721 , \29625 , \29626 );
nand \U$43407 ( \43722 , \43720 , \43721 );
and \U$43408 ( \43723 , \30119 , \43722 );
nand \U$43409 ( \43724 , \29873 , \29874 );
or \U$43410 ( \43725 , \30118 , \43724 );
nand \U$43411 ( \43726 , \30116 , \30117 );
nand \U$43412 ( \43727 , \43725 , \43726 );
nor \U$43413 ( \43728 , \43723 , \43727 );
or \U$43414 ( \43729 , \31044 , \43728 );
nand \U$43415 ( \43730 , \30357 , \30358 );
or \U$43416 ( \43731 , \30590 , \43730 );
nand \U$43417 ( \43732 , \30588 , \30589 );
nand \U$43418 ( \43733 , \43731 , \43732 );
and \U$43419 ( \43734 , \31043 , \43733 );
nand \U$43420 ( \43735 , \30818 , \30819 );
or \U$43421 ( \43736 , \31042 , \43735 );
nand \U$43422 ( \43737 , \31040 , \31041 );
nand \U$43423 ( \43738 , \43736 , \43737 );
nor \U$43424 ( \43739 , \43734 , \43738 );
nand \U$43425 ( \43740 , \43729 , \43739 );
and \U$43426 ( \43741 , \32640 , \43740 );
nand \U$43427 ( \43742 , \31261 , \31262 );
or \U$43428 ( \43743 , \31474 , \43742 );
nand \U$43429 ( \43744 , \31472 , \31473 );
nand \U$43430 ( \43745 , \43743 , \43744 );
and \U$43431 ( \43746 , \31882 , \43745 );
nand \U$43432 ( \43747 , \31680 , \31681 );
or \U$43433 ( \43748 , \31881 , \43747 );
nand \U$43434 ( \43749 , \31879 , \31880 );
nand \U$43435 ( \43750 , \43748 , \43749 );
nor \U$43436 ( \43751 , \43746 , \43750 );
or \U$43437 ( \43752 , \32639 , \43751 );
nand \U$43438 ( \43753 , \32078 , \32079 );
or \U$43439 ( \43754 , \32269 , \43753 );
nand \U$43440 ( \43755 , \32267 , \32268 );
nand \U$43441 ( \43756 , \43754 , \43755 );
and \U$43442 ( \43757 , \32638 , \43756 );
nand \U$43443 ( \43758 , \32452 , \32456 );
or \U$43444 ( \43759 , \32637 , \43758 );
nand \U$43445 ( \43760 , \32632 , \32636 );
nand \U$43446 ( \43761 , \43759 , \43760 );
nor \U$43447 ( \43762 , \43757 , \43761 );
nand \U$43448 ( \43763 , \43752 , \43762 );
nor \U$43449 ( \43764 , \43741 , \43763 );
nand \U$43450 ( \43765 , \43718 , \43764 );
and \U$43451 ( \43766 , \35779 , \43765 );
nand \U$43452 ( \43767 , \32812 , \32816 );
or \U$43453 ( \43768 , \32984 , \43767 );
nand \U$43454 ( \43769 , \32982 , \32983 );
nand \U$43455 ( \43770 , \43768 , \43769 );
and \U$43456 ( \43771 , \33309 , \43770 );
nand \U$43457 ( \43772 , \33147 , \33148 );
or \U$43458 ( \43773 , \33308 , \43772 );
nand \U$43459 ( \43774 , \33306 , \33307 );
nand \U$43460 ( \43775 , \43773 , \43774 );
nor \U$43461 ( \43776 , \43771 , \43775 );
or \U$43462 ( \43777 , \33914 , \43776 );
nand \U$43463 ( \43778 , \33465 , \33466 );
or \U$43464 ( \43779 , \33620 , \43778 );
nand \U$43465 ( \43780 , \33618 , \33619 );
nand \U$43466 ( \43781 , \43779 , \43780 );
and \U$43467 ( \43782 , \33913 , \43781 );
nand \U$43468 ( \43783 , \33768 , \33769 );
or \U$43469 ( \43784 , \33912 , \43783 );
nand \U$43470 ( \43785 , \33910 , \33911 );
nand \U$43471 ( \43786 , \43784 , \43785 );
nor \U$43472 ( \43787 , \43782 , \43786 );
nand \U$43473 ( \43788 , \43777 , \43787 );
and \U$43474 ( \43789 , \34867 , \43788 );
nand \U$43475 ( \43790 , \34050 , \34051 );
or \U$43476 ( \43791 , \34181 , \43790 );
nand \U$43477 ( \43792 , \34179 , \34180 );
nand \U$43478 ( \43793 , \43791 , \43792 );
and \U$43479 ( \43794 , \34432 , \43793 );
nand \U$43480 ( \43795 , \34308 , \34309 );
or \U$43481 ( \43796 , \34431 , \43795 );
nand \U$43482 ( \43797 , \34429 , \34430 );
nand \U$43483 ( \43798 , \43796 , \43797 );
nor \U$43484 ( \43799 , \43794 , \43798 );
or \U$43485 ( \43800 , \34866 , \43799 );
nand \U$43486 ( \43801 , \34545 , \34549 );
or \U$43487 ( \43802 , \34660 , \43801 );
nand \U$43488 ( \43803 , \34655 , \34659 );
nand \U$43489 ( \43804 , \43802 , \43803 );
and \U$43490 ( \43805 , \34865 , \43804 );
nand \U$43491 ( \43806 , \34763 , \34764 );
or \U$43492 ( \43807 , \34864 , \43806 );
nand \U$43493 ( \43808 , \34862 , \34863 );
nand \U$43494 ( \43809 , \43807 , \43808 );
nor \U$43495 ( \43810 , \43805 , \43809 );
nand \U$43496 ( \43811 , \43800 , \43810 );
nor \U$43497 ( \43812 , \43789 , \43811 );
or \U$43498 ( \43813 , \35778 , \43812 );
nand \U$43499 ( \43814 , \34963 , \34964 );
or \U$43500 ( \43815 , \35054 , \43814 );
nand \U$43501 ( \43816 , \35052 , \35053 );
nand \U$43502 ( \43817 , \43815 , \43816 );
and \U$43503 ( \43818 , \35222 , \43817 );
nand \U$43504 ( \43819 , \35140 , \35141 );
or \U$43505 ( \43820 , \35221 , \43819 );
nand \U$43506 ( \43821 , \35219 , \35220 );
nand \U$43507 ( \43822 , \43820 , \43821 );
nor \U$43508 ( \43823 , \43818 , \43822 );
or \U$43509 ( \43824 , \35499 , \43823 );
nand \U$43510 ( \43825 , \35298 , \35299 );
or \U$43511 ( \43826 , \35370 , \43825 );
nand \U$43512 ( \43827 , \35365 , \35369 );
nand \U$43513 ( \43828 , \43826 , \43827 );
and \U$43514 ( \43829 , \35498 , \43828 );
nand \U$43515 ( \43830 , \35434 , \35435 );
or \U$43516 ( \43831 , \35497 , \43830 );
nand \U$43517 ( \43832 , \35495 , \35496 );
nand \U$43518 ( \43833 , \43831 , \43832 );
nor \U$43519 ( \43834 , \43829 , \43833 );
nand \U$43520 ( \43835 , \43824 , \43834 );
and \U$43521 ( \43836 , \35777 , \43835 );
nand \U$43522 ( \43837 , \35555 , \35556 );
or \U$43523 ( \43838 , \35606 , \43837 );
nand \U$43524 ( \43839 , \35604 , \35605 );
nand \U$43525 ( \43840 , \43838 , \43839 );
and \U$43526 ( \43841 , \35695 , \43840 );
nand \U$43527 ( \43842 , \35652 , \35653 );
or \U$43528 ( \43843 , \35694 , \43842 );
nand \U$43529 ( \43844 , \35689 , \35693 );
nand \U$43530 ( \43845 , \43843 , \43844 );
nor \U$43531 ( \43846 , \43841 , \43845 );
or \U$43532 ( \43847 , \35776 , \43846 );
nand \U$43533 ( \43848 , \35729 , \35730 );
or \U$43534 ( \43849 , \35753 , \43848 );
nand \U$43535 ( \43850 , \35751 , \35752 );
nand \U$43536 ( \43851 , \43849 , \43850 );
and \U$43537 ( \43852 , \35775 , \43851 );
nand \U$43538 ( \43853 , \35765 , \35766 );
or \U$43539 ( \43854 , \35774 , \43853 );
nand \U$43540 ( \43855 , \35769 , \35773 );
nand \U$43541 ( \43856 , \43854 , \43855 );
nor \U$43542 ( \43857 , \43852 , \43856 );
nand \U$43543 ( \43858 , \43847 , \43857 );
nor \U$43544 ( \43859 , \43836 , \43858 );
nand \U$43545 ( \43860 , \43813 , \43859 );
nor \U$43546 ( \43861 , \43766 , \43860 );
nand \U$43547 ( \43862 , \43671 , \43861 );
not \U$43548 ( \43863 , \43862 );
xor \U$43549 ( \43864 , \22062 , \43863 );
buf \U$43550 ( \43865 , \43864 );
_HMUX rb622 ( \43866_nRb622 , \21589 , \43865 , RIc0c97c8_1 );
buf \U$43551 ( \43867 , \43866_nRb622 );
xor \U$43552 ( \43868 , \402 , \21585 );
buf \U$43553 ( \43869 , \43868 );
not \U$43554 ( \43870 , \35774 );
nand \U$43555 ( \43871 , \43855 , \43870 );
nor \U$43556 ( \43872 , \41857 , \24724 );
nor \U$43557 ( \43873 , \25038 , \25353 );
nand \U$43558 ( \43874 , \43872 , \43873 );
nor \U$43559 ( \43875 , \25668 , \25981 );
nor \U$43560 ( \43876 , \26291 , \26597 );
nand \U$43561 ( \43877 , \43875 , \43876 );
nor \U$43562 ( \43878 , \43874 , \43877 );
nor \U$43563 ( \43879 , \26898 , \27198 );
nor \U$43564 ( \43880 , \27488 , \27774 );
nand \U$43565 ( \43881 , \43879 , \43880 );
nor \U$43566 ( \43882 , \28051 , \28328 );
nor \U$43567 ( \43883 , \28595 , \28860 );
nand \U$43568 ( \43884 , \43882 , \43883 );
nor \U$43569 ( \43885 , \43881 , \43884 );
nand \U$43570 ( \43886 , \43878 , \43885 );
nor \U$43571 ( \43887 , \29120 , \29378 );
nor \U$43572 ( \43888 , \29627 , \29875 );
nand \U$43573 ( \43889 , \43887 , \43888 );
nor \U$43574 ( \43890 , \30118 , \30359 );
nor \U$43575 ( \43891 , \30590 , \30820 );
nand \U$43576 ( \43892 , \43890 , \43891 );
nor \U$43577 ( \43893 , \43889 , \43892 );
nor \U$43578 ( \43894 , \31042 , \31263 );
nor \U$43579 ( \43895 , \31474 , \31682 );
nand \U$43580 ( \43896 , \43894 , \43895 );
nor \U$43581 ( \43897 , \31881 , \32080 );
nor \U$43582 ( \43898 , \32269 , \32457 );
nand \U$43583 ( \43899 , \43897 , \43898 );
nor \U$43584 ( \43900 , \43896 , \43899 );
nand \U$43585 ( \43901 , \43893 , \43900 );
nor \U$43586 ( \43902 , \43886 , \43901 );
nor \U$43587 ( \43903 , \32637 , \32817 );
nor \U$43588 ( \43904 , \32984 , \33149 );
nand \U$43589 ( \43905 , \43903 , \43904 );
nor \U$43590 ( \43906 , \33308 , \33467 );
nor \U$43591 ( \43907 , \33620 , \33770 );
nand \U$43592 ( \43908 , \43906 , \43907 );
nor \U$43593 ( \43909 , \43905 , \43908 );
nor \U$43594 ( \43910 , \33912 , \34052 );
nor \U$43595 ( \43911 , \34181 , \34310 );
nand \U$43596 ( \43912 , \43910 , \43911 );
nor \U$43597 ( \43913 , \34431 , \34550 );
nor \U$43598 ( \43914 , \34660 , \34765 );
nand \U$43599 ( \43915 , \43913 , \43914 );
nor \U$43600 ( \43916 , \43912 , \43915 );
nand \U$43601 ( \43917 , \43909 , \43916 );
nor \U$43602 ( \43918 , \34864 , \34965 );
nor \U$43603 ( \43919 , \35054 , \35142 );
nand \U$43604 ( \43920 , \43918 , \43919 );
nor \U$43605 ( \43921 , \35221 , \35300 );
nor \U$43606 ( \43922 , \35370 , \35436 );
nand \U$43607 ( \43923 , \43921 , \43922 );
nor \U$43608 ( \43924 , \43920 , \43923 );
nor \U$43609 ( \43925 , \35497 , \35557 );
nor \U$43610 ( \43926 , \35606 , \35654 );
nand \U$43611 ( \43927 , \43925 , \43926 );
nor \U$43612 ( \43928 , \35694 , \35731 );
nor \U$43613 ( \43929 , \35753 , \35767 );
nand \U$43614 ( \43930 , \43928 , \43929 );
nor \U$43615 ( \43931 , \43927 , \43930 );
nand \U$43616 ( \43932 , \43924 , \43931 );
nor \U$43617 ( \43933 , \43917 , \43932 );
nand \U$43618 ( \43934 , \43902 , \43933 );
nor \U$43619 ( \43935 , \43170 , \36532 );
nor \U$43620 ( \43936 , \36687 , \36849 );
nand \U$43621 ( \43937 , \43935 , \43936 );
nor \U$43622 ( \43938 , \37014 , \37187 );
nor \U$43623 ( \43939 , \37362 , \37544 );
nand \U$43624 ( \43940 , \43938 , \43939 );
nor \U$43625 ( \43941 , \43937 , \43940 );
nor \U$43626 ( \43942 , \37729 , \37923 );
nor \U$43627 ( \43943 , \38118 , \38320 );
nand \U$43628 ( \43944 , \43942 , \43943 );
nor \U$43629 ( \43945 , \38525 , \38737 );
nor \U$43630 ( \43946 , \38955 , \39177 );
nand \U$43631 ( \43947 , \43945 , \43946 );
nor \U$43632 ( \43948 , \43944 , \43947 );
nand \U$43633 ( \43949 , \43941 , \43948 );
nor \U$43634 ( \43950 , \39402 , \39637 );
nor \U$43635 ( \43951 , \39872 , \40114 );
nand \U$43636 ( \43952 , \43950 , \43951 );
nor \U$43637 ( \43953 , \40359 , \40612 );
nor \U$43638 ( \43954 , \40867 , \41129 );
nand \U$43639 ( \43955 , \43953 , \43954 );
nor \U$43640 ( \43956 , \43952 , \43955 );
nor \U$43641 ( \43957 , \41394 , \41560 );
nor \U$43642 ( \43958 , \41667 , \41739 );
nand \U$43643 ( \43959 , \43957 , \43958 );
nor \U$43644 ( \43960 , \41784 , \41819 );
nor \U$43645 ( \43961 , \41841 , \41854 );
nand \U$43646 ( \43962 , \43960 , \43961 );
nor \U$43647 ( \43963 , \43959 , \43962 );
nand \U$43648 ( \43964 , \43956 , \43963 );
nor \U$43649 ( \43965 , \43949 , \43964 );
nor \U$43650 ( \43966 , \43425 , \42103 );
nor \U$43651 ( \43967 , \42178 , \42260 );
nand \U$43652 ( \43968 , \43966 , \43967 );
nor \U$43653 ( \43969 , \42345 , \42438 );
nor \U$43654 ( \43970 , \42533 , \42635 );
nand \U$43655 ( \43971 , \43969 , \43970 );
nor \U$43656 ( \43972 , \43968 , \43971 );
nor \U$43657 ( \43973 , \42740 , \42854 );
nor \U$43658 ( \43974 , \42969 , \43043 );
nand \U$43659 ( \43975 , \43973 , \43974 );
nor \U$43660 ( \43976 , \43088 , \43123 );
nor \U$43661 ( \43977 , \43148 , \43163 );
nand \U$43662 ( \43978 , \43976 , \43977 );
nor \U$43663 ( \43979 , \43975 , \43978 );
nand \U$43664 ( \43980 , \43972 , \43979 );
nor \U$43665 ( \43981 , \43472 , \43238 );
nor \U$43666 ( \43982 , \43273 , \43315 );
nand \U$43667 ( \43983 , \43981 , \43982 );
nor \U$43668 ( \43984 , \43360 , \43389 );
nor \U$43669 ( \43985 , \43406 , \43418 );
nand \U$43670 ( \43986 , \43984 , \43985 );
nor \U$43671 ( \43987 , \43983 , \43986 );
nor \U$43672 ( \43988 , \43478 , \43443 );
nor \U$43673 ( \43989 , \43458 , \43468 );
nand \U$43674 ( \43990 , \43988 , \43989 );
or \U$43675 ( \43991 , \43990 , \43486 );
or \U$43676 ( \43992 , \43443 , \43488 );
nand \U$43677 ( \43993 , \43992 , \43492 );
and \U$43678 ( \43994 , \43989 , \43993 );
or \U$43679 ( \43995 , \43468 , \43494 );
nand \U$43680 ( \43996 , \43995 , \43497 );
nor \U$43681 ( \43997 , \43994 , \43996 );
nand \U$43682 ( \43998 , \43991 , \43997 );
and \U$43683 ( \43999 , \43987 , \43998 );
or \U$43684 ( \44000 , \43238 , \43499 );
nand \U$43685 ( \44001 , \44000 , \43504 );
and \U$43686 ( \44002 , \43982 , \44001 );
or \U$43687 ( \44003 , \43315 , \43506 );
nand \U$43688 ( \44004 , \44003 , \43509 );
nor \U$43689 ( \44005 , \44002 , \44004 );
or \U$43690 ( \44006 , \43986 , \44005 );
or \U$43691 ( \44007 , \43389 , \43511 );
nand \U$43692 ( \44008 , \44007 , \43515 );
and \U$43693 ( \44009 , \43985 , \44008 );
or \U$43694 ( \44010 , \43418 , \43517 );
nand \U$43695 ( \44011 , \44010 , \43520 );
nor \U$43696 ( \44012 , \44009 , \44011 );
nand \U$43697 ( \44013 , \44006 , \44012 );
nor \U$43698 ( \44014 , \43999 , \44013 );
or \U$43699 ( \44015 , \43980 , \44014 );
or \U$43700 ( \44016 , \42103 , \43522 );
nand \U$43701 ( \44017 , \44016 , \43528 );
and \U$43702 ( \44018 , \43967 , \44017 );
or \U$43703 ( \44019 , \42260 , \43530 );
nand \U$43704 ( \44020 , \44019 , \43533 );
nor \U$43705 ( \44021 , \44018 , \44020 );
or \U$43706 ( \44022 , \43971 , \44021 );
or \U$43707 ( \44023 , \42438 , \43535 );
nand \U$43708 ( \44024 , \44023 , \43539 );
and \U$43709 ( \44025 , \43970 , \44024 );
or \U$43710 ( \44026 , \42635 , \43541 );
nand \U$43711 ( \44027 , \44026 , \43544 );
nor \U$43712 ( \44028 , \44025 , \44027 );
nand \U$43713 ( \44029 , \44022 , \44028 );
and \U$43714 ( \44030 , \43979 , \44029 );
or \U$43715 ( \44031 , \42854 , \43546 );
nand \U$43716 ( \44032 , \44031 , \43551 );
and \U$43717 ( \44033 , \43974 , \44032 );
or \U$43718 ( \44034 , \43043 , \43553 );
nand \U$43719 ( \44035 , \44034 , \43556 );
nor \U$43720 ( \44036 , \44033 , \44035 );
or \U$43721 ( \44037 , \43978 , \44036 );
or \U$43722 ( \44038 , \43123 , \43558 );
nand \U$43723 ( \44039 , \44038 , \43562 );
and \U$43724 ( \44040 , \43977 , \44039 );
or \U$43725 ( \44041 , \43163 , \43564 );
nand \U$43726 ( \44042 , \44041 , \43567 );
nor \U$43727 ( \44043 , \44040 , \44042 );
nand \U$43728 ( \44044 , \44037 , \44043 );
nor \U$43729 ( \44045 , \44030 , \44044 );
nand \U$43730 ( \44046 , \44015 , \44045 );
and \U$43731 ( \44047 , \43965 , \44046 );
or \U$43732 ( \44048 , \36532 , \43569 );
nand \U$43733 ( \44049 , \44048 , \43576 );
and \U$43734 ( \44050 , \43936 , \44049 );
or \U$43735 ( \44051 , \36849 , \43578 );
nand \U$43736 ( \44052 , \44051 , \43581 );
nor \U$43737 ( \44053 , \44050 , \44052 );
or \U$43738 ( \44054 , \43940 , \44053 );
or \U$43739 ( \44055 , \37187 , \43583 );
nand \U$43740 ( \44056 , \44055 , \43587 );
and \U$43741 ( \44057 , \43939 , \44056 );
or \U$43742 ( \44058 , \37544 , \43589 );
nand \U$43743 ( \44059 , \44058 , \43592 );
nor \U$43744 ( \44060 , \44057 , \44059 );
nand \U$43745 ( \44061 , \44054 , \44060 );
and \U$43746 ( \44062 , \43948 , \44061 );
or \U$43747 ( \44063 , \37923 , \43594 );
nand \U$43748 ( \44064 , \44063 , \43599 );
and \U$43749 ( \44065 , \43943 , \44064 );
or \U$43750 ( \44066 , \38320 , \43601 );
nand \U$43751 ( \44067 , \44066 , \43604 );
nor \U$43752 ( \44068 , \44065 , \44067 );
or \U$43753 ( \44069 , \43947 , \44068 );
or \U$43754 ( \44070 , \38737 , \43606 );
nand \U$43755 ( \44071 , \44070 , \43610 );
and \U$43756 ( \44072 , \43946 , \44071 );
or \U$43757 ( \44073 , \39177 , \43612 );
nand \U$43758 ( \44074 , \44073 , \43615 );
nor \U$43759 ( \44075 , \44072 , \44074 );
nand \U$43760 ( \44076 , \44069 , \44075 );
nor \U$43761 ( \44077 , \44062 , \44076 );
or \U$43762 ( \44078 , \43964 , \44077 );
or \U$43763 ( \44079 , \39637 , \43617 );
nand \U$43764 ( \44080 , \44079 , \43623 );
and \U$43765 ( \44081 , \43951 , \44080 );
or \U$43766 ( \44082 , \40114 , \43625 );
nand \U$43767 ( \44083 , \44082 , \43628 );
nor \U$43768 ( \44084 , \44081 , \44083 );
or \U$43769 ( \44085 , \43955 , \44084 );
or \U$43770 ( \44086 , \40612 , \43630 );
nand \U$43771 ( \44087 , \44086 , \43634 );
and \U$43772 ( \44088 , \43954 , \44087 );
or \U$43773 ( \44089 , \41129 , \43636 );
nand \U$43774 ( \44090 , \44089 , \43639 );
nor \U$43775 ( \44091 , \44088 , \44090 );
nand \U$43776 ( \44092 , \44085 , \44091 );
and \U$43777 ( \44093 , \43963 , \44092 );
or \U$43778 ( \44094 , \41560 , \43641 );
nand \U$43779 ( \44095 , \44094 , \43646 );
and \U$43780 ( \44096 , \43958 , \44095 );
or \U$43781 ( \44097 , \41739 , \43648 );
nand \U$43782 ( \44098 , \44097 , \43651 );
nor \U$43783 ( \44099 , \44096 , \44098 );
or \U$43784 ( \44100 , \43962 , \44099 );
or \U$43785 ( \44101 , \41819 , \43653 );
nand \U$43786 ( \44102 , \44101 , \43657 );
and \U$43787 ( \44103 , \43961 , \44102 );
or \U$43788 ( \44104 , \41854 , \43659 );
nand \U$43789 ( \44105 , \44104 , \43662 );
nor \U$43790 ( \44106 , \44103 , \44105 );
nand \U$43791 ( \44107 , \44100 , \44106 );
nor \U$43792 ( \44108 , \44093 , \44107 );
nand \U$43793 ( \44109 , \44078 , \44108 );
nor \U$43794 ( \44110 , \44047 , \44109 );
or \U$43795 ( \44111 , \43934 , \44110 );
or \U$43796 ( \44112 , \24724 , \43664 );
nand \U$43797 ( \44113 , \44112 , \43672 );
and \U$43798 ( \44114 , \43873 , \44113 );
or \U$43799 ( \44115 , \25353 , \43674 );
nand \U$43800 ( \44116 , \44115 , \43677 );
nor \U$43801 ( \44117 , \44114 , \44116 );
or \U$43802 ( \44118 , \43877 , \44117 );
or \U$43803 ( \44119 , \25981 , \43679 );
nand \U$43804 ( \44120 , \44119 , \43683 );
and \U$43805 ( \44121 , \43876 , \44120 );
or \U$43806 ( \44122 , \26597 , \43685 );
nand \U$43807 ( \44123 , \44122 , \43688 );
nor \U$43808 ( \44124 , \44121 , \44123 );
nand \U$43809 ( \44125 , \44118 , \44124 );
and \U$43810 ( \44126 , \43885 , \44125 );
or \U$43811 ( \44127 , \27198 , \43690 );
nand \U$43812 ( \44128 , \44127 , \43695 );
and \U$43813 ( \44129 , \43880 , \44128 );
or \U$43814 ( \44130 , \27774 , \43697 );
nand \U$43815 ( \44131 , \44130 , \43700 );
nor \U$43816 ( \44132 , \44129 , \44131 );
or \U$43817 ( \44133 , \43884 , \44132 );
or \U$43818 ( \44134 , \28328 , \43702 );
nand \U$43819 ( \44135 , \44134 , \43706 );
and \U$43820 ( \44136 , \43883 , \44135 );
or \U$43821 ( \44137 , \28860 , \43708 );
nand \U$43822 ( \44138 , \44137 , \43711 );
nor \U$43823 ( \44139 , \44136 , \44138 );
nand \U$43824 ( \44140 , \44133 , \44139 );
nor \U$43825 ( \44141 , \44126 , \44140 );
or \U$43826 ( \44142 , \43901 , \44141 );
or \U$43827 ( \44143 , \29378 , \43713 );
nand \U$43828 ( \44144 , \44143 , \43719 );
and \U$43829 ( \44145 , \43888 , \44144 );
or \U$43830 ( \44146 , \29875 , \43721 );
nand \U$43831 ( \44147 , \44146 , \43724 );
nor \U$43832 ( \44148 , \44145 , \44147 );
or \U$43833 ( \44149 , \43892 , \44148 );
or \U$43834 ( \44150 , \30359 , \43726 );
nand \U$43835 ( \44151 , \44150 , \43730 );
and \U$43836 ( \44152 , \43891 , \44151 );
or \U$43837 ( \44153 , \30820 , \43732 );
nand \U$43838 ( \44154 , \44153 , \43735 );
nor \U$43839 ( \44155 , \44152 , \44154 );
nand \U$43840 ( \44156 , \44149 , \44155 );
and \U$43841 ( \44157 , \43900 , \44156 );
or \U$43842 ( \44158 , \31263 , \43737 );
nand \U$43843 ( \44159 , \44158 , \43742 );
and \U$43844 ( \44160 , \43895 , \44159 );
or \U$43845 ( \44161 , \31682 , \43744 );
nand \U$43846 ( \44162 , \44161 , \43747 );
nor \U$43847 ( \44163 , \44160 , \44162 );
or \U$43848 ( \44164 , \43899 , \44163 );
or \U$43849 ( \44165 , \32080 , \43749 );
nand \U$43850 ( \44166 , \44165 , \43753 );
and \U$43851 ( \44167 , \43898 , \44166 );
or \U$43852 ( \44168 , \32457 , \43755 );
nand \U$43853 ( \44169 , \44168 , \43758 );
nor \U$43854 ( \44170 , \44167 , \44169 );
nand \U$43855 ( \44171 , \44164 , \44170 );
nor \U$43856 ( \44172 , \44157 , \44171 );
nand \U$43857 ( \44173 , \44142 , \44172 );
and \U$43858 ( \44174 , \43933 , \44173 );
or \U$43859 ( \44175 , \32817 , \43760 );
nand \U$43860 ( \44176 , \44175 , \43767 );
and \U$43861 ( \44177 , \43904 , \44176 );
or \U$43862 ( \44178 , \33149 , \43769 );
nand \U$43863 ( \44179 , \44178 , \43772 );
nor \U$43864 ( \44180 , \44177 , \44179 );
or \U$43865 ( \44181 , \43908 , \44180 );
or \U$43866 ( \44182 , \33467 , \43774 );
nand \U$43867 ( \44183 , \44182 , \43778 );
and \U$43868 ( \44184 , \43907 , \44183 );
or \U$43869 ( \44185 , \33770 , \43780 );
nand \U$43870 ( \44186 , \44185 , \43783 );
nor \U$43871 ( \44187 , \44184 , \44186 );
nand \U$43872 ( \44188 , \44181 , \44187 );
and \U$43873 ( \44189 , \43916 , \44188 );
or \U$43874 ( \44190 , \34052 , \43785 );
nand \U$43875 ( \44191 , \44190 , \43790 );
and \U$43876 ( \44192 , \43911 , \44191 );
or \U$43877 ( \44193 , \34310 , \43792 );
nand \U$43878 ( \44194 , \44193 , \43795 );
nor \U$43879 ( \44195 , \44192 , \44194 );
or \U$43880 ( \44196 , \43915 , \44195 );
or \U$43881 ( \44197 , \34550 , \43797 );
nand \U$43882 ( \44198 , \44197 , \43801 );
and \U$43883 ( \44199 , \43914 , \44198 );
or \U$43884 ( \44200 , \34765 , \43803 );
nand \U$43885 ( \44201 , \44200 , \43806 );
nor \U$43886 ( \44202 , \44199 , \44201 );
nand \U$43887 ( \44203 , \44196 , \44202 );
nor \U$43888 ( \44204 , \44189 , \44203 );
or \U$43889 ( \44205 , \43932 , \44204 );
or \U$43890 ( \44206 , \34965 , \43808 );
nand \U$43891 ( \44207 , \44206 , \43814 );
and \U$43892 ( \44208 , \43919 , \44207 );
or \U$43893 ( \44209 , \35142 , \43816 );
nand \U$43894 ( \44210 , \44209 , \43819 );
nor \U$43895 ( \44211 , \44208 , \44210 );
or \U$43896 ( \44212 , \43923 , \44211 );
or \U$43897 ( \44213 , \35300 , \43821 );
nand \U$43898 ( \44214 , \44213 , \43825 );
and \U$43899 ( \44215 , \43922 , \44214 );
or \U$43900 ( \44216 , \35436 , \43827 );
nand \U$43901 ( \44217 , \44216 , \43830 );
nor \U$43902 ( \44218 , \44215 , \44217 );
nand \U$43903 ( \44219 , \44212 , \44218 );
and \U$43904 ( \44220 , \43931 , \44219 );
or \U$43905 ( \44221 , \35557 , \43832 );
nand \U$43906 ( \44222 , \44221 , \43837 );
and \U$43907 ( \44223 , \43926 , \44222 );
or \U$43908 ( \44224 , \35654 , \43839 );
nand \U$43909 ( \44225 , \44224 , \43842 );
nor \U$43910 ( \44226 , \44223 , \44225 );
or \U$43911 ( \44227 , \43930 , \44226 );
or \U$43912 ( \44228 , \35731 , \43844 );
nand \U$43913 ( \44229 , \44228 , \43848 );
and \U$43914 ( \44230 , \43929 , \44229 );
or \U$43915 ( \44231 , \35767 , \43850 );
nand \U$43916 ( \44232 , \44231 , \43853 );
nor \U$43917 ( \44233 , \44230 , \44232 );
nand \U$43918 ( \44234 , \44227 , \44233 );
nor \U$43919 ( \44235 , \44220 , \44234 );
nand \U$43920 ( \44236 , \44205 , \44235 );
nor \U$43921 ( \44237 , \44174 , \44236 );
nand \U$43922 ( \44238 , \44111 , \44237 );
not \U$43923 ( \44239 , \44238 );
xor \U$43924 ( \44240 , \43871 , \44239 );
buf \U$43925 ( \44241 , \44240 );
_HMUX rb5ec ( \44242_nRb5ec , \43869 , \44241 , RIc0c97c8_1 );
buf \U$43926 ( \44243 , \44242_nRb5ec );
xor \U$43927 ( \44244 , \472 , \21583 );
buf \U$43928 ( \44245 , \44244 );
not \U$43929 ( \44246 , \35767 );
nand \U$43930 ( \44247 , \43853 , \44246 );
nand \U$43931 ( \44248 , \41858 , \25039 );
nand \U$43932 ( \44249 , \25669 , \26292 );
nor \U$43933 ( \44250 , \44248 , \44249 );
nand \U$43934 ( \44251 , \26899 , \27489 );
nand \U$43935 ( \44252 , \28052 , \28596 );
nor \U$43936 ( \44253 , \44251 , \44252 );
nand \U$43937 ( \44254 , \44250 , \44253 );
nand \U$43938 ( \44255 , \29121 , \29628 );
nand \U$43939 ( \44256 , \30119 , \30591 );
nor \U$43940 ( \44257 , \44255 , \44256 );
nand \U$43941 ( \44258 , \31043 , \31475 );
nand \U$43942 ( \44259 , \31882 , \32270 );
nor \U$43943 ( \44260 , \44258 , \44259 );
nand \U$43944 ( \44261 , \44257 , \44260 );
nor \U$43945 ( \44262 , \44254 , \44261 );
nand \U$43946 ( \44263 , \32638 , \32985 );
nand \U$43947 ( \44264 , \33309 , \33621 );
nor \U$43948 ( \44265 , \44263 , \44264 );
nand \U$43949 ( \44266 , \33913 , \34182 );
nand \U$43950 ( \44267 , \34432 , \34661 );
nor \U$43951 ( \44268 , \44266 , \44267 );
nand \U$43952 ( \44269 , \44265 , \44268 );
nand \U$43953 ( \44270 , \34865 , \35055 );
nand \U$43954 ( \44271 , \35222 , \35371 );
nor \U$43955 ( \44272 , \44270 , \44271 );
nand \U$43956 ( \44273 , \35498 , \35607 );
nand \U$43957 ( \44274 , \35695 , \35754 );
nor \U$43958 ( \44275 , \44273 , \44274 );
nand \U$43959 ( \44276 , \44272 , \44275 );
nor \U$43960 ( \44277 , \44269 , \44276 );
nand \U$43961 ( \44278 , \44262 , \44277 );
nand \U$43962 ( \44279 , \43171 , \36688 );
nand \U$43963 ( \44280 , \37015 , \37363 );
nor \U$43964 ( \44281 , \44279 , \44280 );
nand \U$43965 ( \44282 , \37730 , \38119 );
nand \U$43966 ( \44283 , \38526 , \38956 );
nor \U$43967 ( \44284 , \44282 , \44283 );
nand \U$43968 ( \44285 , \44281 , \44284 );
nand \U$43969 ( \44286 , \39403 , \39873 );
nand \U$43970 ( \44287 , \40360 , \40868 );
nor \U$43971 ( \44288 , \44286 , \44287 );
nand \U$43972 ( \44289 , \41395 , \41668 );
nand \U$43973 ( \44290 , \41785 , \41842 );
nor \U$43974 ( \44291 , \44289 , \44290 );
nand \U$43975 ( \44292 , \44288 , \44291 );
nor \U$43976 ( \44293 , \44285 , \44292 );
nand \U$43977 ( \44294 , \43426 , \42179 );
nand \U$43978 ( \44295 , \42346 , \42534 );
nor \U$43979 ( \44296 , \44294 , \44295 );
nand \U$43980 ( \44297 , \42741 , \42970 );
nand \U$43981 ( \44298 , \43089 , \43149 );
nor \U$43982 ( \44299 , \44297 , \44298 );
nand \U$43983 ( \44300 , \44296 , \44299 );
nand \U$43984 ( \44301 , \43473 , \43274 );
nand \U$43985 ( \44302 , \43361 , \43407 );
nor \U$43986 ( \44303 , \44301 , \44302 );
and \U$43987 ( \44304 , \43459 , \43489 );
nor \U$43988 ( \44305 , \44304 , \43495 );
not \U$43989 ( \44306 , \44305 );
and \U$43990 ( \44307 , \44303 , \44306 );
and \U$43991 ( \44308 , \43274 , \43500 );
nor \U$43992 ( \44309 , \44308 , \43507 );
or \U$43993 ( \44310 , \44302 , \44309 );
and \U$43994 ( \44311 , \43407 , \43512 );
nor \U$43995 ( \44312 , \44311 , \43518 );
nand \U$43996 ( \44313 , \44310 , \44312 );
nor \U$43997 ( \44314 , \44307 , \44313 );
or \U$43998 ( \44315 , \44300 , \44314 );
and \U$43999 ( \44316 , \42179 , \43523 );
nor \U$44000 ( \44317 , \44316 , \43531 );
or \U$44001 ( \44318 , \44295 , \44317 );
and \U$44002 ( \44319 , \42534 , \43536 );
nor \U$44003 ( \44320 , \44319 , \43542 );
nand \U$44004 ( \44321 , \44318 , \44320 );
and \U$44005 ( \44322 , \44299 , \44321 );
and \U$44006 ( \44323 , \42970 , \43547 );
nor \U$44007 ( \44324 , \44323 , \43554 );
or \U$44008 ( \44325 , \44298 , \44324 );
and \U$44009 ( \44326 , \43149 , \43559 );
nor \U$44010 ( \44327 , \44326 , \43565 );
nand \U$44011 ( \44328 , \44325 , \44327 );
nor \U$44012 ( \44329 , \44322 , \44328 );
nand \U$44013 ( \44330 , \44315 , \44329 );
and \U$44014 ( \44331 , \44293 , \44330 );
and \U$44015 ( \44332 , \36688 , \43570 );
nor \U$44016 ( \44333 , \44332 , \43579 );
or \U$44017 ( \44334 , \44280 , \44333 );
and \U$44018 ( \44335 , \37363 , \43584 );
nor \U$44019 ( \44336 , \44335 , \43590 );
nand \U$44020 ( \44337 , \44334 , \44336 );
and \U$44021 ( \44338 , \44284 , \44337 );
and \U$44022 ( \44339 , \38119 , \43595 );
nor \U$44023 ( \44340 , \44339 , \43602 );
or \U$44024 ( \44341 , \44283 , \44340 );
and \U$44025 ( \44342 , \38956 , \43607 );
nor \U$44026 ( \44343 , \44342 , \43613 );
nand \U$44027 ( \44344 , \44341 , \44343 );
nor \U$44028 ( \44345 , \44338 , \44344 );
or \U$44029 ( \44346 , \44292 , \44345 );
and \U$44030 ( \44347 , \39873 , \43618 );
nor \U$44031 ( \44348 , \44347 , \43626 );
or \U$44032 ( \44349 , \44287 , \44348 );
and \U$44033 ( \44350 , \40868 , \43631 );
nor \U$44034 ( \44351 , \44350 , \43637 );
nand \U$44035 ( \44352 , \44349 , \44351 );
and \U$44036 ( \44353 , \44291 , \44352 );
and \U$44037 ( \44354 , \41668 , \43642 );
nor \U$44038 ( \44355 , \44354 , \43649 );
or \U$44039 ( \44356 , \44290 , \44355 );
and \U$44040 ( \44357 , \41842 , \43654 );
nor \U$44041 ( \44358 , \44357 , \43660 );
nand \U$44042 ( \44359 , \44356 , \44358 );
nor \U$44043 ( \44360 , \44353 , \44359 );
nand \U$44044 ( \44361 , \44346 , \44360 );
nor \U$44045 ( \44362 , \44331 , \44361 );
or \U$44046 ( \44363 , \44278 , \44362 );
and \U$44047 ( \44364 , \25039 , \43665 );
nor \U$44048 ( \44365 , \44364 , \43675 );
or \U$44049 ( \44366 , \44249 , \44365 );
and \U$44050 ( \44367 , \26292 , \43680 );
nor \U$44051 ( \44368 , \44367 , \43686 );
nand \U$44052 ( \44369 , \44366 , \44368 );
and \U$44053 ( \44370 , \44253 , \44369 );
and \U$44054 ( \44371 , \27489 , \43691 );
nor \U$44055 ( \44372 , \44371 , \43698 );
or \U$44056 ( \44373 , \44252 , \44372 );
and \U$44057 ( \44374 , \28596 , \43703 );
nor \U$44058 ( \44375 , \44374 , \43709 );
nand \U$44059 ( \44376 , \44373 , \44375 );
nor \U$44060 ( \44377 , \44370 , \44376 );
or \U$44061 ( \44378 , \44261 , \44377 );
and \U$44062 ( \44379 , \29628 , \43714 );
nor \U$44063 ( \44380 , \44379 , \43722 );
or \U$44064 ( \44381 , \44256 , \44380 );
and \U$44065 ( \44382 , \30591 , \43727 );
nor \U$44066 ( \44383 , \44382 , \43733 );
nand \U$44067 ( \44384 , \44381 , \44383 );
and \U$44068 ( \44385 , \44260 , \44384 );
and \U$44069 ( \44386 , \31475 , \43738 );
nor \U$44070 ( \44387 , \44386 , \43745 );
or \U$44071 ( \44388 , \44259 , \44387 );
and \U$44072 ( \44389 , \32270 , \43750 );
nor \U$44073 ( \44390 , \44389 , \43756 );
nand \U$44074 ( \44391 , \44388 , \44390 );
nor \U$44075 ( \44392 , \44385 , \44391 );
nand \U$44076 ( \44393 , \44378 , \44392 );
and \U$44077 ( \44394 , \44277 , \44393 );
and \U$44078 ( \44395 , \32985 , \43761 );
nor \U$44079 ( \44396 , \44395 , \43770 );
or \U$44080 ( \44397 , \44264 , \44396 );
and \U$44081 ( \44398 , \33621 , \43775 );
nor \U$44082 ( \44399 , \44398 , \43781 );
nand \U$44083 ( \44400 , \44397 , \44399 );
and \U$44084 ( \44401 , \44268 , \44400 );
and \U$44085 ( \44402 , \34182 , \43786 );
nor \U$44086 ( \44403 , \44402 , \43793 );
or \U$44087 ( \44404 , \44267 , \44403 );
and \U$44088 ( \44405 , \34661 , \43798 );
nor \U$44089 ( \44406 , \44405 , \43804 );
nand \U$44090 ( \44407 , \44404 , \44406 );
nor \U$44091 ( \44408 , \44401 , \44407 );
or \U$44092 ( \44409 , \44276 , \44408 );
and \U$44093 ( \44410 , \35055 , \43809 );
nor \U$44094 ( \44411 , \44410 , \43817 );
or \U$44095 ( \44412 , \44271 , \44411 );
and \U$44096 ( \44413 , \35371 , \43822 );
nor \U$44097 ( \44414 , \44413 , \43828 );
nand \U$44098 ( \44415 , \44412 , \44414 );
and \U$44099 ( \44416 , \44275 , \44415 );
and \U$44100 ( \44417 , \35607 , \43833 );
nor \U$44101 ( \44418 , \44417 , \43840 );
or \U$44102 ( \44419 , \44274 , \44418 );
and \U$44103 ( \44420 , \35754 , \43845 );
nor \U$44104 ( \44421 , \44420 , \43851 );
nand \U$44105 ( \44422 , \44419 , \44421 );
nor \U$44106 ( \44423 , \44416 , \44422 );
nand \U$44107 ( \44424 , \44409 , \44423 );
nor \U$44108 ( \44425 , \44394 , \44424 );
nand \U$44109 ( \44426 , \44363 , \44425 );
not \U$44110 ( \44427 , \44426 );
xor \U$44111 ( \44428 , \44247 , \44427 );
buf \U$44112 ( \44429 , \44428 );
_HMUX rb5a9 ( \44430_nRb5a9 , \44245 , \44429 , RIc0c97c8_1 );
buf \U$44113 ( \44431 , \44430_nRb5a9 );
xor \U$44114 ( \44432 , \524 , \21581 );
buf \U$44115 ( \44433 , \44432 );
not \U$44116 ( \44434 , \35753 );
nand \U$44117 ( \44435 , \43850 , \44434 );
nand \U$44118 ( \44436 , \43961 , \43872 );
nand \U$44119 ( \44437 , \43873 , \43875 );
nor \U$44120 ( \44438 , \44436 , \44437 );
nand \U$44121 ( \44439 , \43876 , \43879 );
nand \U$44122 ( \44440 , \43880 , \43882 );
nor \U$44123 ( \44441 , \44439 , \44440 );
nand \U$44124 ( \44442 , \44438 , \44441 );
nand \U$44125 ( \44443 , \43883 , \43887 );
nand \U$44126 ( \44444 , \43888 , \43890 );
nor \U$44127 ( \44445 , \44443 , \44444 );
nand \U$44128 ( \44446 , \43891 , \43894 );
nand \U$44129 ( \44447 , \43895 , \43897 );
nor \U$44130 ( \44448 , \44446 , \44447 );
nand \U$44131 ( \44449 , \44445 , \44448 );
nor \U$44132 ( \44450 , \44442 , \44449 );
nand \U$44133 ( \44451 , \43898 , \43903 );
nand \U$44134 ( \44452 , \43904 , \43906 );
nor \U$44135 ( \44453 , \44451 , \44452 );
nand \U$44136 ( \44454 , \43907 , \43910 );
nand \U$44137 ( \44455 , \43911 , \43913 );
nor \U$44138 ( \44456 , \44454 , \44455 );
nand \U$44139 ( \44457 , \44453 , \44456 );
nand \U$44140 ( \44458 , \43914 , \43918 );
nand \U$44141 ( \44459 , \43919 , \43921 );
nor \U$44142 ( \44460 , \44458 , \44459 );
nand \U$44143 ( \44461 , \43922 , \43925 );
nand \U$44144 ( \44462 , \43926 , \43928 );
nor \U$44145 ( \44463 , \44461 , \44462 );
nand \U$44146 ( \44464 , \44460 , \44463 );
nor \U$44147 ( \44465 , \44457 , \44464 );
nand \U$44148 ( \44466 , \44450 , \44465 );
nand \U$44149 ( \44467 , \43977 , \43935 );
nand \U$44150 ( \44468 , \43936 , \43938 );
nor \U$44151 ( \44469 , \44467 , \44468 );
nand \U$44152 ( \44470 , \43939 , \43942 );
nand \U$44153 ( \44471 , \43943 , \43945 );
nor \U$44154 ( \44472 , \44470 , \44471 );
nand \U$44155 ( \44473 , \44469 , \44472 );
nand \U$44156 ( \44474 , \43946 , \43950 );
nand \U$44157 ( \44475 , \43951 , \43953 );
nor \U$44158 ( \44476 , \44474 , \44475 );
nand \U$44159 ( \44477 , \43954 , \43957 );
nand \U$44160 ( \44478 , \43958 , \43960 );
nor \U$44161 ( \44479 , \44477 , \44478 );
nand \U$44162 ( \44480 , \44476 , \44479 );
nor \U$44163 ( \44481 , \44473 , \44480 );
nand \U$44164 ( \44482 , \43985 , \43966 );
nand \U$44165 ( \44483 , \43967 , \43969 );
nor \U$44166 ( \44484 , \44482 , \44483 );
nand \U$44167 ( \44485 , \43970 , \43973 );
nand \U$44168 ( \44486 , \43974 , \43976 );
nor \U$44169 ( \44487 , \44485 , \44486 );
nand \U$44170 ( \44488 , \44484 , \44487 );
nand \U$44171 ( \44489 , \43989 , \43981 );
nand \U$44172 ( \44490 , \43982 , \43984 );
nor \U$44173 ( \44491 , \44489 , \44490 );
not \U$44174 ( \44492 , \43486 );
and \U$44175 ( \44493 , \43988 , \44492 );
nor \U$44176 ( \44494 , \44493 , \43993 );
not \U$44177 ( \44495 , \44494 );
and \U$44178 ( \44496 , \44491 , \44495 );
and \U$44179 ( \44497 , \43981 , \43996 );
nor \U$44180 ( \44498 , \44497 , \44001 );
or \U$44181 ( \44499 , \44490 , \44498 );
and \U$44182 ( \44500 , \43984 , \44004 );
nor \U$44183 ( \44501 , \44500 , \44008 );
nand \U$44184 ( \44502 , \44499 , \44501 );
nor \U$44185 ( \44503 , \44496 , \44502 );
or \U$44186 ( \44504 , \44488 , \44503 );
and \U$44187 ( \44505 , \43966 , \44011 );
nor \U$44188 ( \44506 , \44505 , \44017 );
or \U$44189 ( \44507 , \44483 , \44506 );
and \U$44190 ( \44508 , \43969 , \44020 );
nor \U$44191 ( \44509 , \44508 , \44024 );
nand \U$44192 ( \44510 , \44507 , \44509 );
and \U$44193 ( \44511 , \44487 , \44510 );
and \U$44194 ( \44512 , \43973 , \44027 );
nor \U$44195 ( \44513 , \44512 , \44032 );
or \U$44196 ( \44514 , \44486 , \44513 );
and \U$44197 ( \44515 , \43976 , \44035 );
nor \U$44198 ( \44516 , \44515 , \44039 );
nand \U$44199 ( \44517 , \44514 , \44516 );
nor \U$44200 ( \44518 , \44511 , \44517 );
nand \U$44201 ( \44519 , \44504 , \44518 );
and \U$44202 ( \44520 , \44481 , \44519 );
and \U$44203 ( \44521 , \43935 , \44042 );
nor \U$44204 ( \44522 , \44521 , \44049 );
or \U$44205 ( \44523 , \44468 , \44522 );
and \U$44206 ( \44524 , \43938 , \44052 );
nor \U$44207 ( \44525 , \44524 , \44056 );
nand \U$44208 ( \44526 , \44523 , \44525 );
and \U$44209 ( \44527 , \44472 , \44526 );
and \U$44210 ( \44528 , \43942 , \44059 );
nor \U$44211 ( \44529 , \44528 , \44064 );
or \U$44212 ( \44530 , \44471 , \44529 );
and \U$44213 ( \44531 , \43945 , \44067 );
nor \U$44214 ( \44532 , \44531 , \44071 );
nand \U$44215 ( \44533 , \44530 , \44532 );
nor \U$44216 ( \44534 , \44527 , \44533 );
or \U$44217 ( \44535 , \44480 , \44534 );
and \U$44218 ( \44536 , \43950 , \44074 );
nor \U$44219 ( \44537 , \44536 , \44080 );
or \U$44220 ( \44538 , \44475 , \44537 );
and \U$44221 ( \44539 , \43953 , \44083 );
nor \U$44222 ( \44540 , \44539 , \44087 );
nand \U$44223 ( \44541 , \44538 , \44540 );
and \U$44224 ( \44542 , \44479 , \44541 );
and \U$44225 ( \44543 , \43957 , \44090 );
nor \U$44226 ( \44544 , \44543 , \44095 );
or \U$44227 ( \44545 , \44478 , \44544 );
and \U$44228 ( \44546 , \43960 , \44098 );
nor \U$44229 ( \44547 , \44546 , \44102 );
nand \U$44230 ( \44548 , \44545 , \44547 );
nor \U$44231 ( \44549 , \44542 , \44548 );
nand \U$44232 ( \44550 , \44535 , \44549 );
nor \U$44233 ( \44551 , \44520 , \44550 );
or \U$44234 ( \44552 , \44466 , \44551 );
and \U$44235 ( \44553 , \43872 , \44105 );
nor \U$44236 ( \44554 , \44553 , \44113 );
or \U$44237 ( \44555 , \44437 , \44554 );
and \U$44238 ( \44556 , \43875 , \44116 );
nor \U$44239 ( \44557 , \44556 , \44120 );
nand \U$44240 ( \44558 , \44555 , \44557 );
and \U$44241 ( \44559 , \44441 , \44558 );
and \U$44242 ( \44560 , \43879 , \44123 );
nor \U$44243 ( \44561 , \44560 , \44128 );
or \U$44244 ( \44562 , \44440 , \44561 );
and \U$44245 ( \44563 , \43882 , \44131 );
nor \U$44246 ( \44564 , \44563 , \44135 );
nand \U$44247 ( \44565 , \44562 , \44564 );
nor \U$44248 ( \44566 , \44559 , \44565 );
or \U$44249 ( \44567 , \44449 , \44566 );
and \U$44250 ( \44568 , \43887 , \44138 );
nor \U$44251 ( \44569 , \44568 , \44144 );
or \U$44252 ( \44570 , \44444 , \44569 );
and \U$44253 ( \44571 , \43890 , \44147 );
nor \U$44254 ( \44572 , \44571 , \44151 );
nand \U$44255 ( \44573 , \44570 , \44572 );
and \U$44256 ( \44574 , \44448 , \44573 );
and \U$44257 ( \44575 , \43894 , \44154 );
nor \U$44258 ( \44576 , \44575 , \44159 );
or \U$44259 ( \44577 , \44447 , \44576 );
and \U$44260 ( \44578 , \43897 , \44162 );
nor \U$44261 ( \44579 , \44578 , \44166 );
nand \U$44262 ( \44580 , \44577 , \44579 );
nor \U$44263 ( \44581 , \44574 , \44580 );
nand \U$44264 ( \44582 , \44567 , \44581 );
and \U$44265 ( \44583 , \44465 , \44582 );
and \U$44266 ( \44584 , \43903 , \44169 );
nor \U$44267 ( \44585 , \44584 , \44176 );
or \U$44268 ( \44586 , \44452 , \44585 );
and \U$44269 ( \44587 , \43906 , \44179 );
nor \U$44270 ( \44588 , \44587 , \44183 );
nand \U$44271 ( \44589 , \44586 , \44588 );
and \U$44272 ( \44590 , \44456 , \44589 );
and \U$44273 ( \44591 , \43910 , \44186 );
nor \U$44274 ( \44592 , \44591 , \44191 );
or \U$44275 ( \44593 , \44455 , \44592 );
and \U$44276 ( \44594 , \43913 , \44194 );
nor \U$44277 ( \44595 , \44594 , \44198 );
nand \U$44278 ( \44596 , \44593 , \44595 );
nor \U$44279 ( \44597 , \44590 , \44596 );
or \U$44280 ( \44598 , \44464 , \44597 );
and \U$44281 ( \44599 , \43918 , \44201 );
nor \U$44282 ( \44600 , \44599 , \44207 );
or \U$44283 ( \44601 , \44459 , \44600 );
and \U$44284 ( \44602 , \43921 , \44210 );
nor \U$44285 ( \44603 , \44602 , \44214 );
nand \U$44286 ( \44604 , \44601 , \44603 );
and \U$44287 ( \44605 , \44463 , \44604 );
and \U$44288 ( \44606 , \43925 , \44217 );
nor \U$44289 ( \44607 , \44606 , \44222 );
or \U$44290 ( \44608 , \44462 , \44607 );
and \U$44291 ( \44609 , \43928 , \44225 );
nor \U$44292 ( \44610 , \44609 , \44229 );
nand \U$44293 ( \44611 , \44608 , \44610 );
nor \U$44294 ( \44612 , \44605 , \44611 );
nand \U$44295 ( \44613 , \44598 , \44612 );
nor \U$44296 ( \44614 , \44583 , \44613 );
nand \U$44297 ( \44615 , \44552 , \44614 );
not \U$44298 ( \44616 , \44615 );
xor \U$44299 ( \44617 , \44435 , \44616 );
buf \U$44300 ( \44618 , \44617 );
_HMUX rb55a ( \44619_nRb55a , \44433 , \44618 , RIc0c97c8_1 );
buf \U$44301 ( \44620 , \44619_nRb55a );
xor \U$44302 ( \44621 , \574 , \21579 );
buf \U$44303 ( \44622 , \44621 );
not \U$44304 ( \44623 , \35731 );
nand \U$44305 ( \44624 , \43848 , \44623 );
nor \U$44306 ( \44625 , \41859 , \25670 );
nor \U$44307 ( \44626 , \26900 , \28053 );
nand \U$44308 ( \44627 , \44625 , \44626 );
nor \U$44309 ( \44628 , \29122 , \30120 );
nor \U$44310 ( \44629 , \31044 , \31883 );
nand \U$44311 ( \44630 , \44628 , \44629 );
nor \U$44312 ( \44631 , \44627 , \44630 );
nor \U$44313 ( \44632 , \32639 , \33310 );
nor \U$44314 ( \44633 , \33914 , \34433 );
nand \U$44315 ( \44634 , \44632 , \44633 );
nor \U$44316 ( \44635 , \34866 , \35223 );
nor \U$44317 ( \44636 , \35499 , \35696 );
nand \U$44318 ( \44637 , \44635 , \44636 );
nor \U$44319 ( \44638 , \44634 , \44637 );
nand \U$44320 ( \44639 , \44631 , \44638 );
nor \U$44321 ( \44640 , \43172 , \37016 );
nor \U$44322 ( \44641 , \37731 , \38527 );
nand \U$44323 ( \44642 , \44640 , \44641 );
nor \U$44324 ( \44643 , \39404 , \40361 );
nor \U$44325 ( \44644 , \41396 , \41786 );
nand \U$44326 ( \44645 , \44643 , \44644 );
nor \U$44327 ( \44646 , \44642 , \44645 );
nor \U$44328 ( \44647 , \43427 , \42347 );
nor \U$44329 ( \44648 , \42742 , \43090 );
nand \U$44330 ( \44649 , \44647 , \44648 );
nor \U$44331 ( \44650 , \43474 , \43362 );
and \U$44332 ( \44651 , \44650 , \43489 );
or \U$44333 ( \44652 , \43362 , \43501 );
nand \U$44334 ( \44653 , \44652 , \43513 );
nor \U$44335 ( \44654 , \44651 , \44653 );
or \U$44336 ( \44655 , \44649 , \44654 );
or \U$44337 ( \44656 , \42347 , \43524 );
nand \U$44338 ( \44657 , \44656 , \43537 );
and \U$44339 ( \44658 , \44648 , \44657 );
or \U$44340 ( \44659 , \43090 , \43548 );
nand \U$44341 ( \44660 , \44659 , \43560 );
nor \U$44342 ( \44661 , \44658 , \44660 );
nand \U$44343 ( \44662 , \44655 , \44661 );
and \U$44344 ( \44663 , \44646 , \44662 );
or \U$44345 ( \44664 , \37016 , \43571 );
nand \U$44346 ( \44665 , \44664 , \43585 );
and \U$44347 ( \44666 , \44641 , \44665 );
or \U$44348 ( \44667 , \38527 , \43596 );
nand \U$44349 ( \44668 , \44667 , \43608 );
nor \U$44350 ( \44669 , \44666 , \44668 );
or \U$44351 ( \44670 , \44645 , \44669 );
or \U$44352 ( \44671 , \40361 , \43619 );
nand \U$44353 ( \44672 , \44671 , \43632 );
and \U$44354 ( \44673 , \44644 , \44672 );
or \U$44355 ( \44674 , \41786 , \43643 );
nand \U$44356 ( \44675 , \44674 , \43655 );
nor \U$44357 ( \44676 , \44673 , \44675 );
nand \U$44358 ( \44677 , \44670 , \44676 );
nor \U$44359 ( \44678 , \44663 , \44677 );
or \U$44360 ( \44679 , \44639 , \44678 );
or \U$44361 ( \44680 , \25670 , \43666 );
nand \U$44362 ( \44681 , \44680 , \43681 );
and \U$44363 ( \44682 , \44626 , \44681 );
or \U$44364 ( \44683 , \28053 , \43692 );
nand \U$44365 ( \44684 , \44683 , \43704 );
nor \U$44366 ( \44685 , \44682 , \44684 );
or \U$44367 ( \44686 , \44630 , \44685 );
or \U$44368 ( \44687 , \30120 , \43715 );
nand \U$44369 ( \44688 , \44687 , \43728 );
and \U$44370 ( \44689 , \44629 , \44688 );
or \U$44371 ( \44690 , \31883 , \43739 );
nand \U$44372 ( \44691 , \44690 , \43751 );
nor \U$44373 ( \44692 , \44689 , \44691 );
nand \U$44374 ( \44693 , \44686 , \44692 );
and \U$44375 ( \44694 , \44638 , \44693 );
or \U$44376 ( \44695 , \33310 , \43762 );
nand \U$44377 ( \44696 , \44695 , \43776 );
and \U$44378 ( \44697 , \44633 , \44696 );
or \U$44379 ( \44698 , \34433 , \43787 );
nand \U$44380 ( \44699 , \44698 , \43799 );
nor \U$44381 ( \44700 , \44697 , \44699 );
or \U$44382 ( \44701 , \44637 , \44700 );
or \U$44383 ( \44702 , \35223 , \43810 );
nand \U$44384 ( \44703 , \44702 , \43823 );
and \U$44385 ( \44704 , \44636 , \44703 );
or \U$44386 ( \44705 , \35696 , \43834 );
nand \U$44387 ( \44706 , \44705 , \43846 );
nor \U$44388 ( \44707 , \44704 , \44706 );
nand \U$44389 ( \44708 , \44701 , \44707 );
nor \U$44390 ( \44709 , \44694 , \44708 );
nand \U$44391 ( \44710 , \44679 , \44709 );
not \U$44392 ( \44711 , \44710 );
xor \U$44393 ( \44712 , \44624 , \44711 );
buf \U$44394 ( \44713 , \44712 );
_HMUX rb500 ( \44714_nRb500 , \44622 , \44713 , RIc0c97c8_1 );
buf \U$44395 ( \44715 , \44714_nRb500 );
xor \U$44396 ( \44716 , \627 , \21577 );
buf \U$44397 ( \44717 , \44716 );
not \U$44398 ( \44718 , \35694 );
nand \U$44399 ( \44719 , \43844 , \44718 );
nor \U$44400 ( \44720 , \43962 , \43874 );
nor \U$44401 ( \44721 , \43877 , \43881 );
nand \U$44402 ( \44722 , \44720 , \44721 );
nor \U$44403 ( \44723 , \43884 , \43889 );
nor \U$44404 ( \44724 , \43892 , \43896 );
nand \U$44405 ( \44725 , \44723 , \44724 );
nor \U$44406 ( \44726 , \44722 , \44725 );
nor \U$44407 ( \44727 , \43899 , \43905 );
nor \U$44408 ( \44728 , \43908 , \43912 );
nand \U$44409 ( \44729 , \44727 , \44728 );
nor \U$44410 ( \44730 , \43915 , \43920 );
nor \U$44411 ( \44731 , \43923 , \43927 );
nand \U$44412 ( \44732 , \44730 , \44731 );
nor \U$44413 ( \44733 , \44729 , \44732 );
nand \U$44414 ( \44734 , \44726 , \44733 );
nor \U$44415 ( \44735 , \43978 , \43937 );
nor \U$44416 ( \44736 , \43940 , \43944 );
nand \U$44417 ( \44737 , \44735 , \44736 );
nor \U$44418 ( \44738 , \43947 , \43952 );
nor \U$44419 ( \44739 , \43955 , \43959 );
nand \U$44420 ( \44740 , \44738 , \44739 );
nor \U$44421 ( \44741 , \44737 , \44740 );
nor \U$44422 ( \44742 , \43986 , \43968 );
nor \U$44423 ( \44743 , \43971 , \43975 );
nand \U$44424 ( \44744 , \44742 , \44743 );
nor \U$44425 ( \44745 , \43990 , \43983 );
and \U$44426 ( \44746 , \44745 , \44492 );
or \U$44427 ( \44747 , \43983 , \43997 );
nand \U$44428 ( \44748 , \44747 , \44005 );
nor \U$44429 ( \44749 , \44746 , \44748 );
or \U$44430 ( \44750 , \44744 , \44749 );
or \U$44431 ( \44751 , \43968 , \44012 );
nand \U$44432 ( \44752 , \44751 , \44021 );
and \U$44433 ( \44753 , \44743 , \44752 );
or \U$44434 ( \44754 , \43975 , \44028 );
nand \U$44435 ( \44755 , \44754 , \44036 );
nor \U$44436 ( \44756 , \44753 , \44755 );
nand \U$44437 ( \44757 , \44750 , \44756 );
and \U$44438 ( \44758 , \44741 , \44757 );
or \U$44439 ( \44759 , \43937 , \44043 );
nand \U$44440 ( \44760 , \44759 , \44053 );
and \U$44441 ( \44761 , \44736 , \44760 );
or \U$44442 ( \44762 , \43944 , \44060 );
nand \U$44443 ( \44763 , \44762 , \44068 );
nor \U$44444 ( \44764 , \44761 , \44763 );
or \U$44445 ( \44765 , \44740 , \44764 );
or \U$44446 ( \44766 , \43952 , \44075 );
nand \U$44447 ( \44767 , \44766 , \44084 );
and \U$44448 ( \44768 , \44739 , \44767 );
or \U$44449 ( \44769 , \43959 , \44091 );
nand \U$44450 ( \44770 , \44769 , \44099 );
nor \U$44451 ( \44771 , \44768 , \44770 );
nand \U$44452 ( \44772 , \44765 , \44771 );
nor \U$44453 ( \44773 , \44758 , \44772 );
or \U$44454 ( \44774 , \44734 , \44773 );
or \U$44455 ( \44775 , \43874 , \44106 );
nand \U$44456 ( \44776 , \44775 , \44117 );
and \U$44457 ( \44777 , \44721 , \44776 );
or \U$44458 ( \44778 , \43881 , \44124 );
nand \U$44459 ( \44779 , \44778 , \44132 );
nor \U$44460 ( \44780 , \44777 , \44779 );
or \U$44461 ( \44781 , \44725 , \44780 );
or \U$44462 ( \44782 , \43889 , \44139 );
nand \U$44463 ( \44783 , \44782 , \44148 );
and \U$44464 ( \44784 , \44724 , \44783 );
or \U$44465 ( \44785 , \43896 , \44155 );
nand \U$44466 ( \44786 , \44785 , \44163 );
nor \U$44467 ( \44787 , \44784 , \44786 );
nand \U$44468 ( \44788 , \44781 , \44787 );
and \U$44469 ( \44789 , \44733 , \44788 );
or \U$44470 ( \44790 , \43905 , \44170 );
nand \U$44471 ( \44791 , \44790 , \44180 );
and \U$44472 ( \44792 , \44728 , \44791 );
or \U$44473 ( \44793 , \43912 , \44187 );
nand \U$44474 ( \44794 , \44793 , \44195 );
nor \U$44475 ( \44795 , \44792 , \44794 );
or \U$44476 ( \44796 , \44732 , \44795 );
or \U$44477 ( \44797 , \43920 , \44202 );
nand \U$44478 ( \44798 , \44797 , \44211 );
and \U$44479 ( \44799 , \44731 , \44798 );
or \U$44480 ( \44800 , \43927 , \44218 );
nand \U$44481 ( \44801 , \44800 , \44226 );
nor \U$44482 ( \44802 , \44799 , \44801 );
nand \U$44483 ( \44803 , \44796 , \44802 );
nor \U$44484 ( \44804 , \44789 , \44803 );
nand \U$44485 ( \44805 , \44774 , \44804 );
not \U$44486 ( \44806 , \44805 );
xor \U$44487 ( \44807 , \44719 , \44806 );
buf \U$44488 ( \44808 , \44807 );
_HMUX rb49d ( \44809_nRb49d , \44717 , \44808 , RIc0c97c8_1 );
buf \U$44489 ( \44810 , \44809_nRb49d );
xor \U$44490 ( \44811 , \747 , \21575 );
buf \U$44491 ( \44812 , \44811 );
not \U$44492 ( \44813 , \35654 );
nand \U$44493 ( \44814 , \43842 , \44813 );
nor \U$44494 ( \44815 , \44290 , \44248 );
nor \U$44495 ( \44816 , \44249 , \44251 );
nand \U$44496 ( \44817 , \44815 , \44816 );
nor \U$44497 ( \44818 , \44252 , \44255 );
nor \U$44498 ( \44819 , \44256 , \44258 );
nand \U$44499 ( \44820 , \44818 , \44819 );
nor \U$44500 ( \44821 , \44817 , \44820 );
nor \U$44501 ( \44822 , \44259 , \44263 );
nor \U$44502 ( \44823 , \44264 , \44266 );
nand \U$44503 ( \44824 , \44822 , \44823 );
nor \U$44504 ( \44825 , \44267 , \44270 );
nor \U$44505 ( \44826 , \44271 , \44273 );
nand \U$44506 ( \44827 , \44825 , \44826 );
nor \U$44507 ( \44828 , \44824 , \44827 );
nand \U$44508 ( \44829 , \44821 , \44828 );
nor \U$44509 ( \44830 , \44298 , \44279 );
nor \U$44510 ( \44831 , \44280 , \44282 );
nand \U$44511 ( \44832 , \44830 , \44831 );
nor \U$44512 ( \44833 , \44283 , \44286 );
nor \U$44513 ( \44834 , \44287 , \44289 );
nand \U$44514 ( \44835 , \44833 , \44834 );
nor \U$44515 ( \44836 , \44832 , \44835 );
nor \U$44516 ( \44837 , \44302 , \44294 );
nor \U$44517 ( \44838 , \44295 , \44297 );
nand \U$44518 ( \44839 , \44837 , \44838 );
or \U$44519 ( \44840 , \44301 , \44305 );
nand \U$44520 ( \44841 , \44840 , \44309 );
not \U$44521 ( \44842 , \44841 );
or \U$44522 ( \44843 , \44839 , \44842 );
or \U$44523 ( \44844 , \44294 , \44312 );
nand \U$44524 ( \44845 , \44844 , \44317 );
and \U$44525 ( \44846 , \44838 , \44845 );
or \U$44526 ( \44847 , \44297 , \44320 );
nand \U$44527 ( \44848 , \44847 , \44324 );
nor \U$44528 ( \44849 , \44846 , \44848 );
nand \U$44529 ( \44850 , \44843 , \44849 );
and \U$44530 ( \44851 , \44836 , \44850 );
or \U$44531 ( \44852 , \44279 , \44327 );
nand \U$44532 ( \44853 , \44852 , \44333 );
and \U$44533 ( \44854 , \44831 , \44853 );
or \U$44534 ( \44855 , \44282 , \44336 );
nand \U$44535 ( \44856 , \44855 , \44340 );
nor \U$44536 ( \44857 , \44854 , \44856 );
or \U$44537 ( \44858 , \44835 , \44857 );
or \U$44538 ( \44859 , \44286 , \44343 );
nand \U$44539 ( \44860 , \44859 , \44348 );
and \U$44540 ( \44861 , \44834 , \44860 );
or \U$44541 ( \44862 , \44289 , \44351 );
nand \U$44542 ( \44863 , \44862 , \44355 );
nor \U$44543 ( \44864 , \44861 , \44863 );
nand \U$44544 ( \44865 , \44858 , \44864 );
nor \U$44545 ( \44866 , \44851 , \44865 );
or \U$44546 ( \44867 , \44829 , \44866 );
or \U$44547 ( \44868 , \44248 , \44358 );
nand \U$44548 ( \44869 , \44868 , \44365 );
and \U$44549 ( \44870 , \44816 , \44869 );
or \U$44550 ( \44871 , \44251 , \44368 );
nand \U$44551 ( \44872 , \44871 , \44372 );
nor \U$44552 ( \44873 , \44870 , \44872 );
or \U$44553 ( \44874 , \44820 , \44873 );
or \U$44554 ( \44875 , \44255 , \44375 );
nand \U$44555 ( \44876 , \44875 , \44380 );
and \U$44556 ( \44877 , \44819 , \44876 );
or \U$44557 ( \44878 , \44258 , \44383 );
nand \U$44558 ( \44879 , \44878 , \44387 );
nor \U$44559 ( \44880 , \44877 , \44879 );
nand \U$44560 ( \44881 , \44874 , \44880 );
and \U$44561 ( \44882 , \44828 , \44881 );
or \U$44562 ( \44883 , \44263 , \44390 );
nand \U$44563 ( \44884 , \44883 , \44396 );
and \U$44564 ( \44885 , \44823 , \44884 );
or \U$44565 ( \44886 , \44266 , \44399 );
nand \U$44566 ( \44887 , \44886 , \44403 );
nor \U$44567 ( \44888 , \44885 , \44887 );
or \U$44568 ( \44889 , \44827 , \44888 );
or \U$44569 ( \44890 , \44270 , \44406 );
nand \U$44570 ( \44891 , \44890 , \44411 );
and \U$44571 ( \44892 , \44826 , \44891 );
or \U$44572 ( \44893 , \44273 , \44414 );
nand \U$44573 ( \44894 , \44893 , \44418 );
nor \U$44574 ( \44895 , \44892 , \44894 );
nand \U$44575 ( \44896 , \44889 , \44895 );
nor \U$44576 ( \44897 , \44882 , \44896 );
nand \U$44577 ( \44898 , \44867 , \44897 );
not \U$44578 ( \44899 , \44898 );
xor \U$44579 ( \44900 , \44814 , \44899 );
buf \U$44580 ( \44901 , \44900 );
_HMUX rb432 ( \44902_nRb432 , \44812 , \44901 , RIc0c97c8_1 );
buf \U$44581 ( \44903 , \44902_nRb432 );
xor \U$44582 ( \44904 , \821 , \21573 );
buf \U$44583 ( \44905 , \44904 );
not \U$44584 ( \44906 , \35606 );
nand \U$44585 ( \44907 , \43839 , \44906 );
nor \U$44586 ( \44908 , \44478 , \44436 );
nor \U$44587 ( \44909 , \44437 , \44439 );
nand \U$44588 ( \44910 , \44908 , \44909 );
nor \U$44589 ( \44911 , \44440 , \44443 );
nor \U$44590 ( \44912 , \44444 , \44446 );
nand \U$44591 ( \44913 , \44911 , \44912 );
nor \U$44592 ( \44914 , \44910 , \44913 );
nor \U$44593 ( \44915 , \44447 , \44451 );
nor \U$44594 ( \44916 , \44452 , \44454 );
nand \U$44595 ( \44917 , \44915 , \44916 );
nor \U$44596 ( \44918 , \44455 , \44458 );
nor \U$44597 ( \44919 , \44459 , \44461 );
nand \U$44598 ( \44920 , \44918 , \44919 );
nor \U$44599 ( \44921 , \44917 , \44920 );
nand \U$44600 ( \44922 , \44914 , \44921 );
nor \U$44601 ( \44923 , \44486 , \44467 );
nor \U$44602 ( \44924 , \44468 , \44470 );
nand \U$44603 ( \44925 , \44923 , \44924 );
nor \U$44604 ( \44926 , \44471 , \44474 );
nor \U$44605 ( \44927 , \44475 , \44477 );
nand \U$44606 ( \44928 , \44926 , \44927 );
nor \U$44607 ( \44929 , \44925 , \44928 );
nor \U$44608 ( \44930 , \44490 , \44482 );
nor \U$44609 ( \44931 , \44483 , \44485 );
nand \U$44610 ( \44932 , \44930 , \44931 );
or \U$44611 ( \44933 , \44489 , \44494 );
nand \U$44612 ( \44934 , \44933 , \44498 );
not \U$44613 ( \44935 , \44934 );
or \U$44614 ( \44936 , \44932 , \44935 );
or \U$44615 ( \44937 , \44482 , \44501 );
nand \U$44616 ( \44938 , \44937 , \44506 );
and \U$44617 ( \44939 , \44931 , \44938 );
or \U$44618 ( \44940 , \44485 , \44509 );
nand \U$44619 ( \44941 , \44940 , \44513 );
nor \U$44620 ( \44942 , \44939 , \44941 );
nand \U$44621 ( \44943 , \44936 , \44942 );
and \U$44622 ( \44944 , \44929 , \44943 );
or \U$44623 ( \44945 , \44467 , \44516 );
nand \U$44624 ( \44946 , \44945 , \44522 );
and \U$44625 ( \44947 , \44924 , \44946 );
or \U$44626 ( \44948 , \44470 , \44525 );
nand \U$44627 ( \44949 , \44948 , \44529 );
nor \U$44628 ( \44950 , \44947 , \44949 );
or \U$44629 ( \44951 , \44928 , \44950 );
or \U$44630 ( \44952 , \44474 , \44532 );
nand \U$44631 ( \44953 , \44952 , \44537 );
and \U$44632 ( \44954 , \44927 , \44953 );
or \U$44633 ( \44955 , \44477 , \44540 );
nand \U$44634 ( \44956 , \44955 , \44544 );
nor \U$44635 ( \44957 , \44954 , \44956 );
nand \U$44636 ( \44958 , \44951 , \44957 );
nor \U$44637 ( \44959 , \44944 , \44958 );
or \U$44638 ( \44960 , \44922 , \44959 );
or \U$44639 ( \44961 , \44436 , \44547 );
nand \U$44640 ( \44962 , \44961 , \44554 );
and \U$44641 ( \44963 , \44909 , \44962 );
or \U$44642 ( \44964 , \44439 , \44557 );
nand \U$44643 ( \44965 , \44964 , \44561 );
nor \U$44644 ( \44966 , \44963 , \44965 );
or \U$44645 ( \44967 , \44913 , \44966 );
or \U$44646 ( \44968 , \44443 , \44564 );
nand \U$44647 ( \44969 , \44968 , \44569 );
and \U$44648 ( \44970 , \44912 , \44969 );
or \U$44649 ( \44971 , \44446 , \44572 );
nand \U$44650 ( \44972 , \44971 , \44576 );
nor \U$44651 ( \44973 , \44970 , \44972 );
nand \U$44652 ( \44974 , \44967 , \44973 );
and \U$44653 ( \44975 , \44921 , \44974 );
or \U$44654 ( \44976 , \44451 , \44579 );
nand \U$44655 ( \44977 , \44976 , \44585 );
and \U$44656 ( \44978 , \44916 , \44977 );
or \U$44657 ( \44979 , \44454 , \44588 );
nand \U$44658 ( \44980 , \44979 , \44592 );
nor \U$44659 ( \44981 , \44978 , \44980 );
or \U$44660 ( \44982 , \44920 , \44981 );
or \U$44661 ( \44983 , \44458 , \44595 );
nand \U$44662 ( \44984 , \44983 , \44600 );
and \U$44663 ( \44985 , \44919 , \44984 );
or \U$44664 ( \44986 , \44461 , \44603 );
nand \U$44665 ( \44987 , \44986 , \44607 );
nor \U$44666 ( \44988 , \44985 , \44987 );
nand \U$44667 ( \44989 , \44982 , \44988 );
nor \U$44668 ( \44990 , \44975 , \44989 );
nand \U$44669 ( \44991 , \44960 , \44990 );
not \U$44670 ( \44992 , \44991 );
xor \U$44671 ( \44993 , \44907 , \44992 );
buf \U$44672 ( \44994 , \44993 );
_HMUX rb3bb ( \44995_nRb3bb , \44905 , \44994 , RIc0c97c8_1 );
buf \U$44673 ( \44996 , \44995_nRb3bb );
xor \U$44674 ( \44997 , \896 , \21571 );
buf \U$44675 ( \44998 , \44997 );
not \U$44676 ( \44999 , \35557 );
nand \U$44677 ( \45000 , \43837 , \44999 );
nand \U$44678 ( \45001 , \41860 , \26901 );
nand \U$44679 ( \45002 , \29123 , \31045 );
nor \U$44680 ( \45003 , \45001 , \45002 );
nand \U$44681 ( \45004 , \32640 , \33915 );
nand \U$44682 ( \45005 , \34867 , \35500 );
nor \U$44683 ( \45006 , \45004 , \45005 );
nand \U$44684 ( \45007 , \45003 , \45006 );
nand \U$44685 ( \45008 , \43173 , \37732 );
nand \U$44686 ( \45009 , \39405 , \41397 );
nor \U$44687 ( \45010 , \45008 , \45009 );
nand \U$44688 ( \45011 , \43428 , \42743 );
not \U$44689 ( \45012 , \43502 );
or \U$44690 ( \45013 , \45011 , \45012 );
and \U$44691 ( \45014 , \42743 , \43525 );
nor \U$44692 ( \45015 , \45014 , \43549 );
nand \U$44693 ( \45016 , \45013 , \45015 );
and \U$44694 ( \45017 , \45010 , \45016 );
and \U$44695 ( \45018 , \37732 , \43572 );
nor \U$44696 ( \45019 , \45018 , \43597 );
or \U$44697 ( \45020 , \45009 , \45019 );
and \U$44698 ( \45021 , \41397 , \43620 );
nor \U$44699 ( \45022 , \45021 , \43644 );
nand \U$44700 ( \45023 , \45020 , \45022 );
nor \U$44701 ( \45024 , \45017 , \45023 );
or \U$44702 ( \45025 , \45007 , \45024 );
and \U$44703 ( \45026 , \26901 , \43667 );
nor \U$44704 ( \45027 , \45026 , \43693 );
or \U$44705 ( \45028 , \45002 , \45027 );
and \U$44706 ( \45029 , \31045 , \43716 );
nor \U$44707 ( \45030 , \45029 , \43740 );
nand \U$44708 ( \45031 , \45028 , \45030 );
and \U$44709 ( \45032 , \45006 , \45031 );
and \U$44710 ( \45033 , \33915 , \43763 );
nor \U$44711 ( \45034 , \45033 , \43788 );
or \U$44712 ( \45035 , \45005 , \45034 );
and \U$44713 ( \45036 , \35500 , \43811 );
nor \U$44714 ( \45037 , \45036 , \43835 );
nand \U$44715 ( \45038 , \45035 , \45037 );
nor \U$44716 ( \45039 , \45032 , \45038 );
nand \U$44717 ( \45040 , \45025 , \45039 );
not \U$44718 ( \45041 , \45040 );
xor \U$44719 ( \45042 , \45000 , \45041 );
buf \U$44720 ( \45043 , \45042 );
_HMUX rb33b ( \45044_nRb33b , \44998 , \45043 , RIc0c97c8_1 );
buf \U$44721 ( \45045 , \45044_nRb33b );
xor \U$44722 ( \45046 , \977 , \21569 );
buf \U$44723 ( \45047 , \45046 );
not \U$44724 ( \45048 , \35497 );
nand \U$44725 ( \45049 , \43832 , \45048 );
nand \U$44726 ( \45050 , \43963 , \43878 );
nand \U$44727 ( \45051 , \43885 , \43893 );
nor \U$44728 ( \45052 , \45050 , \45051 );
nand \U$44729 ( \45053 , \43900 , \43909 );
nand \U$44730 ( \45054 , \43916 , \43924 );
nor \U$44731 ( \45055 , \45053 , \45054 );
nand \U$44732 ( \45056 , \45052 , \45055 );
nand \U$44733 ( \45057 , \43979 , \43941 );
nand \U$44734 ( \45058 , \43948 , \43956 );
nor \U$44735 ( \45059 , \45057 , \45058 );
nand \U$44736 ( \45060 , \43987 , \43972 );
not \U$44737 ( \45061 , \43998 );
or \U$44738 ( \45062 , \45060 , \45061 );
and \U$44739 ( \45063 , \43972 , \44013 );
nor \U$44740 ( \45064 , \45063 , \44029 );
nand \U$44741 ( \45065 , \45062 , \45064 );
and \U$44742 ( \45066 , \45059 , \45065 );
and \U$44743 ( \45067 , \43941 , \44044 );
nor \U$44744 ( \45068 , \45067 , \44061 );
or \U$44745 ( \45069 , \45058 , \45068 );
and \U$44746 ( \45070 , \43956 , \44076 );
nor \U$44747 ( \45071 , \45070 , \44092 );
nand \U$44748 ( \45072 , \45069 , \45071 );
nor \U$44749 ( \45073 , \45066 , \45072 );
or \U$44750 ( \45074 , \45056 , \45073 );
and \U$44751 ( \45075 , \43878 , \44107 );
nor \U$44752 ( \45076 , \45075 , \44125 );
or \U$44753 ( \45077 , \45051 , \45076 );
and \U$44754 ( \45078 , \43893 , \44140 );
nor \U$44755 ( \45079 , \45078 , \44156 );
nand \U$44756 ( \45080 , \45077 , \45079 );
and \U$44757 ( \45081 , \45055 , \45080 );
and \U$44758 ( \45082 , \43909 , \44171 );
nor \U$44759 ( \45083 , \45082 , \44188 );
or \U$44760 ( \45084 , \45054 , \45083 );
and \U$44761 ( \45085 , \43924 , \44203 );
nor \U$44762 ( \45086 , \45085 , \44219 );
nand \U$44763 ( \45087 , \45084 , \45086 );
nor \U$44764 ( \45088 , \45081 , \45087 );
nand \U$44765 ( \45089 , \45074 , \45088 );
not \U$44766 ( \45090 , \45089 );
xor \U$44767 ( \45091 , \45049 , \45090 );
buf \U$44768 ( \45092 , \45091 );
_HMUX rb2b1 ( \45093_nRb2b1 , \45047 , \45092 , RIc0c97c8_1 );
buf \U$44769 ( \45094 , \45093_nRb2b1 );
xor \U$44770 ( \45095 , \1060 , \21567 );
buf \U$44771 ( \45096 , \45095 );
not \U$44772 ( \45097 , \35436 );
nand \U$44773 ( \45098 , \43830 , \45097 );
nand \U$44774 ( \45099 , \44291 , \44250 );
nand \U$44775 ( \45100 , \44253 , \44257 );
nor \U$44776 ( \45101 , \45099 , \45100 );
nand \U$44777 ( \45102 , \44260 , \44265 );
nand \U$44778 ( \45103 , \44268 , \44272 );
nor \U$44779 ( \45104 , \45102 , \45103 );
nand \U$44780 ( \45105 , \45101 , \45104 );
nand \U$44781 ( \45106 , \44299 , \44281 );
nand \U$44782 ( \45107 , \44284 , \44288 );
nor \U$44783 ( \45108 , \45106 , \45107 );
nand \U$44784 ( \45109 , \44303 , \44296 );
or \U$44785 ( \45110 , \45109 , \44305 );
and \U$44786 ( \45111 , \44296 , \44313 );
nor \U$44787 ( \45112 , \45111 , \44321 );
nand \U$44788 ( \45113 , \45110 , \45112 );
and \U$44789 ( \45114 , \45108 , \45113 );
and \U$44790 ( \45115 , \44281 , \44328 );
nor \U$44791 ( \45116 , \45115 , \44337 );
or \U$44792 ( \45117 , \45107 , \45116 );
and \U$44793 ( \45118 , \44288 , \44344 );
nor \U$44794 ( \45119 , \45118 , \44352 );
nand \U$44795 ( \45120 , \45117 , \45119 );
nor \U$44796 ( \45121 , \45114 , \45120 );
or \U$44797 ( \45122 , \45105 , \45121 );
and \U$44798 ( \45123 , \44250 , \44359 );
nor \U$44799 ( \45124 , \45123 , \44369 );
or \U$44800 ( \45125 , \45100 , \45124 );
and \U$44801 ( \45126 , \44257 , \44376 );
nor \U$44802 ( \45127 , \45126 , \44384 );
nand \U$44803 ( \45128 , \45125 , \45127 );
and \U$44804 ( \45129 , \45104 , \45128 );
and \U$44805 ( \45130 , \44265 , \44391 );
nor \U$44806 ( \45131 , \45130 , \44400 );
or \U$44807 ( \45132 , \45103 , \45131 );
and \U$44808 ( \45133 , \44272 , \44407 );
nor \U$44809 ( \45134 , \45133 , \44415 );
nand \U$44810 ( \45135 , \45132 , \45134 );
nor \U$44811 ( \45136 , \45129 , \45135 );
nand \U$44812 ( \45137 , \45122 , \45136 );
not \U$44813 ( \45138 , \45137 );
xor \U$44814 ( \45139 , \45098 , \45138 );
buf \U$44815 ( \45140 , \45139 );
_HMUX rb21b ( \45141_nRb21b , \45096 , \45140 , RIc0c97c8_1 );
buf \U$44816 ( \45142 , \45141_nRb21b );
xor \U$44817 ( \45143 , \1139 , \21565 );
buf \U$44818 ( \45144 , \45143 );
not \U$44819 ( \45145 , \35370 );
nand \U$44820 ( \45146 , \43827 , \45145 );
nand \U$44821 ( \45147 , \44479 , \44438 );
nand \U$44822 ( \45148 , \44441 , \44445 );
nor \U$44823 ( \45149 , \45147 , \45148 );
nand \U$44824 ( \45150 , \44448 , \44453 );
nand \U$44825 ( \45151 , \44456 , \44460 );
nor \U$44826 ( \45152 , \45150 , \45151 );
nand \U$44827 ( \45153 , \45149 , \45152 );
nand \U$44828 ( \45154 , \44487 , \44469 );
nand \U$44829 ( \45155 , \44472 , \44476 );
nor \U$44830 ( \45156 , \45154 , \45155 );
nand \U$44831 ( \45157 , \44491 , \44484 );
or \U$44832 ( \45158 , \45157 , \44494 );
and \U$44833 ( \45159 , \44484 , \44502 );
nor \U$44834 ( \45160 , \45159 , \44510 );
nand \U$44835 ( \45161 , \45158 , \45160 );
and \U$44836 ( \45162 , \45156 , \45161 );
and \U$44837 ( \45163 , \44469 , \44517 );
nor \U$44838 ( \45164 , \45163 , \44526 );
or \U$44839 ( \45165 , \45155 , \45164 );
and \U$44840 ( \45166 , \44476 , \44533 );
nor \U$44841 ( \45167 , \45166 , \44541 );
nand \U$44842 ( \45168 , \45165 , \45167 );
nor \U$44843 ( \45169 , \45162 , \45168 );
or \U$44844 ( \45170 , \45153 , \45169 );
and \U$44845 ( \45171 , \44438 , \44548 );
nor \U$44846 ( \45172 , \45171 , \44558 );
or \U$44847 ( \45173 , \45148 , \45172 );
and \U$44848 ( \45174 , \44445 , \44565 );
nor \U$44849 ( \45175 , \45174 , \44573 );
nand \U$44850 ( \45176 , \45173 , \45175 );
and \U$44851 ( \45177 , \45152 , \45176 );
and \U$44852 ( \45178 , \44453 , \44580 );
nor \U$44853 ( \45179 , \45178 , \44589 );
or \U$44854 ( \45180 , \45151 , \45179 );
and \U$44855 ( \45181 , \44460 , \44596 );
nor \U$44856 ( \45182 , \45181 , \44604 );
nand \U$44857 ( \45183 , \45180 , \45182 );
nor \U$44858 ( \45184 , \45177 , \45183 );
nand \U$44859 ( \45185 , \45170 , \45184 );
not \U$44860 ( \45186 , \45185 );
xor \U$44861 ( \45187 , \45146 , \45186 );
buf \U$44862 ( \45188 , \45187 );
_HMUX rb17c ( \45189_nRb17c , \45144 , \45188 , RIc0c97c8_1 );
buf \U$44863 ( \45190 , \45189_nRb17c );
xor \U$44864 ( \45191 , \1321 , \21563 );
buf \U$44865 ( \45192 , \45191 );
not \U$44866 ( \45193 , \35300 );
nand \U$44867 ( \45194 , \43825 , \45193 );
nand \U$44868 ( \45195 , \44644 , \44625 );
nand \U$44869 ( \45196 , \44626 , \44628 );
nor \U$44870 ( \45197 , \45195 , \45196 );
nand \U$44871 ( \45198 , \44629 , \44632 );
nand \U$44872 ( \45199 , \44633 , \44635 );
nor \U$44873 ( \45200 , \45198 , \45199 );
nand \U$44874 ( \45201 , \45197 , \45200 );
nand \U$44875 ( \45202 , \44648 , \44640 );
nand \U$44876 ( \45203 , \44641 , \44643 );
nor \U$44877 ( \45204 , \45202 , \45203 );
nand \U$44878 ( \45205 , \44650 , \44647 );
or \U$44879 ( \45206 , \45205 , \43490 );
and \U$44880 ( \45207 , \44647 , \44653 );
nor \U$44881 ( \45208 , \45207 , \44657 );
nand \U$44882 ( \45209 , \45206 , \45208 );
and \U$44883 ( \45210 , \45204 , \45209 );
and \U$44884 ( \45211 , \44640 , \44660 );
nor \U$44885 ( \45212 , \45211 , \44665 );
or \U$44886 ( \45213 , \45203 , \45212 );
and \U$44887 ( \45214 , \44643 , \44668 );
nor \U$44888 ( \45215 , \45214 , \44672 );
nand \U$44889 ( \45216 , \45213 , \45215 );
nor \U$44890 ( \45217 , \45210 , \45216 );
or \U$44891 ( \45218 , \45201 , \45217 );
and \U$44892 ( \45219 , \44625 , \44675 );
nor \U$44893 ( \45220 , \45219 , \44681 );
or \U$44894 ( \45221 , \45196 , \45220 );
and \U$44895 ( \45222 , \44628 , \44684 );
nor \U$44896 ( \45223 , \45222 , \44688 );
nand \U$44897 ( \45224 , \45221 , \45223 );
and \U$44898 ( \45225 , \45200 , \45224 );
and \U$44899 ( \45226 , \44632 , \44691 );
nor \U$44900 ( \45227 , \45226 , \44696 );
or \U$44901 ( \45228 , \45199 , \45227 );
and \U$44902 ( \45229 , \44635 , \44699 );
nor \U$44903 ( \45230 , \45229 , \44703 );
nand \U$44904 ( \45231 , \45228 , \45230 );
nor \U$44905 ( \45232 , \45225 , \45231 );
nand \U$44906 ( \45233 , \45218 , \45232 );
not \U$44907 ( \45234 , \45233 );
xor \U$44908 ( \45235 , \45194 , \45234 );
buf \U$44909 ( \45236 , \45235 );
_HMUX rb0d5 ( \45237_nRb0d5 , \45192 , \45236 , RIc0c97c8_1 );
buf \U$44910 ( \45238 , \45237_nRb0d5 );
xor \U$44911 ( \45239 , \1435 , \21561 );
buf \U$44912 ( \45240 , \45239 );
not \U$44913 ( \45241 , \35221 );
nand \U$44914 ( \45242 , \43821 , \45241 );
nand \U$44915 ( \45243 , \44739 , \44720 );
nand \U$44916 ( \45244 , \44721 , \44723 );
nor \U$44917 ( \45245 , \45243 , \45244 );
nand \U$44918 ( \45246 , \44724 , \44727 );
nand \U$44919 ( \45247 , \44728 , \44730 );
nor \U$44920 ( \45248 , \45246 , \45247 );
nand \U$44921 ( \45249 , \45245 , \45248 );
nand \U$44922 ( \45250 , \44743 , \44735 );
nand \U$44923 ( \45251 , \44736 , \44738 );
nor \U$44924 ( \45252 , \45250 , \45251 );
nand \U$44925 ( \45253 , \44745 , \44742 );
or \U$44926 ( \45254 , \45253 , \43486 );
and \U$44927 ( \45255 , \44742 , \44748 );
nor \U$44928 ( \45256 , \45255 , \44752 );
nand \U$44929 ( \45257 , \45254 , \45256 );
and \U$44930 ( \45258 , \45252 , \45257 );
and \U$44931 ( \45259 , \44735 , \44755 );
nor \U$44932 ( \45260 , \45259 , \44760 );
or \U$44933 ( \45261 , \45251 , \45260 );
and \U$44934 ( \45262 , \44738 , \44763 );
nor \U$44935 ( \45263 , \45262 , \44767 );
nand \U$44936 ( \45264 , \45261 , \45263 );
nor \U$44937 ( \45265 , \45258 , \45264 );
or \U$44938 ( \45266 , \45249 , \45265 );
and \U$44939 ( \45267 , \44720 , \44770 );
nor \U$44940 ( \45268 , \45267 , \44776 );
or \U$44941 ( \45269 , \45244 , \45268 );
and \U$44942 ( \45270 , \44723 , \44779 );
nor \U$44943 ( \45271 , \45270 , \44783 );
nand \U$44944 ( \45272 , \45269 , \45271 );
and \U$44945 ( \45273 , \45248 , \45272 );
and \U$44946 ( \45274 , \44727 , \44786 );
nor \U$44947 ( \45275 , \45274 , \44791 );
or \U$44948 ( \45276 , \45247 , \45275 );
and \U$44949 ( \45277 , \44730 , \44794 );
nor \U$44950 ( \45278 , \45277 , \44798 );
nand \U$44951 ( \45279 , \45276 , \45278 );
nor \U$44952 ( \45280 , \45273 , \45279 );
nand \U$44953 ( \45281 , \45266 , \45280 );
not \U$44954 ( \45282 , \45281 );
xor \U$44955 ( \45283 , \45242 , \45282 );
buf \U$44956 ( \45284 , \45283 );
_HMUX rb022 ( \45285_nRb022 , \45240 , \45284 , RIc0c97c8_1 );
buf \U$44957 ( \45286 , \45285_nRb022 );
xor \U$44958 ( \45287 , \1549 , \21559 );
buf \U$44959 ( \45288 , \45287 );
not \U$44960 ( \45289 , \35142 );
nand \U$44961 ( \45290 , \43819 , \45289 );
nand \U$44962 ( \45291 , \44834 , \44815 );
nand \U$44963 ( \45292 , \44816 , \44818 );
nor \U$44964 ( \45293 , \45291 , \45292 );
nand \U$44965 ( \45294 , \44819 , \44822 );
nand \U$44966 ( \45295 , \44823 , \44825 );
nor \U$44967 ( \45296 , \45294 , \45295 );
nand \U$44968 ( \45297 , \45293 , \45296 );
nand \U$44969 ( \45298 , \44838 , \44830 );
nand \U$44970 ( \45299 , \44831 , \44833 );
nor \U$44971 ( \45300 , \45298 , \45299 );
and \U$44972 ( \45301 , \44837 , \44841 );
nor \U$44973 ( \45302 , \45301 , \44845 );
not \U$44974 ( \45303 , \45302 );
and \U$44975 ( \45304 , \45300 , \45303 );
and \U$44976 ( \45305 , \44830 , \44848 );
nor \U$44977 ( \45306 , \45305 , \44853 );
or \U$44978 ( \45307 , \45299 , \45306 );
and \U$44979 ( \45308 , \44833 , \44856 );
nor \U$44980 ( \45309 , \45308 , \44860 );
nand \U$44981 ( \45310 , \45307 , \45309 );
nor \U$44982 ( \45311 , \45304 , \45310 );
or \U$44983 ( \45312 , \45297 , \45311 );
and \U$44984 ( \45313 , \44815 , \44863 );
nor \U$44985 ( \45314 , \45313 , \44869 );
or \U$44986 ( \45315 , \45292 , \45314 );
and \U$44987 ( \45316 , \44818 , \44872 );
nor \U$44988 ( \45317 , \45316 , \44876 );
nand \U$44989 ( \45318 , \45315 , \45317 );
and \U$44990 ( \45319 , \45296 , \45318 );
and \U$44991 ( \45320 , \44822 , \44879 );
nor \U$44992 ( \45321 , \45320 , \44884 );
or \U$44993 ( \45322 , \45295 , \45321 );
and \U$44994 ( \45323 , \44825 , \44887 );
nor \U$44995 ( \45324 , \45323 , \44891 );
nand \U$44996 ( \45325 , \45322 , \45324 );
nor \U$44997 ( \45326 , \45319 , \45325 );
nand \U$44998 ( \45327 , \45312 , \45326 );
not \U$44999 ( \45328 , \45327 );
xor \U$45000 ( \45329 , \45290 , \45328 );
buf \U$45001 ( \45330 , \45329 );
_HMUX raf66 ( \45331_nRaf66 , \45288 , \45330 , RIc0c97c8_1 );
buf \U$45002 ( \45332 , \45331_nRaf66 );
xor \U$45003 ( \45333 , \1664 , \21557 );
buf \U$45004 ( \45334 , \45333 );
not \U$45005 ( \45335 , \35054 );
nand \U$45006 ( \45336 , \43816 , \45335 );
nand \U$45007 ( \45337 , \44927 , \44908 );
nand \U$45008 ( \45338 , \44909 , \44911 );
nor \U$45009 ( \45339 , \45337 , \45338 );
nand \U$45010 ( \45340 , \44912 , \44915 );
nand \U$45011 ( \45341 , \44916 , \44918 );
nor \U$45012 ( \45342 , \45340 , \45341 );
nand \U$45013 ( \45343 , \45339 , \45342 );
nand \U$45014 ( \45344 , \44931 , \44923 );
nand \U$45015 ( \45345 , \44924 , \44926 );
nor \U$45016 ( \45346 , \45344 , \45345 );
and \U$45017 ( \45347 , \44930 , \44934 );
nor \U$45018 ( \45348 , \45347 , \44938 );
not \U$45019 ( \45349 , \45348 );
and \U$45020 ( \45350 , \45346 , \45349 );
and \U$45021 ( \45351 , \44923 , \44941 );
nor \U$45022 ( \45352 , \45351 , \44946 );
or \U$45023 ( \45353 , \45345 , \45352 );
and \U$45024 ( \45354 , \44926 , \44949 );
nor \U$45025 ( \45355 , \45354 , \44953 );
nand \U$45026 ( \45356 , \45353 , \45355 );
nor \U$45027 ( \45357 , \45350 , \45356 );
or \U$45028 ( \45358 , \45343 , \45357 );
and \U$45029 ( \45359 , \44908 , \44956 );
nor \U$45030 ( \45360 , \45359 , \44962 );
or \U$45031 ( \45361 , \45338 , \45360 );
and \U$45032 ( \45362 , \44911 , \44965 );
nor \U$45033 ( \45363 , \45362 , \44969 );
nand \U$45034 ( \45364 , \45361 , \45363 );
and \U$45035 ( \45365 , \45342 , \45364 );
and \U$45036 ( \45366 , \44915 , \44972 );
nor \U$45037 ( \45367 , \45366 , \44977 );
or \U$45038 ( \45368 , \45341 , \45367 );
and \U$45039 ( \45369 , \44918 , \44980 );
nor \U$45040 ( \45370 , \45369 , \44984 );
nand \U$45041 ( \45371 , \45368 , \45370 );
nor \U$45042 ( \45372 , \45365 , \45371 );
nand \U$45043 ( \45373 , \45358 , \45372 );
not \U$45044 ( \45374 , \45373 );
xor \U$45045 ( \45375 , \45336 , \45374 );
buf \U$45046 ( \45376 , \45375 );
_HMUX raea0 ( \45377_nRaea0 , \45334 , \45376 , RIc0c97c8_1 );
buf \U$45047 ( \45378 , \45377_nRaea0 );
xor \U$45048 ( \45379 , \1780 , \21555 );
buf \U$45049 ( \45380 , \45379 );
not \U$45050 ( \45381 , \34965 );
nand \U$45051 ( \45382 , \43814 , \45381 );
nor \U$45052 ( \45383 , \41861 , \29124 );
nor \U$45053 ( \45384 , \32641 , \34868 );
nand \U$45054 ( \45385 , \45383 , \45384 );
nor \U$45055 ( \45386 , \43174 , \39406 );
not \U$45056 ( \45387 , \43526 );
and \U$45057 ( \45388 , \45386 , \45387 );
or \U$45058 ( \45389 , \39406 , \43573 );
nand \U$45059 ( \45390 , \45389 , \43621 );
nor \U$45060 ( \45391 , \45388 , \45390 );
or \U$45061 ( \45392 , \45385 , \45391 );
or \U$45062 ( \45393 , \29124 , \43668 );
nand \U$45063 ( \45394 , \45393 , \43717 );
and \U$45064 ( \45395 , \45384 , \45394 );
or \U$45065 ( \45396 , \34868 , \43764 );
nand \U$45066 ( \45397 , \45396 , \43812 );
nor \U$45067 ( \45398 , \45395 , \45397 );
nand \U$45068 ( \45399 , \45392 , \45398 );
not \U$45069 ( \45400 , \45399 );
xor \U$45070 ( \45401 , \45382 , \45400 );
buf \U$45071 ( \45402 , \45401 );
_HMUX radd0 ( \45403_nRadd0 , \45380 , \45402 , RIc0c97c8_1 );
buf \U$45072 ( \45404 , \45403_nRadd0 );
xor \U$45073 ( \45405 , \1903 , \21553 );
buf \U$45074 ( \45406 , \45405 );
not \U$45075 ( \45407 , \34864 );
nand \U$45076 ( \45408 , \43808 , \45407 );
nor \U$45077 ( \45409 , \43964 , \43886 );
nor \U$45078 ( \45410 , \43901 , \43917 );
nand \U$45079 ( \45411 , \45409 , \45410 );
nor \U$45080 ( \45412 , \43980 , \43949 );
not \U$45081 ( \45413 , \44014 );
and \U$45082 ( \45414 , \45412 , \45413 );
or \U$45083 ( \45415 , \43949 , \44045 );
nand \U$45084 ( \45416 , \45415 , \44077 );
nor \U$45085 ( \45417 , \45414 , \45416 );
or \U$45086 ( \45418 , \45411 , \45417 );
or \U$45087 ( \45419 , \43886 , \44108 );
nand \U$45088 ( \45420 , \45419 , \44141 );
and \U$45089 ( \45421 , \45410 , \45420 );
or \U$45090 ( \45422 , \43917 , \44172 );
nand \U$45091 ( \45423 , \45422 , \44204 );
nor \U$45092 ( \45424 , \45421 , \45423 );
nand \U$45093 ( \45425 , \45418 , \45424 );
not \U$45094 ( \45426 , \45425 );
xor \U$45095 ( \45427 , \45408 , \45426 );
buf \U$45096 ( \45428 , \45427 );
_HMUX racf6 ( \45429_nRacf6 , \45406 , \45428 , RIc0c97c8_1 );
buf \U$45097 ( \45430 , \45429_nRacf6 );
xor \U$45098 ( \45431 , \2024 , \21551 );
buf \U$45099 ( \45432 , \45431 );
not \U$45100 ( \45433 , \34765 );
nand \U$45101 ( \45434 , \43806 , \45433 );
nor \U$45102 ( \45435 , \44292 , \44254 );
nor \U$45103 ( \45436 , \44261 , \44269 );
nand \U$45104 ( \45437 , \45435 , \45436 );
nor \U$45105 ( \45438 , \44300 , \44285 );
not \U$45106 ( \45439 , \44314 );
and \U$45107 ( \45440 , \45438 , \45439 );
or \U$45108 ( \45441 , \44285 , \44329 );
nand \U$45109 ( \45442 , \45441 , \44345 );
nor \U$45110 ( \45443 , \45440 , \45442 );
or \U$45111 ( \45444 , \45437 , \45443 );
or \U$45112 ( \45445 , \44254 , \44360 );
nand \U$45113 ( \45446 , \45445 , \44377 );
and \U$45114 ( \45447 , \45436 , \45446 );
or \U$45115 ( \45448 , \44269 , \44392 );
nand \U$45116 ( \45449 , \45448 , \44408 );
nor \U$45117 ( \45450 , \45447 , \45449 );
nand \U$45118 ( \45451 , \45444 , \45450 );
not \U$45119 ( \45452 , \45451 );
xor \U$45120 ( \45453 , \45434 , \45452 );
buf \U$45121 ( \45454 , \45453 );
_HMUX rac12 ( \45455_nRac12 , \45432 , \45454 , RIc0c97c8_1 );
buf \U$45122 ( \45456 , \45455_nRac12 );
xor \U$45123 ( \45457 , \2157 , \21549 );
buf \U$45124 ( \45458 , \45457 );
not \U$45125 ( \45459 , \34660 );
nand \U$45126 ( \45460 , \43803 , \45459 );
nor \U$45127 ( \45461 , \44480 , \44442 );
nor \U$45128 ( \45462 , \44449 , \44457 );
nand \U$45129 ( \45463 , \45461 , \45462 );
nor \U$45130 ( \45464 , \44488 , \44473 );
not \U$45131 ( \45465 , \44503 );
and \U$45132 ( \45466 , \45464 , \45465 );
or \U$45133 ( \45467 , \44473 , \44518 );
nand \U$45134 ( \45468 , \45467 , \44534 );
nor \U$45135 ( \45469 , \45466 , \45468 );
or \U$45136 ( \45470 , \45463 , \45469 );
or \U$45137 ( \45471 , \44442 , \44549 );
nand \U$45138 ( \45472 , \45471 , \44566 );
and \U$45139 ( \45473 , \45462 , \45472 );
or \U$45140 ( \45474 , \44457 , \44581 );
nand \U$45141 ( \45475 , \45474 , \44597 );
nor \U$45142 ( \45476 , \45473 , \45475 );
nand \U$45143 ( \45477 , \45470 , \45476 );
not \U$45144 ( \45478 , \45477 );
xor \U$45145 ( \45479 , \45460 , \45478 );
buf \U$45146 ( \45480 , \45479 );
_HMUX rab27 ( \45481_nRab27 , \45458 , \45480 , RIc0c97c8_1 );
buf \U$45147 ( \45482 , \45481_nRab27 );
xor \U$45148 ( \45483 , \2294 , \21547 );
buf \U$45149 ( \45484 , \45483 );
not \U$45150 ( \45485 , \34550 );
nand \U$45151 ( \45486 , \43801 , \45485 );
nor \U$45152 ( \45487 , \44645 , \44627 );
nor \U$45153 ( \45488 , \44630 , \44634 );
nand \U$45154 ( \45489 , \45487 , \45488 );
nor \U$45155 ( \45490 , \44649 , \44642 );
not \U$45156 ( \45491 , \44654 );
and \U$45157 ( \45492 , \45490 , \45491 );
or \U$45158 ( \45493 , \44642 , \44661 );
nand \U$45159 ( \45494 , \45493 , \44669 );
nor \U$45160 ( \45495 , \45492 , \45494 );
or \U$45161 ( \45496 , \45489 , \45495 );
or \U$45162 ( \45497 , \44627 , \44676 );
nand \U$45163 ( \45498 , \45497 , \44685 );
and \U$45164 ( \45499 , \45488 , \45498 );
or \U$45165 ( \45500 , \44634 , \44692 );
nand \U$45166 ( \45501 , \45500 , \44700 );
nor \U$45167 ( \45502 , \45499 , \45501 );
nand \U$45168 ( \45503 , \45496 , \45502 );
not \U$45169 ( \45504 , \45503 );
xor \U$45170 ( \45505 , \45486 , \45504 );
buf \U$45171 ( \45506 , \45505 );
_HMUX raa31 ( \45507_nRaa31 , \45484 , \45506 , RIc0c97c8_1 );
buf \U$45172 ( \45508 , \45507_nRaa31 );
xor \U$45173 ( \45509 , \2574 , \21545 );
buf \U$45174 ( \45510 , \45509 );
not \U$45175 ( \45511 , \34431 );
nand \U$45176 ( \45512 , \43797 , \45511 );
nor \U$45177 ( \45513 , \44740 , \44722 );
nor \U$45178 ( \45514 , \44725 , \44729 );
nand \U$45179 ( \45515 , \45513 , \45514 );
nor \U$45180 ( \45516 , \44744 , \44737 );
not \U$45181 ( \45517 , \44749 );
and \U$45182 ( \45518 , \45516 , \45517 );
or \U$45183 ( \45519 , \44737 , \44756 );
nand \U$45184 ( \45520 , \45519 , \44764 );
nor \U$45185 ( \45521 , \45518 , \45520 );
or \U$45186 ( \45522 , \45515 , \45521 );
or \U$45187 ( \45523 , \44722 , \44771 );
nand \U$45188 ( \45524 , \45523 , \44780 );
and \U$45189 ( \45525 , \45514 , \45524 );
or \U$45190 ( \45526 , \44729 , \44787 );
nand \U$45191 ( \45527 , \45526 , \44795 );
nor \U$45192 ( \45528 , \45525 , \45527 );
nand \U$45193 ( \45529 , \45522 , \45528 );
not \U$45194 ( \45530 , \45529 );
xor \U$45195 ( \45531 , \45512 , \45530 );
buf \U$45196 ( \45532 , \45531 );
_HMUX ra92e ( \45533_nRa92e , \45510 , \45532 , RIc0c97c8_1 );
buf \U$45197 ( \45534 , \45533_nRa92e );
xor \U$45198 ( \45535 , \2747 , \21543 );
buf \U$45199 ( \45536 , \45535 );
not \U$45200 ( \45537 , \34310 );
nand \U$45201 ( \45538 , \43795 , \45537 );
nor \U$45202 ( \45539 , \44835 , \44817 );
nor \U$45203 ( \45540 , \44820 , \44824 );
nand \U$45204 ( \45541 , \45539 , \45540 );
nor \U$45205 ( \45542 , \44839 , \44832 );
and \U$45206 ( \45543 , \45542 , \44841 );
or \U$45207 ( \45544 , \44832 , \44849 );
nand \U$45208 ( \45545 , \45544 , \44857 );
nor \U$45209 ( \45546 , \45543 , \45545 );
or \U$45210 ( \45547 , \45541 , \45546 );
or \U$45211 ( \45548 , \44817 , \44864 );
nand \U$45212 ( \45549 , \45548 , \44873 );
and \U$45213 ( \45550 , \45540 , \45549 );
or \U$45214 ( \45551 , \44824 , \44880 );
nand \U$45215 ( \45552 , \45551 , \44888 );
nor \U$45216 ( \45553 , \45550 , \45552 );
nand \U$45217 ( \45554 , \45547 , \45553 );
not \U$45218 ( \45555 , \45554 );
xor \U$45219 ( \45556 , \45538 , \45555 );
buf \U$45220 ( \45557 , \45556 );
_HMUX ra820 ( \45558_nRa820 , \45536 , \45557 , RIc0c97c8_1 );
buf \U$45221 ( \45559 , \45558_nRa820 );
xor \U$45222 ( \45560 , \2913 , \21541 );
buf \U$45223 ( \45561 , \45560 );
not \U$45224 ( \45562 , \34181 );
nand \U$45225 ( \45563 , \43792 , \45562 );
nor \U$45226 ( \45564 , \44928 , \44910 );
nor \U$45227 ( \45565 , \44913 , \44917 );
nand \U$45228 ( \45566 , \45564 , \45565 );
nor \U$45229 ( \45567 , \44932 , \44925 );
and \U$45230 ( \45568 , \45567 , \44934 );
or \U$45231 ( \45569 , \44925 , \44942 );
nand \U$45232 ( \45570 , \45569 , \44950 );
nor \U$45233 ( \45571 , \45568 , \45570 );
or \U$45234 ( \45572 , \45566 , \45571 );
or \U$45235 ( \45573 , \44910 , \44957 );
nand \U$45236 ( \45574 , \45573 , \44966 );
and \U$45237 ( \45575 , \45565 , \45574 );
or \U$45238 ( \45576 , \44917 , \44973 );
nand \U$45239 ( \45577 , \45576 , \44981 );
nor \U$45240 ( \45578 , \45575 , \45577 );
nand \U$45241 ( \45579 , \45572 , \45578 );
not \U$45242 ( \45580 , \45579 );
xor \U$45243 ( \45581 , \45563 , \45580 );
buf \U$45244 ( \45582 , \45581 );
_HMUX ra706 ( \45583_nRa706 , \45561 , \45582 , RIc0c97c8_1 );
buf \U$45245 ( \45584 , \45583_nRa706 );
xor \U$45246 ( \45585 , \3080 , \21539 );
buf \U$45247 ( \45586 , \45585 );
not \U$45248 ( \45587 , \34052 );
nand \U$45249 ( \45588 , \43790 , \45587 );
nor \U$45250 ( \45589 , \45009 , \45001 );
nor \U$45251 ( \45590 , \45002 , \45004 );
nand \U$45252 ( \45591 , \45589 , \45590 );
nor \U$45253 ( \45592 , \45011 , \45008 );
and \U$45254 ( \45593 , \45592 , \43502 );
or \U$45255 ( \45594 , \45008 , \45015 );
nand \U$45256 ( \45595 , \45594 , \45019 );
nor \U$45257 ( \45596 , \45593 , \45595 );
or \U$45258 ( \45597 , \45591 , \45596 );
or \U$45259 ( \45598 , \45001 , \45022 );
nand \U$45260 ( \45599 , \45598 , \45027 );
and \U$45261 ( \45600 , \45590 , \45599 );
or \U$45262 ( \45601 , \45004 , \45030 );
nand \U$45263 ( \45602 , \45601 , \45034 );
nor \U$45264 ( \45603 , \45600 , \45602 );
nand \U$45265 ( \45604 , \45597 , \45603 );
not \U$45266 ( \45605 , \45604 );
xor \U$45267 ( \45606 , \45588 , \45605 );
buf \U$45268 ( \45607 , \45606 );
_HMUX ra5e5 ( \45608_nRa5e5 , \45586 , \45607 , RIc0c97c8_1 );
buf \U$45269 ( \45609 , \45608_nRa5e5 );
xor \U$45270 ( \45610 , \3253 , \21537 );
buf \U$45271 ( \45611 , \45610 );
not \U$45272 ( \45612 , \33912 );
nand \U$45273 ( \45613 , \43785 , \45612 );
nor \U$45274 ( \45614 , \45058 , \45050 );
nor \U$45275 ( \45615 , \45051 , \45053 );
nand \U$45276 ( \45616 , \45614 , \45615 );
nor \U$45277 ( \45617 , \45060 , \45057 );
and \U$45278 ( \45618 , \45617 , \43998 );
or \U$45279 ( \45619 , \45057 , \45064 );
nand \U$45280 ( \45620 , \45619 , \45068 );
nor \U$45281 ( \45621 , \45618 , \45620 );
or \U$45282 ( \45622 , \45616 , \45621 );
or \U$45283 ( \45623 , \45050 , \45071 );
nand \U$45284 ( \45624 , \45623 , \45076 );
and \U$45285 ( \45625 , \45615 , \45624 );
or \U$45286 ( \45626 , \45053 , \45079 );
nand \U$45287 ( \45627 , \45626 , \45083 );
nor \U$45288 ( \45628 , \45625 , \45627 );
nand \U$45289 ( \45629 , \45622 , \45628 );
not \U$45290 ( \45630 , \45629 );
xor \U$45291 ( \45631 , \45613 , \45630 );
buf \U$45292 ( \45632 , \45631 );
_HMUX ra4bb ( \45633_nRa4bb , \45611 , \45632 , RIc0c97c8_1 );
buf \U$45293 ( \45634 , \45633_nRa4bb );
xor \U$45294 ( \45635 , \3428 , \21535 );
buf \U$45295 ( \45636 , \45635 );
not \U$45296 ( \45637 , \33770 );
nand \U$45297 ( \45638 , \43783 , \45637 );
nor \U$45298 ( \45639 , \45107 , \45099 );
nor \U$45299 ( \45640 , \45100 , \45102 );
nand \U$45300 ( \45641 , \45639 , \45640 );
nor \U$45301 ( \45642 , \45109 , \45106 );
and \U$45302 ( \45643 , \45642 , \44306 );
or \U$45303 ( \45644 , \45106 , \45112 );
nand \U$45304 ( \45645 , \45644 , \45116 );
nor \U$45305 ( \45646 , \45643 , \45645 );
or \U$45306 ( \45647 , \45641 , \45646 );
or \U$45307 ( \45648 , \45099 , \45119 );
nand \U$45308 ( \45649 , \45648 , \45124 );
and \U$45309 ( \45650 , \45640 , \45649 );
or \U$45310 ( \45651 , \45102 , \45127 );
nand \U$45311 ( \45652 , \45651 , \45131 );
nor \U$45312 ( \45653 , \45650 , \45652 );
nand \U$45313 ( \45654 , \45647 , \45653 );
not \U$45314 ( \45655 , \45654 );
xor \U$45315 ( \45656 , \45638 , \45655 );
buf \U$45316 ( \45657 , \45656 );
_HMUX ra384 ( \45658_nRa384 , \45636 , \45657 , RIc0c97c8_1 );
buf \U$45317 ( \45659 , \45658_nRa384 );
xor \U$45318 ( \45660 , \3599 , \21533 );
buf \U$45319 ( \45661 , \45660 );
not \U$45320 ( \45662 , \33620 );
nand \U$45321 ( \45663 , \43780 , \45662 );
nor \U$45322 ( \45664 , \45155 , \45147 );
nor \U$45323 ( \45665 , \45148 , \45150 );
nand \U$45324 ( \45666 , \45664 , \45665 );
nor \U$45325 ( \45667 , \45157 , \45154 );
and \U$45326 ( \45668 , \45667 , \44495 );
or \U$45327 ( \45669 , \45154 , \45160 );
nand \U$45328 ( \45670 , \45669 , \45164 );
nor \U$45329 ( \45671 , \45668 , \45670 );
or \U$45330 ( \45672 , \45666 , \45671 );
or \U$45331 ( \45673 , \45147 , \45167 );
nand \U$45332 ( \45674 , \45673 , \45172 );
and \U$45333 ( \45675 , \45665 , \45674 );
or \U$45334 ( \45676 , \45150 , \45175 );
nand \U$45335 ( \45677 , \45676 , \45179 );
nor \U$45336 ( \45678 , \45675 , \45677 );
nand \U$45337 ( \45679 , \45672 , \45678 );
not \U$45338 ( \45680 , \45679 );
xor \U$45339 ( \45681 , \45663 , \45680 );
buf \U$45340 ( \45682 , \45681 );
_HMUX ra241 ( \45683_nRa241 , \45661 , \45682 , RIc0c97c8_1 );
buf \U$45341 ( \45684 , \45683_nRa241 );
xor \U$45342 ( \45685 , \3780 , \21531 );
buf \U$45343 ( \45686 , \45685 );
not \U$45344 ( \45687 , \33467 );
nand \U$45345 ( \45688 , \43778 , \45687 );
nor \U$45346 ( \45689 , \45203 , \45195 );
nor \U$45347 ( \45690 , \45196 , \45198 );
nand \U$45348 ( \45691 , \45689 , \45690 );
nor \U$45349 ( \45692 , \45205 , \45202 );
and \U$45350 ( \45693 , \45692 , \43489 );
or \U$45351 ( \45694 , \45202 , \45208 );
nand \U$45352 ( \45695 , \45694 , \45212 );
nor \U$45353 ( \45696 , \45693 , \45695 );
or \U$45354 ( \45697 , \45691 , \45696 );
or \U$45355 ( \45698 , \45195 , \45215 );
nand \U$45356 ( \45699 , \45698 , \45220 );
and \U$45357 ( \45700 , \45690 , \45699 );
or \U$45358 ( \45701 , \45198 , \45223 );
nand \U$45359 ( \45702 , \45701 , \45227 );
nor \U$45360 ( \45703 , \45700 , \45702 );
nand \U$45361 ( \45704 , \45697 , \45703 );
not \U$45362 ( \45705 , \45704 );
xor \U$45363 ( \45706 , \45688 , \45705 );
buf \U$45364 ( \45707 , \45706 );
_HMUX ra0f3 ( \45708_nRa0f3 , \45686 , \45707 , RIc0c97c8_1 );
buf \U$45365 ( \45709 , \45708_nRa0f3 );
xor \U$45366 ( \45710 , \3957 , \21529 );
buf \U$45367 ( \45711 , \45710 );
not \U$45368 ( \45712 , \33308 );
nand \U$45369 ( \45713 , \43774 , \45712 );
nor \U$45370 ( \45714 , \45251 , \45243 );
nor \U$45371 ( \45715 , \45244 , \45246 );
nand \U$45372 ( \45716 , \45714 , \45715 );
nor \U$45373 ( \45717 , \45253 , \45250 );
and \U$45374 ( \45718 , \45717 , \44492 );
or \U$45375 ( \45719 , \45250 , \45256 );
nand \U$45376 ( \45720 , \45719 , \45260 );
nor \U$45377 ( \45721 , \45718 , \45720 );
or \U$45378 ( \45722 , \45716 , \45721 );
or \U$45379 ( \45723 , \45243 , \45263 );
nand \U$45380 ( \45724 , \45723 , \45268 );
and \U$45381 ( \45725 , \45715 , \45724 );
or \U$45382 ( \45726 , \45246 , \45271 );
nand \U$45383 ( \45727 , \45726 , \45275 );
nor \U$45384 ( \45728 , \45725 , \45727 );
nand \U$45385 ( \45729 , \45722 , \45728 );
not \U$45386 ( \45730 , \45729 );
xor \U$45387 ( \45731 , \45713 , \45730 );
buf \U$45388 ( \45732 , \45731 );
_HMUX r9f9c ( \45733_nR9f9c , \45711 , \45732 , RIc0c97c8_1 );
buf \U$45389 ( \45734 , \45733_nR9f9c );
xor \U$45390 ( \45735 , \4154 , \21527 );
buf \U$45391 ( \45736 , \45735 );
not \U$45392 ( \45737 , \33149 );
nand \U$45393 ( \45738 , \43772 , \45737 );
nor \U$45394 ( \45739 , \45299 , \45291 );
nor \U$45395 ( \45740 , \45292 , \45294 );
nand \U$45396 ( \45741 , \45739 , \45740 );
or \U$45397 ( \45742 , \45298 , \45302 );
nand \U$45398 ( \45743 , \45742 , \45306 );
not \U$45399 ( \45744 , \45743 );
or \U$45400 ( \45745 , \45741 , \45744 );
or \U$45401 ( \45746 , \45291 , \45309 );
nand \U$45402 ( \45747 , \45746 , \45314 );
and \U$45403 ( \45748 , \45740 , \45747 );
or \U$45404 ( \45749 , \45294 , \45317 );
nand \U$45405 ( \45750 , \45749 , \45321 );
nor \U$45406 ( \45751 , \45748 , \45750 );
nand \U$45407 ( \45752 , \45745 , \45751 );
not \U$45408 ( \45753 , \45752 );
xor \U$45409 ( \45754 , \45738 , \45753 );
buf \U$45410 ( \45755 , \45754 );
_HMUX r9e40 ( \45756_nR9e40 , \45736 , \45755 , RIc0c97c8_1 );
buf \U$45411 ( \45757 , \45756_nR9e40 );
xor \U$45412 ( \45758 , \4350 , \21525 );
buf \U$45413 ( \45759 , \45758 );
not \U$45414 ( \45760 , \32984 );
nand \U$45415 ( \45761 , \43769 , \45760 );
nor \U$45416 ( \45762 , \45345 , \45337 );
nor \U$45417 ( \45763 , \45338 , \45340 );
nand \U$45418 ( \45764 , \45762 , \45763 );
or \U$45419 ( \45765 , \45344 , \45348 );
nand \U$45420 ( \45766 , \45765 , \45352 );
not \U$45421 ( \45767 , \45766 );
or \U$45422 ( \45768 , \45764 , \45767 );
or \U$45423 ( \45769 , \45337 , \45355 );
nand \U$45424 ( \45770 , \45769 , \45360 );
and \U$45425 ( \45771 , \45763 , \45770 );
or \U$45426 ( \45772 , \45340 , \45363 );
nand \U$45427 ( \45773 , \45772 , \45367 );
nor \U$45428 ( \45774 , \45771 , \45773 );
nand \U$45429 ( \45775 , \45768 , \45774 );
not \U$45430 ( \45776 , \45775 );
xor \U$45431 ( \45777 , \45761 , \45776 );
buf \U$45432 ( \45778 , \45777 );
_HMUX r9cdd ( \45779_nR9cdd , \45759 , \45778 , RIc0c97c8_1 );
buf \U$45433 ( \45780 , \45779_nR9cdd );
xor \U$45434 ( \45781 , \4552 , \21523 );
buf \U$45435 ( \45782 , \45781 );
not \U$45436 ( \45783 , \32817 );
nand \U$45437 ( \45784 , \43767 , \45783 );
nand \U$45438 ( \45785 , \41862 , \32642 );
not \U$45439 ( \45786 , \43574 );
or \U$45440 ( \45787 , \45785 , \45786 );
and \U$45441 ( \45788 , \32642 , \43669 );
nor \U$45442 ( \45789 , \45788 , \43765 );
nand \U$45443 ( \45790 , \45787 , \45789 );
not \U$45444 ( \45791 , \45790 );
xor \U$45445 ( \45792 , \45784 , \45791 );
buf \U$45446 ( \45793 , \45792 );
_HMUX r9b72 ( \45794_nR9b72 , \45782 , \45793 , RIc0c97c8_1 );
buf \U$45447 ( \45795 , \45794_nR9b72 );
xor \U$45448 ( \45796 , \4759 , \21521 );
buf \U$45449 ( \45797 , \45796 );
not \U$45450 ( \45798 , \32637 );
nand \U$45451 ( \45799 , \43760 , \45798 );
nand \U$45452 ( \45800 , \43965 , \43902 );
not \U$45453 ( \45801 , \44046 );
or \U$45454 ( \45802 , \45800 , \45801 );
and \U$45455 ( \45803 , \43902 , \44109 );
nor \U$45456 ( \45804 , \45803 , \44173 );
nand \U$45457 ( \45805 , \45802 , \45804 );
not \U$45458 ( \45806 , \45805 );
xor \U$45459 ( \45807 , \45799 , \45806 );
buf \U$45460 ( \45808 , \45807 );
_HMUX r99fc ( \45809_nR99fc , \45797 , \45808 , RIc0c97c8_1 );
buf \U$45461 ( \45810 , \45809_nR99fc );
xor \U$45462 ( \45811 , \4969 , \21519 );
buf \U$45463 ( \45812 , \45811 );
not \U$45464 ( \45813 , \32457 );
nand \U$45465 ( \45814 , \43758 , \45813 );
nand \U$45466 ( \45815 , \44293 , \44262 );
not \U$45467 ( \45816 , \44330 );
or \U$45468 ( \45817 , \45815 , \45816 );
and \U$45469 ( \45818 , \44262 , \44361 );
nor \U$45470 ( \45819 , \45818 , \44393 );
nand \U$45471 ( \45820 , \45817 , \45819 );
not \U$45472 ( \45821 , \45820 );
xor \U$45473 ( \45822 , \45814 , \45821 );
buf \U$45474 ( \45823 , \45822 );
_HMUX r9879 ( \45824_nR9879 , \45812 , \45823 , RIc0c97c8_1 );
buf \U$45475 ( \45825 , \45824_nR9879 );
xor \U$45476 ( \45826 , \5398 , \21517 );
buf \U$45477 ( \45827 , \45826 );
not \U$45478 ( \45828 , \32269 );
nand \U$45479 ( \45829 , \43755 , \45828 );
nand \U$45480 ( \45830 , \44481 , \44450 );
not \U$45481 ( \45831 , \44519 );
or \U$45482 ( \45832 , \45830 , \45831 );
and \U$45483 ( \45833 , \44450 , \44550 );
nor \U$45484 ( \45834 , \45833 , \44582 );
nand \U$45485 ( \45835 , \45832 , \45834 );
not \U$45486 ( \45836 , \45835 );
xor \U$45487 ( \45837 , \45829 , \45836 );
buf \U$45488 ( \45838 , \45837 );
_HMUX r96ea ( \45839_nR96ea , \45827 , \45838 , RIc0c97c8_1 );
buf \U$45489 ( \45840 , \45839_nR96ea );
xor \U$45490 ( \45841 , \5641 , \21515 );
buf \U$45491 ( \45842 , \45841 );
not \U$45492 ( \45843 , \32080 );
nand \U$45493 ( \45844 , \43753 , \45843 );
nand \U$45494 ( \45845 , \44646 , \44631 );
not \U$45495 ( \45846 , \44662 );
or \U$45496 ( \45847 , \45845 , \45846 );
and \U$45497 ( \45848 , \44631 , \44677 );
nor \U$45498 ( \45849 , \45848 , \44693 );
nand \U$45499 ( \45850 , \45847 , \45849 );
not \U$45500 ( \45851 , \45850 );
xor \U$45501 ( \45852 , \45844 , \45851 );
buf \U$45502 ( \45853 , \45852 );
_HMUX r9552 ( \45854_nR9552 , \45842 , \45853 , RIc0c97c8_1 );
buf \U$45503 ( \45855 , \45854_nR9552 );
xor \U$45504 ( \45856 , \5873 , \21513 );
buf \U$45505 ( \45857 , \45856 );
not \U$45506 ( \45858 , \31881 );
nand \U$45507 ( \45859 , \43749 , \45858 );
nand \U$45508 ( \45860 , \44741 , \44726 );
not \U$45509 ( \45861 , \44757 );
or \U$45510 ( \45862 , \45860 , \45861 );
and \U$45511 ( \45863 , \44726 , \44772 );
nor \U$45512 ( \45864 , \45863 , \44788 );
nand \U$45513 ( \45865 , \45862 , \45864 );
not \U$45514 ( \45866 , \45865 );
xor \U$45515 ( \45867 , \45859 , \45866 );
buf \U$45516 ( \45868 , \45867 );
_HMUX r93b0 ( \45869_nR93b0 , \45857 , \45868 , RIc0c97c8_1 );
buf \U$45517 ( \45870 , \45869_nR93b0 );
xor \U$45518 ( \45871 , \6121 , \21511 );
buf \U$45519 ( \45872 , \45871 );
not \U$45520 ( \45873 , \31682 );
nand \U$45521 ( \45874 , \43747 , \45873 );
nand \U$45522 ( \45875 , \44836 , \44821 );
not \U$45523 ( \45876 , \44850 );
or \U$45524 ( \45877 , \45875 , \45876 );
and \U$45525 ( \45878 , \44821 , \44865 );
nor \U$45526 ( \45879 , \45878 , \44881 );
nand \U$45527 ( \45880 , \45877 , \45879 );
not \U$45528 ( \45881 , \45880 );
xor \U$45529 ( \45882 , \45874 , \45881 );
buf \U$45530 ( \45883 , \45882 );
_HMUX r9204 ( \45884_nR9204 , \45872 , \45883 , RIc0c97c8_1 );
buf \U$45531 ( \45885 , \45884_nR9204 );
xor \U$45532 ( \45886 , \6374 , \21509 );
buf \U$45533 ( \45887 , \45886 );
not \U$45534 ( \45888 , \31474 );
nand \U$45535 ( \45889 , \43744 , \45888 );
nand \U$45536 ( \45890 , \44929 , \44914 );
not \U$45537 ( \45891 , \44943 );
or \U$45538 ( \45892 , \45890 , \45891 );
and \U$45539 ( \45893 , \44914 , \44958 );
nor \U$45540 ( \45894 , \45893 , \44974 );
nand \U$45541 ( \45895 , \45892 , \45894 );
not \U$45542 ( \45896 , \45895 );
xor \U$45543 ( \45897 , \45889 , \45896 );
buf \U$45544 ( \45898 , \45897 );
_HMUX r904e ( \45899_nR904e , \45887 , \45898 , RIc0c97c8_1 );
buf \U$45545 ( \45900 , \45899_nR904e );
xor \U$45546 ( \45901 , \6630 , \21507 );
buf \U$45547 ( \45902 , \45901 );
not \U$45548 ( \45903 , \31263 );
nand \U$45549 ( \45904 , \43742 , \45903 );
nand \U$45550 ( \45905 , \45010 , \45003 );
not \U$45551 ( \45906 , \45016 );
or \U$45552 ( \45907 , \45905 , \45906 );
and \U$45553 ( \45908 , \45003 , \45023 );
nor \U$45554 ( \45909 , \45908 , \45031 );
nand \U$45555 ( \45910 , \45907 , \45909 );
not \U$45556 ( \45911 , \45910 );
xor \U$45557 ( \45912 , \45904 , \45911 );
buf \U$45558 ( \45913 , \45912 );
_HMUX r8e8c ( \45914_nR8e8c , \45902 , \45913 , RIc0c97c8_1 );
buf \U$45559 ( \45915 , \45914_nR8e8c );
xor \U$45560 ( \45916 , \6887 , \21505 );
buf \U$45561 ( \45917 , \45916 );
not \U$45562 ( \45918 , \31042 );
nand \U$45563 ( \45919 , \43737 , \45918 );
nand \U$45564 ( \45920 , \45059 , \45052 );
not \U$45565 ( \45921 , \45065 );
or \U$45566 ( \45922 , \45920 , \45921 );
and \U$45567 ( \45923 , \45052 , \45072 );
nor \U$45568 ( \45924 , \45923 , \45080 );
nand \U$45569 ( \45925 , \45922 , \45924 );
not \U$45570 ( \45926 , \45925 );
xor \U$45571 ( \45927 , \45919 , \45926 );
buf \U$45572 ( \45928 , \45927 );
_HMUX r8cbe ( \45929_nR8cbe , \45917 , \45928 , RIc0c97c8_1 );
buf \U$45573 ( \45930 , \45929_nR8cbe );
xor \U$45574 ( \45931 , \7150 , \21503 );
buf \U$45575 ( \45932 , \45931 );
not \U$45576 ( \45933 , \30820 );
nand \U$45577 ( \45934 , \43735 , \45933 );
nand \U$45578 ( \45935 , \45108 , \45101 );
not \U$45579 ( \45936 , \45113 );
or \U$45580 ( \45937 , \45935 , \45936 );
and \U$45581 ( \45938 , \45101 , \45120 );
nor \U$45582 ( \45939 , \45938 , \45128 );
nand \U$45583 ( \45940 , \45937 , \45939 );
not \U$45584 ( \45941 , \45940 );
xor \U$45585 ( \45942 , \45934 , \45941 );
buf \U$45586 ( \45943 , \45942 );
_HMUX r8ae6 ( \45944_nR8ae6 , \45932 , \45943 , RIc0c97c8_1 );
buf \U$45587 ( \45945 , \45944_nR8ae6 );
xor \U$45588 ( \45946 , \7415 , \21501 );
buf \U$45589 ( \45947 , \45946 );
not \U$45590 ( \45948 , \30590 );
nand \U$45591 ( \45949 , \43732 , \45948 );
nand \U$45592 ( \45950 , \45156 , \45149 );
not \U$45593 ( \45951 , \45161 );
or \U$45594 ( \45952 , \45950 , \45951 );
and \U$45595 ( \45953 , \45149 , \45168 );
nor \U$45596 ( \45954 , \45953 , \45176 );
nand \U$45597 ( \45955 , \45952 , \45954 );
not \U$45598 ( \45956 , \45955 );
xor \U$45599 ( \45957 , \45949 , \45956 );
buf \U$45600 ( \45958 , \45957 );
_HMUX r8903 ( \45959_nR8903 , \45947 , \45958 , RIc0c97c8_1 );
buf \U$45601 ( \45960 , \45959_nR8903 );
xor \U$45602 ( \45961 , \7676 , \21499 );
buf \U$45603 ( \45962 , \45961 );
not \U$45604 ( \45963 , \30359 );
nand \U$45605 ( \45964 , \43730 , \45963 );
nand \U$45606 ( \45965 , \45204 , \45197 );
not \U$45607 ( \45966 , \45209 );
or \U$45608 ( \45967 , \45965 , \45966 );
and \U$45609 ( \45968 , \45197 , \45216 );
nor \U$45610 ( \45969 , \45968 , \45224 );
nand \U$45611 ( \45970 , \45967 , \45969 );
not \U$45612 ( \45971 , \45970 );
xor \U$45613 ( \45972 , \45964 , \45971 );
buf \U$45614 ( \45973 , \45972 );
_HMUX r8717 ( \45974_nR8717 , \45962 , \45973 , RIc0c97c8_1 );
buf \U$45615 ( \45975 , \45974_nR8717 );
xor \U$45616 ( \45976 , \7942 , \21497 );
buf \U$45617 ( \45977 , \45976 );
not \U$45618 ( \45978 , \30118 );
nand \U$45619 ( \45979 , \43726 , \45978 );
nand \U$45620 ( \45980 , \45252 , \45245 );
not \U$45621 ( \45981 , \45257 );
or \U$45622 ( \45982 , \45980 , \45981 );
and \U$45623 ( \45983 , \45245 , \45264 );
nor \U$45624 ( \45984 , \45983 , \45272 );
nand \U$45625 ( \45985 , \45982 , \45984 );
not \U$45626 ( \45986 , \45985 );
xor \U$45627 ( \45987 , \45979 , \45986 );
buf \U$45628 ( \45988 , \45987 );
_HMUX r8521 ( \45989_nR8521 , \45977 , \45988 , RIc0c97c8_1 );
buf \U$45629 ( \45990 , \45989_nR8521 );
xor \U$45630 ( \45991 , \8208 , \21495 );
buf \U$45631 ( \45992 , \45991 );
not \U$45632 ( \45993 , \29875 );
nand \U$45633 ( \45994 , \43724 , \45993 );
nand \U$45634 ( \45995 , \45300 , \45293 );
or \U$45635 ( \45996 , \45995 , \45302 );
and \U$45636 ( \45997 , \45293 , \45310 );
nor \U$45637 ( \45998 , \45997 , \45318 );
nand \U$45638 ( \45999 , \45996 , \45998 );
not \U$45639 ( \46000 , \45999 );
xor \U$45640 ( \46001 , \45994 , \46000 );
buf \U$45641 ( \46002 , \46001 );
_HMUX r831f ( \46003_nR831f , \45992 , \46002 , RIc0c97c8_1 );
buf \U$45642 ( \46004 , \46003_nR831f );
xor \U$45643 ( \46005 , \8503 , \21493 );
buf \U$45644 ( \46006 , \46005 );
not \U$45645 ( \46007 , \29627 );
nand \U$45646 ( \46008 , \43721 , \46007 );
nand \U$45647 ( \46009 , \45346 , \45339 );
or \U$45648 ( \46010 , \46009 , \45348 );
and \U$45649 ( \46011 , \45339 , \45356 );
nor \U$45650 ( \46012 , \46011 , \45364 );
nand \U$45651 ( \46013 , \46010 , \46012 );
not \U$45652 ( \46014 , \46013 );
xor \U$45653 ( \46015 , \46008 , \46014 );
buf \U$45654 ( \46016 , \46015 );
_HMUX r8114 ( \46017_nR8114 , \46006 , \46016 , RIc0c97c8_1 );
buf \U$45655 ( \46018 , \46017_nR8114 );
xor \U$45656 ( \46019 , \8786 , \21491 );
buf \U$45657 ( \46020 , \46019 );
not \U$45658 ( \46021 , \29378 );
nand \U$45659 ( \46022 , \43719 , \46021 );
nand \U$45660 ( \46023 , \45386 , \45383 );
or \U$45661 ( \46024 , \46023 , \43526 );
and \U$45662 ( \46025 , \45383 , \45390 );
nor \U$45663 ( \46026 , \46025 , \45394 );
nand \U$45664 ( \46027 , \46024 , \46026 );
not \U$45665 ( \46028 , \46027 );
xor \U$45666 ( \46029 , \46022 , \46028 );
buf \U$45667 ( \46030 , \46029 );
_HMUX r7f04 ( \46031_nR7f04 , \46020 , \46030 , RIc0c97c8_1 );
buf \U$45668 ( \46032 , \46031_nR7f04 );
xor \U$45669 ( \46033 , \9074 , \21489 );
buf \U$45670 ( \46034 , \46033 );
not \U$45671 ( \46035 , \29120 );
nand \U$45672 ( \46036 , \43713 , \46035 );
nand \U$45673 ( \46037 , \45412 , \45409 );
or \U$45674 ( \46038 , \46037 , \44014 );
and \U$45675 ( \46039 , \45409 , \45416 );
nor \U$45676 ( \46040 , \46039 , \45420 );
nand \U$45677 ( \46041 , \46038 , \46040 );
not \U$45678 ( \46042 , \46041 );
xor \U$45679 ( \46043 , \46036 , \46042 );
buf \U$45680 ( \46044 , \46043 );
_HMUX r7ced ( \46045_nR7ced , \46034 , \46044 , RIc0c97c8_1 );
buf \U$45681 ( \46046 , \46045_nR7ced );
xor \U$45682 ( \46047 , \9375 , \21487 );
buf \U$45683 ( \46048 , \46047 );
not \U$45684 ( \46049 , \28860 );
nand \U$45685 ( \46050 , \43711 , \46049 );
nand \U$45686 ( \46051 , \45438 , \45435 );
or \U$45687 ( \46052 , \46051 , \44314 );
and \U$45688 ( \46053 , \45435 , \45442 );
nor \U$45689 ( \46054 , \46053 , \45446 );
nand \U$45690 ( \46055 , \46052 , \46054 );
not \U$45691 ( \46056 , \46055 );
xor \U$45692 ( \46057 , \46050 , \46056 );
buf \U$45693 ( \46058 , \46057 );
_HMUX r7acb ( \46059_nR7acb , \46048 , \46058 , RIc0c97c8_1 );
buf \U$45694 ( \46060 , \46059_nR7acb );
xor \U$45695 ( \46061 , \9671 , \21485 );
buf \U$45696 ( \46062 , \46061 );
not \U$45697 ( \46063 , \28595 );
nand \U$45698 ( \46064 , \43708 , \46063 );
nand \U$45699 ( \46065 , \45464 , \45461 );
or \U$45700 ( \46066 , \46065 , \44503 );
and \U$45701 ( \46067 , \45461 , \45468 );
nor \U$45702 ( \46068 , \46067 , \45472 );
nand \U$45703 ( \46069 , \46066 , \46068 );
not \U$45704 ( \46070 , \46069 );
xor \U$45705 ( \46071 , \46064 , \46070 );
buf \U$45706 ( \46072 , \46071 );
_HMUX r789f ( \46073_nR789f , \46062 , \46072 , RIc0c97c8_1 );
buf \U$45707 ( \46074 , \46073_nR789f );
xor \U$45708 ( \46075 , \9980 , \21483 );
buf \U$45709 ( \46076 , \46075 );
not \U$45710 ( \46077 , \28328 );
nand \U$45711 ( \46078 , \43706 , \46077 );
nand \U$45712 ( \46079 , \45490 , \45487 );
or \U$45713 ( \46080 , \46079 , \44654 );
and \U$45714 ( \46081 , \45487 , \45494 );
nor \U$45715 ( \46082 , \46081 , \45498 );
nand \U$45716 ( \46083 , \46080 , \46082 );
not \U$45717 ( \46084 , \46083 );
xor \U$45718 ( \46085 , \46078 , \46084 );
buf \U$45719 ( \46086 , \46085 );
_HMUX r766c ( \46087_nR766c , \46076 , \46086 , RIc0c97c8_1 );
buf \U$45720 ( \46088 , \46087_nR766c );
xor \U$45721 ( \46089 , \10298 , \21481 );
buf \U$45722 ( \46090 , \46089 );
not \U$45723 ( \46091 , \28051 );
nand \U$45724 ( \46092 , \43702 , \46091 );
nand \U$45725 ( \46093 , \45516 , \45513 );
or \U$45726 ( \46094 , \46093 , \44749 );
and \U$45727 ( \46095 , \45513 , \45520 );
nor \U$45728 ( \46096 , \46095 , \45524 );
nand \U$45729 ( \46097 , \46094 , \46096 );
not \U$45730 ( \46098 , \46097 );
xor \U$45731 ( \46099 , \46092 , \46098 );
buf \U$45732 ( \46100 , \46099 );
_HMUX r742e ( \46101_nR742e , \46090 , \46100 , RIc0c97c8_1 );
buf \U$45733 ( \46102 , \46101_nR742e );
xor \U$45734 ( \46103 , \10614 , \21479 );
buf \U$45735 ( \46104 , \46103 );
not \U$45736 ( \46105 , \27774 );
nand \U$45737 ( \46106 , \43700 , \46105 );
nand \U$45738 ( \46107 , \45542 , \45539 );
or \U$45739 ( \46108 , \46107 , \44842 );
and \U$45740 ( \46109 , \45539 , \45545 );
nor \U$45741 ( \46110 , \46109 , \45549 );
nand \U$45742 ( \46111 , \46108 , \46110 );
not \U$45743 ( \46112 , \46111 );
xor \U$45744 ( \46113 , \46106 , \46112 );
buf \U$45745 ( \46114 , \46113 );
_HMUX r71e6 ( \46115_nR71e6 , \46104 , \46114 , RIc0c97c8_1 );
buf \U$45746 ( \46116 , \46115_nR71e6 );
xor \U$45747 ( \46117 , \10927 , \21477 );
buf \U$45748 ( \46118 , \46117 );
not \U$45749 ( \46119 , \27488 );
nand \U$45750 ( \46120 , \43697 , \46119 );
nand \U$45751 ( \46121 , \45567 , \45564 );
or \U$45752 ( \46122 , \46121 , \44935 );
and \U$45753 ( \46123 , \45564 , \45570 );
nor \U$45754 ( \46124 , \46123 , \45574 );
nand \U$45755 ( \46125 , \46122 , \46124 );
not \U$45756 ( \46126 , \46125 );
xor \U$45757 ( \46127 , \46120 , \46126 );
buf \U$45758 ( \46128 , \46127 );
_HMUX r6f94 ( \46129_nR6f94 , \46118 , \46128 , RIc0c97c8_1 );
buf \U$45759 ( \46130 , \46129_nR6f94 );
xor \U$45760 ( \46131 , \11238 , \21475 );
buf \U$45761 ( \46132 , \46131 );
not \U$45762 ( \46133 , \27198 );
nand \U$45763 ( \46134 , \43695 , \46133 );
nand \U$45764 ( \46135 , \45592 , \45589 );
or \U$45765 ( \46136 , \46135 , \45012 );
and \U$45766 ( \46137 , \45589 , \45595 );
nor \U$45767 ( \46138 , \46137 , \45599 );
nand \U$45768 ( \46139 , \46136 , \46138 );
not \U$45769 ( \46140 , \46139 );
xor \U$45770 ( \46141 , \46134 , \46140 );
buf \U$45771 ( \46142 , \46141 );
_HMUX r6d35 ( \46143_nR6d35 , \46132 , \46142 , RIc0c97c8_1 );
buf \U$45772 ( \46144 , \46143_nR6d35 );
xor \U$45773 ( \46145 , \11556 , \21473 );
buf \U$45774 ( \46146 , \46145 );
not \U$45775 ( \46147 , \26898 );
nand \U$45776 ( \46148 , \43690 , \46147 );
nand \U$45777 ( \46149 , \45617 , \45614 );
or \U$45778 ( \46150 , \46149 , \45061 );
and \U$45779 ( \46151 , \45614 , \45620 );
nor \U$45780 ( \46152 , \46151 , \45624 );
nand \U$45781 ( \46153 , \46150 , \46152 );
not \U$45782 ( \46154 , \46153 );
xor \U$45783 ( \46155 , \46148 , \46154 );
buf \U$45784 ( \46156 , \46155 );
_HMUX r6aca ( \46157_nR6aca , \46146 , \46156 , RIc0c97c8_1 );
buf \U$45785 ( \46158 , \46157_nR6aca );
xor \U$45786 ( \46159 , \11872 , \21471 );
buf \U$45787 ( \46160 , \46159 );
not \U$45788 ( \46161 , \26597 );
nand \U$45789 ( \46162 , \43688 , \46161 );
nand \U$45790 ( \46163 , \45642 , \45639 );
or \U$45791 ( \46164 , \46163 , \44305 );
and \U$45792 ( \46165 , \45639 , \45645 );
nor \U$45793 ( \46166 , \46165 , \45649 );
nand \U$45794 ( \46167 , \46164 , \46166 );
not \U$45795 ( \46168 , \46167 );
xor \U$45796 ( \46169 , \46162 , \46168 );
buf \U$45797 ( \46170 , \46169 );
_HMUX r6854 ( \46171_nR6854 , \46160 , \46170 , RIc0c97c8_1 );
buf \U$45798 ( \46172 , \46171_nR6854 );
xor \U$45799 ( \46173 , \12172 , \21469 );
buf \U$45800 ( \46174 , \46173 );
not \U$45801 ( \46175 , \26291 );
nand \U$45802 ( \46176 , \43685 , \46175 );
nand \U$45803 ( \46177 , \45667 , \45664 );
or \U$45804 ( \46178 , \46177 , \44494 );
and \U$45805 ( \46179 , \45664 , \45670 );
nor \U$45806 ( \46180 , \46179 , \45674 );
nand \U$45807 ( \46181 , \46178 , \46180 );
not \U$45808 ( \46182 , \46181 );
xor \U$45809 ( \46183 , \46176 , \46182 );
buf \U$45810 ( \46184 , \46183 );
_HMUX r65d5 ( \46185_nR65d5 , \46174 , \46184 , RIc0c97c8_1 );
buf \U$45811 ( \46186 , \46185_nR65d5 );
xor \U$45812 ( \46187 , \12488 , \21467 );
buf \U$45813 ( \46188 , \46187 );
not \U$45814 ( \46189 , \25981 );
nand \U$45815 ( \46190 , \43683 , \46189 );
nand \U$45816 ( \46191 , \45692 , \45689 );
or \U$45817 ( \46192 , \46191 , \43490 );
and \U$45818 ( \46193 , \45689 , \45695 );
nor \U$45819 ( \46194 , \46193 , \45699 );
nand \U$45820 ( \46195 , \46192 , \46194 );
not \U$45821 ( \46196 , \46195 );
xor \U$45822 ( \46197 , \46190 , \46196 );
buf \U$45823 ( \46198 , \46197 );
_HMUX r634e ( \46199_nR634e , \46188 , \46198 , RIc0c97c8_1 );
buf \U$45824 ( \46200 , \46199_nR634e );
xor \U$45825 ( \46201 , \12773 , \21465 );
buf \U$45826 ( \46202 , \46201 );
not \U$45827 ( \46203 , \25668 );
nand \U$45828 ( \46204 , \43679 , \46203 );
nand \U$45829 ( \46205 , \45717 , \45714 );
or \U$45830 ( \46206 , \46205 , \43486 );
and \U$45831 ( \46207 , \45714 , \45720 );
nor \U$45832 ( \46208 , \46207 , \45724 );
nand \U$45833 ( \46209 , \46206 , \46208 );
not \U$45834 ( \46210 , \46209 );
xor \U$45835 ( \46211 , \46204 , \46210 );
buf \U$45836 ( \46212 , \46211 );
_HMUX r60c1 ( \46213_nR60c1 , \46202 , \46212 , RIc0c97c8_1 );
buf \U$45837 ( \46214 , \46213_nR60c1 );
xor \U$45838 ( \46215 , \13052 , \21463 );
buf \U$45839 ( \46216 , \46215 );
not \U$45840 ( \46217 , \25353 );
nand \U$45841 ( \46218 , \43677 , \46217 );
and \U$45842 ( \46219 , \45739 , \45743 );
nor \U$45843 ( \46220 , \46219 , \45747 );
xor \U$45844 ( \46221 , \46218 , \46220 );
buf \U$45845 ( \46222 , \46221 );
_HMUX r5e2f ( \46223_nR5e2f , \46216 , \46222 , RIc0c97c8_1 );
buf \U$45846 ( \46224 , \46223_nR5e2f );
xor \U$45847 ( \46225 , \13355 , \21461 );
buf \U$45848 ( \46226 , \46225 );
not \U$45849 ( \46227 , \25038 );
nand \U$45850 ( \46228 , \43674 , \46227 );
and \U$45851 ( \46229 , \45762 , \45766 );
nor \U$45852 ( \46230 , \46229 , \45770 );
xor \U$45853 ( \46231 , \46228 , \46230 );
buf \U$45854 ( \46232 , \46231 );
_HMUX r5ba1 ( \46233_nR5ba1 , \46226 , \46232 , RIc0c97c8_1 );
buf \U$45855 ( \46234 , \46233_nR5ba1 );
xor \U$45856 ( \46235 , \13626 , \21459 );
buf \U$45857 ( \46236 , \46235 );
not \U$45858 ( \46237 , \24724 );
nand \U$45859 ( \46238 , \43672 , \46237 );
xor \U$45860 ( \46239 , \46238 , \43670 );
buf \U$45861 ( \46240 , \46239 );
_HMUX r590c ( \46241_nR590c , \46236 , \46240 , RIc0c97c8_1 );
buf \U$45862 ( \46242 , \46241_nR590c );
xor \U$45863 ( \46243 , \13902 , \21457 );
buf \U$45864 ( \46244 , \46243 );
not \U$45865 ( \46245 , \41857 );
nand \U$45866 ( \46246 , \43664 , \46245 );
xor \U$45867 ( \46247 , \46246 , \44110 );
buf \U$45868 ( \46248 , \46247 );
_HMUX r5671 ( \46249_nR5671 , \46244 , \46248 , RIc0c97c8_1 );
buf \U$45869 ( \46250 , \46249_nR5671 );
xor \U$45870 ( \46251 , \14179 , \21455 );
buf \U$45871 ( \46252 , \46251 );
not \U$45872 ( \46253 , \41854 );
nand \U$45873 ( \46254 , \43662 , \46253 );
xor \U$45874 ( \46255 , \46254 , \44362 );
buf \U$45875 ( \46256 , \46255 );
_HMUX r53dc ( \46257_nR53dc , \46252 , \46256 , RIc0c97c8_1 );
buf \U$45876 ( \46258 , \46257_nR53dc );
xor \U$45877 ( \46259 , \14449 , \21453 );
buf \U$45878 ( \46260 , \46259 );
not \U$45879 ( \46261 , \41841 );
nand \U$45880 ( \46262 , \43659 , \46261 );
xor \U$45881 ( \46263 , \46262 , \44551 );
buf \U$45882 ( \46264 , \46263 );
_HMUX r5155 ( \46265_nR5155 , \46260 , \46264 , RIc0c97c8_1 );
buf \U$45883 ( \46266 , \46265_nR5155 );
xor \U$45884 ( \46267 , \14711 , \21451 );
buf \U$45885 ( \46268 , \46267 );
not \U$45886 ( \46269 , \41819 );
nand \U$45887 ( \46270 , \43657 , \46269 );
xor \U$45888 ( \46271 , \46270 , \44678 );
buf \U$45889 ( \46272 , \46271 );
_HMUX r4ed4 ( \46273_nR4ed4 , \46268 , \46272 , RIc0c97c8_1 );
buf \U$45890 ( \46274 , \46273_nR4ed4 );
xor \U$45891 ( \46275 , \14972 , \21449 );
buf \U$45892 ( \46276 , \46275 );
not \U$45893 ( \46277 , \41784 );
nand \U$45894 ( \46278 , \43653 , \46277 );
xor \U$45895 ( \46279 , \46278 , \44773 );
buf \U$45896 ( \46280 , \46279 );
_HMUX r4c61 ( \46281_nR4c61 , \46276 , \46280 , RIc0c97c8_1 );
buf \U$45897 ( \46282 , \46281_nR4c61 );
xor \U$45898 ( \46283 , \14980 , \21447 );
buf \U$45899 ( \46284 , \46283 );
not \U$45900 ( \46285 , \41739 );
nand \U$45901 ( \46286 , \43651 , \46285 );
xor \U$45902 ( \46287 , \46286 , \44866 );
buf \U$45903 ( \46288 , \46287 );
_HMUX r49f4 ( \46289_nR49f4 , \46284 , \46288 , RIc0c97c8_1 );
buf \U$45904 ( \46290 , \46289_nR49f4 );
xor \U$45905 ( \46291 , \15226 , \21445 );
buf \U$45906 ( \46292 , \46291 );
not \U$45907 ( \46293 , \41667 );
nand \U$45908 ( \46294 , \43648 , \46293 );
xor \U$45909 ( \46295 , \46294 , \44959 );
buf \U$45910 ( \46296 , \46295 );
_HMUX r4795 ( \46297_nR4795 , \46292 , \46296 , RIc0c97c8_1 );
buf \U$45911 ( \46298 , \46297_nR4795 );
xor \U$45912 ( \46299 , \15456 , \21443 );
buf \U$45913 ( \46300 , \46299 );
not \U$45914 ( \46301 , \41560 );
nand \U$45915 ( \46302 , \43646 , \46301 );
xor \U$45916 ( \46303 , \46302 , \45024 );
buf \U$45917 ( \46304 , \46303 );
_HMUX r453c ( \46305_nR453c , \46300 , \46304 , RIc0c97c8_1 );
buf \U$45918 ( \46306 , \46305_nR453c );
xor \U$45919 ( \46307 , \15706 , \21441 );
buf \U$45920 ( \46308 , \46307 );
not \U$45921 ( \46309 , \41394 );
nand \U$45922 ( \46310 , \43641 , \46309 );
xor \U$45923 ( \46311 , \46310 , \45073 );
buf \U$45924 ( \46312 , \46311 );
_HMUX r42f1 ( \46313_nR42f1 , \46308 , \46312 , RIc0c97c8_1 );
buf \U$45925 ( \46314 , \46313_nR42f1 );
xor \U$45926 ( \46315 , \15931 , \21439 );
buf \U$45927 ( \46316 , \46315 );
not \U$45928 ( \46317 , \41129 );
nand \U$45929 ( \46318 , \43639 , \46317 );
xor \U$45930 ( \46319 , \46318 , \45121 );
buf \U$45931 ( \46320 , \46319 );
_HMUX r40ac ( \46321_nR40ac , \46316 , \46320 , RIc0c97c8_1 );
buf \U$45932 ( \46322 , \46321_nR40ac );
xor \U$45933 ( \46323 , \16150 , \21437 );
buf \U$45934 ( \46324 , \46323 );
not \U$45935 ( \46325 , \40867 );
nand \U$45936 ( \46326 , \43636 , \46325 );
xor \U$45937 ( \46327 , \46326 , \45169 );
buf \U$45938 ( \46328 , \46327 );
_HMUX r3e75 ( \46329_nR3e75 , \46324 , \46328 , RIc0c97c8_1 );
buf \U$45939 ( \46330 , \46329_nR3e75 );
xor \U$45940 ( \46331 , \16380 , \21435 );
buf \U$45941 ( \46332 , \46331 );
not \U$45942 ( \46333 , \40612 );
nand \U$45943 ( \46334 , \43634 , \46333 );
xor \U$45944 ( \46335 , \46334 , \45217 );
buf \U$45945 ( \46336 , \46335 );
_HMUX r3c44 ( \46337_nR3c44 , \46332 , \46336 , RIc0c97c8_1 );
buf \U$45946 ( \46338 , \46337_nR3c44 );
xor \U$45947 ( \46339 , \16611 , \21433 );
buf \U$45948 ( \46340 , \46339 );
not \U$45949 ( \46341 , \40359 );
nand \U$45950 ( \46342 , \43630 , \46341 );
xor \U$45951 ( \46343 , \46342 , \45265 );
buf \U$45952 ( \46344 , \46343 );
_HMUX r3a21 ( \46345_nR3a21 , \46340 , \46344 , RIc0c97c8_1 );
buf \U$45953 ( \46346 , \46345_nR3a21 );
xor \U$45954 ( \46347 , \16822 , \21431 );
buf \U$45955 ( \46348 , \46347 );
not \U$45956 ( \46349 , \40114 );
nand \U$45957 ( \46350 , \43628 , \46349 );
xor \U$45958 ( \46351 , \46350 , \45311 );
buf \U$45959 ( \46352 , \46351 );
_HMUX r3804 ( \46353_nR3804 , \46348 , \46352 , RIc0c97c8_1 );
buf \U$45960 ( \46354 , \46353_nR3804 );
xor \U$45961 ( \46355 , \17035 , \21429 );
buf \U$45962 ( \46356 , \46355 );
not \U$45963 ( \46357 , \39872 );
nand \U$45964 ( \46358 , \43625 , \46357 );
xor \U$45965 ( \46359 , \46358 , \45357 );
buf \U$45966 ( \46360 , \46359 );
_HMUX r35f4 ( \46361_nR35f4 , \46356 , \46360 , RIc0c97c8_1 );
buf \U$45967 ( \46362 , \46361_nR35f4 );
xor \U$45968 ( \46363 , \17232 , \21427 );
buf \U$45969 ( \46364 , \46363 );
not \U$45970 ( \46365 , \39637 );
nand \U$45971 ( \46366 , \43623 , \46365 );
xor \U$45972 ( \46367 , \46366 , \45391 );
buf \U$45973 ( \46368 , \46367 );
_HMUX r33ea ( \46369_nR33ea , \46364 , \46368 , RIc0c97c8_1 );
buf \U$45974 ( \46370 , \46369_nR33ea );
xor \U$45975 ( \46371 , \17428 , \21425 );
buf \U$45976 ( \46372 , \46371 );
not \U$45977 ( \46373 , \39402 );
nand \U$45978 ( \46374 , \43617 , \46373 );
xor \U$45979 ( \46375 , \46374 , \45417 );
buf \U$45980 ( \46376 , \46375 );
_HMUX r31ee ( \46377_nR31ee , \46372 , \46376 , RIc0c97c8_1 );
buf \U$45981 ( \46378 , \46377_nR31ee );
xor \U$45982 ( \46379 , \17636 , \21423 );
buf \U$45983 ( \46380 , \46379 );
not \U$45984 ( \46381 , \39177 );
nand \U$45985 ( \46382 , \43615 , \46381 );
xor \U$45986 ( \46383 , \46382 , \45443 );
buf \U$45987 ( \46384 , \46383 );
_HMUX r2ff8 ( \46385_nR2ff8 , \46380 , \46384 , RIc0c97c8_1 );
buf \U$45988 ( \46386 , \46385_nR2ff8 );
xor \U$45989 ( \46387 , \17821 , \21421 );
buf \U$45990 ( \46388 , \46387 );
not \U$45991 ( \46389 , \38955 );
nand \U$45992 ( \46390 , \43612 , \46389 );
xor \U$45993 ( \46391 , \46390 , \45469 );
buf \U$45994 ( \46392 , \46391 );
_HMUX r2e10 ( \46393_nR2e10 , \46388 , \46392 , RIc0c97c8_1 );
buf \U$45995 ( \46394 , \46393_nR2e10 );
xor \U$45996 ( \46395 , \18008 , \21419 );
buf \U$45997 ( \46396 , \46395 );
not \U$45998 ( \46397 , \38737 );
nand \U$45999 ( \46398 , \43610 , \46397 );
xor \U$46000 ( \46399 , \46398 , \45495 );
buf \U$46001 ( \46400 , \46399 );
_HMUX r2c28 ( \46401_nR2c28 , \46396 , \46400 , RIc0c97c8_1 );
buf \U$46002 ( \46402 , \46401_nR2c28 );
xor \U$46003 ( \46403 , \18198 , \21417 );
buf \U$46004 ( \46404 , \46403 );
not \U$46005 ( \46405 , \38525 );
nand \U$46006 ( \46406 , \43606 , \46405 );
xor \U$46007 ( \46407 , \46406 , \45521 );
buf \U$46008 ( \46408 , \46407 );
_HMUX r2a56 ( \46409_nR2a56 , \46404 , \46408 , RIc0c97c8_1 );
buf \U$46009 ( \46410 , \46409_nR2a56 );
xor \U$46010 ( \46411 , \18374 , \21415 );
buf \U$46011 ( \46412 , \46411 );
not \U$46012 ( \46413 , \38320 );
nand \U$46013 ( \46414 , \43604 , \46413 );
xor \U$46014 ( \46415 , \46414 , \45546 );
buf \U$46015 ( \46416 , \46415 );
_HMUX r2888 ( \46417_nR2888 , \46412 , \46416 , RIc0c97c8_1 );
buf \U$46016 ( \46418 , \46417_nR2888 );
xor \U$46017 ( \46419 , \18545 , \21413 );
buf \U$46018 ( \46420 , \46419 );
not \U$46019 ( \46421 , \38118 );
nand \U$46020 ( \46422 , \43601 , \46421 );
xor \U$46021 ( \46423 , \46422 , \45571 );
buf \U$46022 ( \46424 , \46423 );
_HMUX r26c9 ( \46425_nR26c9 , \46420 , \46424 , RIc0c97c8_1 );
buf \U$46023 ( \46426 , \46425_nR26c9 );
xor \U$46024 ( \46427 , \18553 , \21411 );
buf \U$46025 ( \46428 , \46427 );
not \U$46026 ( \46429 , \37923 );
nand \U$46027 ( \46430 , \43599 , \46429 );
xor \U$46028 ( \46431 , \46430 , \45596 );
buf \U$46029 ( \46432 , \46431 );
_HMUX r2510 ( \46433_nR2510 , \46428 , \46432 , RIc0c97c8_1 );
buf \U$46030 ( \46434 , \46433_nR2510 );
xor \U$46031 ( \46435 , \18721 , \21409 );
buf \U$46032 ( \46436 , \46435 );
not \U$46033 ( \46437 , \37729 );
nand \U$46034 ( \46438 , \43594 , \46437 );
xor \U$46035 ( \46439 , \46438 , \45621 );
buf \U$46036 ( \46440 , \46439 );
_HMUX r2365 ( \46441_nR2365 , \46436 , \46440 , RIc0c97c8_1 );
buf \U$46037 ( \46442 , \46441_nR2365 );
xor \U$46038 ( \46443 , \18861 , \21407 );
buf \U$46039 ( \46444 , \46443 );
not \U$46040 ( \46445 , \37544 );
nand \U$46041 ( \46446 , \43592 , \46445 );
xor \U$46042 ( \46447 , \46446 , \45646 );
buf \U$46043 ( \46448 , \46447 );
_HMUX r21c0 ( \46449_nR21c0 , \46444 , \46448 , RIc0c97c8_1 );
buf \U$46044 ( \46450 , \46449_nR21c0 );
xor \U$46045 ( \46451 , \19013 , \21405 );
buf \U$46046 ( \46452 , \46451 );
not \U$46047 ( \46453 , \37362 );
nand \U$46048 ( \46454 , \43589 , \46453 );
xor \U$46049 ( \46455 , \46454 , \45671 );
buf \U$46050 ( \46456 , \46455 );
_HMUX r2029 ( \46457_nR2029 , \46452 , \46456 , RIc0c97c8_1 );
buf \U$46051 ( \46458 , \46457_nR2029 );
xor \U$46052 ( \46459 , \19177 , \21403 );
buf \U$46053 ( \46460 , \46459 );
not \U$46054 ( \46461 , \37187 );
nand \U$46055 ( \46462 , \43587 , \46461 );
xor \U$46056 ( \46463 , \46462 , \45696 );
buf \U$46057 ( \46464 , \46463 );
_HMUX r1e98 ( \46465_nR1e98 , \46460 , \46464 , RIc0c97c8_1 );
buf \U$46058 ( \46466 , \46465_nR1e98 );
xor \U$46059 ( \46467 , \19316 , \21401 );
buf \U$46060 ( \46468 , \46467 );
not \U$46061 ( \46469 , \37014 );
nand \U$46062 ( \46470 , \43583 , \46469 );
xor \U$46063 ( \46471 , \46470 , \45721 );
buf \U$46064 ( \46472 , \46471 );
_HMUX r1d15 ( \46473_nR1d15 , \46468 , \46472 , RIc0c97c8_1 );
buf \U$46065 ( \46474 , \46473_nR1d15 );
xor \U$46066 ( \46475 , \19441 , \21399 );
buf \U$46067 ( \46476 , \46475 );
not \U$46068 ( \46477 , \36849 );
nand \U$46069 ( \46478 , \43581 , \46477 );
xor \U$46070 ( \46479 , \46478 , \45744 );
buf \U$46071 ( \46480 , \46479 );
_HMUX r1b98 ( \46481_nR1b98 , \46476 , \46480 , RIc0c97c8_1 );
buf \U$46072 ( \46482 , \46481_nR1b98 );
xor \U$46073 ( \46483 , \19585 , \21397 );
buf \U$46074 ( \46484 , \46483 );
not \U$46075 ( \46485 , \36687 );
nand \U$46076 ( \46486 , \43578 , \46485 );
xor \U$46077 ( \46487 , \46486 , \45767 );
buf \U$46078 ( \46488 , \46487 );
_HMUX r1a2b ( \46489_nR1a2b , \46484 , \46488 , RIc0c97c8_1 );
buf \U$46079 ( \46490 , \46489_nR1a2b );
xor \U$46080 ( \46491 , \19709 , \21395 );
buf \U$46081 ( \46492 , \46491 );
not \U$46082 ( \46493 , \36532 );
nand \U$46083 ( \46494 , \43576 , \46493 );
xor \U$46084 ( \46495 , \46494 , \45786 );
buf \U$46085 ( \46496 , \46495 );
_HMUX r18c4 ( \46497_nR18c4 , \46492 , \46496 , RIc0c97c8_1 );
buf \U$46086 ( \46498 , \46497_nR18c4 );
xor \U$46087 ( \46499 , \19849 , \21393 );
buf \U$46088 ( \46500 , \46499 );
not \U$46089 ( \46501 , \43170 );
nand \U$46090 ( \46502 , \43569 , \46501 );
xor \U$46091 ( \46503 , \46502 , \45801 );
buf \U$46092 ( \46504 , \46503 );
_HMUX r176b ( \46505_nR176b , \46500 , \46504 , RIc0c97c8_1 );
buf \U$46093 ( \46506 , \46505_nR176b );
xor \U$46094 ( \46507 , \19973 , \21391 );
buf \U$46095 ( \46508 , \46507 );
not \U$46096 ( \46509 , \43163 );
nand \U$46097 ( \46510 , \43567 , \46509 );
xor \U$46098 ( \46511 , \46510 , \45816 );
buf \U$46099 ( \46512 , \46511 );
_HMUX r1618 ( \46513_nR1618 , \46508 , \46512 , RIc0c97c8_1 );
buf \U$46100 ( \46514 , \46513_nR1618 );
xor \U$46101 ( \46515 , \20088 , \21389 );
buf \U$46102 ( \46516 , \46515 );
not \U$46103 ( \46517 , \43148 );
nand \U$46104 ( \46518 , \43564 , \46517 );
xor \U$46105 ( \46519 , \46518 , \45831 );
buf \U$46106 ( \46520 , \46519 );
_HMUX r14d3 ( \46521_nR14d3 , \46516 , \46520 , RIc0c97c8_1 );
buf \U$46107 ( \46522 , \46521_nR14d3 );
xor \U$46108 ( \46523 , \20096 , \21387 );
buf \U$46109 ( \46524 , \46523 );
not \U$46110 ( \46525 , \43123 );
nand \U$46111 ( \46526 , \43562 , \46525 );
xor \U$46112 ( \46527 , \46526 , \45846 );
buf \U$46113 ( \46528 , \46527 );
_HMUX r1394 ( \46529_nR1394 , \46524 , \46528 , RIc0c97c8_1 );
buf \U$46114 ( \46530 , \46529_nR1394 );
xor \U$46115 ( \46531 , \20192 , \21385 );
buf \U$46116 ( \46532 , \46531 );
not \U$46117 ( \46533 , \43088 );
nand \U$46118 ( \46534 , \43558 , \46533 );
xor \U$46119 ( \46535 , \46534 , \45861 );
buf \U$46120 ( \46536 , \46535 );
_HMUX r1263 ( \46537_nR1263 , \46532 , \46536 , RIc0c97c8_1 );
buf \U$46121 ( \46538 , \46537_nR1263 );
xor \U$46122 ( \46539 , \20307 , \21383 );
buf \U$46123 ( \46540 , \46539 );
not \U$46124 ( \46541 , \43043 );
nand \U$46125 ( \46542 , \43556 , \46541 );
xor \U$46126 ( \46543 , \46542 , \45876 );
buf \U$46127 ( \46544 , \46543 );
_HMUX r1138 ( \46545_nR1138 , \46540 , \46544 , RIc0c97c8_1 );
buf \U$46128 ( \46546 , \46545_nR1138 );
xor \U$46129 ( \46547 , \20395 , \21381 );
buf \U$46130 ( \46548 , \46547 );
not \U$46131 ( \46549 , \42969 );
nand \U$46132 ( \46550 , \43553 , \46549 );
xor \U$46133 ( \46551 , \46550 , \45891 );
buf \U$46134 ( \46552 , \46551 );
_HMUX r101b ( \46553_nR101b , \46548 , \46552 , RIc0c97c8_1 );
buf \U$46135 ( \46554 , \46553_nR101b );
xor \U$46136 ( \46555 , \20487 , \21379 );
buf \U$46137 ( \46556 , \46555 );
not \U$46138 ( \46557 , \42854 );
nand \U$46139 ( \46558 , \43551 , \46557 );
xor \U$46140 ( \46559 , \46558 , \45906 );
buf \U$46141 ( \46560 , \46559 );
_HMUX rf04 ( \46561_nRf04 , \46556 , \46560 , RIc0c97c8_1 );
buf \U$46142 ( \46562 , \46561_nRf04 );
xor \U$46143 ( \46563 , \20575 , \21377 );
buf \U$46144 ( \46564 , \46563 );
not \U$46145 ( \46565 , \42740 );
nand \U$46146 ( \46566 , \43546 , \46565 );
xor \U$46147 ( \46567 , \46566 , \45921 );
buf \U$46148 ( \46568 , \46567 );
_HMUX rdfb ( \46569_nRdfb , \46564 , \46568 , RIc0c97c8_1 );
buf \U$46149 ( \46570 , \46569_nRdfb );
xor \U$46150 ( \46571 , \20670 , \21375 );
buf \U$46151 ( \46572 , \46571 );
not \U$46152 ( \46573 , \42635 );
nand \U$46153 ( \46574 , \43544 , \46573 );
xor \U$46154 ( \46575 , \46574 , \45936 );
buf \U$46155 ( \46576 , \46575 );
_HMUX rcf8 ( \46577_nRcf8 , \46572 , \46576 , RIc0c97c8_1 );
buf \U$46156 ( \46578 , \46577_nRcf8 );
xor \U$46157 ( \46579 , \20750 , \21373 );
buf \U$46158 ( \46580 , \46579 );
not \U$46159 ( \46581 , \42533 );
nand \U$46160 ( \46582 , \43541 , \46581 );
xor \U$46161 ( \46583 , \46582 , \45951 );
buf \U$46162 ( \46584 , \46583 );
_HMUX rc03 ( \46585_nRc03 , \46580 , \46584 , RIc0c97c8_1 );
buf \U$46163 ( \46586 , \46585_nRc03 );
xor \U$46164 ( \46587 , \20829 , \21371 );
buf \U$46165 ( \46588 , \46587 );
not \U$46166 ( \46589 , \42438 );
nand \U$46167 ( \46590 , \43539 , \46589 );
xor \U$46168 ( \46591 , \46590 , \45966 );
buf \U$46169 ( \46592 , \46591 );
_HMUX rb14 ( \46593_nRb14 , \46588 , \46592 , RIc0c97c8_1 );
buf \U$46170 ( \46594 , \46593_nRb14 );
xor \U$46171 ( \46595 , \20837 , \21369 );
buf \U$46172 ( \46596 , \46595 );
not \U$46173 ( \46597 , \42345 );
nand \U$46174 ( \46598 , \43535 , \46597 );
xor \U$46175 ( \46599 , \46598 , \45981 );
buf \U$46176 ( \46600 , \46599 );
_HMUX ra33 ( \46601_nRa33 , \46596 , \46600 , RIc0c97c8_1 );
buf \U$46177 ( \46602 , \46601_nRa33 );
xor \U$46178 ( \46603 , \20896 , \21367 );
buf \U$46179 ( \46604 , \46603 );
not \U$46180 ( \46605 , \42260 );
nand \U$46181 ( \46606 , \43533 , \46605 );
xor \U$46182 ( \46607 , \46606 , \45302 );
buf \U$46183 ( \46608 , \46607 );
_HMUX r958 ( \46609_nR958 , \46604 , \46608 , RIc0c97c8_1 );
buf \U$46184 ( \46610 , \46609_nR958 );
xor \U$46185 ( \46611 , \20951 , \21365 );
buf \U$46186 ( \46612 , \46611 );
not \U$46187 ( \46613 , \42178 );
nand \U$46188 ( \46614 , \43530 , \46613 );
xor \U$46189 ( \46615 , \46614 , \45348 );
buf \U$46190 ( \46616 , \46615 );
_HMUX r88f ( \46617_nR88f , \46612 , \46616 , RIc0c97c8_1 );
buf \U$46191 ( \46618 , \46617_nR88f );
xor \U$46192 ( \46619 , \21022 , \21363 );
buf \U$46193 ( \46620 , \46619 );
not \U$46194 ( \46621 , \42103 );
nand \U$46195 ( \46622 , \43528 , \46621 );
xor \U$46196 ( \46623 , \46622 , \43526 );
buf \U$46197 ( \46624 , \46623 );
_HMUX r7cc ( \46625_nR7cc , \46620 , \46624 , RIc0c97c8_1 );
buf \U$46198 ( \46626 , \46625_nR7cc );
xor \U$46199 ( \46627 , \21075 , \21361 );
buf \U$46200 ( \46628 , \46627 );
not \U$46201 ( \46629 , \43425 );
nand \U$46202 ( \46630 , \43522 , \46629 );
xor \U$46203 ( \46631 , \46630 , \44014 );
buf \U$46204 ( \46632 , \46631 );
_HMUX r717 ( \46633_nR717 , \46628 , \46632 , RIc0c97c8_1 );
buf \U$46205 ( \46634 , \46633_nR717 );
xor \U$46206 ( \46635 , \21114 , \21359 );
buf \U$46207 ( \46636 , \46635 );
not \U$46208 ( \46637 , \43418 );
nand \U$46209 ( \46638 , \43520 , \46637 );
xor \U$46210 ( \46639 , \46638 , \44314 );
buf \U$46211 ( \46640 , \46639 );
_HMUX r668 ( \46641_nR668 , \46636 , \46640 , RIc0c97c8_1 );
buf \U$46212 ( \46642 , \46641_nR668 );
xor \U$46213 ( \46643 , \21167 , \21357 );
buf \U$46214 ( \46644 , \46643 );
not \U$46215 ( \46645 , \43406 );
nand \U$46216 ( \46646 , \43517 , \46645 );
xor \U$46217 ( \46647 , \46646 , \44503 );
buf \U$46218 ( \46648 , \46647 );
_HMUX r5c6 ( \46649_nR5c6 , \46644 , \46648 , RIc0c97c8_1 );
buf \U$46219 ( \46650 , \46649_nR5c6 );
xor \U$46220 ( \46651 , \21175 , \21355 );
buf \U$46221 ( \46652 , \46651 );
not \U$46222 ( \46653 , \43389 );
nand \U$46223 ( \46654 , \43515 , \46653 );
xor \U$46224 ( \46655 , \46654 , \44654 );
buf \U$46225 ( \46656 , \46655 );
_HMUX r52a ( \46657_nR52a , \46652 , \46656 , RIc0c97c8_1 );
buf \U$46226 ( \46658 , \46657_nR52a );
xor \U$46227 ( \46659 , \21209 , \21353 );
buf \U$46228 ( \46660 , \46659 );
not \U$46229 ( \46661 , \43360 );
nand \U$46230 ( \46662 , \43511 , \46661 );
xor \U$46231 ( \46663 , \46662 , \44749 );
buf \U$46232 ( \46664 , \46663 );
_HMUX r49d ( \46665_nR49d , \46660 , \46664 , RIc0c97c8_1 );
buf \U$46233 ( \46666 , \46665_nR49d );
xor \U$46234 ( \46667 , \21243 , \21351 );
buf \U$46235 ( \46668 , \46667 );
not \U$46236 ( \46669 , \43315 );
nand \U$46237 ( \46670 , \43509 , \46669 );
xor \U$46238 ( \46671 , \46670 , \44842 );
buf \U$46239 ( \46672 , \46671 );
_HMUX r416 ( \46673_nR416 , \46668 , \46672 , RIc0c97c8_1 );
buf \U$46240 ( \46674 , \46673_nR416 );
xor \U$46241 ( \46675 , \21251 , \21349 );
buf \U$46242 ( \46676 , \46675 );
not \U$46243 ( \46677 , \43273 );
nand \U$46244 ( \46678 , \43506 , \46677 );
xor \U$46245 ( \46679 , \46678 , \44935 );
buf \U$46246 ( \46680 , \46679 );
_HMUX r39f ( \46681_nR39f , \46676 , \46680 , RIc0c97c8_1 );
buf \U$46247 ( \46682 , \46681_nR39f );
endmodule

