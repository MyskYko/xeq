//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RI2b5e785ebcf0_2,RI2b5e785ebc78_3,RI2b5e785ebc00_4,RI2b5e785ebb88_5,RI2b5e785ebb10_6,RI2b5e785eba98_7,RI2b5e785eba20_8,RI2b5e785eb9a8_9,RI2b5e785eb930_10,
        RI2b5e785eb8b8_11,RI2b5e785eb840_12,RI2b5e785daa40_28,RI2b5e785ae9b8_600,RI2b5e785aea30_599,RI2b5e785aeaa8_598,RI2b5e785aeb20_597,RI2b5e785aeb98_596,RI2b5e785aec10_595,RI2b5e785aec88_594,
        RI2b5e785aed00_593,RI2b5e785aed78_592,RI2b5e785aedf0_591,RI2b5e785aee68_590,RI2b5e785aeee0_589,RI2b5e785aef58_588,RI2b5e78549540_41,RI2b5e785388a8_54,RI2b5e784a6330_67,RI2b5e78495698_80,
        RI2b5e78495080_93,RI2b5e78403b80_106,RI2b5e775b1e60_119,RI2b5e7750bdf8_132,RI2b5e774ff5d0_145,RI2b5e774f65e8_158,RI2b5e774eabd0_171,RI2b5e774de3a8_184,RI2b5e774d53c0_197,RI2b5e785f4300_210,
        RI2b5e785f3ce8_223,RI2b5e785eb0c0_236,RI2b5e785da9c8_29,RI2b5e785494c8_42,RI2b5e78538830_55,RI2b5e784a62b8_68,RI2b5e78495620_81,RI2b5e78495008_94,RI2b5e78403b08_107,RI2b5e775b1de8_120,
        RI2b5e7750bd80_133,RI2b5e774ff558_146,RI2b5e774f6570_159,RI2b5e774eab58_172,RI2b5e774de330_185,RI2b5e774d5348_198,RI2b5e785f4288_211,RI2b5e785f3658_224,RI2b5e785eb048_237,RI2b5e785da950_30,
        RI2b5e78549450_43,RI2b5e785387b8_56,RI2b5e784a6240_69,RI2b5e784955a8_82,RI2b5e78494f90_95,RI2b5e78403a90_108,RI2b5e775b1d70_121,RI2b5e7750bd08_134,RI2b5e774ff4e0_147,RI2b5e774f64f8_160,
        RI2b5e774eaae0_173,RI2b5e774de2b8_186,RI2b5e774d52d0_199,RI2b5e785f4210_212,RI2b5e785eb5e8_225,RI2b5e785e6c50_238,RI2b5e785da8d8_31,RI2b5e785493d8_44,RI2b5e78538740_57,RI2b5e784a61c8_70,
        RI2b5e78495530_83,RI2b5e78494f18_96,RI2b5e78403a18_109,RI2b5e775b1cf8_122,RI2b5e7750bc90_135,RI2b5e774ff468_148,RI2b5e774f6480_161,RI2b5e774eaa68_174,RI2b5e774de240_187,RI2b5e774d5258_200,
        RI2b5e785f4198_213,RI2b5e785eb570_226,RI2b5e785e6bd8_239,RI2b5e785da860_32,RI2b5e78549360_45,RI2b5e785386c8_58,RI2b5e784a6150_71,RI2b5e784954b8_84,RI2b5e78494ea0_97,RI2b5e784039a0_110,
        RI2b5e775b1c80_123,RI2b5e7750bc18_136,RI2b5e774ff3f0_149,RI2b5e774f6408_162,RI2b5e774ea9f0_175,RI2b5e774de1c8_188,RI2b5e774d51e0_201,RI2b5e785f4120_214,RI2b5e785eb4f8_227,RI2b5e785e64d0_240,
        RI2b5e78549900_33,RI2b5e78538c68_46,RI2b5e78538650_59,RI2b5e784a60d8_72,RI2b5e78495440_85,RI2b5e78494e28_98,RI2b5e78403928_111,RI2b5e775b1c08_124,RI2b5e7750bba0_137,RI2b5e774ff378_150,
        RI2b5e774f6390_163,RI2b5e774ea978_176,RI2b5e774de150_189,RI2b5e774d5168_202,RI2b5e785f40a8_215,RI2b5e785eb480_228,RI2b5e785da608_241,RI2b5e78549888_34,RI2b5e78538bf0_47,RI2b5e785385d8_60,
        RI2b5e784a6060_73,RI2b5e784953c8_86,RI2b5e78403ec8_99,RI2b5e775b21a8_112,RI2b5e775b1b90_125,RI2b5e7750bb28_138,RI2b5e774ff300_151,RI2b5e774f6318_164,RI2b5e774ea900_177,RI2b5e774de0d8_190,
        RI2b5e774d50f0_203,RI2b5e785f4030_216,RI2b5e785eb408_229,RI2b5e785da590_242,RI2b5e78549810_35,RI2b5e78538b78_48,RI2b5e78538560_61,RI2b5e784a5fe8_74,RI2b5e78495350_87,RI2b5e78403e50_100,
        RI2b5e775b2130_113,RI2b5e775b1b18_126,RI2b5e7750bab0_139,RI2b5e774ff288_152,RI2b5e774f62a0_165,RI2b5e774ea888_178,RI2b5e774de060_191,RI2b5e774d5078_204,RI2b5e785f3fb8_217,RI2b5e785eb390_230,
        RI2b5e785da518_243,RI2b5e78549798_36,RI2b5e78538b00_49,RI2b5e785384e8_62,RI2b5e784a5f70_75,RI2b5e784952d8_88,RI2b5e78403dd8_101,RI2b5e775b20b8_114,RI2b5e775b1aa0_127,RI2b5e7750ba38_140,
        RI2b5e774ff210_153,RI2b5e774f6228_166,RI2b5e774ea810_179,RI2b5e774ddfe8_192,RI2b5e774d5000_205,RI2b5e785f3f40_218,RI2b5e785eb318_231,RI2b5e785da4a0_244,RI2b5e78549720_37,RI2b5e78538a88_50,
        RI2b5e78538470_63,RI2b5e784a5ef8_76,RI2b5e78495260_89,RI2b5e78403d60_102,RI2b5e775b2040_115,RI2b5e775b1a28_128,RI2b5e7750b9c0_141,RI2b5e774ff198_154,RI2b5e774f61b0_167,RI2b5e774ea798_180,
        RI2b5e774ddf70_193,RI2b5e774d4f88_206,RI2b5e785f3ec8_219,RI2b5e785eb2a0_232,RI2b5e785da428_245,RI2b5e785496a8_38,RI2b5e78538a10_51,RI2b5e785383f8_64,RI2b5e784a5e80_77,RI2b5e784951e8_90,
        RI2b5e78403ce8_103,RI2b5e775b1fc8_116,RI2b5e775b19b0_129,RI2b5e7750b948_142,RI2b5e774ff120_155,RI2b5e774f6138_168,RI2b5e774ea720_181,RI2b5e774ddef8_194,RI2b5e774d4f10_207,RI2b5e785f3e50_220,
        RI2b5e785eb228_233,RI2b5e785da3b0_246,RI2b5e785db148_13,RI2b5e78549630_39,RI2b5e78538998_52,RI2b5e78538380_65,RI2b5e784a5e08_78,RI2b5e78495170_91,RI2b5e78403c70_104,RI2b5e775b1f50_117,
        RI2b5e775b1938_130,RI2b5e7750b8d0_143,RI2b5e774ff0a8_156,RI2b5e774f60c0_169,RI2b5e774ea6a8_182,RI2b5e774dde80_195,RI2b5e774d4e98_208,RI2b5e785f3dd8_221,RI2b5e785eb1b0_234,RI2b5e785da338_247,
        RI2b5e785da248_249,RI2b5e785be750_269,RI2b5e785bc4a0_289,RI2b5e785bbb40_309,RI2b5e785b9c50_329,RI2b5e785b8120_349,RI2b5e785b77c0_369,RI2b5e785b6e60_389,RI2b5e785b56f0_409,RI2b5e785b4d90_429,
        RI2b5e785b39e0_449,RI2b5e785b3080_469,RI2b5e785b2720_489,RI2b5e785b1730_509,RI2b5e785b0dd0_529,RI2b5e785b0470_549,RI2b5e785af840_569,RI2b5e785ebd68_1,RI2b5e785daab8_27,RI2b5e785495b8_40,
        RI2b5e78538920_53,RI2b5e784a63a8_66,RI2b5e78495710_79,RI2b5e784950f8_92,RI2b5e78403bf8_105,RI2b5e775b1ed8_118,RI2b5e775b18c0_131,RI2b5e7750b858_144,RI2b5e774ff030_157,RI2b5e774f6048_170,
        RI2b5e774ea630_183,RI2b5e774dde08_196,RI2b5e774d4e20_209,RI2b5e785f3d60_222,RI2b5e785eb138_235,RI2b5e785da2c0_248,RI2b5e785be7c8_268,RI2b5e785bc518_288,RI2b5e785bbbb8_308,RI2b5e785b9cc8_328,
        RI2b5e785b9368_348,RI2b5e785b7838_368,RI2b5e785b6ed8_388,RI2b5e785b5768_408,RI2b5e785b4e08_428,RI2b5e785b3a58_448,RI2b5e785b30f8_468,RI2b5e785b2798_488,RI2b5e785b17a8_508,RI2b5e785b0e48_528,
        RI2b5e785b04e8_548,RI2b5e785afb88_568,RI2b5e785da1d0_250,RI2b5e785be6d8_270,RI2b5e785bc428_290,RI2b5e785bbac8_310,RI2b5e785b9bd8_330,RI2b5e785b80a8_350,RI2b5e785b7748_370,RI2b5e785b6de8_390,
        RI2b5e785b5678_410,RI2b5e785b4d18_430,RI2b5e785b3968_450,RI2b5e785b3008_470,RI2b5e785b26a8_490,RI2b5e785b16b8_510,RI2b5e785b0d58_530,RI2b5e785b03f8_550,RI2b5e785af7c8_570,RI2b5e785da0e0_252,
        RI2b5e785be5e8_272,RI2b5e785bc338_292,RI2b5e785bb9d8_312,RI2b5e785b9ae8_332,RI2b5e785b7fb8_352,RI2b5e785b7658_372,RI2b5e785b5ee8_392,RI2b5e785b5588_412,RI2b5e785b4c28_432,RI2b5e785b3878_452,
        RI2b5e785b2f18_472,RI2b5e785b25b8_492,RI2b5e785b15c8_512,RI2b5e785b0c68_532,RI2b5e785b0308_552,RI2b5e785af6d8_572,RI2b5e785da158_251,RI2b5e785be660_271,RI2b5e785bc3b0_291,RI2b5e785bba50_311,
        RI2b5e785b9b60_331,RI2b5e785b8030_351,RI2b5e785b76d0_371,RI2b5e785b6d70_391,RI2b5e785b5600_411,RI2b5e785b4ca0_431,RI2b5e785b38f0_451,RI2b5e785b2f90_471,RI2b5e785b2630_491,RI2b5e785b1640_511,
        RI2b5e785b0ce0_531,RI2b5e785b0380_551,RI2b5e785af750_571,RI2b5e785da068_253,RI2b5e785be570_273,RI2b5e785bc2c0_293,RI2b5e785bb960_313,RI2b5e785b9a70_333,RI2b5e785b7f40_353,RI2b5e785b75e0_373,
        RI2b5e785b5e70_393,RI2b5e785b5510_413,RI2b5e785b4bb0_433,RI2b5e785b3800_453,RI2b5e785b2ea0_473,RI2b5e785b2540_493,RI2b5e785b1550_513,RI2b5e785b0bf0_533,RI2b5e785b0290_553,RI2b5e785af660_573,
        RI2b5e785c2bc0_255,RI2b5e785be480_275,RI2b5e785bc1d0_295,RI2b5e785ba2e0_315,RI2b5e785b9980_335,RI2b5e785b7e50_355,RI2b5e785b74f0_375,RI2b5e785b5d80_395,RI2b5e785b5420_415,RI2b5e785b4ac0_435,
        RI2b5e785b3710_455,RI2b5e785b2db0_475,RI2b5e785b2450_495,RI2b5e785b1460_515,RI2b5e785b0b00_535,RI2b5e785b01a0_555,RI2b5e785af570_575,RI2b5e785c2c38_254,RI2b5e785be4f8_274,RI2b5e785bc248_294,
        RI2b5e785ba358_314,RI2b5e785b99f8_334,RI2b5e785b7ec8_354,RI2b5e785b7568_374,RI2b5e785b5df8_394,RI2b5e785b5498_414,RI2b5e785b4b38_434,RI2b5e785b3788_454,RI2b5e785b2e28_474,RI2b5e785b24c8_494,
        RI2b5e785b14d8_514,RI2b5e785b0b78_534,RI2b5e785b0218_554,RI2b5e785af5e8_574,RI2b5e785c0a00_257,RI2b5e785be390_277,RI2b5e785bc0e0_297,RI2b5e785ba1f0_317,RI2b5e785b9890_337,RI2b5e785b7d60_357,
        RI2b5e785b7400_377,RI2b5e785b5c90_397,RI2b5e785b5330_417,RI2b5e785b49d0_437,RI2b5e785b3620_457,RI2b5e785b2cc0_477,RI2b5e785b2360_497,RI2b5e785b1370_517,RI2b5e785b0a10_537,RI2b5e785b00b0_557,
        RI2b5e785af480_577,RI2b5e785c2b48_256,RI2b5e785be408_276,RI2b5e785bc158_296,RI2b5e785ba268_316,RI2b5e785b9908_336,RI2b5e785b7dd8_356,RI2b5e785b7478_376,RI2b5e785b5d08_396,RI2b5e785b53a8_416,
        RI2b5e785b4a48_436,RI2b5e785b3698_456,RI2b5e785b2d38_476,RI2b5e785b23d8_496,RI2b5e785b13e8_516,RI2b5e785b0a88_536,RI2b5e785b0128_556,RI2b5e785af4f8_576,RI2b5e785c0910_259,RI2b5e785be2a0_279,
        RI2b5e785bbff0_299,RI2b5e785ba100_319,RI2b5e785b97a0_339,RI2b5e785b7c70_359,RI2b5e785b7310_379,RI2b5e785b5ba0_399,RI2b5e785b5240_419,RI2b5e785b48e0_439,RI2b5e785b3530_459,RI2b5e785b2bd0_479,
        RI2b5e785b2270_499,RI2b5e785b1280_519,RI2b5e785b0920_539,RI2b5e785affc0_559,RI2b5e785af390_579,RI2b5e785c0988_258,RI2b5e785be318_278,RI2b5e785bc068_298,RI2b5e785ba178_318,RI2b5e785b9818_338,
        RI2b5e785b7ce8_358,RI2b5e785b7388_378,RI2b5e785b5c18_398,RI2b5e785b52b8_418,RI2b5e785b4958_438,RI2b5e785b35a8_458,RI2b5e785b2c48_478,RI2b5e785b22e8_498,RI2b5e785b12f8_518,RI2b5e785b0998_538,
        RI2b5e785b0038_558,RI2b5e785af408_578,RI2b5e785c0820_261,RI2b5e785be1b0_281,RI2b5e785bbf00_301,RI2b5e785ba010_321,RI2b5e785b96b0_341,RI2b5e785b7b80_361,RI2b5e785b7220_381,RI2b5e785b5ab0_401,
        RI2b5e785b5150_421,RI2b5e785b47f0_441,RI2b5e785b3440_461,RI2b5e785b2ae0_481,RI2b5e785b2180_501,RI2b5e785b1190_521,RI2b5e785b0830_541,RI2b5e785afed0_561,RI2b5e785af2a0_581,RI2b5e785c0898_260,
        RI2b5e785be228_280,RI2b5e785bbf78_300,RI2b5e785ba088_320,RI2b5e785b9728_340,RI2b5e785b7bf8_360,RI2b5e785b7298_380,RI2b5e785b5b28_400,RI2b5e785b51c8_420,RI2b5e785b4868_440,RI2b5e785b34b8_460,
        RI2b5e785b2b58_480,RI2b5e785b21f8_500,RI2b5e785b1208_520,RI2b5e785b08a8_540,RI2b5e785aff48_560,RI2b5e785af318_580,RI2b5e785c0730_263,RI2b5e785be0c0_283,RI2b5e785bbe10_303,RI2b5e785b9f20_323,
        RI2b5e785b95c0_343,RI2b5e785b7a90_363,RI2b5e785b7130_383,RI2b5e785b59c0_403,RI2b5e785b5060_423,RI2b5e785b3cb0_443,RI2b5e785b3350_463,RI2b5e785b29f0_483,RI2b5e785b1a00_503,RI2b5e785b10a0_523,
        RI2b5e785b0740_543,RI2b5e785afde0_563,RI2b5e785af1b0_583,RI2b5e785c07a8_262,RI2b5e785be138_282,RI2b5e785bbe88_302,RI2b5e785b9f98_322,RI2b5e785b9638_342,RI2b5e785b7b08_362,RI2b5e785b71a8_382,
        RI2b5e785b5a38_402,RI2b5e785b50d8_422,RI2b5e785b4778_442,RI2b5e785b33c8_462,RI2b5e785b2a68_482,RI2b5e785b1a78_502,RI2b5e785b1118_522,RI2b5e785b07b8_542,RI2b5e785afe58_562,RI2b5e785af228_582,
        RI2b5e785c0640_265,RI2b5e785bdfd0_285,RI2b5e785bbd20_305,RI2b5e785b9e30_325,RI2b5e785b94d0_345,RI2b5e785b79a0_365,RI2b5e785b7040_385,RI2b5e785b58d0_405,RI2b5e785b4f70_425,RI2b5e785b3bc0_445,
        RI2b5e785b3260_465,RI2b5e785b2900_485,RI2b5e785b1910_505,RI2b5e785b0fb0_525,RI2b5e785b0650_545,RI2b5e785afcf0_565,RI2b5e785af0c0_585,RI2b5e785c06b8_264,RI2b5e785be048_284,RI2b5e785bbd98_304,
        RI2b5e785b9ea8_324,RI2b5e785b9548_344,RI2b5e785b7a18_364,RI2b5e785b70b8_384,RI2b5e785b5948_404,RI2b5e785b4fe8_424,RI2b5e785b3c38_444,RI2b5e785b32d8_464,RI2b5e785b2978_484,RI2b5e785b1988_504,
        RI2b5e785b1028_524,RI2b5e785b06c8_544,RI2b5e785afd68_564,RI2b5e785af138_584,RI2b5e785c05c8_266,RI2b5e785bdf58_286,RI2b5e785bbca8_306,RI2b5e785b9db8_326,RI2b5e785b9458_346,RI2b5e785b7928_366,
        RI2b5e785b6fc8_386,RI2b5e785b5858_406,RI2b5e785b4ef8_426,RI2b5e785b3b48_446,RI2b5e785b31e8_466,RI2b5e785b2888_486,RI2b5e785b1898_506,RI2b5e785b0f38_526,RI2b5e785b05d8_546,RI2b5e785afc78_566,
        RI2b5e785af048_586,RI2b5e785c0550_267,RI2b5e785bc590_287,RI2b5e785bbc30_307,RI2b5e785b9d40_327,RI2b5e785b93e0_347,RI2b5e785b78b0_367,RI2b5e785b6f50_387,RI2b5e785b57e0_407,RI2b5e785b4e80_427,
        RI2b5e785b3ad0_447,RI2b5e785b3170_467,RI2b5e785b2810_487,RI2b5e785b1820_507,RI2b5e785b0ec0_527,RI2b5e785b0560_547,RI2b5e785afc00_567,RI2b5e785aefd0_587,RI2b5e785ae328_614,RI2b5e785db058_15,
        RI2b5e785dafe0_16,RI2b5e785daf68_17,RI2b5e785daef0_18,RI2b5e785dae78_19,RI2b5e785dae00_20,RI2b5e785dad88_21,RI2b5e785dad10_22,RI2b5e785dac98_23,RI2b5e785dac20_24,RI2b5e785daba8_25,
        RI2b5e785ae3a0_613,RI2b5e785ae418_612,RI2b5e785ae490_611,RI2b5e785ae508_610,RI2b5e785ae580_609,RI2b5e785ae5f8_608,RI2b5e785ae670_607,RI2b5e785ae6e8_606,RI2b5e785ae760_605,RI2b5e785ae7d8_604,
        RI2b5e785ae850_603,RI2b5e785ae8c8_602,RI2b5e785ae940_601,RI2b5e785dab30_26,RI2b5e785db0d0_14,R_267_b04ddc8,R_268_b04de70,R_269_b04df18,R_26a_b04dfc0,R_26b_b04e068,
        R_26c_b04e110,R_26d_b04e1b8,R_26e_b04e260,R_26f_b04e308,R_270_b04e3b0,R_271_b04e458,R_272_b04e500,R_273_b04e5a8,R_274_b04e650,R_275_b04e6f8,
        R_276_b04e7a0,R_277_b04e848,R_278_b04e8f0,R_279_b04e998,R_27a_b04ea40,R_27b_b04eae8,R_27c_b04eb90,R_27d_b04ec38,R_27e_b04ece0,R_27f_b04ed88,
        R_280_b04ee30,R_281_b04eed8,R_282_b04ef80,R_283_b04f028,R_284_b04f0d0,R_285_b04f178,R_286_b04f220,R_287_b04f2c8,R_288_b04f370,R_289_b04f418,
        R_28a_b04f4c0,R_28b_b04f568,R_28c_b04f610,R_28d_b04f6b8,R_28e_b04f760,R_28f_b04f808,R_290_b04f8b0,R_291_b04f958,R_292_b04fa00,R_293_b04faa8,
        R_294_b04fb50,R_295_b04fbf8,R_296_b04fca0,R_297_b04fd48,R_298_b04fdf0,R_299_b04fe98,R_29a_b04ff40,R_29b_b04ffe8,R_29c_b050090,R_29d_b050138,
        R_29e_b0501e0,R_29f_b050288,R_2a0_b050330,R_2a1_b0503d8,R_2a2_b050480,R_2a3_b050528,R_2a4_b0505d0,R_2a5_b050678,R_2a6_b050720,R_2a7_b0507c8,
        R_2a8_b050870,R_2a9_b050918,R_2aa_b0509c0);
input RI2b5e785ebcf0_2,RI2b5e785ebc78_3,RI2b5e785ebc00_4,RI2b5e785ebb88_5,RI2b5e785ebb10_6,RI2b5e785eba98_7,RI2b5e785eba20_8,RI2b5e785eb9a8_9,RI2b5e785eb930_10,
        RI2b5e785eb8b8_11,RI2b5e785eb840_12,RI2b5e785daa40_28,RI2b5e785ae9b8_600,RI2b5e785aea30_599,RI2b5e785aeaa8_598,RI2b5e785aeb20_597,RI2b5e785aeb98_596,RI2b5e785aec10_595,RI2b5e785aec88_594,
        RI2b5e785aed00_593,RI2b5e785aed78_592,RI2b5e785aedf0_591,RI2b5e785aee68_590,RI2b5e785aeee0_589,RI2b5e785aef58_588,RI2b5e78549540_41,RI2b5e785388a8_54,RI2b5e784a6330_67,RI2b5e78495698_80,
        RI2b5e78495080_93,RI2b5e78403b80_106,RI2b5e775b1e60_119,RI2b5e7750bdf8_132,RI2b5e774ff5d0_145,RI2b5e774f65e8_158,RI2b5e774eabd0_171,RI2b5e774de3a8_184,RI2b5e774d53c0_197,RI2b5e785f4300_210,
        RI2b5e785f3ce8_223,RI2b5e785eb0c0_236,RI2b5e785da9c8_29,RI2b5e785494c8_42,RI2b5e78538830_55,RI2b5e784a62b8_68,RI2b5e78495620_81,RI2b5e78495008_94,RI2b5e78403b08_107,RI2b5e775b1de8_120,
        RI2b5e7750bd80_133,RI2b5e774ff558_146,RI2b5e774f6570_159,RI2b5e774eab58_172,RI2b5e774de330_185,RI2b5e774d5348_198,RI2b5e785f4288_211,RI2b5e785f3658_224,RI2b5e785eb048_237,RI2b5e785da950_30,
        RI2b5e78549450_43,RI2b5e785387b8_56,RI2b5e784a6240_69,RI2b5e784955a8_82,RI2b5e78494f90_95,RI2b5e78403a90_108,RI2b5e775b1d70_121,RI2b5e7750bd08_134,RI2b5e774ff4e0_147,RI2b5e774f64f8_160,
        RI2b5e774eaae0_173,RI2b5e774de2b8_186,RI2b5e774d52d0_199,RI2b5e785f4210_212,RI2b5e785eb5e8_225,RI2b5e785e6c50_238,RI2b5e785da8d8_31,RI2b5e785493d8_44,RI2b5e78538740_57,RI2b5e784a61c8_70,
        RI2b5e78495530_83,RI2b5e78494f18_96,RI2b5e78403a18_109,RI2b5e775b1cf8_122,RI2b5e7750bc90_135,RI2b5e774ff468_148,RI2b5e774f6480_161,RI2b5e774eaa68_174,RI2b5e774de240_187,RI2b5e774d5258_200,
        RI2b5e785f4198_213,RI2b5e785eb570_226,RI2b5e785e6bd8_239,RI2b5e785da860_32,RI2b5e78549360_45,RI2b5e785386c8_58,RI2b5e784a6150_71,RI2b5e784954b8_84,RI2b5e78494ea0_97,RI2b5e784039a0_110,
        RI2b5e775b1c80_123,RI2b5e7750bc18_136,RI2b5e774ff3f0_149,RI2b5e774f6408_162,RI2b5e774ea9f0_175,RI2b5e774de1c8_188,RI2b5e774d51e0_201,RI2b5e785f4120_214,RI2b5e785eb4f8_227,RI2b5e785e64d0_240,
        RI2b5e78549900_33,RI2b5e78538c68_46,RI2b5e78538650_59,RI2b5e784a60d8_72,RI2b5e78495440_85,RI2b5e78494e28_98,RI2b5e78403928_111,RI2b5e775b1c08_124,RI2b5e7750bba0_137,RI2b5e774ff378_150,
        RI2b5e774f6390_163,RI2b5e774ea978_176,RI2b5e774de150_189,RI2b5e774d5168_202,RI2b5e785f40a8_215,RI2b5e785eb480_228,RI2b5e785da608_241,RI2b5e78549888_34,RI2b5e78538bf0_47,RI2b5e785385d8_60,
        RI2b5e784a6060_73,RI2b5e784953c8_86,RI2b5e78403ec8_99,RI2b5e775b21a8_112,RI2b5e775b1b90_125,RI2b5e7750bb28_138,RI2b5e774ff300_151,RI2b5e774f6318_164,RI2b5e774ea900_177,RI2b5e774de0d8_190,
        RI2b5e774d50f0_203,RI2b5e785f4030_216,RI2b5e785eb408_229,RI2b5e785da590_242,RI2b5e78549810_35,RI2b5e78538b78_48,RI2b5e78538560_61,RI2b5e784a5fe8_74,RI2b5e78495350_87,RI2b5e78403e50_100,
        RI2b5e775b2130_113,RI2b5e775b1b18_126,RI2b5e7750bab0_139,RI2b5e774ff288_152,RI2b5e774f62a0_165,RI2b5e774ea888_178,RI2b5e774de060_191,RI2b5e774d5078_204,RI2b5e785f3fb8_217,RI2b5e785eb390_230,
        RI2b5e785da518_243,RI2b5e78549798_36,RI2b5e78538b00_49,RI2b5e785384e8_62,RI2b5e784a5f70_75,RI2b5e784952d8_88,RI2b5e78403dd8_101,RI2b5e775b20b8_114,RI2b5e775b1aa0_127,RI2b5e7750ba38_140,
        RI2b5e774ff210_153,RI2b5e774f6228_166,RI2b5e774ea810_179,RI2b5e774ddfe8_192,RI2b5e774d5000_205,RI2b5e785f3f40_218,RI2b5e785eb318_231,RI2b5e785da4a0_244,RI2b5e78549720_37,RI2b5e78538a88_50,
        RI2b5e78538470_63,RI2b5e784a5ef8_76,RI2b5e78495260_89,RI2b5e78403d60_102,RI2b5e775b2040_115,RI2b5e775b1a28_128,RI2b5e7750b9c0_141,RI2b5e774ff198_154,RI2b5e774f61b0_167,RI2b5e774ea798_180,
        RI2b5e774ddf70_193,RI2b5e774d4f88_206,RI2b5e785f3ec8_219,RI2b5e785eb2a0_232,RI2b5e785da428_245,RI2b5e785496a8_38,RI2b5e78538a10_51,RI2b5e785383f8_64,RI2b5e784a5e80_77,RI2b5e784951e8_90,
        RI2b5e78403ce8_103,RI2b5e775b1fc8_116,RI2b5e775b19b0_129,RI2b5e7750b948_142,RI2b5e774ff120_155,RI2b5e774f6138_168,RI2b5e774ea720_181,RI2b5e774ddef8_194,RI2b5e774d4f10_207,RI2b5e785f3e50_220,
        RI2b5e785eb228_233,RI2b5e785da3b0_246,RI2b5e785db148_13,RI2b5e78549630_39,RI2b5e78538998_52,RI2b5e78538380_65,RI2b5e784a5e08_78,RI2b5e78495170_91,RI2b5e78403c70_104,RI2b5e775b1f50_117,
        RI2b5e775b1938_130,RI2b5e7750b8d0_143,RI2b5e774ff0a8_156,RI2b5e774f60c0_169,RI2b5e774ea6a8_182,RI2b5e774dde80_195,RI2b5e774d4e98_208,RI2b5e785f3dd8_221,RI2b5e785eb1b0_234,RI2b5e785da338_247,
        RI2b5e785da248_249,RI2b5e785be750_269,RI2b5e785bc4a0_289,RI2b5e785bbb40_309,RI2b5e785b9c50_329,RI2b5e785b8120_349,RI2b5e785b77c0_369,RI2b5e785b6e60_389,RI2b5e785b56f0_409,RI2b5e785b4d90_429,
        RI2b5e785b39e0_449,RI2b5e785b3080_469,RI2b5e785b2720_489,RI2b5e785b1730_509,RI2b5e785b0dd0_529,RI2b5e785b0470_549,RI2b5e785af840_569,RI2b5e785ebd68_1,RI2b5e785daab8_27,RI2b5e785495b8_40,
        RI2b5e78538920_53,RI2b5e784a63a8_66,RI2b5e78495710_79,RI2b5e784950f8_92,RI2b5e78403bf8_105,RI2b5e775b1ed8_118,RI2b5e775b18c0_131,RI2b5e7750b858_144,RI2b5e774ff030_157,RI2b5e774f6048_170,
        RI2b5e774ea630_183,RI2b5e774dde08_196,RI2b5e774d4e20_209,RI2b5e785f3d60_222,RI2b5e785eb138_235,RI2b5e785da2c0_248,RI2b5e785be7c8_268,RI2b5e785bc518_288,RI2b5e785bbbb8_308,RI2b5e785b9cc8_328,
        RI2b5e785b9368_348,RI2b5e785b7838_368,RI2b5e785b6ed8_388,RI2b5e785b5768_408,RI2b5e785b4e08_428,RI2b5e785b3a58_448,RI2b5e785b30f8_468,RI2b5e785b2798_488,RI2b5e785b17a8_508,RI2b5e785b0e48_528,
        RI2b5e785b04e8_548,RI2b5e785afb88_568,RI2b5e785da1d0_250,RI2b5e785be6d8_270,RI2b5e785bc428_290,RI2b5e785bbac8_310,RI2b5e785b9bd8_330,RI2b5e785b80a8_350,RI2b5e785b7748_370,RI2b5e785b6de8_390,
        RI2b5e785b5678_410,RI2b5e785b4d18_430,RI2b5e785b3968_450,RI2b5e785b3008_470,RI2b5e785b26a8_490,RI2b5e785b16b8_510,RI2b5e785b0d58_530,RI2b5e785b03f8_550,RI2b5e785af7c8_570,RI2b5e785da0e0_252,
        RI2b5e785be5e8_272,RI2b5e785bc338_292,RI2b5e785bb9d8_312,RI2b5e785b9ae8_332,RI2b5e785b7fb8_352,RI2b5e785b7658_372,RI2b5e785b5ee8_392,RI2b5e785b5588_412,RI2b5e785b4c28_432,RI2b5e785b3878_452,
        RI2b5e785b2f18_472,RI2b5e785b25b8_492,RI2b5e785b15c8_512,RI2b5e785b0c68_532,RI2b5e785b0308_552,RI2b5e785af6d8_572,RI2b5e785da158_251,RI2b5e785be660_271,RI2b5e785bc3b0_291,RI2b5e785bba50_311,
        RI2b5e785b9b60_331,RI2b5e785b8030_351,RI2b5e785b76d0_371,RI2b5e785b6d70_391,RI2b5e785b5600_411,RI2b5e785b4ca0_431,RI2b5e785b38f0_451,RI2b5e785b2f90_471,RI2b5e785b2630_491,RI2b5e785b1640_511,
        RI2b5e785b0ce0_531,RI2b5e785b0380_551,RI2b5e785af750_571,RI2b5e785da068_253,RI2b5e785be570_273,RI2b5e785bc2c0_293,RI2b5e785bb960_313,RI2b5e785b9a70_333,RI2b5e785b7f40_353,RI2b5e785b75e0_373,
        RI2b5e785b5e70_393,RI2b5e785b5510_413,RI2b5e785b4bb0_433,RI2b5e785b3800_453,RI2b5e785b2ea0_473,RI2b5e785b2540_493,RI2b5e785b1550_513,RI2b5e785b0bf0_533,RI2b5e785b0290_553,RI2b5e785af660_573,
        RI2b5e785c2bc0_255,RI2b5e785be480_275,RI2b5e785bc1d0_295,RI2b5e785ba2e0_315,RI2b5e785b9980_335,RI2b5e785b7e50_355,RI2b5e785b74f0_375,RI2b5e785b5d80_395,RI2b5e785b5420_415,RI2b5e785b4ac0_435,
        RI2b5e785b3710_455,RI2b5e785b2db0_475,RI2b5e785b2450_495,RI2b5e785b1460_515,RI2b5e785b0b00_535,RI2b5e785b01a0_555,RI2b5e785af570_575,RI2b5e785c2c38_254,RI2b5e785be4f8_274,RI2b5e785bc248_294,
        RI2b5e785ba358_314,RI2b5e785b99f8_334,RI2b5e785b7ec8_354,RI2b5e785b7568_374,RI2b5e785b5df8_394,RI2b5e785b5498_414,RI2b5e785b4b38_434,RI2b5e785b3788_454,RI2b5e785b2e28_474,RI2b5e785b24c8_494,
        RI2b5e785b14d8_514,RI2b5e785b0b78_534,RI2b5e785b0218_554,RI2b5e785af5e8_574,RI2b5e785c0a00_257,RI2b5e785be390_277,RI2b5e785bc0e0_297,RI2b5e785ba1f0_317,RI2b5e785b9890_337,RI2b5e785b7d60_357,
        RI2b5e785b7400_377,RI2b5e785b5c90_397,RI2b5e785b5330_417,RI2b5e785b49d0_437,RI2b5e785b3620_457,RI2b5e785b2cc0_477,RI2b5e785b2360_497,RI2b5e785b1370_517,RI2b5e785b0a10_537,RI2b5e785b00b0_557,
        RI2b5e785af480_577,RI2b5e785c2b48_256,RI2b5e785be408_276,RI2b5e785bc158_296,RI2b5e785ba268_316,RI2b5e785b9908_336,RI2b5e785b7dd8_356,RI2b5e785b7478_376,RI2b5e785b5d08_396,RI2b5e785b53a8_416,
        RI2b5e785b4a48_436,RI2b5e785b3698_456,RI2b5e785b2d38_476,RI2b5e785b23d8_496,RI2b5e785b13e8_516,RI2b5e785b0a88_536,RI2b5e785b0128_556,RI2b5e785af4f8_576,RI2b5e785c0910_259,RI2b5e785be2a0_279,
        RI2b5e785bbff0_299,RI2b5e785ba100_319,RI2b5e785b97a0_339,RI2b5e785b7c70_359,RI2b5e785b7310_379,RI2b5e785b5ba0_399,RI2b5e785b5240_419,RI2b5e785b48e0_439,RI2b5e785b3530_459,RI2b5e785b2bd0_479,
        RI2b5e785b2270_499,RI2b5e785b1280_519,RI2b5e785b0920_539,RI2b5e785affc0_559,RI2b5e785af390_579,RI2b5e785c0988_258,RI2b5e785be318_278,RI2b5e785bc068_298,RI2b5e785ba178_318,RI2b5e785b9818_338,
        RI2b5e785b7ce8_358,RI2b5e785b7388_378,RI2b5e785b5c18_398,RI2b5e785b52b8_418,RI2b5e785b4958_438,RI2b5e785b35a8_458,RI2b5e785b2c48_478,RI2b5e785b22e8_498,RI2b5e785b12f8_518,RI2b5e785b0998_538,
        RI2b5e785b0038_558,RI2b5e785af408_578,RI2b5e785c0820_261,RI2b5e785be1b0_281,RI2b5e785bbf00_301,RI2b5e785ba010_321,RI2b5e785b96b0_341,RI2b5e785b7b80_361,RI2b5e785b7220_381,RI2b5e785b5ab0_401,
        RI2b5e785b5150_421,RI2b5e785b47f0_441,RI2b5e785b3440_461,RI2b5e785b2ae0_481,RI2b5e785b2180_501,RI2b5e785b1190_521,RI2b5e785b0830_541,RI2b5e785afed0_561,RI2b5e785af2a0_581,RI2b5e785c0898_260,
        RI2b5e785be228_280,RI2b5e785bbf78_300,RI2b5e785ba088_320,RI2b5e785b9728_340,RI2b5e785b7bf8_360,RI2b5e785b7298_380,RI2b5e785b5b28_400,RI2b5e785b51c8_420,RI2b5e785b4868_440,RI2b5e785b34b8_460,
        RI2b5e785b2b58_480,RI2b5e785b21f8_500,RI2b5e785b1208_520,RI2b5e785b08a8_540,RI2b5e785aff48_560,RI2b5e785af318_580,RI2b5e785c0730_263,RI2b5e785be0c0_283,RI2b5e785bbe10_303,RI2b5e785b9f20_323,
        RI2b5e785b95c0_343,RI2b5e785b7a90_363,RI2b5e785b7130_383,RI2b5e785b59c0_403,RI2b5e785b5060_423,RI2b5e785b3cb0_443,RI2b5e785b3350_463,RI2b5e785b29f0_483,RI2b5e785b1a00_503,RI2b5e785b10a0_523,
        RI2b5e785b0740_543,RI2b5e785afde0_563,RI2b5e785af1b0_583,RI2b5e785c07a8_262,RI2b5e785be138_282,RI2b5e785bbe88_302,RI2b5e785b9f98_322,RI2b5e785b9638_342,RI2b5e785b7b08_362,RI2b5e785b71a8_382,
        RI2b5e785b5a38_402,RI2b5e785b50d8_422,RI2b5e785b4778_442,RI2b5e785b33c8_462,RI2b5e785b2a68_482,RI2b5e785b1a78_502,RI2b5e785b1118_522,RI2b5e785b07b8_542,RI2b5e785afe58_562,RI2b5e785af228_582,
        RI2b5e785c0640_265,RI2b5e785bdfd0_285,RI2b5e785bbd20_305,RI2b5e785b9e30_325,RI2b5e785b94d0_345,RI2b5e785b79a0_365,RI2b5e785b7040_385,RI2b5e785b58d0_405,RI2b5e785b4f70_425,RI2b5e785b3bc0_445,
        RI2b5e785b3260_465,RI2b5e785b2900_485,RI2b5e785b1910_505,RI2b5e785b0fb0_525,RI2b5e785b0650_545,RI2b5e785afcf0_565,RI2b5e785af0c0_585,RI2b5e785c06b8_264,RI2b5e785be048_284,RI2b5e785bbd98_304,
        RI2b5e785b9ea8_324,RI2b5e785b9548_344,RI2b5e785b7a18_364,RI2b5e785b70b8_384,RI2b5e785b5948_404,RI2b5e785b4fe8_424,RI2b5e785b3c38_444,RI2b5e785b32d8_464,RI2b5e785b2978_484,RI2b5e785b1988_504,
        RI2b5e785b1028_524,RI2b5e785b06c8_544,RI2b5e785afd68_564,RI2b5e785af138_584,RI2b5e785c05c8_266,RI2b5e785bdf58_286,RI2b5e785bbca8_306,RI2b5e785b9db8_326,RI2b5e785b9458_346,RI2b5e785b7928_366,
        RI2b5e785b6fc8_386,RI2b5e785b5858_406,RI2b5e785b4ef8_426,RI2b5e785b3b48_446,RI2b5e785b31e8_466,RI2b5e785b2888_486,RI2b5e785b1898_506,RI2b5e785b0f38_526,RI2b5e785b05d8_546,RI2b5e785afc78_566,
        RI2b5e785af048_586,RI2b5e785c0550_267,RI2b5e785bc590_287,RI2b5e785bbc30_307,RI2b5e785b9d40_327,RI2b5e785b93e0_347,RI2b5e785b78b0_367,RI2b5e785b6f50_387,RI2b5e785b57e0_407,RI2b5e785b4e80_427,
        RI2b5e785b3ad0_447,RI2b5e785b3170_467,RI2b5e785b2810_487,RI2b5e785b1820_507,RI2b5e785b0ec0_527,RI2b5e785b0560_547,RI2b5e785afc00_567,RI2b5e785aefd0_587,RI2b5e785ae328_614,RI2b5e785db058_15,
        RI2b5e785dafe0_16,RI2b5e785daf68_17,RI2b5e785daef0_18,RI2b5e785dae78_19,RI2b5e785dae00_20,RI2b5e785dad88_21,RI2b5e785dad10_22,RI2b5e785dac98_23,RI2b5e785dac20_24,RI2b5e785daba8_25,
        RI2b5e785ae3a0_613,RI2b5e785ae418_612,RI2b5e785ae490_611,RI2b5e785ae508_610,RI2b5e785ae580_609,RI2b5e785ae5f8_608,RI2b5e785ae670_607,RI2b5e785ae6e8_606,RI2b5e785ae760_605,RI2b5e785ae7d8_604,
        RI2b5e785ae850_603,RI2b5e785ae8c8_602,RI2b5e785ae940_601,RI2b5e785dab30_26,RI2b5e785db0d0_14;
output R_267_b04ddc8,R_268_b04de70,R_269_b04df18,R_26a_b04dfc0,R_26b_b04e068,R_26c_b04e110,R_26d_b04e1b8,R_26e_b04e260,R_26f_b04e308,
        R_270_b04e3b0,R_271_b04e458,R_272_b04e500,R_273_b04e5a8,R_274_b04e650,R_275_b04e6f8,R_276_b04e7a0,R_277_b04e848,R_278_b04e8f0,R_279_b04e998,
        R_27a_b04ea40,R_27b_b04eae8,R_27c_b04eb90,R_27d_b04ec38,R_27e_b04ece0,R_27f_b04ed88,R_280_b04ee30,R_281_b04eed8,R_282_b04ef80,R_283_b04f028,
        R_284_b04f0d0,R_285_b04f178,R_286_b04f220,R_287_b04f2c8,R_288_b04f370,R_289_b04f418,R_28a_b04f4c0,R_28b_b04f568,R_28c_b04f610,R_28d_b04f6b8,
        R_28e_b04f760,R_28f_b04f808,R_290_b04f8b0,R_291_b04f958,R_292_b04fa00,R_293_b04faa8,R_294_b04fb50,R_295_b04fbf8,R_296_b04fca0,R_297_b04fd48,
        R_298_b04fdf0,R_299_b04fe98,R_29a_b04ff40,R_29b_b04ffe8,R_29c_b050090,R_29d_b050138,R_29e_b0501e0,R_29f_b050288,R_2a0_b050330,R_2a1_b0503d8,
        R_2a2_b050480,R_2a3_b050528,R_2a4_b0505d0,R_2a5_b050678,R_2a6_b050720,R_2a7_b0507c8,R_2a8_b050870,R_2a9_b050918,R_2aa_b0509c0;

wire \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 ,
         \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 ,
         \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 ,
         \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 ,
         \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 ,
         \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 ,
         \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 ,
         \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 ,
         \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 ,
         \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 ,
         \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 ,
         \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 ,
         \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 ,
         \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 ,
         \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 ,
         \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 ,
         \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 ,
         \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 ,
         \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 ,
         \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 ,
         \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 ,
         \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 ,
         \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 ,
         \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 ,
         \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 ,
         \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 ,
         \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 ,
         \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 ,
         \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 ,
         \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 ,
         \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 ,
         \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 ,
         \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 ,
         \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 ,
         \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 ,
         \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 ,
         \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 ,
         \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 ,
         \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 ,
         \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 ,
         \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 ,
         \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 ,
         \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 ,
         \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 ,
         \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 ,
         \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 ,
         \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 ,
         \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 ,
         \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 ,
         \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 ,
         \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 ,
         \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 ,
         \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 ,
         \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 ,
         \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 ,
         \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 ,
         \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 ,
         \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 ,
         \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 ,
         \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 ,
         \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 ,
         \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 ,
         \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 ,
         \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 ,
         \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 ,
         \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
         \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 ,
         \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 ,
         \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 ,
         \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 ,
         \1382 , \1383 , \1384 , \1385 , \1386 , \1387_N$1 , \1388_N$2 , \1389_N$3 , \1390_N$4 , \1391_N$5 ,
         \1392_N$6 , \1393_N$7 , \1394_N$8 , \1395_N$9 , \1396_N$10 , \1397_N$11 , \1398_N$12 , \1399_N$13 , \1400_N$14 , \1401_N$15 ,
         \1402_N$16 , \1403_N$17 , \1404_N$18 , \1405_N$20 , \1406_N$21 , \1407_N$22 , \1408_N$23 , \1409_N$24 , \1410_N$25 , \1411_N$26 ,
         \1412_N$27 , \1413_N$28 , \1414_N$29 , \1415_N$30 , \1416_N$31 , \1417_N$32 , \1418_N$33 , \1419_N$34 , \1420_N$35 , \1421_N$36 ,
         \1422_N$37 , \1423_N$38 , \1424_N$39 , \1425_N$40 , \1426_N$41 , \1427_N$42 , \1428_N$43 , \1429_N$45 , \1430_N$46 , \1431_N$47 ,
         \1432_N$48 , \1433_N$49 , \1434_N$50 , \1435_N$51 , \1436_N$52 , \1437_N$53 , \1438_N$54 , \1439_N$55 , \1440_N$56 , \1441_N$57 ,
         \1442_N$58 , \1443_N$59 , \1444_N$60 , \1445_N$61 , \1446_N$62 , \1447_N$63 , \1448_N$64 , \1449_N$65 , \1450_N$66 , \1451_N$67 ,
         \1452_N$68 , \1453_N$69 , \1454_N$70 , \1455_N$71 , \1456_N$72 , \1457_N$73 , \1458_N$74 , \1459_N$75 , \1460_N$76 , \1461_N$77 ,
         \1462_N$78 , \1463_N$79 , \1464_N$80 , \1465_N$81 , \1466_N$82 , \1467_N$83 , \1468_N$85 , \1469_N$86 , \1470_N$87 , \1471_N$88 ,
         \1472_N$90 , \1473_N$91 , \1474_N$92 , \1475_N$93 , \1476_N$94 , \1477_N$95 , \1478_N$96 , \1479_N$98 , \1480_N$99 , \1481_N$100 ,
         \1482_N$101 , \1483_N$102 , \1484_N$103 , \1485_N$104 , \1486_N$105 , \1487_N$106 , \1488_N$107 , \1489_N$108 , \1490_N$109 , \1491_N$110 ,
         \1492_N$111 , \1493_N$112 , \1494_N$113 , \1495_N$114 , \1496_N$115 , \1497_N$116 , \1498_N$117 , \1499_N$118 , \1500_N$119 , \1501_N$120 ,
         \1502_N$121 , \1503_N$122 , \1504_N$123 , \1505_N$124 , \1506_N$125 , \1507_N$126 , \1508_N$127 , \1509_N$128 , \1510_N$129 , \1511_N$130 ,
         \1512_N$131 , \1513_N$132 , \1514_N$133 , \1515_N$134 , \1516_N$135 , \1517_N$137 , \1518_N$138 , \1519_N$139 , \1520_N$140 , \1521_N$141 ,
         \1522_N$142 , \1523_N$143 , \1524_N$144 , \1525_N$145 , \1526_N$146 , \1527_N$147 , \1528_N$148 , \1529_N$149 , \1530_N$150 , \1531_N$151 ,
         \1532_N$152 , \1533_N$153 , \1534_N$154 , \1535_N$155 , \1536_N$156 , \1537_N$157 , \1538_N$158 , \1539_N$159 , \1540_N$160 , \1541_N$161 ,
         \1542_N$162 , \1543_N$163 , \1544_N$164 , \1545_N$165 , \1546_N$166 , \1547_N$167 , \1548_N$168 , \1549_N$169 , \1550_N$171 , \1551_N$172 ,
         \1552_N$173 , \1553_N$174 , \1554_N$175 , \1555_N$176 , \1556_N$177 , \1557_N$178 , \1558_N$179 , \1559_N$180 , \1560_N$181 , \1561_N$182 ,
         \1562_N$183 , \1563_N$184 , \1564_N$185 , \1565_N$186 , \1566_N$187 , \1567_N$188 , \1568_N$189 , \1569_N$190 , \1570_N$191 , \1571_N$192 ,
         \1572_N$193 , \1573_N$194 , \1574_N$195 , \1575_N$196 , \1576_N$197 , \1577_N$198 , \1578_N$199 , \1579_N$200 , \1580_N$201 , \1581_N$203 ,
         \1582_N$204 , \1583_N$205 , \1584_N$206 , \1585_N$207 , \1586_N$208 , \1587_N$209 , \1588_N$210 , \1589_N$211 , \1590_N$212 , \1591_N$213 ,
         \1592_N$214 , \1593_N$215 , \1594_N$216 , \1595_N$217 , \1596_N$218 , \1597_N$219 , \1598_N$220 , \1599_N$221 , \1600_N$222 , \1601_N$223 ,
         \1602_N$224 , \1603_N$225 , \1604_N$226 , \1605_N$228 , \1606_N$229 , \1607_N$230 , \1608_N$231 , \1609_N$232 , \1610_N$233 , \1611_N$234 ,
         \1612_N$235 , \1613_N$236 , \1614_N$237 , \1615_N$238 , \1616_N$239 , \1617_N$240 , \1618_N$241 , \1619_N$242 , \1620_N$243 , \1621_N$244 ,
         \1622_N$245 , \1623_N$246 , \1624_N$247 , \1625_N$248 , \1626_N$249 , \1627_N$250 , \1628_N$251 , \1629_N$252 , \1630_N$253 , \1631_N$254 ,
         \1632_N$255 , \1633_N$256 , \1634_N$257 , \1635_N$258 , \1636_N$259 , \1637_N$260 , \1638_N$261 , \1639_N$262 , \1640_N$263 , \1641_N$264 ,
         \1642_N$265 , \1643_N$266 , \1644_N$268 , \1645_N$269 , \1646_N$270 , \1647_N$271 , \1648_N$273 , \1649_N$274 , \1650_N$275 , \1651_N$276 ,
         \1652_N$277 , \1653_N$278 , \1654_N$279 , \1655_N$281 , \1656_N$282 , \1657_N$283 , \1658_N$284 , \1659_N$285 , \1660_N$286 , \1661_N$287 ,
         \1662_N$288 , \1663_N$289 , \1664_N$290 , \1665_N$291 , \1666_N$292 , \1667_N$293 , \1668_N$294 , \1669_N$295 , \1670_N$296 , \1671_N$297 ,
         \1672_N$298 , \1673_N$299 , \1674_N$300 , \1675_N$301 , \1676_N$302 , \1677_N$303 , \1678_N$304 , \1679_N$305 , \1680_N$306 , \1681_N$307 ,
         \1682_N$308 , \1683_N$309 , \1684_N$310 , \1685_N$311 , \1686_N$312 , \1687_N$313 , \1688_N$314 , \1689_N$315 , \1690_N$316 , \1691_N$317 ,
         \1692_N$318 , \1693_N$320 , \1694_N$321 , \1695_N$322 , \1696_N$323 , \1697_N$324 , \1698_N$325 , \1699_N$326 , \1700_N$327 , \1701_N$328 ,
         \1702_N$329 , \1703_N$330 , \1704_N$331 , \1705_N$332 , \1706_N$333 , \1707_N$334 , \1708_N$335 , \1709_N$336 , \1710_N$337 , \1711_N$338 ,
         \1712_N$339 , \1713_N$340 , \1714_N$341 , \1715_N$342 , \1716_N$343 , \1717_N$344 , \1718_N$345 , \1719_N$346 , \1720_N$347 , \1721_N$348 ,
         \1722_N$349 , \1723_N$350 , \1724_N$351 , \1725_N$352 , \1726_N$354 , \1727_N$355 , \1728_N$356 , \1729_N$357 , \1730_N$358 , \1731_N$359 ,
         \1732_N$360 , \1733_N$361 , \1734_N$362 , \1735_N$363 , \1736_N$364 , \1737_N$365 , \1738_N$366 , \1739_N$367 , \1740_N$368 , \1741_N$369 ,
         \1742_N$370 , \1743_N$371 , \1744_N$372 , \1745_N$373 , \1746_N$374 , \1747_N$375 , \1748_N$376 , \1749_N$377 , \1750_N$378 , \1751_N$379 ,
         \1752_N$380 , \1753_N$381 , \1754_N$382 , \1755_N$383 , \1756_N$384 , \1757_N$386 , \1758_N$387 , \1759_N$388 , \1760_N$389 , \1761_N$390 ,
         \1762_N$391 , \1763_N$392 , \1764_N$393 , \1765_N$394 , \1766_N$395 , \1767_N$396 , \1768_N$397 , \1769_N$398 , \1770_N$399 , \1771_N$400 ,
         \1772_N$401 , \1773_N$402 , \1774_N$403 , \1775_N$404 , \1776_N$405 , \1777_N$406 , \1778_N$407 , \1779_N$408 , \1780_N$409 , \1781_N$411 ,
         \1782_N$412 , \1783_N$413 , \1784_N$414 , \1785_N$415 , \1786_N$416 , \1787_N$417 , \1788_N$418 , \1789_N$419 , \1790_N$420 , \1791_N$421 ,
         \1792_N$422 , \1793_N$423 , \1794_N$424 , \1795_N$425 , \1796_N$426 , \1797_N$427 , \1798_N$428 , \1799_N$429 , \1800_N$430 , \1801_N$431 ,
         \1802_N$432 , \1803_N$433 , \1804_N$434 , \1805_N$435 , \1806_N$436 , \1807_N$437 , \1808_N$438 , \1809_N$439 , \1810_N$440 , \1811_N$441 ,
         \1812_N$442 , \1813_N$443 , \1814_N$444 , \1815_N$445 , \1816_N$446 , \1817_N$447 , \1818_N$448 , \1819_N$449 , \1820_N$451 , \1821_N$452 ,
         \1822_N$453 , \1823_N$454 , \1824_N$456 , \1825_N$457 , \1826_N$458 , \1827_N$459 , \1828_N$460 , \1829_N$461 , \1830_N$462 , \1831_N$464 ,
         \1832_N$465 , \1833_N$466 , \1834_N$467 , \1835_N$468 , \1836_N$469 , \1837_N$470 , \1838_N$471 , \1839_N$472 , \1840_N$473 , \1841_N$474 ,
         \1842_N$475 , \1843_N$476 , \1844_N$477 , \1845_N$478 , \1846_N$479 , \1847_N$480 , \1848_N$481 , \1849_N$482 , \1850_N$483 , \1851_N$484 ,
         \1852_N$485 , \1853_N$486 , \1854_N$487 , \1855_N$488 , \1856_N$489 , \1857_N$490 , \1858_N$491 , \1859_N$492 , \1860_N$493 , \1861_N$494 ,
         \1862_N$495 , \1863_N$496 , \1864_N$497 , \1865_N$498 , \1866_N$499 , \1867_N$500 , \1868_N$501 , \1869_N$503 , \1870_N$504 , \1871_N$505 ,
         \1872_N$506 , \1873_N$507 , \1874_N$508 , \1875_N$509 , \1876_N$510 , \1877_N$511 , \1878_N$512 , \1879_N$513 , \1880_N$514 , \1881_N$515 ,
         \1882_N$516 , \1883_N$517 , \1884_N$518 , \1885_N$519 , \1886_N$520 , \1887_N$521 , \1888_N$522 , \1889_N$523 , \1890_N$524 , \1891_N$525 ,
         \1892_N$526 , \1893_N$527 , \1894_N$528 , \1895_N$529 , \1896_N$530 , \1897_N$531 , \1898_N$532 , \1899_N$533 , \1900_N$534 , \1901_N$535 ,
         \1902_N$537 , \1903_N$538 , \1904_N$539 , \1905_N$540 , \1906_N$541 , \1907_N$542 , \1908_N$543 , \1909_N$544 , \1910_N$545 , \1911_N$546 ,
         \1912_N$547 , \1913_N$548 , \1914_N$549 , \1915_N$550 , \1916_N$551 , \1917_N$552 , \1918_N$553 , \1919_N$554 , \1920_N$555 , \1921_N$556 ,
         \1922_N$557 , \1923_N$558 , \1924_N$559 , \1925_N$560 , \1926_N$561 , \1927_N$562 , \1928_N$563 , \1929_N$564 , \1930_N$565 , \1931_N$566 ,
         \1932_N$567 , \1933_N$569 , \1934_N$570 , \1935_N$571 , \1936_N$572 , \1937_N$573 , \1938_N$574 , \1939_N$575 , \1940_N$576 , \1941_N$577 ,
         \1942_N$578 , \1943_N$579 , \1944_N$580 , \1945_N$581 , \1946_N$582 , \1947_N$583 , \1948_N$584 , \1949_N$585 , \1950_N$586 , \1951_N$587 ,
         \1952_N$588 , \1953_N$589 , \1954_N$590 , \1955_N$591 , \1956_N$592 , \1957_N$594 , \1958_N$595 , \1959_N$596 , \1960_N$597 , \1961_N$598 ,
         \1962_N$599 , \1963_N$600 , \1964_N$601 , \1965_N$602 , \1966_N$603 , \1967_N$604 , \1968_N$605 , \1969_N$606 , \1970_N$607 , \1971_N$608 ,
         \1972_N$609 , \1973_N$610 , \1974_N$611 , \1975_N$612 , \1976_N$613 , \1977_N$614 , \1978_N$615 , \1979_N$616 , \1980_N$617 , \1981_N$618 ,
         \1982_N$619 , \1983_N$620 , \1984_N$621 , \1985_N$622 , \1986_N$623 , \1987_N$624 , \1988_N$625 , \1989_N$626 , \1990_N$627 , \1991_N$628 ,
         \1992_N$629 , \1993_N$630 , \1994_N$631 , \1995_N$632 , \1996_N$634 , \1997_N$635 , \1998_N$636 , \1999_N$637 , \2000_N$639 , \2001_N$640 ,
         \2002_N$641 , \2003_N$642 , \2004_N$643 , \2005_N$644 , \2006_N$645 , \2007_N$647 , \2008_N$648 , \2009_N$649 , \2010_N$650 , \2011_N$651 ,
         \2012_N$652 , \2013_N$653 , \2014_N$654 , \2015_N$655 , \2016_N$656 , \2017_N$657 , \2018_N$658 , \2019_N$659 , \2020_N$660 , \2021_N$661 ,
         \2022_N$662 , \2023_N$663 , \2024_N$664 , \2025_N$665 , \2026_N$666 , \2027_N$667 , \2028_N$668 , \2029_N$669 , \2030_N$670 , \2031_N$671 ,
         \2032_N$672 , \2033_N$673 , \2034_N$674 , \2035_N$675 , \2036_N$676 , \2037_N$677 , \2038_N$678 , \2039_N$679 , \2040_N$680 , \2041_N$681 ,
         \2042_N$682 , \2043_N$683 , \2044_N$684 , \2045_N$686 , \2046_N$687 , \2047_N$688 , \2048_N$689 , \2049_N$690 , \2050_N$691 , \2051_N$692 ,
         \2052_N$693 , \2053_N$694 , \2054_N$695 , \2055_N$696 , \2056_N$697 , \2057_N$698 , \2058_N$699 , \2059_N$700 , \2060_N$701 , \2061_N$702 ,
         \2062_N$703 , \2063_N$704 , \2064_N$705 , \2065_N$706 , \2066_N$707 , \2067_N$708 , \2068_N$709 , \2069_N$710 , \2070_N$711 , \2071_N$712 ,
         \2072_N$713 , \2073_N$714 , \2074_N$715 , \2075_N$716 , \2076_N$717 , \2077_N$718 , \2078_N$720 , \2079_N$721 , \2080_N$722 , \2081_N$723 ,
         \2082_N$724 , \2083_N$725 , \2084_N$726 , \2085_N$727 , \2086_N$728 , \2087_N$729 , \2088_N$730 , \2089_N$731 , \2090_N$732 , \2091_ZERO ,
         \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 ,
         \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 ,
         \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120_N$19 , \2121_N$44 ,
         \2122_N$84 , \2123_N$89 , \2124_N$97 , \2125_N$136 , \2126_N$170 , \2127_N$202 , \2128_N$227 , \2129_N$267 , \2130_N$272 , \2131_N$280 ,
         \2132_N$319 , \2133_N$353 , \2134_N$385 , \2135_N$410 , \2136_N$450 , \2137_N$455 , \2138_N$463 , \2139_N$502 , \2140_N$536 , \2141_N$568 ,
         \2142_N$593 , \2143_N$633 , \2144_N$638 , \2145_N$646 , \2146_N$685 , \2147_N$719 , \2148_ONE , \2149 , \2150 , \2151 ,
         \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 ,
         \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 ,
         \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 ,
         \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 ,
         \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 ,
         \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 ,
         \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 ,
         \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229_nG2199 , \2230 , \2231 ,
         \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 ,
         \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 ,
         \2252 , \2253 , \2254_nG2175 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 ,
         \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 ,
         \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279_nG1fee , \2280 , \2281 ,
         \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 ,
         \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 ,
         \2302 , \2303 , \2304_nG1fca , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 ,
         \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 ,
         \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329_nG1e55 , \2330 , \2331 ,
         \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 ,
         \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 ,
         \2352 , \2353 , \2354_nG1e31 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 ,
         \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 ,
         \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379_nG1cf3 , \2380 , \2381 ,
         \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 ,
         \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 ,
         \2402 , \2403 , \2404_nG1ccf , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 ,
         \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 ,
         \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429_nG1bc2 , \2430 , \2431 ,
         \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 ,
         \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 ,
         \2452 , \2453 , \2454_nG1bdb , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 ,
         \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 ,
         \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479_nG1aa5 , \2480 , \2481 ,
         \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 ,
         \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 ,
         \2502 , \2503_nG1a89 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 ,
         \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 ,
         \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 ,
         \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538_nG21a2 , \2539 , \2540 , \2541 ,
         \2542_nG217e , \2543 , \2544 , \2545 , \2546_nG1ff7 , \2547 , \2548 , \2549 , \2550 , \2551 ,
         \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 ,
         \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 ,
         \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 ,
         \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 ,
         \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 ,
         \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 ,
         \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 ,
         \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 ,
         \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 ,
         \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 ,
         \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 ,
         \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 ,
         \2672_nG2899 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 ,
         \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 ,
         \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700_nG2361 , \2701 ,
         \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 ,
         \2712_nG2376 , \2713 , \2714 , \2715 , \2716_nG236a , \2717 , \2718 , \2719 , \2720 , \2721 ,
         \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 ,
         \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741_nG298d ,
         \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 ,
         \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 ,
         \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768_nG27d7 , \2769 , \2770 , \2771 ,
         \2772_nG2572 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 ,
         \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 ,
         \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 ,
         \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 ,
         \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 ,
         \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 ,
         \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839_nG1fd3 , \2840 , \2841 ,
         \2842 , \2843 , \2844_nG1e5e , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 ,
         \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 ,
         \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 ,
         \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879_nG263c , \2880 , \2881 ,
         \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 ,
         \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900_nG2716 , \2901 ,
         \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 ,
         \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 ,
         \2922 , \2923_nG2551 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 ,
         \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 ,
         \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 ,
         \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 ,
         \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 ,
         \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 ,
         \2982 , \2983 , \2984 , \2985 , \2986_nG1aac , \2987 , \2988 , \2989_nG1a8c , \2990 , \2991 ,
         \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 ,
         \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 ,
         \3012 , \3013 , \3014 , \3015 , \3016_nG239e , \3017 , \3018 , \3019 , \3020_nG1be7 , \3021 ,
         \3022 , \3023 , \3024_nG1beb , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 ,
         \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 ,
         \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049_nG2472 , \3050 , \3051 ,
         \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 ,
         \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 ,
         \3072 , \3073 , \3074 , \3075 , \3076_nG21d1 , \3077 , \3078 , \3079 , \3080_nG1cfc , \3081 ,
         \3082 , \3083 , \3084_nG1cd8 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 ,
         \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 ,
         \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109_nG22a8 , \3110 , \3111 ,
         \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 ,
         \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 ,
         \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138_nG2012 , \3139 , \3140 , \3141 ,
         \3142_nG1e3a , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 ,
         \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 ,
         \3162 , \3163 , \3164 , \3165 , \3166 , \3167_nG20db , \3168 , \3169 , \3170 , \3171 ,
         \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 ,
         \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 ,
         \3192 , \3193_nG1e79 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 ,
         \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 ,
         \3212 , \3213 , \3214_nG1f2c , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 ,
         \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 ,
         \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238_nG1d15 , \3239 , \3240 , \3241 ,
         \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 ,
         \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259_nG1dbc , \3260 , \3261 ,
         \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 ,
         \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 ,
         \3282 , \3283 , \3284 , \3285 , \3286_nG1ba5 , \3287 , \3288 , \3289 , \3290 , \3291 ,
         \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 ,
         \3302 , \3303 , \3304 , \3305 , \3306 , \3307_nG1c76 , \3308 , \3309 , \3310 , \3311 ,
         \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 ,
         \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330_nG1b63 , \3331 ,
         \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 ,
         \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 ,
         \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 ,
         \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 ,
         \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 ,
         \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 ,
         \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 ,
         \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 ,
         \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 ,
         \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 ,
         \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 ,
         \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 ,
         \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 ,
         \3462 , \3463_nG1a4f , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 ,
         \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 ,
         \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 ,
         \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 ,
         \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 ,
         \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 ,
         \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 ,
         \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 ,
         \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 ,
         \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 ,
         \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 ,
         \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 ,
         \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 ,
         \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 ,
         \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 ,
         \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 ,
         \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 ,
         \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 ,
         \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 ,
         \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 ,
         \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 ,
         \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 ,
         \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 ,
         \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 ,
         \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 ,
         \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 ,
         \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 ,
         \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 ,
         \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 ,
         \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 ,
         \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 ,
         \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 ,
         \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 ,
         \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 ,
         \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 ,
         \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 ,
         \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 ,
         \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 ,
         \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 ,
         \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 ,
         \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 ,
         \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 ,
         \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 ,
         \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 ,
         \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 ,
         \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 ,
         \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 ,
         \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 ,
         \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 ,
         \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 ,
         \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 ,
         \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 ,
         \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 ,
         \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 ,
         \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 ,
         \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 ,
         \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 ,
         \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 ,
         \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 ,
         \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 ,
         \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 ,
         \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 ,
         \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 ,
         \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 ,
         \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 ,
         \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 ,
         \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 ,
         \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 ,
         \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 ,
         \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 ,
         \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 ,
         \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 ,
         \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 ,
         \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 ,
         \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 ,
         \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 ,
         \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 ,
         \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 ,
         \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 ,
         \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 ,
         \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 ,
         \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 ,
         \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 ,
         \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 ,
         \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 ,
         \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 ,
         \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 ,
         \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 ,
         \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 ,
         \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 ,
         \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 ,
         \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 ,
         \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 ,
         \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 ,
         \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 ,
         \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 ,
         \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 ,
         \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 ,
         \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 ,
         \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 ,
         \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 ,
         \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 ,
         \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 ,
         \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 ,
         \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 ,
         \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 ,
         \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 ,
         \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 ,
         \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 ,
         \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 ,
         \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 ,
         \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 ,
         \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 ,
         \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 ,
         \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 ,
         \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 ,
         \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 ,
         \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 ,
         \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 ,
         \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 ,
         \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 ,
         \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 ,
         \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 ,
         \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 ,
         \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 ,
         \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 ,
         \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 ,
         \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 ,
         \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 ,
         \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 ,
         \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 ,
         \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 ,
         \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 ,
         \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 ,
         \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 ,
         \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 ,
         \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 ,
         \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 ,
         \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 ,
         \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 ,
         \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 ,
         \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 ,
         \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 ,
         \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 ,
         \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 ,
         \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 ,
         \4922 , \4923 , \4924 , \4925 , \4926_nG3284 , \4927 , \4928 , \4929 , \4930 , \4931 ,
         \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 ,
         \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 ,
         \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 ,
         \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 ,
         \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 ,
         \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 ,
         \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 ,
         \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 ,
         \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 ,
         \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 ,
         \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 ,
         \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 ,
         \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 ,
         \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 ,
         \5072 , \5073 , \5074 , \5075_nG2232 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 ,
         \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 ,
         \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100_nG220e , \5101 ,
         \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 ,
         \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 ,
         \5122 , \5123 , \5124 , \5125_nG207b , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 ,
         \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 ,
         \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150_nG2057 , \5151 ,
         \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 ,
         \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 ,
         \5172 , \5173 , \5174 , \5175_nG1ed8 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 ,
         \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 ,
         \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200_nG1eb4 , \5201 ,
         \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 ,
         \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 ,
         \5222 , \5223 , \5224 , \5225_nG1d69 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 ,
         \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 ,
         \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250_nG1d45 , \5251 ,
         \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 ,
         \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 ,
         \5272 , \5273 , \5274 , \5275_nG1c2a , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 ,
         \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 ,
         \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300_nG1c43 , \5301 ,
         \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 ,
         \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 ,
         \5322 , \5323 , \5324 , \5325_nG1b40 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 ,
         \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 ,
         \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349_nG1b24 , \5350 , \5351 ,
         \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 ,
         \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 ,
         \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 ,
         \5382 , \5383 , \5384_nG223b , \5385 , \5386 , \5387 , \5388_nG2217 , \5389 , \5390 , \5391 ,
         \5392_nG2084 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 ,
         \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 ,
         \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 ,
         \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 ,
         \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 ,
         \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 ,
         \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 ,
         \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 ,
         \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 ,
         \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 ,
         \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 ,
         \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 ,
         \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518_nG290c , \5519 , \5520 , \5521 ,
         \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 ,
         \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 ,
         \5542 , \5543 , \5544 , \5545 , \5546_nG23ed , \5547 , \5548 , \5549 , \5550 , \5551 ,
         \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558_nG2402 , \5559 , \5560 , \5561 ,
         \5562_nG23f6 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 ,
         \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 ,
         \5582 , \5583 , \5584 , \5585 , \5586 , \5587_nG2a01 , \5588 , \5589 , \5590 , \5591 ,
         \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 ,
         \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 ,
         \5612 , \5613 , \5614_nG2843 , \5615 , \5616 , \5617 , \5618_nG25dc , \5619 , \5620 , \5621 ,
         \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 ,
         \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 ,
         \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 ,
         \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 ,
         \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 ,
         \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 ,
         \5682 , \5683 , \5684 , \5685_nG2060 , \5686 , \5687 , \5688 , \5689 , \5690_nG1ee1 , \5691 ,
         \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 ,
         \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 ,
         \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 ,
         \5722 , \5723 , \5724 , \5725_nG26a4 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 ,
         \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 ,
         \5742 , \5743 , \5744 , \5745 , \5746_nG2782 , \5747 , \5748 , \5749 , \5750 , \5751 ,
         \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 ,
         \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769_nG25bb , \5770 , \5771 ,
         \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 ,
         \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 ,
         \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 ,
         \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 ,
         \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 ,
         \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 ,
         \5832_nG1b47 , \5833 , \5834 , \5835_nG1b27 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 ,
         \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 ,
         \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 ,
         \5862_nG242a , \5863 , \5864 , \5865 , \5866_nG1c4f , \5867 , \5868 , \5869 , \5870_nG1c53 , \5871 ,
         \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 ,
         \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 ,
         \5892 , \5893 , \5894 , \5895_nG24d7 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 ,
         \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 ,
         \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 ,
         \5922_nG226a , \5923 , \5924 , \5925 , \5926_nG1d72 , \5927 , \5928 , \5929 , \5930_nG1d4e , \5931 ,
         \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 ,
         \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 ,
         \5952 , \5953 , \5954 , \5955_nG2302 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 ,
         \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 ,
         \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 ,
         \5982 , \5983 , \5984_nG209f , \5985 , \5986 , \5987 , \5988_nG1ebd , \5989 , \5990 , \5991 ,
         \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 ,
         \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 ,
         \6012 , \6013_nG2129 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 ,
         \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 ,
         \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039_nG1efc , \6040 , \6041 ,
         \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 ,
         \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060_nG1f70 , \6061 ,
         \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 ,
         \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 ,
         \6082 , \6083 , \6084_nG1d8b , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 ,
         \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 ,
         \6102 , \6103 , \6104 , \6105_nG1df2 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 ,
         \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 ,
         \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 ,
         \6132_nG1c0d , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 ,
         \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 ,
         \6152 , \6153_nG1ca0 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 ,
         \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 ,
         \6172 , \6173 , \6174 , \6175 , \6176_nG1b85 , \6177 , \6178 , \6179 , \6180 , \6181 ,
         \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 ,
         \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 ,
         \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 ,
         \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 ,
         \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 ,
         \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 ,
         \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 ,
         \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 ,
         \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 ,
         \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 ,
         \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 ,
         \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 ,
         \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309_nG1aea , \6310 , \6311 ,
         \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 ,
         \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 ,
         \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 ,
         \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 ,
         \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 ,
         \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 ,
         \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 ,
         \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 ,
         \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 ,
         \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 ,
         \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 ,
         \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 ,
         \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 ,
         \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 ,
         \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 ,
         \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 ,
         \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 ,
         \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 ,
         \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 ,
         \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 ,
         \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 ,
         \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 ,
         \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 ,
         \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 ,
         \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 ,
         \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 ,
         \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 ,
         \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 ,
         \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 ,
         \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 ,
         \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 ,
         \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 ,
         \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 ,
         \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 ,
         \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 ,
         \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 ,
         \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 ,
         \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 ,
         \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 ,
         \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 ,
         \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 ,
         \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 ,
         \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 ,
         \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 ,
         \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 ,
         \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 ,
         \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 ,
         \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 ,
         \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 ,
         \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 ,
         \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 ,
         \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 ,
         \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 ,
         \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 ,
         \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 ,
         \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 ,
         \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 ,
         \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 ,
         \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 ,
         \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 ,
         \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 ,
         \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 ,
         \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 ,
         \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 ,
         \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 ,
         \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 ,
         \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 ,
         \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 ,
         \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 ,
         \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 ,
         \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 ,
         \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 ,
         \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 ,
         \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 ,
         \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 ,
         \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 ,
         \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 ,
         \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 ,
         \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 ,
         \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 ,
         \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 ,
         \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 ,
         \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 ,
         \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 ,
         \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 ,
         \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 ,
         \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 ,
         \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 ,
         \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 ,
         \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 ,
         \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 ,
         \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 ,
         \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 ,
         \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 ,
         \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 ,
         \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 ,
         \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 ,
         \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 ,
         \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 ,
         \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 ,
         \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 ,
         \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 ,
         \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 ,
         \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 ,
         \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 ,
         \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 ,
         \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 ,
         \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 ,
         \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 ,
         \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 ,
         \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 ,
         \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 ,
         \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 ,
         \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 ,
         \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 ,
         \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 ,
         \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 ,
         \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 ,
         \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 ,
         \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 ,
         \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
         \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 ,
         \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 ,
         \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 ,
         \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 ,
         \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 ,
         \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 ,
         \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 ,
         \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 ,
         \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 ,
         \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 ,
         \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 ,
         \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 ,
         \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 ,
         \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 ,
         \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 ,
         \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 ,
         \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 ,
         \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 ,
         \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 ,
         \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 ,
         \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 ,
         \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 ,
         \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 ,
         \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 ,
         \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 ,
         \7772_nG32b2 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 ,
         \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 ,
         \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 ,
         \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 ,
         \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 ,
         \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 ,
         \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 ,
         \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 ,
         \7852 , \7853 , \7854_nG1080 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 ,
         \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 ,
         \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879_nG1099 , \7880 , \7881 ,
         \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 ,
         \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 ,
         \7902 , \7903 , \7904_nG10b2 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 ,
         \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 ,
         \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929_nG10cb , \7930 , \7931 ,
         \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 ,
         \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 ,
         \7952 , \7953 , \7954_nG10e4 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 ,
         \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 ,
         \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979_nG10fd , \7980 , \7981 ,
         \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 ,
         \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 ,
         \8002 , \8003 , \8004_nG1116 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 ,
         \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 ,
         \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029_nG112f , \8030 , \8031 ,
         \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 ,
         \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 ,
         \8052 , \8053 , \8054_nG1148 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 ,
         \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 ,
         \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079_nG1161 , \8080 , \8081 ,
         \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 ,
         \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 ,
         \8102 , \8103 , \8104_nG117a , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 ,
         \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 ,
         \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129_nG1193 , \8130 , \8131 ,
         \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 ,
         \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 ,
         \8152 , \8153_nG11ad , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 ,
         \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 ,
         \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 ,
         \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 ,
         \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 ,
         \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 ,
         \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 ,
         \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 ,
         \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 ,
         \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 ,
         \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 ,
         \8262 , \8263_nG1220 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 ,
         \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 ,
         \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 ,
         \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 ,
         \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 ,
         \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318_nG1257 , \8319 , \8320 , \8321 ,
         \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 ,
         \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339_nG126c , \8340 , \8341 ,
         \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 ,
         \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360_nG1281 , \8361 ,
         \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 ,
         \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381_nG1296 ,
         \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 ,
         \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 ,
         \8402_nG12ab , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 ,
         \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 ,
         \8422 , \8423_nG12c0 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 ,
         \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 ,
         \8442 , \8443 , \8444_nG12d5 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 ,
         \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 ,
         \8462 , \8463 , \8464 , \8465_nG12ea , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 ,
         \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 ,
         \8482 , \8483 , \8484 , \8485 , \8486_nG12ff , \8487 , \8488 , \8489 , \8490 , \8491 ,
         \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 ,
         \8502 , \8503 , \8504 , \8505 , \8506 , \8507_nG1314 , \8508 , \8509 , \8510 , \8511 ,
         \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 ,
         \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528_nG1329 , \8529 , \8530 , \8531 ,
         \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 ,
         \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549_nG133e , \8550 , \8551 ,
         \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 ,
         \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570_nG1353 , \8571 ,
         \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 ,
         \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591_nG1368 ,
         \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 ,
         \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 ,
         \8612_nG137d , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 ,
         \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 ,
         \8632 , \8633_nG1392 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 ,
         \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 ,
         \8652 , \8653 , \8654_nG13a7 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 ,
         \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 ,
         \8672 , \8673 , \8674 , \8675_nG13bc , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 ,
         \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 ,
         \8692 , \8693 , \8694 , \8695 , \8696_nG13d1 , \8697 , \8698 , \8699 , \8700 , \8701 ,
         \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 ,
         \8712 , \8713 , \8714 , \8715 , \8716 , \8717_nG13e6 , \8718 , \8719 , \8720 , \8721 ,
         \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 ,
         \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738_nG13fb , \8739 , \8740 , \8741 ,
         \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 ,
         \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759_nG1410 , \8760 , \8761 ,
         \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 ,
         \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780_nG1425 , \8781 ,
         \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 ,
         \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801_nG143a ,
         \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 ,
         \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 ,
         \8822_nG144f , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 ,
         \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 ,
         \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 ,
         \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 ,
         \8862 , \8863_nG32b3 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 ,
         \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 ,
         \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 ,
         \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 ,
         \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 ,
         \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 ,
         \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 ,
         \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 ,
         \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 ,
         \8952 , \8953 , \8954 , \8955 , \8956_nG3221 , \8957 , \8958 , \8959 , \8960 , \8961 ,
         \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 ,
         \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 ,
         \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 ,
         \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 ,
         \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 ,
         \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 ,
         \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 ,
         \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 ,
         \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048_nG3255 , \9049_nG3256 , \9050 , \9051 ,
         \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 ,
         \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 ,
         \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 ,
         \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 ,
         \9092 , \9093 , \9094 , \9095_nG31b2 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 ,
         \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 ,
         \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 ,
         \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 ,
         \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140_nG31ec , \9141_nG31ed ,
         \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 ,
         \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 ,
         \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 ,
         \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 ,
         \9182 , \9183 , \9184 , \9185 , \9186_nG3135 , \9187 , \9188 , \9189 , \9190 , \9191 ,
         \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 ,
         \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 ,
         \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 ,
         \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230_nG3177 , \9231_nG3178 ,
         \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 ,
         \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 ,
         \9252 , \9253 , \9254_nG30ac , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 ,
         \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 ,
         \9272 , \9273 , \9274 , \9275 , \9276_nG30f2 , \9277_nG30f3 , \9278 , \9279 , \9280 , \9281 ,
         \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 ,
         \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300_nG301d , \9301 ,
         \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 ,
         \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 ,
         \9322_nG3065 , \9323_nG3066 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 ,
         \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 ,
         \9342 , \9343 , \9344 , \9345_nG2f88 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 ,
         \9352 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 ,
         \9362 , \9363 , \9364 , \9365 , \9366_nG2fd4 , \9367_nG2fd5 , \9368 , \9369 , \9370 , \9371 ,
         \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 ,
         \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389_nG2eeb , \9390 , \9391 ,
         \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 ,
         \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410_nG2f3b , \9411_nG2f3c ,
         \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 ,
         \9422 , \9423_nG2e49 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 ,
         \9432 , \9433 , \9434_nG2e9a , \9435_nG2e9b , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 ,
         \9442 , \9443 , \9444 , \9445 , \9446 , \9447_nG2d9e , \9448 , \9449 , \9450 , \9451 ,
         \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458_nG2df7 , \9459_nG2df8 , \9460 , \9461 ,
         \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471_nG2ce8 ,
         \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 ,
         \9482_nG2d44 , \9483_nG2d45 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 ,
         \9492 , \9493 , \9494 , \9495_nG2c2b , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 ,
         \9502 , \9503 , \9504 , \9505 , \9506_nG2c8b , \9507_nG2c8c , \9508 , \9509 , \9510 , \9511 ,
         \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518_nG2b6b , \9519 , \9520 , \9521 ,
         \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528_nG2bca , \9529_nG2bcb , \9530 , \9531 ,
         \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540_nG2aac , \9541 ,
         \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550_nG2b0b , \9551_nG2b0c ,
         \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 ,
         \9562_nG29d8 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 ,
         \9572_nG2a4c , \9573_nG2a4d , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 ,
         \9582 , \9583 , \9584_nG28f0 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 ,
         \9592 , \9593 , \9594_nG2963 , \9595_nG2964 , \9596 , \9597 , \9598 , \9599 , \9600_nG2810 , \9601 ,
         \9602 , \9603 , \9604_nG287c , \9605_nG287d , \9606 , \9607 , \9608 , \9609 , \9610_nG2737 , \9611 ,
         \9612 , \9613 , \9614_nG27a3 , \9615_nG27a4 , \9616 , \9617 , \9618 , \9619 , \9620_nG2662 , \9621 ,
         \9622 , \9623 , \9624_nG26ca , \9625_nG26cb , \9626 , \9627 , \9628 , \9629 , \9630_nG258f , \9631 ,
         \9632 , \9633 , \9634_nG25f9 , \9635_nG25fa , \9636 , \9637 , \9638 , \9639 , \9640_nG24bf , \9641 ,
         \9642 , \9643 , \9644_nG2524 , \9645_nG2525 , \9646 , \9647 , \9648 , \9649 , \9650_nG23cd , \9651 ,
         \9652 , \9653 , \9654_nG2459 , \9655_nG245a , \9656 , \9657 , \9658 , \9659 , \9660_nG22e6 , \9661 ,
         \9662 , \9663 , \9664_nG2340 , \9665_nG2341 , \9666 , \9667 , \9668 , \9669 , \9670_nG21f2 , \9671 ,
         \9672 , \9673 , \9674_nG228b , \9675_nG228c , \9676 , \9677 , \9678 , \9679 , \9680_nG210a , \9681 ,
         \9682 , \9683 , \9684_nG2158 , \9685_nG2159 , \9686 , \9687 , \9688 , \9689 , \9690_nG202e , \9691 ,
         \9692 , \9693 , \9694_nG20bb , \9695_nG20bc , \9696 , \9697 , \9698 , \9699 , \9700_nG1f5c , \9701 ,
         \9702 , \9703 , \9704_nG1fa0 , \9705_nG1fa1 , \9706 , \9707 , \9708 , \9709 , \9710_nG1e94 , \9711 ,
         \9712 , \9713 , \9714_nG1f17 , \9715_nG1f18 , \9716 , \9717 , \9718 , \9719 , \9720_nG1dda , \9721 ,
         \9722 , \9723 , \9724_nG1e10 , \9725_nG1e11 , \9726 , \9727 , \9728 , \9729 , \9730_nG1d2d , \9731 ,
         \9732 , \9733 , \9734_nG1da3 , \9735_nG1da4 , \9736 , \9737 , \9738 , \9739 , \9740_nG1c8c , \9741 ,
         \9742 , \9743 , \9744_nG1cb6 , \9745_nG1cb7 , \9746 , \9747 , \9748 , \9749 , \9750_nG1bf9 , \9751 ,
         \9752 , \9753 , \9754_nG1c61 , \9755_nG1c62 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761_nG1b6e ,
         \9762 , \9763 , \9764 , \9765 , \9766_nG1b90 , \9767_nG1b91 , \9768 , \9769 , \9770_nG1ab0 , \9771 ,
         \9772_nG1b4b , \9773_nG1b4c , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 ,
         \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 ,
         \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 ,
         \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 ,
         \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 ,
         \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 ,
         \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 ,
         \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 ,
         \9852 , \9853 , \9854 , \9855_nG3a87 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 ,
         \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 ,
         \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880_nG3a63 , \9881 ,
         \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 ,
         \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 ,
         \9902 , \9903 , \9904 , \9905_nG38dc , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 ,
         \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 ,
         \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930_nG38b8 , \9931 ,
         \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 ,
         \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 ,
         \9952 , \9953 , \9954 , \9955_nG3743 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 ,
         \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 ,
         \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980_nG371f , \9981 ,
         \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 ,
         \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 ,
         \10002 , \10003 , \10004 , \10005_nG35e1 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 ,
         \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 ,
         \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030_nG35bd , \10031 ,
         \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 ,
         \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 ,
         \10052 , \10053 , \10054 , \10055_nG34b0 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 ,
         \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 ,
         \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080_nG34c9 , \10081 ,
         \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 ,
         \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 ,
         \10102 , \10103 , \10104 , \10105_nG3393 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 ,
         \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 ,
         \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129_nG3377 , \10130 , \10131 ,
         \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 ,
         \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 ,
         \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 ,
         \10162 , \10163 , \10164_nG3a90 , \10165 , \10166 , \10167 , \10168_nG3a6c , \10169 , \10170 , \10171 ,
         \10172_nG38e5 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 ,
         \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 ,
         \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 ,
         \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 ,
         \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 ,
         \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 ,
         \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 ,
         \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 ,
         \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 ,
         \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 ,
         \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 ,
         \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 ,
         \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298_nG4187 , \10299 , \10300 , \10301 ,
         \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 ,
         \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 ,
         \10322 , \10323 , \10324 , \10325 , \10326_nG3c4f , \10327 , \10328 , \10329 , \10330 , \10331 ,
         \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338_nG3c64 , \10339 , \10340 , \10341 ,
         \10342_nG3c58 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 ,
         \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 ,
         \10362 , \10363 , \10364 , \10365 , \10366 , \10367_nG427b , \10368 , \10369 , \10370 , \10371 ,
         \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 ,
         \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 ,
         \10392 , \10393 , \10394_nG40c5 , \10395 , \10396 , \10397 , \10398_nG3e60 , \10399 , \10400 , \10401 ,
         \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 ,
         \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 ,
         \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 ,
         \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 ,
         \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 ,
         \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 ,
         \10462 , \10463 , \10464 , \10465_nG38c1 , \10466 , \10467 , \10468 , \10469 , \10470_nG374c , \10471 ,
         \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 ,
         \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 ,
         \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 ,
         \10502 , \10503 , \10504 , \10505_nG3f2a , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 ,
         \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 ,
         \10522 , \10523 , \10524 , \10525 , \10526_nG4004 , \10527 , \10528 , \10529 , \10530 , \10531 ,
         \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 ,
         \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549_nG3e3f , \10550 , \10551 ,
         \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 ,
         \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 ,
         \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 ,
         \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 ,
         \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 ,
         \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 ,
         \10612_nG339a , \10613 , \10614 , \10615_nG337a , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 ,
         \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 ,
         \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 ,
         \10642_nG3c8c , \10643 , \10644 , \10645 , \10646_nG34d5 , \10647 , \10648 , \10649 , \10650_nG34d9 , \10651 ,
         \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 ,
         \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 ,
         \10672 , \10673 , \10674 , \10675_nG3d60 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 ,
         \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 ,
         \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 ,
         \10702_nG3abf , \10703 , \10704 , \10705 , \10706_nG35ea , \10707 , \10708 , \10709 , \10710_nG35c6 , \10711 ,
         \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 ,
         \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 ,
         \10732 , \10733 , \10734 , \10735_nG3b96 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 ,
         \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 ,
         \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 ,
         \10762 , \10763 , \10764_nG3900 , \10765 , \10766 , \10767 , \10768_nG3728 , \10769 , \10770 , \10771 ,
         \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 ,
         \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 ,
         \10792 , \10793_nG39c9 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 ,
         \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 ,
         \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819_nG3767 , \10820 , \10821 ,
         \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 ,
         \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840_nG381a , \10841 ,
         \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 ,
         \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 ,
         \10862 , \10863 , \10864_nG3603 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 ,
         \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 ,
         \10882 , \10883 , \10884 , \10885_nG36aa , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 ,
         \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 ,
         \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 ,
         \10912_nG3493 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 ,
         \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 ,
         \10932 , \10933_nG3564 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 ,
         \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 ,
         \10952 , \10953 , \10954 , \10955 , \10956_nG3451 , \10957 , \10958 , \10959 , \10960 , \10961 ,
         \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 ,
         \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 ,
         \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 ,
         \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 ,
         \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 ,
         \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 ,
         \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 ,
         \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 ,
         \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 ,
         \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 ,
         \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 ,
         \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 ,
         \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089_nG333d , \11090 , \11091 ,
         \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 ,
         \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 ,
         \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 ,
         \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 ,
         \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 ,
         \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 ,
         \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 ,
         \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 ,
         \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 ,
         \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 ,
         \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 ,
         \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 ,
         \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 ,
         \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 ,
         \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 ,
         \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 ,
         \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 ,
         \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 ,
         \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 ,
         \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 ,
         \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 ,
         \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 ,
         \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 ,
         \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 ,
         \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 ,
         \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 ,
         \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 ,
         \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 ,
         \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 ,
         \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 ,
         \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 ,
         \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 ,
         \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 ,
         \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 ,
         \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 ,
         \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 ,
         \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 ,
         \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 ,
         \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 ,
         \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 ,
         \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 ,
         \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 ,
         \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 ,
         \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 ,
         \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 ,
         \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 ,
         \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 ,
         \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 ,
         \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 ,
         \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 ,
         \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 ,
         \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 ,
         \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 ,
         \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 ,
         \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 ,
         \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 ,
         \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 ,
         \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 ,
         \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 ,
         \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 ,
         \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 ,
         \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 ,
         \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 ,
         \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 ,
         \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 ,
         \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 ,
         \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 ,
         \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 ,
         \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 ,
         \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 ,
         \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 ,
         \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 ,
         \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 ,
         \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 ,
         \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 ,
         \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 ,
         \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 ,
         \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 ,
         \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 ,
         \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 ,
         \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 ,
         \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 ,
         \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 ,
         \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 ,
         \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 ,
         \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 ,
         \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 ,
         \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 ,
         \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 ,
         \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 ,
         \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 ,
         \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 ,
         \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 ,
         \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 ,
         \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 ,
         \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 ,
         \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 ,
         \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 ,
         \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 ,
         \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 ,
         \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 ,
         \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 ,
         \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 ,
         \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 ,
         \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 ,
         \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 ,
         \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 ,
         \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 ,
         \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 ,
         \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 ,
         \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 ,
         \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 ,
         \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 ,
         \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 ,
         \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 ,
         \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 ,
         \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 ,
         \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 ,
         \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 ,
         \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 ,
         \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 ,
         \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 ,
         \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 ,
         \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 ,
         \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 ,
         \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 ,
         \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 ,
         \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 ,
         \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 ,
         \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 ,
         \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 ,
         \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 ,
         \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 ,
         \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 ,
         \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 ,
         \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 ,
         \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 ,
         \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 ,
         \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 ,
         \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 ,
         \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 ,
         \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 ,
         \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 ,
         \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 ,
         \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 ,
         \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 ,
         \12552_nG4b72 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 ,
         \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 ,
         \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 ,
         \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 ,
         \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 ,
         \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 ,
         \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 ,
         \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 ,
         \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 ,
         \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 ,
         \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 ,
         \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 ,
         \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 ,
         \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 ,
         \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701_nG3b20 ,
         \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 ,
         \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 ,
         \12722 , \12723 , \12724 , \12725 , \12726_nG3afc , \12727 , \12728 , \12729 , \12730 , \12731 ,
         \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 ,
         \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751_nG3969 ,
         \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 ,
         \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 ,
         \12772 , \12773 , \12774 , \12775 , \12776_nG3945 , \12777 , \12778 , \12779 , \12780 , \12781 ,
         \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 ,
         \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801_nG37c6 ,
         \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 ,
         \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 ,
         \12822 , \12823 , \12824 , \12825 , \12826_nG37a2 , \12827 , \12828 , \12829 , \12830 , \12831 ,
         \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 ,
         \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851_nG3657 ,
         \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 ,
         \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 ,
         \12872 , \12873 , \12874 , \12875 , \12876_nG3633 , \12877 , \12878 , \12879 , \12880 , \12881 ,
         \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 ,
         \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901_nG3518 ,
         \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 ,
         \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 ,
         \12922 , \12923 , \12924 , \12925 , \12926_nG3531 , \12927 , \12928 , \12929 , \12930 , \12931 ,
         \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 ,
         \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951_nG342e ,
         \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 ,
         \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 ,
         \12972 , \12973 , \12974 , \12975_nG3412 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 ,
         \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 ,
         \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 ,
         \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010_nG3b29 , \13011 ,
         \13012 , \13013 , \13014_nG3b05 , \13015 , \13016 , \13017 , \13018_nG3972 , \13019 , \13020 , \13021 ,
         \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 ,
         \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 ,
         \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 ,
         \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 ,
         \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 ,
         \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 ,
         \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 ,
         \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 ,
         \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 ,
         \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 ,
         \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 ,
         \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 ,
         \13142 , \13143 , \13144_nG41fa , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 ,
         \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 ,
         \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 ,
         \13172_nG3cdb , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 ,
         \13182 , \13183 , \13184_nG3cf0 , \13185 , \13186 , \13187 , \13188_nG3ce4 , \13189 , \13190 , \13191 ,
         \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 ,
         \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 ,
         \13212 , \13213_nG42ef , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 ,
         \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 ,
         \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240_nG4131 , \13241 ,
         \13242 , \13243 , \13244_nG3eca , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 ,
         \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 ,
         \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 ,
         \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 ,
         \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 ,
         \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 ,
         \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311_nG394e ,
         \13312 , \13313 , \13314 , \13315 , \13316_nG37cf , \13317 , \13318 , \13319 , \13320 , \13321 ,
         \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 ,
         \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 ,
         \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351_nG3f92 ,
         \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 ,
         \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 ,
         \13372_nG4070 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 ,
         \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 ,
         \13392 , \13393 , \13394 , \13395_nG3ea9 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 ,
         \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 ,
         \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 ,
         \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 ,
         \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 ,
         \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 ,
         \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458_nG3435 , \13459 , \13460 , \13461_nG3415 ,
         \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 ,
         \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 ,
         \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488_nG3d18 , \13489 , \13490 , \13491 ,
         \13492_nG353d , \13493 , \13494 , \13495 , \13496_nG3541 , \13497 , \13498 , \13499 , \13500 , \13501 ,
         \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 ,
         \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521_nG3dc5 ,
         \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 ,
         \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 ,
         \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548_nG3b58 , \13549 , \13550 , \13551 ,
         \13552_nG3660 , \13553 , \13554 , \13555 , \13556_nG363c , \13557 , \13558 , \13559 , \13560 , \13561 ,
         \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 ,
         \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581_nG3bf0 ,
         \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 ,
         \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 ,
         \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610_nG398d , \13611 ,
         \13612 , \13613 , \13614_nG37ab , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 ,
         \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 ,
         \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639_nG3a17 , \13640 , \13641 ,
         \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 ,
         \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 ,
         \13662 , \13663 , \13664 , \13665_nG37ea , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 ,
         \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 ,
         \13682 , \13683 , \13684 , \13685 , \13686_nG385e , \13687 , \13688 , \13689 , \13690 , \13691 ,
         \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 ,
         \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710_nG3679 , \13711 ,
         \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 ,
         \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731_nG36e0 ,
         \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 ,
         \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 ,
         \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758_nG34fb , \13759 , \13760 , \13761 ,
         \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 ,
         \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779_nG358e , \13780 , \13781 ,
         \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 ,
         \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 ,
         \13802_nG3473 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 ,
         \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 ,
         \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 ,
         \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 ,
         \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 ,
         \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 ,
         \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 ,
         \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 ,
         \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 ,
         \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 ,
         \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 ,
         \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 ,
         \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 ,
         \13932 , \13933 , \13934 , \13935_nG33d8 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 ,
         \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 ,
         \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 ,
         \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 ,
         \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 ,
         \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 ,
         \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 ,
         \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 ,
         \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 ,
         \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 ,
         \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 ,
         \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 ,
         \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 ,
         \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 ,
         \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 ,
         \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 ,
         \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 ,
         \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 ,
         \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 ,
         \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 ,
         \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 ,
         \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 ,
         \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 ,
         \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 ,
         \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 ,
         \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 ,
         \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 ,
         \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 ,
         \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 ,
         \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 ,
         \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 ,
         \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 ,
         \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 ,
         \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 ,
         \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 ,
         \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 ,
         \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 ,
         \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 ,
         \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 ,
         \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 ,
         \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 ,
         \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 ,
         \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 ,
         \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 ,
         \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 ,
         \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 ,
         \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 ,
         \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 ,
         \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 ,
         \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 ,
         \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 ,
         \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 ,
         \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 ,
         \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 ,
         \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 ,
         \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 ,
         \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 ,
         \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 ,
         \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 ,
         \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 ,
         \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 ,
         \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 ,
         \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 ,
         \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 ,
         \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 ,
         \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 ,
         \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 ,
         \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 ,
         \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 ,
         \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 ,
         \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 ,
         \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 ,
         \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 ,
         \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 ,
         \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 ,
         \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 ,
         \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 ,
         \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 ,
         \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 ,
         \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 ,
         \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 ,
         \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 ,
         \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 ,
         \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 ,
         \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 ,
         \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 ,
         \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 ,
         \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 ,
         \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 ,
         \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 ,
         \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 ,
         \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 ,
         \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 ,
         \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 ,
         \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 ,
         \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 ,
         \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 ,
         \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 ,
         \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 ,
         \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 ,
         \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 ,
         \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 ,
         \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 ,
         \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 ,
         \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 ,
         \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 ,
         \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 ,
         \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 ,
         \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 ,
         \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 ,
         \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 ,
         \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 ,
         \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 ,
         \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 ,
         \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 ,
         \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 ,
         \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 ,
         \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 ,
         \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 ,
         \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 ,
         \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 ,
         \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 ,
         \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 ,
         \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 ,
         \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 ,
         \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 ,
         \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 ,
         \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 ,
         \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 ,
         \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 ,
         \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 ,
         \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 ,
         \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 ,
         \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 ,
         \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 ,
         \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 ,
         \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 ,
         \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 ,
         \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 ,
         \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 ,
         \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 ,
         \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 ,
         \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 ,
         \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 ,
         \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 ,
         \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 ,
         \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398_nG4ba0 , \15399 , \15400 , \15401 ,
         \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 ,
         \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 ,
         \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 ,
         \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 ,
         \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 ,
         \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 ,
         \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 ,
         \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480_nG1512 , \15481 ,
         \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 ,
         \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 ,
         \15502 , \15503 , \15504 , \15505_nG152b , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 ,
         \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 ,
         \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530_nG1544 , \15531 ,
         \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 ,
         \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 ,
         \15552 , \15553 , \15554 , \15555_nG155d , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 ,
         \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 ,
         \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580_nG1576 , \15581 ,
         \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 ,
         \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 ,
         \15602 , \15603 , \15604 , \15605_nG158f , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 ,
         \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 ,
         \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630_nG15a8 , \15631 ,
         \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 ,
         \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 ,
         \15652 , \15653 , \15654 , \15655_nG15c1 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 ,
         \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 ,
         \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680_nG15da , \15681 ,
         \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 ,
         \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 ,
         \15702 , \15703 , \15704 , \15705_nG15f3 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 ,
         \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 ,
         \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730_nG160c , \15731 ,
         \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 ,
         \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 ,
         \15752 , \15753 , \15754 , \15755_nG1625 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 ,
         \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 ,
         \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779_nG163f , \15780 , \15781 ,
         \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 ,
         \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 ,
         \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 ,
         \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 ,
         \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 ,
         \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 ,
         \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 ,
         \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 ,
         \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 ,
         \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 ,
         \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889_nG16b2 , \15890 , \15891 ,
         \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 ,
         \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 ,
         \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 ,
         \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 ,
         \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 ,
         \15942 , \15943 , \15944_nG16e9 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 ,
         \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 ,
         \15962 , \15963 , \15964 , \15965_nG16fe , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 ,
         \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 ,
         \15982 , \15983 , \15984 , \15985 , \15986_nG1713 , \15987 , \15988 , \15989 , \15990 , \15991 ,
         \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 ,
         \16002 , \16003 , \16004 , \16005 , \16006 , \16007_nG1728 , \16008 , \16009 , \16010 , \16011 ,
         \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 ,
         \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028_nG173d , \16029 , \16030 , \16031 ,
         \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 ,
         \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049_nG1752 , \16050 , \16051 ,
         \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 ,
         \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070_nG1767 , \16071 ,
         \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 ,
         \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091_nG177c ,
         \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 ,
         \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 ,
         \16112_nG1791 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 ,
         \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 ,
         \16132 , \16133_nG17a6 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 ,
         \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 ,
         \16152 , \16153 , \16154_nG17bb , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 ,
         \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 ,
         \16172 , \16173 , \16174 , \16175_nG17d0 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 ,
         \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 ,
         \16192 , \16193 , \16194 , \16195 , \16196_nG17e5 , \16197 , \16198 , \16199 , \16200 , \16201 ,
         \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 ,
         \16212 , \16213 , \16214 , \16215 , \16216 , \16217_nG17fa , \16218 , \16219 , \16220 , \16221 ,
         \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 ,
         \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238_nG180f , \16239 , \16240 , \16241 ,
         \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 ,
         \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259_nG1824 , \16260 , \16261 ,
         \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 ,
         \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280_nG1839 , \16281 ,
         \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 ,
         \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301_nG184e ,
         \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 ,
         \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 ,
         \16322_nG1863 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 ,
         \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 ,
         \16342 , \16343_nG1878 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 ,
         \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 ,
         \16362 , \16363 , \16364_nG188d , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 ,
         \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 ,
         \16382 , \16383 , \16384 , \16385_nG18a2 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 ,
         \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 ,
         \16402 , \16403 , \16404 , \16405 , \16406_nG18b7 , \16407 , \16408 , \16409 , \16410 , \16411 ,
         \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 ,
         \16422 , \16423 , \16424 , \16425 , \16426 , \16427_nG18cc , \16428 , \16429 , \16430 , \16431 ,
         \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 ,
         \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448_nG18e1 , \16449 , \16450 , \16451 ,
         \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 ,
         \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 ,
         \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 ,
         \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489_nG4ba1 , \16490 , \16491 ,
         \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 ,
         \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 ,
         \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 ,
         \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 ,
         \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 ,
         \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 ,
         \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 ,
         \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 ,
         \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 ,
         \16582_nG4b0f , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 ,
         \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 ,
         \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 ,
         \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 ,
         \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 ,
         \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 ,
         \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 ,
         \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 ,
         \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 ,
         \16672 , \16673 , \16674_nG4b43 , \16675_nG4b44 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 ,
         \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 ,
         \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 ,
         \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 ,
         \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721_nG4aa0 ,
         \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 ,
         \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 ,
         \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 ,
         \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 ,
         \16762 , \16763 , \16764 , \16765 , \16766_nG4ada , \16767_nG4adb , \16768 , \16769 , \16770 , \16771 ,
         \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 ,
         \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 ,
         \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 ,
         \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 ,
         \16812_nG4a23 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 ,
         \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 ,
         \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 ,
         \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 ,
         \16852 , \16853 , \16854 , \16855 , \16856_nG4a65 , \16857_nG4a66 , \16858 , \16859 , \16860 , \16861 ,
         \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 ,
         \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880_nG499a , \16881 ,
         \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 ,
         \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 ,
         \16902_nG49e0 , \16903_nG49e1 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 ,
         \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 ,
         \16922 , \16923 , \16924 , \16925 , \16926_nG490b , \16927 , \16928 , \16929 , \16930 , \16931 ,
         \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 ,
         \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948_nG4953 , \16949_nG4954 , \16950 , \16951 ,
         \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 ,
         \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971_nG4876 ,
         \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 ,
         \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 ,
         \16992_nG48c2 , \16993_nG48c3 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 ,
         \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 ,
         \17012 , \17013 , \17014 , \17015_nG47d9 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 ,
         \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 ,
         \17032 , \17033 , \17034 , \17035 , \17036_nG4829 , \17037_nG482a , \17038 , \17039 , \17040 , \17041 ,
         \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049_nG4737 , \17050 , \17051 ,
         \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060_nG4788 , \17061_nG4789 ,
         \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 ,
         \17072 , \17073_nG468c , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 ,
         \17082 , \17083 , \17084_nG46e5 , \17085_nG46e6 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 ,
         \17092 , \17093 , \17094 , \17095 , \17096 , \17097_nG45d6 , \17098 , \17099 , \17100 , \17101 ,
         \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108_nG4632 , \17109_nG4633 , \17110 , \17111 ,
         \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121_nG4519 ,
         \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 ,
         \17132_nG4579 , \17133_nG457a , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 ,
         \17142 , \17143 , \17144_nG4459 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 ,
         \17152 , \17153 , \17154_nG44b8 , \17155_nG44b9 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 ,
         \17162 , \17163 , \17164 , \17165 , \17166_nG439a , \17167 , \17168 , \17169 , \17170 , \17171 ,
         \17172 , \17173 , \17174 , \17175 , \17176_nG43f9 , \17177_nG43fa , \17178 , \17179 , \17180 , \17181 ,
         \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188_nG42c6 , \17189 , \17190 , \17191 ,
         \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198_nG433a , \17199_nG433b , \17200 , \17201 ,
         \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210_nG41de , \17211 ,
         \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220_nG4251 , \17221_nG4252 ,
         \17222 , \17223 , \17224 , \17225 , \17226_nG40fe , \17227 , \17228 , \17229 , \17230_nG416a , \17231_nG416b ,
         \17232 , \17233 , \17234 , \17235 , \17236_nG4025 , \17237 , \17238 , \17239 , \17240_nG4091 , \17241_nG4092 ,
         \17242 , \17243 , \17244 , \17245 , \17246_nG3f50 , \17247 , \17248 , \17249 , \17250_nG3fb8 , \17251_nG3fb9 ,
         \17252 , \17253 , \17254 , \17255 , \17256_nG3e7d , \17257 , \17258 , \17259 , \17260_nG3ee7 , \17261_nG3ee8 ,
         \17262 , \17263 , \17264 , \17265 , \17266_nG3dad , \17267 , \17268 , \17269 , \17270_nG3e12 , \17271_nG3e13 ,
         \17272 , \17273 , \17274 , \17275 , \17276_nG3cbb , \17277 , \17278 , \17279 , \17280_nG3d47 , \17281_nG3d48 ,
         \17282 , \17283 , \17284 , \17285 , \17286_nG3bd4 , \17287 , \17288 , \17289 , \17290_nG3c2e , \17291_nG3c2f ,
         \17292 , \17293 , \17294 , \17295 , \17296_nG3ae0 , \17297 , \17298 , \17299 , \17300_nG3b79 , \17301_nG3b7a ,
         \17302 , \17303 , \17304 , \17305 , \17306_nG39f8 , \17307 , \17308 , \17309 , \17310_nG3a46 , \17311_nG3a47 ,
         \17312 , \17313 , \17314 , \17315 , \17316_nG391c , \17317 , \17318 , \17319 , \17320_nG39a9 , \17321_nG39aa ,
         \17322 , \17323 , \17324 , \17325 , \17326_nG384a , \17327 , \17328 , \17329 , \17330_nG388e , \17331_nG388f ,
         \17332 , \17333 , \17334 , \17335 , \17336_nG3782 , \17337 , \17338 , \17339 , \17340_nG3805 , \17341_nG3806 ,
         \17342 , \17343 , \17344 , \17345 , \17346_nG36c8 , \17347 , \17348 , \17349 , \17350_nG36fe , \17351_nG36ff ,
         \17352 , \17353 , \17354 , \17355 , \17356_nG361b , \17357 , \17358 , \17359 , \17360_nG3691 , \17361_nG3692 ,
         \17362 , \17363 , \17364 , \17365 , \17366_nG357a , \17367 , \17368 , \17369 , \17370_nG35a4 , \17371_nG35a5 ,
         \17372 , \17373 , \17374 , \17375 , \17376_nG34e7 , \17377 , \17378 , \17379 , \17380_nG354f , \17381_nG3550 ,
         \17382 , \17383 , \17384 , \17385 , \17386 , \17387_nG345c , \17388 , \17389 , \17390 , \17391 ,
         \17392_nG347e , \17393_nG347f , \17394 , \17395 , \17396_nG339e , \17397 , \17398_nG3439 , \17399_nG343a , \17400 ;
buf \U$labaj1815 ( R_267_b04ddc8, \8864 );
buf \U$labaj1816 ( R_268_b04de70, \9050 );
buf \U$labaj1817 ( R_269_b04df18, \9142 );
buf \U$labaj1818 ( R_26a_b04dfc0, \9232 );
buf \U$labaj1819 ( R_26b_b04e068, \9278 );
buf \U$labaj1820 ( R_26c_b04e110, \9324 );
buf \U$labaj1821 ( R_26d_b04e1b8, \9368 );
buf \U$labaj1822 ( R_26e_b04e260, \9412 );
buf \U$labaj1823 ( R_26f_b04e308, \9436 );
buf \U$labaj1824 ( R_270_b04e3b0, \9460 );
buf \U$labaj1825 ( R_271_b04e458, \9484 );
buf \U$labaj1826 ( R_272_b04e500, \9508 );
buf \U$labaj1827 ( R_273_b04e5a8, \9530 );
buf \U$labaj1828 ( R_274_b04e650, \9552 );
buf \U$labaj1829 ( R_275_b04e6f8, \9574 );
buf \U$labaj1830 ( R_276_b04e7a0, \9596 );
buf \U$labaj1831 ( R_277_b04e848, \9606 );
buf \U$labaj1832 ( R_278_b04e8f0, \9616 );
buf \U$labaj1833 ( R_279_b04e998, \9626 );
buf \U$labaj1834 ( R_27a_b04ea40, \9636 );
buf \U$labaj1835 ( R_27b_b04eae8, \9646 );
buf \U$labaj1836 ( R_27c_b04eb90, \9656 );
buf \U$labaj1837 ( R_27d_b04ec38, \9666 );
buf \U$labaj1838 ( R_27e_b04ece0, \9676 );
buf \U$labaj1839 ( R_27f_b04ed88, \9686 );
buf \U$labaj1840 ( R_280_b04ee30, \9696 );
buf \U$labaj1841 ( R_281_b04eed8, \9706 );
buf \U$labaj1842 ( R_282_b04ef80, \9716 );
buf \U$labaj1843 ( R_283_b04f028, \9726 );
buf \U$labaj1844 ( R_284_b04f0d0, \9736 );
buf \U$labaj1845 ( R_285_b04f178, \9746 );
buf \U$labaj1846 ( R_286_b04f220, \9756 );
buf \U$labaj1847 ( R_287_b04f2c8, \9768 );
buf \U$labaj1848 ( R_288_b04f370, \9774 );
buf \U$labaj1849 ( R_289_b04f418, \16490 );
buf \U$labaj1850 ( R_28a_b04f4c0, \16676 );
buf \U$labaj1851 ( R_28b_b04f568, \16768 );
buf \U$labaj1852 ( R_28c_b04f610, \16858 );
buf \U$labaj1853 ( R_28d_b04f6b8, \16904 );
buf \U$labaj1854 ( R_28e_b04f760, \16950 );
buf \U$labaj1855 ( R_28f_b04f808, \16994 );
buf \U$labaj1856 ( R_290_b04f8b0, \17038 );
buf \U$labaj1857 ( R_291_b04f958, \17062 );
buf \U$labaj1858 ( R_292_b04fa00, \17086 );
buf \U$labaj1859 ( R_293_b04faa8, \17110 );
buf \U$labaj1860 ( R_294_b04fb50, \17134 );
buf \U$labaj1861 ( R_295_b04fbf8, \17156 );
buf \U$labaj1862 ( R_296_b04fca0, \17178 );
buf \U$labaj1863 ( R_297_b04fd48, \17200 );
buf \U$labaj1864 ( R_298_b04fdf0, \17222 );
buf \U$labaj1865 ( R_299_b04fe98, \17232 );
buf \U$labaj1866 ( R_29a_b04ff40, \17242 );
buf \U$labaj1867 ( R_29b_b04ffe8, \17252 );
buf \U$labaj1868 ( R_29c_b050090, \17262 );
buf \U$labaj1869 ( R_29d_b050138, \17272 );
buf \U$labaj1870 ( R_29e_b0501e0, \17282 );
buf \U$labaj1871 ( R_29f_b050288, \17292 );
buf \U$labaj1872 ( R_2a0_b050330, \17302 );
buf \U$labaj1873 ( R_2a1_b0503d8, \17312 );
buf \U$labaj1874 ( R_2a2_b050480, \17322 );
buf \U$labaj1875 ( R_2a3_b050528, \17332 );
buf \U$labaj1876 ( R_2a4_b0505d0, \17342 );
buf \U$labaj1877 ( R_2a5_b050678, \17352 );
buf \U$labaj1878 ( R_2a6_b050720, \17362 );
buf \U$labaj1879 ( R_2a7_b0507c8, \17372 );
buf \U$labaj1880 ( R_2a8_b050870, \17382 );
buf \U$labaj1881 ( R_2a9_b050918, \17394 );
buf \U$labaj1882 ( R_2aa_b0509c0, \17400 );
buf \U$5 ( \2149 , RI2b5e785ebcf0_2);
buf \U$6 ( \2150 , RI2b5e785ebc78_3);
buf \U$7 ( \2151 , RI2b5e785ebc00_4);
buf \U$8 ( \2152 , RI2b5e785ebb88_5);
buf \U$9 ( \2153 , RI2b5e785ebb10_6);
buf \U$10 ( \2154 , RI2b5e785eba98_7);
buf \U$11 ( \2155 , RI2b5e785eba20_8);
buf \U$12 ( \2156 , RI2b5e785eb9a8_9);
buf \U$13 ( \2157 , RI2b5e785eb930_10);
buf \U$14 ( \2158 , RI2b5e785eb8b8_11);
buf \U$15 ( \2159 , RI2b5e785eb840_12);
and \U$16 ( \2160 , \2158 , \2159 );
and \U$17 ( \2161 , \2157 , \2160 );
and \U$18 ( \2162 , \2156 , \2161 );
and \U$19 ( \2163 , \2155 , \2162 );
and \U$20 ( \2164 , \2154 , \2163 );
and \U$21 ( \2165 , \2153 , \2164 );
and \U$22 ( \2166 , \2152 , \2165 );
and \U$23 ( \2167 , \2151 , \2166 );
and \U$24 ( \2168 , \2150 , \2167 );
xor \U$25 ( \2169 , \2149 , \2168 );
buf \U$26 ( \2170 , \2169 );
buf \U$27 ( \2171 , \2170 );
not \U$28 ( \2172 , RI2b5e785aeb98_596);
nor \U$29 ( \2173 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 , RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$30 ( \2174 , RI2b5e785daa40_28, \2173 );
not \U$31 ( \2175 , RI2b5e785ae9b8_600);
not \U$32 ( \2176 , RI2b5e785aea30_599);
not \U$33 ( \2177 , RI2b5e785aeaa8_598);
not \U$34 ( \2178 , RI2b5e785aeb20_597);
nor \U$35 ( \2179 , \2175 , \2176 , \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$36 ( \2180 , RI2b5e78549540_41, \2179 );
nor \U$37 ( \2181 , RI2b5e785ae9b8_600, \2176 , \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$38 ( \2182 , RI2b5e785388a8_54, \2181 );
nor \U$39 ( \2183 , \2175 , RI2b5e785aea30_599, \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$40 ( \2184 , RI2b5e784a6330_67, \2183 );
nor \U$41 ( \2185 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$42 ( \2186 , RI2b5e78495698_80, \2185 );
nor \U$43 ( \2187 , \2175 , \2176 , RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$44 ( \2188 , RI2b5e78495080_93, \2187 );
nor \U$45 ( \2189 , RI2b5e785ae9b8_600, \2176 , RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$46 ( \2190 , RI2b5e78403b80_106, \2189 );
nor \U$47 ( \2191 , \2175 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$48 ( \2192 , RI2b5e775b1e60_119, \2191 );
nor \U$49 ( \2193 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$50 ( \2194 , RI2b5e7750bdf8_132, \2193 );
nor \U$51 ( \2195 , \2175 , \2176 , \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$52 ( \2196 , RI2b5e774ff5d0_145, \2195 );
nor \U$53 ( \2197 , RI2b5e785ae9b8_600, \2176 , \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$54 ( \2198 , RI2b5e774f65e8_158, \2197 );
nor \U$55 ( \2199 , \2175 , RI2b5e785aea30_599, \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$56 ( \2200 , RI2b5e774eabd0_171, \2199 );
nor \U$57 ( \2201 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$58 ( \2202 , RI2b5e774de3a8_184, \2201 );
nor \U$59 ( \2203 , \2175 , \2176 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$60 ( \2204 , RI2b5e774d53c0_197, \2203 );
nor \U$61 ( \2205 , RI2b5e785ae9b8_600, \2176 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$62 ( \2206 , RI2b5e785f4300_210, \2205 );
nor \U$63 ( \2207 , \2175 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$64 ( \2208 , RI2b5e785f3ce8_223, \2207 );
nor \U$65 ( \2209 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$66 ( \2210 , RI2b5e785eb0c0_236, \2209 );
or \U$67 ( \2211 , \2174 , \2180 , \2182 , \2184 , \2186 , \2188 , \2190 , \2192 , \2194 , \2196 , \2198 , \2200 , \2202 , \2204 , \2206 , \2208 , \2210 );
buf \U$68 ( \2212 , RI2b5e785aec10_595);
buf \U$69 ( \2213 , RI2b5e785aec88_594);
buf \U$70 ( \2214 , RI2b5e785aed00_593);
buf \U$71 ( \2215 , RI2b5e785aed78_592);
buf \U$72 ( \2216 , RI2b5e785aedf0_591);
buf \U$73 ( \2217 , RI2b5e785aee68_590);
buf \U$74 ( \2218 , RI2b5e785aeee0_589);
buf \U$75 ( \2219 , RI2b5e785aef58_588);
buf \U$76 ( \2220 , RI2b5e785aeb98_596);
buf \U$77 ( \2221 , RI2b5e785ae9b8_600);
buf \U$78 ( \2222 , RI2b5e785aea30_599);
buf \U$79 ( \2223 , RI2b5e785aeaa8_598);
buf \U$80 ( \2224 , RI2b5e785aeb20_597);
or \U$81 ( \2225 , \2221 , \2222 , \2223 , \2224 );
and \U$82 ( \2226 , \2220 , \2225 );
or \U$83 ( \2227 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2226 );
buf \U$84 ( \2228 , \2227 );
_DC g2199 ( \2229_nG2199 , \2211 , \2228 );
buf \U$85 ( \2230 , \2229_nG2199 );
not \U$86 ( \2231 , \2230 );
xor \U$87 ( \2232 , \2171 , \2231 );
xor \U$88 ( \2233 , \2150 , \2167 );
buf \U$89 ( \2234 , \2233 );
buf \U$90 ( \2235 , \2234 );
and \U$91 ( \2236 , RI2b5e785da9c8_29, \2173 );
and \U$92 ( \2237 , RI2b5e785494c8_42, \2179 );
and \U$93 ( \2238 , RI2b5e78538830_55, \2181 );
and \U$94 ( \2239 , RI2b5e784a62b8_68, \2183 );
and \U$95 ( \2240 , RI2b5e78495620_81, \2185 );
and \U$96 ( \2241 , RI2b5e78495008_94, \2187 );
and \U$97 ( \2242 , RI2b5e78403b08_107, \2189 );
and \U$98 ( \2243 , RI2b5e775b1de8_120, \2191 );
and \U$99 ( \2244 , RI2b5e7750bd80_133, \2193 );
and \U$100 ( \2245 , RI2b5e774ff558_146, \2195 );
and \U$101 ( \2246 , RI2b5e774f6570_159, \2197 );
and \U$102 ( \2247 , RI2b5e774eab58_172, \2199 );
and \U$103 ( \2248 , RI2b5e774de330_185, \2201 );
and \U$104 ( \2249 , RI2b5e774d5348_198, \2203 );
and \U$105 ( \2250 , RI2b5e785f4288_211, \2205 );
and \U$106 ( \2251 , RI2b5e785f3658_224, \2207 );
and \U$107 ( \2252 , RI2b5e785eb048_237, \2209 );
or \U$108 ( \2253 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 );
_DC g2175 ( \2254_nG2175 , \2253 , \2228 );
buf \U$109 ( \2255 , \2254_nG2175 );
not \U$110 ( \2256 , \2255 );
and \U$111 ( \2257 , \2235 , \2256 );
xor \U$112 ( \2258 , \2151 , \2166 );
buf \U$113 ( \2259 , \2258 );
buf \U$114 ( \2260 , \2259 );
and \U$115 ( \2261 , RI2b5e785da950_30, \2173 );
and \U$116 ( \2262 , RI2b5e78549450_43, \2179 );
and \U$117 ( \2263 , RI2b5e785387b8_56, \2181 );
and \U$118 ( \2264 , RI2b5e784a6240_69, \2183 );
and \U$119 ( \2265 , RI2b5e784955a8_82, \2185 );
and \U$120 ( \2266 , RI2b5e78494f90_95, \2187 );
and \U$121 ( \2267 , RI2b5e78403a90_108, \2189 );
and \U$122 ( \2268 , RI2b5e775b1d70_121, \2191 );
and \U$123 ( \2269 , RI2b5e7750bd08_134, \2193 );
and \U$124 ( \2270 , RI2b5e774ff4e0_147, \2195 );
and \U$125 ( \2271 , RI2b5e774f64f8_160, \2197 );
and \U$126 ( \2272 , RI2b5e774eaae0_173, \2199 );
and \U$127 ( \2273 , RI2b5e774de2b8_186, \2201 );
and \U$128 ( \2274 , RI2b5e774d52d0_199, \2203 );
and \U$129 ( \2275 , RI2b5e785f4210_212, \2205 );
and \U$130 ( \2276 , RI2b5e785eb5e8_225, \2207 );
and \U$131 ( \2277 , RI2b5e785e6c50_238, \2209 );
or \U$132 ( \2278 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 );
_DC g1fee ( \2279_nG1fee , \2278 , \2228 );
buf \U$133 ( \2280 , \2279_nG1fee );
not \U$134 ( \2281 , \2280 );
and \U$135 ( \2282 , \2260 , \2281 );
xor \U$136 ( \2283 , \2152 , \2165 );
buf \U$137 ( \2284 , \2283 );
buf \U$138 ( \2285 , \2284 );
and \U$139 ( \2286 , RI2b5e785da8d8_31, \2173 );
and \U$140 ( \2287 , RI2b5e785493d8_44, \2179 );
and \U$141 ( \2288 , RI2b5e78538740_57, \2181 );
and \U$142 ( \2289 , RI2b5e784a61c8_70, \2183 );
and \U$143 ( \2290 , RI2b5e78495530_83, \2185 );
and \U$144 ( \2291 , RI2b5e78494f18_96, \2187 );
and \U$145 ( \2292 , RI2b5e78403a18_109, \2189 );
and \U$146 ( \2293 , RI2b5e775b1cf8_122, \2191 );
and \U$147 ( \2294 , RI2b5e7750bc90_135, \2193 );
and \U$148 ( \2295 , RI2b5e774ff468_148, \2195 );
and \U$149 ( \2296 , RI2b5e774f6480_161, \2197 );
and \U$150 ( \2297 , RI2b5e774eaa68_174, \2199 );
and \U$151 ( \2298 , RI2b5e774de240_187, \2201 );
and \U$152 ( \2299 , RI2b5e774d5258_200, \2203 );
and \U$153 ( \2300 , RI2b5e785f4198_213, \2205 );
and \U$154 ( \2301 , RI2b5e785eb570_226, \2207 );
and \U$155 ( \2302 , RI2b5e785e6bd8_239, \2209 );
or \U$156 ( \2303 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 );
_DC g1fca ( \2304_nG1fca , \2303 , \2228 );
buf \U$157 ( \2305 , \2304_nG1fca );
not \U$158 ( \2306 , \2305 );
and \U$159 ( \2307 , \2285 , \2306 );
xor \U$160 ( \2308 , \2153 , \2164 );
buf \U$161 ( \2309 , \2308 );
buf \U$162 ( \2310 , \2309 );
and \U$163 ( \2311 , RI2b5e785da860_32, \2173 );
and \U$164 ( \2312 , RI2b5e78549360_45, \2179 );
and \U$165 ( \2313 , RI2b5e785386c8_58, \2181 );
and \U$166 ( \2314 , RI2b5e784a6150_71, \2183 );
and \U$167 ( \2315 , RI2b5e784954b8_84, \2185 );
and \U$168 ( \2316 , RI2b5e78494ea0_97, \2187 );
and \U$169 ( \2317 , RI2b5e784039a0_110, \2189 );
and \U$170 ( \2318 , RI2b5e775b1c80_123, \2191 );
and \U$171 ( \2319 , RI2b5e7750bc18_136, \2193 );
and \U$172 ( \2320 , RI2b5e774ff3f0_149, \2195 );
and \U$173 ( \2321 , RI2b5e774f6408_162, \2197 );
and \U$174 ( \2322 , RI2b5e774ea9f0_175, \2199 );
and \U$175 ( \2323 , RI2b5e774de1c8_188, \2201 );
and \U$176 ( \2324 , RI2b5e774d51e0_201, \2203 );
and \U$177 ( \2325 , RI2b5e785f4120_214, \2205 );
and \U$178 ( \2326 , RI2b5e785eb4f8_227, \2207 );
and \U$179 ( \2327 , RI2b5e785e64d0_240, \2209 );
or \U$180 ( \2328 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 );
_DC g1e55 ( \2329_nG1e55 , \2328 , \2228 );
buf \U$181 ( \2330 , \2329_nG1e55 );
not \U$182 ( \2331 , \2330 );
and \U$183 ( \2332 , \2310 , \2331 );
xor \U$184 ( \2333 , \2154 , \2163 );
buf \U$185 ( \2334 , \2333 );
buf \U$186 ( \2335 , \2334 );
and \U$187 ( \2336 , RI2b5e78549900_33, \2173 );
and \U$188 ( \2337 , RI2b5e78538c68_46, \2179 );
and \U$189 ( \2338 , RI2b5e78538650_59, \2181 );
and \U$190 ( \2339 , RI2b5e784a60d8_72, \2183 );
and \U$191 ( \2340 , RI2b5e78495440_85, \2185 );
and \U$192 ( \2341 , RI2b5e78494e28_98, \2187 );
and \U$193 ( \2342 , RI2b5e78403928_111, \2189 );
and \U$194 ( \2343 , RI2b5e775b1c08_124, \2191 );
and \U$195 ( \2344 , RI2b5e7750bba0_137, \2193 );
and \U$196 ( \2345 , RI2b5e774ff378_150, \2195 );
and \U$197 ( \2346 , RI2b5e774f6390_163, \2197 );
and \U$198 ( \2347 , RI2b5e774ea978_176, \2199 );
and \U$199 ( \2348 , RI2b5e774de150_189, \2201 );
and \U$200 ( \2349 , RI2b5e774d5168_202, \2203 );
and \U$201 ( \2350 , RI2b5e785f40a8_215, \2205 );
and \U$202 ( \2351 , RI2b5e785eb480_228, \2207 );
and \U$203 ( \2352 , RI2b5e785da608_241, \2209 );
or \U$204 ( \2353 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 );
_DC g1e31 ( \2354_nG1e31 , \2353 , \2228 );
buf \U$205 ( \2355 , \2354_nG1e31 );
not \U$206 ( \2356 , \2355 );
and \U$207 ( \2357 , \2335 , \2356 );
xor \U$208 ( \2358 , \2155 , \2162 );
buf \U$209 ( \2359 , \2358 );
buf \U$210 ( \2360 , \2359 );
and \U$211 ( \2361 , RI2b5e78549888_34, \2173 );
and \U$212 ( \2362 , RI2b5e78538bf0_47, \2179 );
and \U$213 ( \2363 , RI2b5e785385d8_60, \2181 );
and \U$214 ( \2364 , RI2b5e784a6060_73, \2183 );
and \U$215 ( \2365 , RI2b5e784953c8_86, \2185 );
and \U$216 ( \2366 , RI2b5e78403ec8_99, \2187 );
and \U$217 ( \2367 , RI2b5e775b21a8_112, \2189 );
and \U$218 ( \2368 , RI2b5e775b1b90_125, \2191 );
and \U$219 ( \2369 , RI2b5e7750bb28_138, \2193 );
and \U$220 ( \2370 , RI2b5e774ff300_151, \2195 );
and \U$221 ( \2371 , RI2b5e774f6318_164, \2197 );
and \U$222 ( \2372 , RI2b5e774ea900_177, \2199 );
and \U$223 ( \2373 , RI2b5e774de0d8_190, \2201 );
and \U$224 ( \2374 , RI2b5e774d50f0_203, \2203 );
and \U$225 ( \2375 , RI2b5e785f4030_216, \2205 );
and \U$226 ( \2376 , RI2b5e785eb408_229, \2207 );
and \U$227 ( \2377 , RI2b5e785da590_242, \2209 );
or \U$228 ( \2378 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 );
_DC g1cf3 ( \2379_nG1cf3 , \2378 , \2228 );
buf \U$229 ( \2380 , \2379_nG1cf3 );
not \U$230 ( \2381 , \2380 );
and \U$231 ( \2382 , \2360 , \2381 );
xor \U$232 ( \2383 , \2156 , \2161 );
buf \U$233 ( \2384 , \2383 );
buf \U$234 ( \2385 , \2384 );
and \U$235 ( \2386 , RI2b5e78549810_35, \2173 );
and \U$236 ( \2387 , RI2b5e78538b78_48, \2179 );
and \U$237 ( \2388 , RI2b5e78538560_61, \2181 );
and \U$238 ( \2389 , RI2b5e784a5fe8_74, \2183 );
and \U$239 ( \2390 , RI2b5e78495350_87, \2185 );
and \U$240 ( \2391 , RI2b5e78403e50_100, \2187 );
and \U$241 ( \2392 , RI2b5e775b2130_113, \2189 );
and \U$242 ( \2393 , RI2b5e775b1b18_126, \2191 );
and \U$243 ( \2394 , RI2b5e7750bab0_139, \2193 );
and \U$244 ( \2395 , RI2b5e774ff288_152, \2195 );
and \U$245 ( \2396 , RI2b5e774f62a0_165, \2197 );
and \U$246 ( \2397 , RI2b5e774ea888_178, \2199 );
and \U$247 ( \2398 , RI2b5e774de060_191, \2201 );
and \U$248 ( \2399 , RI2b5e774d5078_204, \2203 );
and \U$249 ( \2400 , RI2b5e785f3fb8_217, \2205 );
and \U$250 ( \2401 , RI2b5e785eb390_230, \2207 );
and \U$251 ( \2402 , RI2b5e785da518_243, \2209 );
or \U$252 ( \2403 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 );
_DC g1ccf ( \2404_nG1ccf , \2403 , \2228 );
buf \U$253 ( \2405 , \2404_nG1ccf );
not \U$254 ( \2406 , \2405 );
and \U$255 ( \2407 , \2385 , \2406 );
xor \U$256 ( \2408 , \2157 , \2160 );
buf \U$257 ( \2409 , \2408 );
buf \U$258 ( \2410 , \2409 );
and \U$259 ( \2411 , RI2b5e78549798_36, \2173 );
and \U$260 ( \2412 , RI2b5e78538b00_49, \2179 );
and \U$261 ( \2413 , RI2b5e785384e8_62, \2181 );
and \U$262 ( \2414 , RI2b5e784a5f70_75, \2183 );
and \U$263 ( \2415 , RI2b5e784952d8_88, \2185 );
and \U$264 ( \2416 , RI2b5e78403dd8_101, \2187 );
and \U$265 ( \2417 , RI2b5e775b20b8_114, \2189 );
and \U$266 ( \2418 , RI2b5e775b1aa0_127, \2191 );
and \U$267 ( \2419 , RI2b5e7750ba38_140, \2193 );
and \U$268 ( \2420 , RI2b5e774ff210_153, \2195 );
and \U$269 ( \2421 , RI2b5e774f6228_166, \2197 );
and \U$270 ( \2422 , RI2b5e774ea810_179, \2199 );
and \U$271 ( \2423 , RI2b5e774ddfe8_192, \2201 );
and \U$272 ( \2424 , RI2b5e774d5000_205, \2203 );
and \U$273 ( \2425 , RI2b5e785f3f40_218, \2205 );
and \U$274 ( \2426 , RI2b5e785eb318_231, \2207 );
and \U$275 ( \2427 , RI2b5e785da4a0_244, \2209 );
or \U$276 ( \2428 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 );
_DC g1bc2 ( \2429_nG1bc2 , \2428 , \2228 );
buf \U$277 ( \2430 , \2429_nG1bc2 );
not \U$278 ( \2431 , \2430 );
and \U$279 ( \2432 , \2410 , \2431 );
xor \U$280 ( \2433 , \2158 , \2159 );
buf \U$281 ( \2434 , \2433 );
buf \U$282 ( \2435 , \2434 );
and \U$283 ( \2436 , RI2b5e78549720_37, \2173 );
and \U$284 ( \2437 , RI2b5e78538a88_50, \2179 );
and \U$285 ( \2438 , RI2b5e78538470_63, \2181 );
and \U$286 ( \2439 , RI2b5e784a5ef8_76, \2183 );
and \U$287 ( \2440 , RI2b5e78495260_89, \2185 );
and \U$288 ( \2441 , RI2b5e78403d60_102, \2187 );
and \U$289 ( \2442 , RI2b5e775b2040_115, \2189 );
and \U$290 ( \2443 , RI2b5e775b1a28_128, \2191 );
and \U$291 ( \2444 , RI2b5e7750b9c0_141, \2193 );
and \U$292 ( \2445 , RI2b5e774ff198_154, \2195 );
and \U$293 ( \2446 , RI2b5e774f61b0_167, \2197 );
and \U$294 ( \2447 , RI2b5e774ea798_180, \2199 );
and \U$295 ( \2448 , RI2b5e774ddf70_193, \2201 );
and \U$296 ( \2449 , RI2b5e774d4f88_206, \2203 );
and \U$297 ( \2450 , RI2b5e785f3ec8_219, \2205 );
and \U$298 ( \2451 , RI2b5e785eb2a0_232, \2207 );
and \U$299 ( \2452 , RI2b5e785da428_245, \2209 );
or \U$300 ( \2453 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 );
_DC g1bdb ( \2454_nG1bdb , \2453 , \2228 );
buf \U$301 ( \2455 , \2454_nG1bdb );
not \U$302 ( \2456 , \2455 );
and \U$303 ( \2457 , \2435 , \2456 );
not \U$304 ( \2458 , \2159 );
buf \U$305 ( \2459 , \2458 );
buf \U$306 ( \2460 , \2459 );
and \U$307 ( \2461 , RI2b5e785496a8_38, \2173 );
and \U$308 ( \2462 , RI2b5e78538a10_51, \2179 );
and \U$309 ( \2463 , RI2b5e785383f8_64, \2181 );
and \U$310 ( \2464 , RI2b5e784a5e80_77, \2183 );
and \U$311 ( \2465 , RI2b5e784951e8_90, \2185 );
and \U$312 ( \2466 , RI2b5e78403ce8_103, \2187 );
and \U$313 ( \2467 , RI2b5e775b1fc8_116, \2189 );
and \U$314 ( \2468 , RI2b5e775b19b0_129, \2191 );
and \U$315 ( \2469 , RI2b5e7750b948_142, \2193 );
and \U$316 ( \2470 , RI2b5e774ff120_155, \2195 );
and \U$317 ( \2471 , RI2b5e774f6138_168, \2197 );
and \U$318 ( \2472 , RI2b5e774ea720_181, \2199 );
and \U$319 ( \2473 , RI2b5e774ddef8_194, \2201 );
and \U$320 ( \2474 , RI2b5e774d4f10_207, \2203 );
and \U$321 ( \2475 , RI2b5e785f3e50_220, \2205 );
and \U$322 ( \2476 , RI2b5e785eb228_233, \2207 );
and \U$323 ( \2477 , RI2b5e785da3b0_246, \2209 );
or \U$324 ( \2478 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 );
_DC g1aa5 ( \2479_nG1aa5 , \2478 , \2228 );
buf \U$325 ( \2480 , \2479_nG1aa5 );
not \U$326 ( \2481 , \2480 );
and \U$327 ( \2482 , \2460 , \2481 );
buf \U$328 ( \2483 , RI2b5e785db148_13);
buf \U$331 ( \2484 , \2483 );
and \U$332 ( \2485 , RI2b5e78549630_39, \2173 );
and \U$333 ( \2486 , RI2b5e78538998_52, \2179 );
and \U$334 ( \2487 , RI2b5e78538380_65, \2181 );
and \U$335 ( \2488 , RI2b5e784a5e08_78, \2183 );
and \U$336 ( \2489 , RI2b5e78495170_91, \2185 );
and \U$337 ( \2490 , RI2b5e78403c70_104, \2187 );
and \U$338 ( \2491 , RI2b5e775b1f50_117, \2189 );
and \U$339 ( \2492 , RI2b5e775b1938_130, \2191 );
and \U$340 ( \2493 , RI2b5e7750b8d0_143, \2193 );
and \U$341 ( \2494 , RI2b5e774ff0a8_156, \2195 );
and \U$342 ( \2495 , RI2b5e774f60c0_169, \2197 );
and \U$343 ( \2496 , RI2b5e774ea6a8_182, \2199 );
and \U$344 ( \2497 , RI2b5e774dde80_195, \2201 );
and \U$345 ( \2498 , RI2b5e774d4e98_208, \2203 );
and \U$346 ( \2499 , RI2b5e785f3dd8_221, \2205 );
and \U$347 ( \2500 , RI2b5e785eb1b0_234, \2207 );
and \U$348 ( \2501 , RI2b5e785da338_247, \2209 );
or \U$349 ( \2502 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 );
_DC g1a89 ( \2503_nG1a89 , \2502 , \2228 );
buf \U$350 ( \2504 , \2503_nG1a89 );
not \U$351 ( \2505 , \2504 );
or \U$352 ( \2506 , \2484 , \2505 );
and \U$353 ( \2507 , \2481 , \2506 );
and \U$354 ( \2508 , \2460 , \2506 );
or \U$355 ( \2509 , \2482 , \2507 , \2508 );
and \U$356 ( \2510 , \2456 , \2509 );
and \U$357 ( \2511 , \2435 , \2509 );
or \U$358 ( \2512 , \2457 , \2510 , \2511 );
and \U$359 ( \2513 , \2431 , \2512 );
and \U$360 ( \2514 , \2410 , \2512 );
or \U$361 ( \2515 , \2432 , \2513 , \2514 );
and \U$362 ( \2516 , \2406 , \2515 );
and \U$363 ( \2517 , \2385 , \2515 );
or \U$364 ( \2518 , \2407 , \2516 , \2517 );
and \U$365 ( \2519 , \2381 , \2518 );
and \U$366 ( \2520 , \2360 , \2518 );
or \U$367 ( \2521 , \2382 , \2519 , \2520 );
and \U$368 ( \2522 , \2356 , \2521 );
and \U$369 ( \2523 , \2335 , \2521 );
or \U$370 ( \2524 , \2357 , \2522 , \2523 );
and \U$371 ( \2525 , \2331 , \2524 );
and \U$372 ( \2526 , \2310 , \2524 );
or \U$373 ( \2527 , \2332 , \2525 , \2526 );
and \U$374 ( \2528 , \2306 , \2527 );
and \U$375 ( \2529 , \2285 , \2527 );
or \U$376 ( \2530 , \2307 , \2528 , \2529 );
and \U$377 ( \2531 , \2281 , \2530 );
and \U$378 ( \2532 , \2260 , \2530 );
or \U$379 ( \2533 , \2282 , \2531 , \2532 );
and \U$380 ( \2534 , \2256 , \2533 );
and \U$381 ( \2535 , \2235 , \2533 );
or \U$382 ( \2536 , \2257 , \2534 , \2535 );
xor \U$383 ( \2537 , \2232 , \2536 );
buf g21a2_GF_PartitionCandidate( \2538_nG21a2 , \2537 );
buf \U$384 ( \2539 , \2538_nG21a2 );
xor \U$385 ( \2540 , \2235 , \2256 );
xor \U$386 ( \2541 , \2540 , \2533 );
buf g217e_GF_PartitionCandidate( \2542_nG217e , \2541 );
buf \U$387 ( \2543 , \2542_nG217e );
xor \U$388 ( \2544 , \2260 , \2281 );
xor \U$389 ( \2545 , \2544 , \2530 );
buf g1ff7_GF_PartitionCandidate( \2546_nG1ff7 , \2545 );
buf \U$390 ( \2547 , \2546_nG1ff7 );
and \U$391 ( \2548 , \2543 , \2547 );
not \U$392 ( \2549 , \2548 );
and \U$393 ( \2550 , \2539 , \2549 );
not \U$394 ( \2551 , \2550 );
buf \U$395 ( \2552 , RI2b5e785ae9b8_600);
buf \U$396 ( \2553 , RI2b5e785aec10_595);
buf \U$397 ( \2554 , RI2b5e785aec88_594);
buf \U$398 ( \2555 , RI2b5e785aed00_593);
buf \U$399 ( \2556 , RI2b5e785aed78_592);
buf \U$400 ( \2557 , RI2b5e785aedf0_591);
buf \U$401 ( \2558 , RI2b5e785aee68_590);
buf \U$402 ( \2559 , RI2b5e785aeee0_589);
buf \U$403 ( \2560 , RI2b5e785aef58_588);
buf \U$404 ( \2561 , RI2b5e785aeb98_596);
nor \U$405 ( \2562 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 );
buf \U$406 ( \2563 , \2562 );
buf \U$407 ( \2564 , \2563 );
xor \U$408 ( \2565 , \2552 , \2564 );
buf \U$409 ( \2566 , \2565 );
buf \U$410 ( \2567 , RI2b5e785aea30_599);
and \U$411 ( \2568 , \2552 , \2564 );
xor \U$412 ( \2569 , \2567 , \2568 );
buf \U$413 ( \2570 , \2569 );
buf \U$414 ( \2571 , RI2b5e785aeaa8_598);
and \U$415 ( \2572 , \2567 , \2568 );
xor \U$416 ( \2573 , \2571 , \2572 );
buf \U$417 ( \2574 , \2573 );
buf \U$418 ( \2575 , RI2b5e785aeb20_597);
and \U$419 ( \2576 , \2571 , \2572 );
xor \U$420 ( \2577 , \2575 , \2576 );
buf \U$421 ( \2578 , \2577 );
buf \U$422 ( \2579 , RI2b5e785aeb98_596);
and \U$423 ( \2580 , \2575 , \2576 );
xor \U$424 ( \2581 , \2579 , \2580 );
buf \U$425 ( \2582 , \2581 );
not \U$426 ( \2583 , \2582 );
buf \U$427 ( \2584 , RI2b5e785aec10_595);
and \U$428 ( \2585 , \2579 , \2580 );
xor \U$429 ( \2586 , \2584 , \2585 );
buf \U$430 ( \2587 , \2586 );
buf \U$431 ( \2588 , RI2b5e785aec88_594);
and \U$432 ( \2589 , \2584 , \2585 );
xor \U$433 ( \2590 , \2588 , \2589 );
buf \U$434 ( \2591 , \2590 );
buf \U$435 ( \2592 , RI2b5e785aed00_593);
and \U$436 ( \2593 , \2588 , \2589 );
xor \U$437 ( \2594 , \2592 , \2593 );
buf \U$438 ( \2595 , \2594 );
buf \U$439 ( \2596 , RI2b5e785aed78_592);
and \U$440 ( \2597 , \2592 , \2593 );
xor \U$441 ( \2598 , \2596 , \2597 );
buf \U$442 ( \2599 , \2598 );
buf \U$443 ( \2600 , RI2b5e785aedf0_591);
and \U$444 ( \2601 , \2596 , \2597 );
xor \U$445 ( \2602 , \2600 , \2601 );
buf \U$446 ( \2603 , \2602 );
buf \U$447 ( \2604 , RI2b5e785aee68_590);
and \U$448 ( \2605 , \2600 , \2601 );
xor \U$449 ( \2606 , \2604 , \2605 );
buf \U$450 ( \2607 , \2606 );
buf \U$451 ( \2608 , RI2b5e785aeee0_589);
and \U$452 ( \2609 , \2604 , \2605 );
xor \U$453 ( \2610 , \2608 , \2609 );
buf \U$454 ( \2611 , \2610 );
buf \U$455 ( \2612 , RI2b5e785aef58_588);
and \U$456 ( \2613 , \2608 , \2609 );
xor \U$457 ( \2614 , \2612 , \2613 );
buf \U$458 ( \2615 , \2614 );
nor \U$459 ( \2616 , \2566 , \2570 , \2574 , \2578 , \2583 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$460 ( \2617 , RI2b5e785da248_249, \2616 );
not \U$461 ( \2618 , \2566 );
not \U$462 ( \2619 , \2570 );
not \U$463 ( \2620 , \2574 );
not \U$464 ( \2621 , \2578 );
nor \U$465 ( \2622 , \2618 , \2619 , \2620 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$466 ( \2623 , RI2b5e785be750_269, \2622 );
nor \U$467 ( \2624 , \2566 , \2619 , \2620 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$468 ( \2625 , RI2b5e785bc4a0_289, \2624 );
nor \U$469 ( \2626 , \2618 , \2570 , \2620 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$470 ( \2627 , RI2b5e785bbb40_309, \2626 );
nor \U$471 ( \2628 , \2566 , \2570 , \2620 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$472 ( \2629 , RI2b5e785b9c50_329, \2628 );
nor \U$473 ( \2630 , \2618 , \2619 , \2574 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$474 ( \2631 , RI2b5e785b8120_349, \2630 );
nor \U$475 ( \2632 , \2566 , \2619 , \2574 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$476 ( \2633 , RI2b5e785b77c0_369, \2632 );
nor \U$477 ( \2634 , \2618 , \2570 , \2574 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$478 ( \2635 , RI2b5e785b6e60_389, \2634 );
nor \U$479 ( \2636 , \2566 , \2570 , \2574 , \2621 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$480 ( \2637 , RI2b5e785b56f0_409, \2636 );
nor \U$481 ( \2638 , \2618 , \2619 , \2620 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$482 ( \2639 , RI2b5e785b4d90_429, \2638 );
nor \U$483 ( \2640 , \2566 , \2619 , \2620 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$484 ( \2641 , RI2b5e785b39e0_449, \2640 );
nor \U$485 ( \2642 , \2618 , \2570 , \2620 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$486 ( \2643 , RI2b5e785b3080_469, \2642 );
nor \U$487 ( \2644 , \2566 , \2570 , \2620 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$488 ( \2645 , RI2b5e785b2720_489, \2644 );
nor \U$489 ( \2646 , \2618 , \2619 , \2574 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$490 ( \2647 , RI2b5e785b1730_509, \2646 );
nor \U$491 ( \2648 , \2566 , \2619 , \2574 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$492 ( \2649 , RI2b5e785b0dd0_529, \2648 );
nor \U$493 ( \2650 , \2618 , \2570 , \2574 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$494 ( \2651 , RI2b5e785b0470_549, \2650 );
nor \U$495 ( \2652 , \2566 , \2570 , \2574 , \2578 , \2582 , \2587 , \2591 , \2595 , \2599 , \2603 , \2607 , \2611 , \2615 );
and \U$496 ( \2653 , RI2b5e785af840_569, \2652 );
or \U$497 ( \2654 , \2617 , \2623 , \2625 , \2627 , \2629 , \2631 , \2633 , \2635 , \2637 , \2639 , \2641 , \2643 , \2645 , \2647 , \2649 , \2651 , \2653 );
buf \U$498 ( \2655 , \2587 );
buf \U$499 ( \2656 , \2591 );
buf \U$500 ( \2657 , \2595 );
buf \U$501 ( \2658 , \2599 );
buf \U$502 ( \2659 , \2603 );
buf \U$503 ( \2660 , \2607 );
buf \U$504 ( \2661 , \2611 );
buf \U$505 ( \2662 , \2615 );
buf \U$506 ( \2663 , \2582 );
buf \U$507 ( \2664 , \2566 );
buf \U$508 ( \2665 , \2570 );
buf \U$509 ( \2666 , \2574 );
buf \U$510 ( \2667 , \2578 );
or \U$511 ( \2668 , \2664 , \2665 , \2666 , \2667 );
and \U$512 ( \2669 , \2663 , \2668 );
or \U$513 ( \2670 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2669 );
buf \U$514 ( \2671 , \2670 );
_DC g2899 ( \2672_nG2899 , \2654 , \2671 );
buf \U$515 ( \2673 , \2672_nG2899 );
buf \U$516 ( \2674 , RI2b5e785ebd68_1);
and \U$517 ( \2675 , \2149 , \2168 );
and \U$518 ( \2676 , \2674 , \2675 );
buf \U$519 ( \2677 , \2676 );
buf \U$520 ( \2678 , \2677 );
xor \U$521 ( \2679 , \2674 , \2675 );
buf \U$522 ( \2680 , \2679 );
buf \U$523 ( \2681 , \2680 );
and \U$524 ( \2682 , RI2b5e785daab8_27, \2173 );
and \U$525 ( \2683 , RI2b5e785495b8_40, \2179 );
and \U$526 ( \2684 , RI2b5e78538920_53, \2181 );
and \U$527 ( \2685 , RI2b5e784a63a8_66, \2183 );
and \U$528 ( \2686 , RI2b5e78495710_79, \2185 );
and \U$529 ( \2687 , RI2b5e784950f8_92, \2187 );
and \U$530 ( \2688 , RI2b5e78403bf8_105, \2189 );
and \U$531 ( \2689 , RI2b5e775b1ed8_118, \2191 );
and \U$532 ( \2690 , RI2b5e775b18c0_131, \2193 );
and \U$533 ( \2691 , RI2b5e7750b858_144, \2195 );
and \U$534 ( \2692 , RI2b5e774ff030_157, \2197 );
and \U$535 ( \2693 , RI2b5e774f6048_170, \2199 );
and \U$536 ( \2694 , RI2b5e774ea630_183, \2201 );
and \U$537 ( \2695 , RI2b5e774dde08_196, \2203 );
and \U$538 ( \2696 , RI2b5e774d4e20_209, \2205 );
and \U$539 ( \2697 , RI2b5e785f3d60_222, \2207 );
and \U$540 ( \2698 , RI2b5e785eb138_235, \2209 );
or \U$541 ( \2699 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 );
_DC g2361 ( \2700_nG2361 , \2699 , \2228 );
buf \U$542 ( \2701 , \2700_nG2361 );
not \U$543 ( \2702 , \2701 );
and \U$544 ( \2703 , \2681 , \2702 );
and \U$545 ( \2704 , \2171 , \2231 );
and \U$546 ( \2705 , \2231 , \2536 );
and \U$547 ( \2706 , \2171 , \2536 );
or \U$548 ( \2707 , \2704 , \2705 , \2706 );
and \U$549 ( \2708 , \2702 , \2707 );
and \U$550 ( \2709 , \2681 , \2707 );
or \U$551 ( \2710 , \2703 , \2708 , \2709 );
xnor \U$552 ( \2711 , \2678 , \2710 );
buf g2376_GF_PartitionCandidate( \2712_nG2376 , \2711 );
buf \U$553 ( \2713 , \2712_nG2376 );
xor \U$554 ( \2714 , \2681 , \2702 );
xor \U$555 ( \2715 , \2714 , \2707 );
buf g236a_GF_PartitionCandidate( \2716_nG236a , \2715 );
buf \U$556 ( \2717 , \2716_nG236a );
xor \U$557 ( \2718 , \2713 , \2717 );
xor \U$558 ( \2719 , \2717 , \2539 );
not \U$559 ( \2720 , \2719 );
and \U$560 ( \2721 , \2718 , \2720 );
and \U$561 ( \2722 , \2673 , \2721 );
and \U$562 ( \2723 , RI2b5e785da2c0_248, \2616 );
and \U$563 ( \2724 , RI2b5e785be7c8_268, \2622 );
and \U$564 ( \2725 , RI2b5e785bc518_288, \2624 );
and \U$565 ( \2726 , RI2b5e785bbbb8_308, \2626 );
and \U$566 ( \2727 , RI2b5e785b9cc8_328, \2628 );
and \U$567 ( \2728 , RI2b5e785b9368_348, \2630 );
and \U$568 ( \2729 , RI2b5e785b7838_368, \2632 );
and \U$569 ( \2730 , RI2b5e785b6ed8_388, \2634 );
and \U$570 ( \2731 , RI2b5e785b5768_408, \2636 );
and \U$571 ( \2732 , RI2b5e785b4e08_428, \2638 );
and \U$572 ( \2733 , RI2b5e785b3a58_448, \2640 );
and \U$573 ( \2734 , RI2b5e785b30f8_468, \2642 );
and \U$574 ( \2735 , RI2b5e785b2798_488, \2644 );
and \U$575 ( \2736 , RI2b5e785b17a8_508, \2646 );
and \U$576 ( \2737 , RI2b5e785b0e48_528, \2648 );
and \U$577 ( \2738 , RI2b5e785b04e8_548, \2650 );
and \U$578 ( \2739 , RI2b5e785afb88_568, \2652 );
or \U$579 ( \2740 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 );
_DC g298d ( \2741_nG298d , \2740 , \2671 );
buf \U$580 ( \2742 , \2741_nG298d );
and \U$581 ( \2743 , \2742 , \2719 );
nor \U$582 ( \2744 , \2722 , \2743 );
and \U$583 ( \2745 , \2717 , \2539 );
not \U$584 ( \2746 , \2745 );
and \U$585 ( \2747 , \2713 , \2746 );
xnor \U$586 ( \2748 , \2744 , \2747 );
xor \U$587 ( \2749 , \2551 , \2748 );
and \U$589 ( \2750 , RI2b5e785da1d0_250, \2616 );
and \U$590 ( \2751 , RI2b5e785be6d8_270, \2622 );
and \U$591 ( \2752 , RI2b5e785bc428_290, \2624 );
and \U$592 ( \2753 , RI2b5e785bbac8_310, \2626 );
and \U$593 ( \2754 , RI2b5e785b9bd8_330, \2628 );
and \U$594 ( \2755 , RI2b5e785b80a8_350, \2630 );
and \U$595 ( \2756 , RI2b5e785b7748_370, \2632 );
and \U$596 ( \2757 , RI2b5e785b6de8_390, \2634 );
and \U$597 ( \2758 , RI2b5e785b5678_410, \2636 );
and \U$598 ( \2759 , RI2b5e785b4d18_430, \2638 );
and \U$599 ( \2760 , RI2b5e785b3968_450, \2640 );
and \U$600 ( \2761 , RI2b5e785b3008_470, \2642 );
and \U$601 ( \2762 , RI2b5e785b26a8_490, \2644 );
and \U$602 ( \2763 , RI2b5e785b16b8_510, \2646 );
and \U$603 ( \2764 , RI2b5e785b0d58_530, \2648 );
and \U$604 ( \2765 , RI2b5e785b03f8_550, \2650 );
and \U$605 ( \2766 , RI2b5e785af7c8_570, \2652 );
or \U$606 ( \2767 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 );
_DC g27d7 ( \2768_nG27d7 , \2767 , \2671 );
buf \U$607 ( \2769 , \2768_nG27d7 );
or \U$608 ( \2770 , \2678 , \2710 );
not \U$609 ( \2771 , \2770 );
buf g2572_GF_PartitionCandidate( \2772_nG2572 , \2771 );
buf \U$610 ( \2773 , \2772_nG2572 );
xor \U$611 ( \2774 , \2773 , \2713 );
and \U$612 ( \2775 , \2769 , \2774 );
nor \U$613 ( \2776 , 1'b0 , \2775 );
xnor \U$615 ( \2777 , \2776 , 1'b0 );
xor \U$616 ( \2778 , \2749 , \2777 );
xor \U$617 ( \2779 , 1'b0 , \2778 );
xor \U$619 ( \2780 , \2539 , \2543 );
xor \U$620 ( \2781 , \2543 , \2547 );
not \U$621 ( \2782 , \2781 );
and \U$622 ( \2783 , \2780 , \2782 );
and \U$623 ( \2784 , \2742 , \2783 );
not \U$624 ( \2785 , \2784 );
xnor \U$625 ( \2786 , \2785 , \2550 );
and \U$626 ( \2787 , \2769 , \2721 );
and \U$627 ( \2788 , \2673 , \2719 );
nor \U$628 ( \2789 , \2787 , \2788 );
xnor \U$629 ( \2790 , \2789 , \2747 );
and \U$630 ( \2791 , \2786 , \2790 );
or \U$632 ( \2792 , 1'b0 , \2791 , 1'b0 );
xor \U$634 ( \2793 , \2792 , 1'b0 );
xor \U$636 ( \2794 , \2793 , 1'b0 );
and \U$637 ( \2795 , \2779 , \2794 );
or \U$638 ( \2796 , 1'b0 , 1'b0 , \2795 );
and \U$641 ( \2797 , \2742 , \2721 );
not \U$642 ( \2798 , \2797 );
xnor \U$643 ( \2799 , \2798 , \2747 );
xor \U$644 ( \2800 , 1'b0 , \2799 );
and \U$646 ( \2801 , \2673 , \2774 );
nor \U$647 ( \2802 , 1'b0 , \2801 );
xnor \U$648 ( \2803 , \2802 , 1'b0 );
xor \U$649 ( \2804 , \2800 , \2803 );
xor \U$650 ( \2805 , 1'b0 , \2804 );
xor \U$652 ( \2806 , \2805 , 1'b1 );
and \U$653 ( \2807 , \2551 , \2748 );
and \U$654 ( \2808 , \2748 , \2777 );
and \U$655 ( \2809 , \2551 , \2777 );
or \U$656 ( \2810 , \2807 , \2808 , \2809 );
xor \U$658 ( \2811 , \2810 , 1'b0 );
xor \U$660 ( \2812 , \2811 , 1'b0 );
xor \U$661 ( \2813 , \2806 , \2812 );
and \U$662 ( \2814 , \2796 , \2813 );
or \U$664 ( \2815 , 1'b0 , \2814 , 1'b0 );
xor \U$666 ( \2816 , \2815 , 1'b0 );
and \U$668 ( \2817 , \2805 , 1'b1 );
and \U$669 ( \2818 , 1'b1 , \2812 );
and \U$670 ( \2819 , \2805 , \2812 );
or \U$671 ( \2820 , \2817 , \2818 , \2819 );
xor \U$672 ( \2821 , 1'b0 , \2820 );
not \U$674 ( \2822 , \2747 );
and \U$676 ( \2823 , \2742 , \2774 );
nor \U$677 ( \2824 , 1'b0 , \2823 );
xnor \U$678 ( \2825 , \2824 , 1'b0 );
xor \U$679 ( \2826 , \2822 , \2825 );
xor \U$681 ( \2827 , \2826 , 1'b0 );
xor \U$682 ( \2828 , 1'b0 , \2827 );
xor \U$684 ( \2829 , \2828 , 1'b0 );
and \U$686 ( \2830 , \2799 , \2803 );
or \U$688 ( \2831 , 1'b0 , \2830 , 1'b0 );
xor \U$690 ( \2832 , \2831 , 1'b0 );
xor \U$692 ( \2833 , \2832 , 1'b0 );
xor \U$693 ( \2834 , \2829 , \2833 );
xor \U$694 ( \2835 , \2821 , \2834 );
xor \U$695 ( \2836 , \2816 , \2835 );
xor \U$701 ( \2837 , \2285 , \2306 );
xor \U$702 ( \2838 , \2837 , \2527 );
buf g1fd3_GF_PartitionCandidate( \2839_nG1fd3 , \2838 );
buf \U$703 ( \2840 , \2839_nG1fd3 );
xor \U$704 ( \2841 , \2547 , \2840 );
xor \U$705 ( \2842 , \2310 , \2331 );
xor \U$706 ( \2843 , \2842 , \2524 );
buf g1e5e_GF_PartitionCandidate( \2844_nG1e5e , \2843 );
buf \U$707 ( \2845 , \2844_nG1e5e );
xor \U$708 ( \2846 , \2840 , \2845 );
not \U$709 ( \2847 , \2846 );
and \U$710 ( \2848 , \2841 , \2847 );
and \U$711 ( \2849 , \2742 , \2848 );
not \U$712 ( \2850 , \2849 );
and \U$713 ( \2851 , \2840 , \2845 );
not \U$714 ( \2852 , \2851 );
and \U$715 ( \2853 , \2547 , \2852 );
xnor \U$716 ( \2854 , \2850 , \2853 );
and \U$717 ( \2855 , \2769 , \2783 );
and \U$718 ( \2856 , \2673 , \2781 );
nor \U$719 ( \2857 , \2855 , \2856 );
xnor \U$720 ( \2858 , \2857 , \2550 );
and \U$721 ( \2859 , \2854 , \2858 );
or \U$723 ( \2860 , 1'b0 , \2859 , 1'b0 );
and \U$724 ( \2861 , RI2b5e785da0e0_252, \2616 );
and \U$725 ( \2862 , RI2b5e785be5e8_272, \2622 );
and \U$726 ( \2863 , RI2b5e785bc338_292, \2624 );
and \U$727 ( \2864 , RI2b5e785bb9d8_312, \2626 );
and \U$728 ( \2865 , RI2b5e785b9ae8_332, \2628 );
and \U$729 ( \2866 , RI2b5e785b7fb8_352, \2630 );
and \U$730 ( \2867 , RI2b5e785b7658_372, \2632 );
and \U$731 ( \2868 , RI2b5e785b5ee8_392, \2634 );
and \U$732 ( \2869 , RI2b5e785b5588_412, \2636 );
and \U$733 ( \2870 , RI2b5e785b4c28_432, \2638 );
and \U$734 ( \2871 , RI2b5e785b3878_452, \2640 );
and \U$735 ( \2872 , RI2b5e785b2f18_472, \2642 );
and \U$736 ( \2873 , RI2b5e785b25b8_492, \2644 );
and \U$737 ( \2874 , RI2b5e785b15c8_512, \2646 );
and \U$738 ( \2875 , RI2b5e785b0c68_532, \2648 );
and \U$739 ( \2876 , RI2b5e785b0308_552, \2650 );
and \U$740 ( \2877 , RI2b5e785af6d8_572, \2652 );
or \U$741 ( \2878 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 );
_DC g263c ( \2879_nG263c , \2878 , \2671 );
buf \U$742 ( \2880 , \2879_nG263c );
and \U$743 ( \2881 , \2880 , \2721 );
and \U$744 ( \2882 , RI2b5e785da158_251, \2616 );
and \U$745 ( \2883 , RI2b5e785be660_271, \2622 );
and \U$746 ( \2884 , RI2b5e785bc3b0_291, \2624 );
and \U$747 ( \2885 , RI2b5e785bba50_311, \2626 );
and \U$748 ( \2886 , RI2b5e785b9b60_331, \2628 );
and \U$749 ( \2887 , RI2b5e785b8030_351, \2630 );
and \U$750 ( \2888 , RI2b5e785b76d0_371, \2632 );
and \U$751 ( \2889 , RI2b5e785b6d70_391, \2634 );
and \U$752 ( \2890 , RI2b5e785b5600_411, \2636 );
and \U$753 ( \2891 , RI2b5e785b4ca0_431, \2638 );
and \U$754 ( \2892 , RI2b5e785b38f0_451, \2640 );
and \U$755 ( \2893 , RI2b5e785b2f90_471, \2642 );
and \U$756 ( \2894 , RI2b5e785b2630_491, \2644 );
and \U$757 ( \2895 , RI2b5e785b1640_511, \2646 );
and \U$758 ( \2896 , RI2b5e785b0ce0_531, \2648 );
and \U$759 ( \2897 , RI2b5e785b0380_551, \2650 );
and \U$760 ( \2898 , RI2b5e785af750_571, \2652 );
or \U$761 ( \2899 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 );
_DC g2716 ( \2900_nG2716 , \2899 , \2671 );
buf \U$762 ( \2901 , \2900_nG2716 );
and \U$763 ( \2902 , \2901 , \2719 );
nor \U$764 ( \2903 , \2881 , \2902 );
xnor \U$765 ( \2904 , \2903 , \2747 );
and \U$767 ( \2905 , RI2b5e785da068_253, \2616 );
and \U$768 ( \2906 , RI2b5e785be570_273, \2622 );
and \U$769 ( \2907 , RI2b5e785bc2c0_293, \2624 );
and \U$770 ( \2908 , RI2b5e785bb960_313, \2626 );
and \U$771 ( \2909 , RI2b5e785b9a70_333, \2628 );
and \U$772 ( \2910 , RI2b5e785b7f40_353, \2630 );
and \U$773 ( \2911 , RI2b5e785b75e0_373, \2632 );
and \U$774 ( \2912 , RI2b5e785b5e70_393, \2634 );
and \U$775 ( \2913 , RI2b5e785b5510_413, \2636 );
and \U$776 ( \2914 , RI2b5e785b4bb0_433, \2638 );
and \U$777 ( \2915 , RI2b5e785b3800_453, \2640 );
and \U$778 ( \2916 , RI2b5e785b2ea0_473, \2642 );
and \U$779 ( \2917 , RI2b5e785b2540_493, \2644 );
and \U$780 ( \2918 , RI2b5e785b1550_513, \2646 );
and \U$781 ( \2919 , RI2b5e785b0bf0_533, \2648 );
and \U$782 ( \2920 , RI2b5e785b0290_553, \2650 );
and \U$783 ( \2921 , RI2b5e785af660_573, \2652 );
or \U$784 ( \2922 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 );
_DC g2551 ( \2923_nG2551 , \2922 , \2671 );
buf \U$785 ( \2924 , \2923_nG2551 );
and \U$786 ( \2925 , \2924 , \2774 );
nor \U$787 ( \2926 , 1'b0 , \2925 );
xnor \U$788 ( \2927 , \2926 , 1'b0 );
and \U$789 ( \2928 , \2904 , \2927 );
or \U$792 ( \2929 , \2928 , 1'b0 , 1'b0 );
and \U$793 ( \2930 , \2860 , \2929 );
or \U$796 ( \2931 , \2930 , 1'b0 , 1'b0 );
and \U$799 ( \2932 , \2880 , \2774 );
nor \U$800 ( \2933 , 1'b0 , \2932 );
xnor \U$801 ( \2934 , \2933 , 1'b0 );
xor \U$803 ( \2935 , \2934 , 1'b0 );
xor \U$805 ( \2936 , \2935 , 1'b0 );
not \U$806 ( \2937 , \2853 );
and \U$807 ( \2938 , \2673 , \2783 );
and \U$808 ( \2939 , \2742 , \2781 );
nor \U$809 ( \2940 , \2938 , \2939 );
xnor \U$810 ( \2941 , \2940 , \2550 );
xor \U$811 ( \2942 , \2937 , \2941 );
and \U$812 ( \2943 , \2901 , \2721 );
and \U$813 ( \2944 , \2769 , \2719 );
nor \U$814 ( \2945 , \2943 , \2944 );
xnor \U$815 ( \2946 , \2945 , \2747 );
xor \U$816 ( \2947 , \2942 , \2946 );
and \U$817 ( \2948 , \2936 , \2947 );
or \U$819 ( \2949 , 1'b0 , \2948 , 1'b0 );
and \U$820 ( \2950 , \2931 , \2949 );
or \U$821 ( \2951 , 1'b0 , 1'b0 , \2950 );
and \U$823 ( \2952 , \2901 , \2774 );
nor \U$824 ( \2953 , 1'b0 , \2952 );
xnor \U$825 ( \2954 , \2953 , 1'b0 );
xor \U$827 ( \2955 , \2954 , 1'b0 );
xor \U$829 ( \2956 , \2955 , 1'b0 );
xor \U$831 ( \2957 , 1'b0 , \2786 );
xor \U$832 ( \2958 , \2957 , \2790 );
xor \U$833 ( \2959 , \2956 , \2958 );
and \U$835 ( \2960 , \2959 , 1'b1 );
and \U$836 ( \2961 , \2937 , \2941 );
and \U$837 ( \2962 , \2941 , \2946 );
and \U$838 ( \2963 , \2937 , \2946 );
or \U$839 ( \2964 , \2961 , \2962 , \2963 );
xor \U$841 ( \2965 , \2964 , 1'b0 );
xor \U$843 ( \2966 , \2965 , 1'b0 );
and \U$844 ( \2967 , 1'b1 , \2966 );
and \U$845 ( \2968 , \2959 , \2966 );
or \U$846 ( \2969 , \2960 , \2967 , \2968 );
and \U$847 ( \2970 , \2951 , \2969 );
xor \U$849 ( \2971 , \2779 , 1'b0 );
xor \U$850 ( \2972 , \2971 , \2794 );
and \U$851 ( \2973 , \2969 , \2972 );
and \U$852 ( \2974 , \2951 , \2972 );
or \U$853 ( \2975 , \2970 , \2973 , \2974 );
xor \U$855 ( \2976 , 1'b0 , \2796 );
xor \U$856 ( \2977 , \2976 , \2813 );
and \U$857 ( \2978 , \2975 , \2977 );
or \U$858 ( \2979 , 1'b0 , 1'b0 , \2978 );
nand \U$859 ( \2980 , \2836 , \2979 );
nor \U$860 ( \2981 , \2836 , \2979 );
not \U$861 ( \2982 , \2981 );
nand \U$862 ( \2983 , \2980 , \2982 );
xor \U$863 ( \2984 , \2460 , \2481 );
xor \U$864 ( \2985 , \2984 , \2506 );
buf g1aac_GF_PartitionCandidate( \2986_nG1aac , \2985 );
buf \U$865 ( \2987 , \2986_nG1aac );
xor \U$866 ( \2988 , \2484 , \2504 );
buf g1a8c_GF_PartitionCandidate( \2989_nG1a8c , \2988 );
buf \U$867 ( \2990 , \2989_nG1a8c );
xor \U$868 ( \2991 , \2987 , \2990 );
not \U$869 ( \2992 , \2990 );
and \U$870 ( \2993 , \2991 , \2992 );
and \U$871 ( \2994 , \2924 , \2993 );
and \U$872 ( \2995 , \2880 , \2990 );
nor \U$873 ( \2996 , \2994 , \2995 );
xnor \U$874 ( \2997 , \2996 , \2987 );
and \U$875 ( \2998 , RI2b5e785c2bc0_255, \2616 );
and \U$876 ( \2999 , RI2b5e785be480_275, \2622 );
and \U$877 ( \3000 , RI2b5e785bc1d0_295, \2624 );
and \U$878 ( \3001 , RI2b5e785ba2e0_315, \2626 );
and \U$879 ( \3002 , RI2b5e785b9980_335, \2628 );
and \U$880 ( \3003 , RI2b5e785b7e50_355, \2630 );
and \U$881 ( \3004 , RI2b5e785b74f0_375, \2632 );
and \U$882 ( \3005 , RI2b5e785b5d80_395, \2634 );
and \U$883 ( \3006 , RI2b5e785b5420_415, \2636 );
and \U$884 ( \3007 , RI2b5e785b4ac0_435, \2638 );
and \U$885 ( \3008 , RI2b5e785b3710_455, \2640 );
and \U$886 ( \3009 , RI2b5e785b2db0_475, \2642 );
and \U$887 ( \3010 , RI2b5e785b2450_495, \2644 );
and \U$888 ( \3011 , RI2b5e785b1460_515, \2646 );
and \U$889 ( \3012 , RI2b5e785b0b00_535, \2648 );
and \U$890 ( \3013 , RI2b5e785b01a0_555, \2650 );
and \U$891 ( \3014 , RI2b5e785af570_575, \2652 );
or \U$892 ( \3015 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 );
_DC g239e ( \3016_nG239e , \3015 , \2671 );
buf \U$893 ( \3017 , \3016_nG239e );
xor \U$894 ( \3018 , \2410 , \2431 );
xor \U$895 ( \3019 , \3018 , \2512 );
buf g1be7_GF_PartitionCandidate( \3020_nG1be7 , \3019 );
buf \U$896 ( \3021 , \3020_nG1be7 );
xor \U$897 ( \3022 , \2435 , \2456 );
xor \U$898 ( \3023 , \3022 , \2509 );
buf g1beb_GF_PartitionCandidate( \3024_nG1beb , \3023 );
buf \U$899 ( \3025 , \3024_nG1beb );
xor \U$900 ( \3026 , \3021 , \3025 );
xor \U$901 ( \3027 , \3025 , \2987 );
not \U$902 ( \3028 , \3027 );
and \U$903 ( \3029 , \3026 , \3028 );
and \U$904 ( \3030 , \3017 , \3029 );
and \U$905 ( \3031 , RI2b5e785c2c38_254, \2616 );
and \U$906 ( \3032 , RI2b5e785be4f8_274, \2622 );
and \U$907 ( \3033 , RI2b5e785bc248_294, \2624 );
and \U$908 ( \3034 , RI2b5e785ba358_314, \2626 );
and \U$909 ( \3035 , RI2b5e785b99f8_334, \2628 );
and \U$910 ( \3036 , RI2b5e785b7ec8_354, \2630 );
and \U$911 ( \3037 , RI2b5e785b7568_374, \2632 );
and \U$912 ( \3038 , RI2b5e785b5df8_394, \2634 );
and \U$913 ( \3039 , RI2b5e785b5498_414, \2636 );
and \U$914 ( \3040 , RI2b5e785b4b38_434, \2638 );
and \U$915 ( \3041 , RI2b5e785b3788_454, \2640 );
and \U$916 ( \3042 , RI2b5e785b2e28_474, \2642 );
and \U$917 ( \3043 , RI2b5e785b24c8_494, \2644 );
and \U$918 ( \3044 , RI2b5e785b14d8_514, \2646 );
and \U$919 ( \3045 , RI2b5e785b0b78_534, \2648 );
and \U$920 ( \3046 , RI2b5e785b0218_554, \2650 );
and \U$921 ( \3047 , RI2b5e785af5e8_574, \2652 );
or \U$922 ( \3048 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 );
_DC g2472 ( \3049_nG2472 , \3048 , \2671 );
buf \U$923 ( \3050 , \3049_nG2472 );
and \U$924 ( \3051 , \3050 , \3027 );
nor \U$925 ( \3052 , \3030 , \3051 );
and \U$926 ( \3053 , \3025 , \2987 );
not \U$927 ( \3054 , \3053 );
and \U$928 ( \3055 , \3021 , \3054 );
xnor \U$929 ( \3056 , \3052 , \3055 );
and \U$930 ( \3057 , \2997 , \3056 );
and \U$931 ( \3058 , RI2b5e785c0a00_257, \2616 );
and \U$932 ( \3059 , RI2b5e785be390_277, \2622 );
and \U$933 ( \3060 , RI2b5e785bc0e0_297, \2624 );
and \U$934 ( \3061 , RI2b5e785ba1f0_317, \2626 );
and \U$935 ( \3062 , RI2b5e785b9890_337, \2628 );
and \U$936 ( \3063 , RI2b5e785b7d60_357, \2630 );
and \U$937 ( \3064 , RI2b5e785b7400_377, \2632 );
and \U$938 ( \3065 , RI2b5e785b5c90_397, \2634 );
and \U$939 ( \3066 , RI2b5e785b5330_417, \2636 );
and \U$940 ( \3067 , RI2b5e785b49d0_437, \2638 );
and \U$941 ( \3068 , RI2b5e785b3620_457, \2640 );
and \U$942 ( \3069 , RI2b5e785b2cc0_477, \2642 );
and \U$943 ( \3070 , RI2b5e785b2360_497, \2644 );
and \U$944 ( \3071 , RI2b5e785b1370_517, \2646 );
and \U$945 ( \3072 , RI2b5e785b0a10_537, \2648 );
and \U$946 ( \3073 , RI2b5e785b00b0_557, \2650 );
and \U$947 ( \3074 , RI2b5e785af480_577, \2652 );
or \U$948 ( \3075 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 );
_DC g21d1 ( \3076_nG21d1 , \3075 , \2671 );
buf \U$949 ( \3077 , \3076_nG21d1 );
xor \U$950 ( \3078 , \2360 , \2381 );
xor \U$951 ( \3079 , \3078 , \2518 );
buf g1cfc_GF_PartitionCandidate( \3080_nG1cfc , \3079 );
buf \U$952 ( \3081 , \3080_nG1cfc );
xor \U$953 ( \3082 , \2385 , \2406 );
xor \U$954 ( \3083 , \3082 , \2515 );
buf g1cd8_GF_PartitionCandidate( \3084_nG1cd8 , \3083 );
buf \U$955 ( \3085 , \3084_nG1cd8 );
xor \U$956 ( \3086 , \3081 , \3085 );
xor \U$957 ( \3087 , \3085 , \3021 );
not \U$958 ( \3088 , \3087 );
and \U$959 ( \3089 , \3086 , \3088 );
and \U$960 ( \3090 , \3077 , \3089 );
and \U$961 ( \3091 , RI2b5e785c2b48_256, \2616 );
and \U$962 ( \3092 , RI2b5e785be408_276, \2622 );
and \U$963 ( \3093 , RI2b5e785bc158_296, \2624 );
and \U$964 ( \3094 , RI2b5e785ba268_316, \2626 );
and \U$965 ( \3095 , RI2b5e785b9908_336, \2628 );
and \U$966 ( \3096 , RI2b5e785b7dd8_356, \2630 );
and \U$967 ( \3097 , RI2b5e785b7478_376, \2632 );
and \U$968 ( \3098 , RI2b5e785b5d08_396, \2634 );
and \U$969 ( \3099 , RI2b5e785b53a8_416, \2636 );
and \U$970 ( \3100 , RI2b5e785b4a48_436, \2638 );
and \U$971 ( \3101 , RI2b5e785b3698_456, \2640 );
and \U$972 ( \3102 , RI2b5e785b2d38_476, \2642 );
and \U$973 ( \3103 , RI2b5e785b23d8_496, \2644 );
and \U$974 ( \3104 , RI2b5e785b13e8_516, \2646 );
and \U$975 ( \3105 , RI2b5e785b0a88_536, \2648 );
and \U$976 ( \3106 , RI2b5e785b0128_556, \2650 );
and \U$977 ( \3107 , RI2b5e785af4f8_576, \2652 );
or \U$978 ( \3108 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 );
_DC g22a8 ( \3109_nG22a8 , \3108 , \2671 );
buf \U$979 ( \3110 , \3109_nG22a8 );
and \U$980 ( \3111 , \3110 , \3087 );
nor \U$981 ( \3112 , \3090 , \3111 );
and \U$982 ( \3113 , \3085 , \3021 );
not \U$983 ( \3114 , \3113 );
and \U$984 ( \3115 , \3081 , \3114 );
xnor \U$985 ( \3116 , \3112 , \3115 );
and \U$986 ( \3117 , \3056 , \3116 );
and \U$987 ( \3118 , \2997 , \3116 );
or \U$988 ( \3119 , \3057 , \3117 , \3118 );
and \U$989 ( \3120 , RI2b5e785c0910_259, \2616 );
and \U$990 ( \3121 , RI2b5e785be2a0_279, \2622 );
and \U$991 ( \3122 , RI2b5e785bbff0_299, \2624 );
and \U$992 ( \3123 , RI2b5e785ba100_319, \2626 );
and \U$993 ( \3124 , RI2b5e785b97a0_339, \2628 );
and \U$994 ( \3125 , RI2b5e785b7c70_359, \2630 );
and \U$995 ( \3126 , RI2b5e785b7310_379, \2632 );
and \U$996 ( \3127 , RI2b5e785b5ba0_399, \2634 );
and \U$997 ( \3128 , RI2b5e785b5240_419, \2636 );
and \U$998 ( \3129 , RI2b5e785b48e0_439, \2638 );
and \U$999 ( \3130 , RI2b5e785b3530_459, \2640 );
and \U$1000 ( \3131 , RI2b5e785b2bd0_479, \2642 );
and \U$1001 ( \3132 , RI2b5e785b2270_499, \2644 );
and \U$1002 ( \3133 , RI2b5e785b1280_519, \2646 );
and \U$1003 ( \3134 , RI2b5e785b0920_539, \2648 );
and \U$1004 ( \3135 , RI2b5e785affc0_559, \2650 );
and \U$1005 ( \3136 , RI2b5e785af390_579, \2652 );
or \U$1006 ( \3137 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 );
_DC g2012 ( \3138_nG2012 , \3137 , \2671 );
buf \U$1007 ( \3139 , \3138_nG2012 );
xor \U$1008 ( \3140 , \2335 , \2356 );
xor \U$1009 ( \3141 , \3140 , \2521 );
buf g1e3a_GF_PartitionCandidate( \3142_nG1e3a , \3141 );
buf \U$1010 ( \3143 , \3142_nG1e3a );
xor \U$1011 ( \3144 , \2845 , \3143 );
xor \U$1012 ( \3145 , \3143 , \3081 );
not \U$1013 ( \3146 , \3145 );
and \U$1014 ( \3147 , \3144 , \3146 );
and \U$1015 ( \3148 , \3139 , \3147 );
and \U$1016 ( \3149 , RI2b5e785c0988_258, \2616 );
and \U$1017 ( \3150 , RI2b5e785be318_278, \2622 );
and \U$1018 ( \3151 , RI2b5e785bc068_298, \2624 );
and \U$1019 ( \3152 , RI2b5e785ba178_318, \2626 );
and \U$1020 ( \3153 , RI2b5e785b9818_338, \2628 );
and \U$1021 ( \3154 , RI2b5e785b7ce8_358, \2630 );
and \U$1022 ( \3155 , RI2b5e785b7388_378, \2632 );
and \U$1023 ( \3156 , RI2b5e785b5c18_398, \2634 );
and \U$1024 ( \3157 , RI2b5e785b52b8_418, \2636 );
and \U$1025 ( \3158 , RI2b5e785b4958_438, \2638 );
and \U$1026 ( \3159 , RI2b5e785b35a8_458, \2640 );
and \U$1027 ( \3160 , RI2b5e785b2c48_478, \2642 );
and \U$1028 ( \3161 , RI2b5e785b22e8_498, \2644 );
and \U$1029 ( \3162 , RI2b5e785b12f8_518, \2646 );
and \U$1030 ( \3163 , RI2b5e785b0998_538, \2648 );
and \U$1031 ( \3164 , RI2b5e785b0038_558, \2650 );
and \U$1032 ( \3165 , RI2b5e785af408_578, \2652 );
or \U$1033 ( \3166 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 );
_DC g20db ( \3167_nG20db , \3166 , \2671 );
buf \U$1034 ( \3168 , \3167_nG20db );
and \U$1035 ( \3169 , \3168 , \3145 );
nor \U$1036 ( \3170 , \3148 , \3169 );
and \U$1037 ( \3171 , \3143 , \3081 );
not \U$1038 ( \3172 , \3171 );
and \U$1039 ( \3173 , \2845 , \3172 );
xnor \U$1040 ( \3174 , \3170 , \3173 );
and \U$1041 ( \3175 , RI2b5e785c0820_261, \2616 );
and \U$1042 ( \3176 , RI2b5e785be1b0_281, \2622 );
and \U$1043 ( \3177 , RI2b5e785bbf00_301, \2624 );
and \U$1044 ( \3178 , RI2b5e785ba010_321, \2626 );
and \U$1045 ( \3179 , RI2b5e785b96b0_341, \2628 );
and \U$1046 ( \3180 , RI2b5e785b7b80_361, \2630 );
and \U$1047 ( \3181 , RI2b5e785b7220_381, \2632 );
and \U$1048 ( \3182 , RI2b5e785b5ab0_401, \2634 );
and \U$1049 ( \3183 , RI2b5e785b5150_421, \2636 );
and \U$1050 ( \3184 , RI2b5e785b47f0_441, \2638 );
and \U$1051 ( \3185 , RI2b5e785b3440_461, \2640 );
and \U$1052 ( \3186 , RI2b5e785b2ae0_481, \2642 );
and \U$1053 ( \3187 , RI2b5e785b2180_501, \2644 );
and \U$1054 ( \3188 , RI2b5e785b1190_521, \2646 );
and \U$1055 ( \3189 , RI2b5e785b0830_541, \2648 );
and \U$1056 ( \3190 , RI2b5e785afed0_561, \2650 );
and \U$1057 ( \3191 , RI2b5e785af2a0_581, \2652 );
or \U$1058 ( \3192 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 );
_DC g1e79 ( \3193_nG1e79 , \3192 , \2671 );
buf \U$1059 ( \3194 , \3193_nG1e79 );
and \U$1060 ( \3195 , \3194 , \2848 );
and \U$1061 ( \3196 , RI2b5e785c0898_260, \2616 );
and \U$1062 ( \3197 , RI2b5e785be228_280, \2622 );
and \U$1063 ( \3198 , RI2b5e785bbf78_300, \2624 );
and \U$1064 ( \3199 , RI2b5e785ba088_320, \2626 );
and \U$1065 ( \3200 , RI2b5e785b9728_340, \2628 );
and \U$1066 ( \3201 , RI2b5e785b7bf8_360, \2630 );
and \U$1067 ( \3202 , RI2b5e785b7298_380, \2632 );
and \U$1068 ( \3203 , RI2b5e785b5b28_400, \2634 );
and \U$1069 ( \3204 , RI2b5e785b51c8_420, \2636 );
and \U$1070 ( \3205 , RI2b5e785b4868_440, \2638 );
and \U$1071 ( \3206 , RI2b5e785b34b8_460, \2640 );
and \U$1072 ( \3207 , RI2b5e785b2b58_480, \2642 );
and \U$1073 ( \3208 , RI2b5e785b21f8_500, \2644 );
and \U$1074 ( \3209 , RI2b5e785b1208_520, \2646 );
and \U$1075 ( \3210 , RI2b5e785b08a8_540, \2648 );
and \U$1076 ( \3211 , RI2b5e785aff48_560, \2650 );
and \U$1077 ( \3212 , RI2b5e785af318_580, \2652 );
or \U$1078 ( \3213 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 );
_DC g1f2c ( \3214_nG1f2c , \3213 , \2671 );
buf \U$1079 ( \3215 , \3214_nG1f2c );
and \U$1080 ( \3216 , \3215 , \2846 );
nor \U$1081 ( \3217 , \3195 , \3216 );
xnor \U$1082 ( \3218 , \3217 , \2853 );
and \U$1083 ( \3219 , \3174 , \3218 );
and \U$1084 ( \3220 , RI2b5e785c0730_263, \2616 );
and \U$1085 ( \3221 , RI2b5e785be0c0_283, \2622 );
and \U$1086 ( \3222 , RI2b5e785bbe10_303, \2624 );
and \U$1087 ( \3223 , RI2b5e785b9f20_323, \2626 );
and \U$1088 ( \3224 , RI2b5e785b95c0_343, \2628 );
and \U$1089 ( \3225 , RI2b5e785b7a90_363, \2630 );
and \U$1090 ( \3226 , RI2b5e785b7130_383, \2632 );
and \U$1091 ( \3227 , RI2b5e785b59c0_403, \2634 );
and \U$1092 ( \3228 , RI2b5e785b5060_423, \2636 );
and \U$1093 ( \3229 , RI2b5e785b3cb0_443, \2638 );
and \U$1094 ( \3230 , RI2b5e785b3350_463, \2640 );
and \U$1095 ( \3231 , RI2b5e785b29f0_483, \2642 );
and \U$1096 ( \3232 , RI2b5e785b1a00_503, \2644 );
and \U$1097 ( \3233 , RI2b5e785b10a0_523, \2646 );
and \U$1098 ( \3234 , RI2b5e785b0740_543, \2648 );
and \U$1099 ( \3235 , RI2b5e785afde0_563, \2650 );
and \U$1100 ( \3236 , RI2b5e785af1b0_583, \2652 );
or \U$1101 ( \3237 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 );
_DC g1d15 ( \3238_nG1d15 , \3237 , \2671 );
buf \U$1102 ( \3239 , \3238_nG1d15 );
and \U$1103 ( \3240 , \3239 , \2783 );
and \U$1104 ( \3241 , RI2b5e785c07a8_262, \2616 );
and \U$1105 ( \3242 , RI2b5e785be138_282, \2622 );
and \U$1106 ( \3243 , RI2b5e785bbe88_302, \2624 );
and \U$1107 ( \3244 , RI2b5e785b9f98_322, \2626 );
and \U$1108 ( \3245 , RI2b5e785b9638_342, \2628 );
and \U$1109 ( \3246 , RI2b5e785b7b08_362, \2630 );
and \U$1110 ( \3247 , RI2b5e785b71a8_382, \2632 );
and \U$1111 ( \3248 , RI2b5e785b5a38_402, \2634 );
and \U$1112 ( \3249 , RI2b5e785b50d8_422, \2636 );
and \U$1113 ( \3250 , RI2b5e785b4778_442, \2638 );
and \U$1114 ( \3251 , RI2b5e785b33c8_462, \2640 );
and \U$1115 ( \3252 , RI2b5e785b2a68_482, \2642 );
and \U$1116 ( \3253 , RI2b5e785b1a78_502, \2644 );
and \U$1117 ( \3254 , RI2b5e785b1118_522, \2646 );
and \U$1118 ( \3255 , RI2b5e785b07b8_542, \2648 );
and \U$1119 ( \3256 , RI2b5e785afe58_562, \2650 );
and \U$1120 ( \3257 , RI2b5e785af228_582, \2652 );
or \U$1121 ( \3258 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 );
_DC g1dbc ( \3259_nG1dbc , \3258 , \2671 );
buf \U$1122 ( \3260 , \3259_nG1dbc );
and \U$1123 ( \3261 , \3260 , \2781 );
nor \U$1124 ( \3262 , \3240 , \3261 );
xnor \U$1125 ( \3263 , \3262 , \2550 );
and \U$1126 ( \3264 , \3218 , \3263 );
and \U$1127 ( \3265 , \3174 , \3263 );
or \U$1128 ( \3266 , \3219 , \3264 , \3265 );
and \U$1129 ( \3267 , \3119 , \3266 );
and \U$1130 ( \3268 , RI2b5e785c0640_265, \2616 );
and \U$1131 ( \3269 , RI2b5e785bdfd0_285, \2622 );
and \U$1132 ( \3270 , RI2b5e785bbd20_305, \2624 );
and \U$1133 ( \3271 , RI2b5e785b9e30_325, \2626 );
and \U$1134 ( \3272 , RI2b5e785b94d0_345, \2628 );
and \U$1135 ( \3273 , RI2b5e785b79a0_365, \2630 );
and \U$1136 ( \3274 , RI2b5e785b7040_385, \2632 );
and \U$1137 ( \3275 , RI2b5e785b58d0_405, \2634 );
and \U$1138 ( \3276 , RI2b5e785b4f70_425, \2636 );
and \U$1139 ( \3277 , RI2b5e785b3bc0_445, \2638 );
and \U$1140 ( \3278 , RI2b5e785b3260_465, \2640 );
and \U$1141 ( \3279 , RI2b5e785b2900_485, \2642 );
and \U$1142 ( \3280 , RI2b5e785b1910_505, \2644 );
and \U$1143 ( \3281 , RI2b5e785b0fb0_525, \2646 );
and \U$1144 ( \3282 , RI2b5e785b0650_545, \2648 );
and \U$1145 ( \3283 , RI2b5e785afcf0_565, \2650 );
and \U$1146 ( \3284 , RI2b5e785af0c0_585, \2652 );
or \U$1147 ( \3285 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 );
_DC g1ba5 ( \3286_nG1ba5 , \3285 , \2671 );
buf \U$1148 ( \3287 , \3286_nG1ba5 );
and \U$1149 ( \3288 , \3287 , \2721 );
and \U$1150 ( \3289 , RI2b5e785c06b8_264, \2616 );
and \U$1151 ( \3290 , RI2b5e785be048_284, \2622 );
and \U$1152 ( \3291 , RI2b5e785bbd98_304, \2624 );
and \U$1153 ( \3292 , RI2b5e785b9ea8_324, \2626 );
and \U$1154 ( \3293 , RI2b5e785b9548_344, \2628 );
and \U$1155 ( \3294 , RI2b5e785b7a18_364, \2630 );
and \U$1156 ( \3295 , RI2b5e785b70b8_384, \2632 );
and \U$1157 ( \3296 , RI2b5e785b5948_404, \2634 );
and \U$1158 ( \3297 , RI2b5e785b4fe8_424, \2636 );
and \U$1159 ( \3298 , RI2b5e785b3c38_444, \2638 );
and \U$1160 ( \3299 , RI2b5e785b32d8_464, \2640 );
and \U$1161 ( \3300 , RI2b5e785b2978_484, \2642 );
and \U$1162 ( \3301 , RI2b5e785b1988_504, \2644 );
and \U$1163 ( \3302 , RI2b5e785b1028_524, \2646 );
and \U$1164 ( \3303 , RI2b5e785b06c8_544, \2648 );
and \U$1165 ( \3304 , RI2b5e785afd68_564, \2650 );
and \U$1166 ( \3305 , RI2b5e785af138_584, \2652 );
or \U$1167 ( \3306 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 );
_DC g1c76 ( \3307_nG1c76 , \3306 , \2671 );
buf \U$1168 ( \3308 , \3307_nG1c76 );
and \U$1169 ( \3309 , \3308 , \2719 );
nor \U$1170 ( \3310 , \3288 , \3309 );
xnor \U$1171 ( \3311 , \3310 , \2747 );
and \U$1173 ( \3312 , RI2b5e785c05c8_266, \2616 );
and \U$1174 ( \3313 , RI2b5e785bdf58_286, \2622 );
and \U$1175 ( \3314 , RI2b5e785bbca8_306, \2624 );
and \U$1176 ( \3315 , RI2b5e785b9db8_326, \2626 );
and \U$1177 ( \3316 , RI2b5e785b9458_346, \2628 );
and \U$1178 ( \3317 , RI2b5e785b7928_366, \2630 );
and \U$1179 ( \3318 , RI2b5e785b6fc8_386, \2632 );
and \U$1180 ( \3319 , RI2b5e785b5858_406, \2634 );
and \U$1181 ( \3320 , RI2b5e785b4ef8_426, \2636 );
and \U$1182 ( \3321 , RI2b5e785b3b48_446, \2638 );
and \U$1183 ( \3322 , RI2b5e785b31e8_466, \2640 );
and \U$1184 ( \3323 , RI2b5e785b2888_486, \2642 );
and \U$1185 ( \3324 , RI2b5e785b1898_506, \2644 );
and \U$1186 ( \3325 , RI2b5e785b0f38_526, \2646 );
and \U$1187 ( \3326 , RI2b5e785b05d8_546, \2648 );
and \U$1188 ( \3327 , RI2b5e785afc78_566, \2650 );
and \U$1189 ( \3328 , RI2b5e785af048_586, \2652 );
or \U$1190 ( \3329 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 );
_DC g1b63 ( \3330_nG1b63 , \3329 , \2671 );
buf \U$1191 ( \3331 , \3330_nG1b63 );
and \U$1192 ( \3332 , \3331 , \2774 );
nor \U$1193 ( \3333 , 1'b0 , \3332 );
xnor \U$1194 ( \3334 , \3333 , 1'b0 );
and \U$1195 ( \3335 , \3311 , \3334 );
and \U$1196 ( \3336 , \3266 , \3335 );
and \U$1197 ( \3337 , \3119 , \3335 );
or \U$1198 ( \3338 , \3267 , \3336 , \3337 );
and \U$1200 ( \3339 , \3260 , \2783 );
and \U$1201 ( \3340 , \3194 , \2781 );
nor \U$1202 ( \3341 , \3339 , \3340 );
xnor \U$1203 ( \3342 , \3341 , \2550 );
and \U$1204 ( \3343 , \3308 , \2721 );
and \U$1205 ( \3344 , \3239 , \2719 );
nor \U$1206 ( \3345 , \3343 , \3344 );
xnor \U$1207 ( \3346 , \3345 , \2747 );
xor \U$1208 ( \3347 , \3342 , \3346 );
and \U$1210 ( \3348 , \3287 , \2774 );
nor \U$1211 ( \3349 , 1'b0 , \3348 );
xnor \U$1212 ( \3350 , \3349 , 1'b0 );
xor \U$1213 ( \3351 , \3347 , \3350 );
and \U$1214 ( \3352 , \3110 , \3089 );
and \U$1215 ( \3353 , \3017 , \3087 );
nor \U$1216 ( \3354 , \3352 , \3353 );
xnor \U$1217 ( \3355 , \3354 , \3115 );
and \U$1218 ( \3356 , \3168 , \3147 );
and \U$1219 ( \3357 , \3077 , \3145 );
nor \U$1220 ( \3358 , \3356 , \3357 );
xnor \U$1221 ( \3359 , \3358 , \3173 );
xor \U$1222 ( \3360 , \3355 , \3359 );
and \U$1223 ( \3361 , \3215 , \2848 );
and \U$1224 ( \3362 , \3139 , \2846 );
nor \U$1225 ( \3363 , \3361 , \3362 );
xnor \U$1226 ( \3364 , \3363 , \2853 );
xor \U$1227 ( \3365 , \3360 , \3364 );
and \U$1228 ( \3366 , \3351 , \3365 );
or \U$1230 ( \3367 , 1'b0 , \3366 , 1'b0 );
xor \U$1231 ( \3368 , \3338 , \3367 );
and \U$1232 ( \3369 , \3239 , \2721 );
and \U$1233 ( \3370 , \3260 , \2719 );
nor \U$1234 ( \3371 , \3369 , \3370 );
xnor \U$1235 ( \3372 , \3371 , \2747 );
and \U$1237 ( \3373 , \3308 , \2774 );
nor \U$1238 ( \3374 , 1'b0 , \3373 );
xnor \U$1239 ( \3375 , \3374 , 1'b0 );
xor \U$1240 ( \3376 , \3372 , \3375 );
xor \U$1242 ( \3377 , \3376 , 1'b0 );
and \U$1243 ( \3378 , \3077 , \3147 );
and \U$1244 ( \3379 , \3110 , \3145 );
nor \U$1245 ( \3380 , \3378 , \3379 );
xnor \U$1246 ( \3381 , \3380 , \3173 );
and \U$1247 ( \3382 , \3139 , \2848 );
and \U$1248 ( \3383 , \3168 , \2846 );
nor \U$1249 ( \3384 , \3382 , \3383 );
xnor \U$1250 ( \3385 , \3384 , \2853 );
xor \U$1251 ( \3386 , \3381 , \3385 );
and \U$1252 ( \3387 , \3194 , \2783 );
and \U$1253 ( \3388 , \3215 , \2781 );
nor \U$1254 ( \3389 , \3387 , \3388 );
xnor \U$1255 ( \3390 , \3389 , \2550 );
xor \U$1256 ( \3391 , \3386 , \3390 );
xor \U$1257 ( \3392 , \3377 , \3391 );
and \U$1258 ( \3393 , \2901 , \2993 );
and \U$1259 ( \3394 , \2769 , \2990 );
nor \U$1260 ( \3395 , \3393 , \3394 );
xnor \U$1261 ( \3396 , \3395 , \2987 );
and \U$1262 ( \3397 , \2924 , \3029 );
and \U$1263 ( \3398 , \2880 , \3027 );
nor \U$1264 ( \3399 , \3397 , \3398 );
xnor \U$1265 ( \3400 , \3399 , \3055 );
xor \U$1266 ( \3401 , \3396 , \3400 );
and \U$1267 ( \3402 , \3017 , \3089 );
and \U$1268 ( \3403 , \3050 , \3087 );
nor \U$1269 ( \3404 , \3402 , \3403 );
xnor \U$1270 ( \3405 , \3404 , \3115 );
xor \U$1271 ( \3406 , \3401 , \3405 );
xor \U$1272 ( \3407 , \3392 , \3406 );
xor \U$1273 ( \3408 , \3368 , \3407 );
and \U$1275 ( \3409 , \3050 , \2993 );
and \U$1276 ( \3410 , \2924 , \2990 );
nor \U$1277 ( \3411 , \3409 , \3410 );
xnor \U$1278 ( \3412 , \3411 , \2987 );
and \U$1279 ( \3413 , \3110 , \3029 );
and \U$1280 ( \3414 , \3017 , \3027 );
nor \U$1281 ( \3415 , \3413 , \3414 );
xnor \U$1282 ( \3416 , \3415 , \3055 );
and \U$1283 ( \3417 , \3412 , \3416 );
or \U$1285 ( \3418 , 1'b0 , \3417 , 1'b0 );
and \U$1286 ( \3419 , \3168 , \3089 );
and \U$1287 ( \3420 , \3077 , \3087 );
nor \U$1288 ( \3421 , \3419 , \3420 );
xnor \U$1289 ( \3422 , \3421 , \3115 );
and \U$1290 ( \3423 , \3215 , \3147 );
and \U$1291 ( \3424 , \3139 , \3145 );
nor \U$1292 ( \3425 , \3423 , \3424 );
xnor \U$1293 ( \3426 , \3425 , \3173 );
and \U$1294 ( \3427 , \3422 , \3426 );
and \U$1295 ( \3428 , \3260 , \2848 );
and \U$1296 ( \3429 , \3194 , \2846 );
nor \U$1297 ( \3430 , \3428 , \3429 );
xnor \U$1298 ( \3431 , \3430 , \2853 );
and \U$1299 ( \3432 , \3426 , \3431 );
and \U$1300 ( \3433 , \3422 , \3431 );
or \U$1301 ( \3434 , \3427 , \3432 , \3433 );
and \U$1302 ( \3435 , \3418 , \3434 );
and \U$1303 ( \3436 , \3308 , \2783 );
and \U$1304 ( \3437 , \3239 , \2781 );
nor \U$1305 ( \3438 , \3436 , \3437 );
xnor \U$1306 ( \3439 , \3438 , \2550 );
and \U$1307 ( \3440 , \3331 , \2721 );
and \U$1308 ( \3441 , \3287 , \2719 );
nor \U$1309 ( \3442 , \3440 , \3441 );
xnor \U$1310 ( \3443 , \3442 , \2747 );
and \U$1311 ( \3444 , \3439 , \3443 );
and \U$1312 ( \3445 , RI2b5e785c0550_267, \2616 );
and \U$1313 ( \3446 , RI2b5e785bc590_287, \2622 );
and \U$1314 ( \3447 , RI2b5e785bbc30_307, \2624 );
and \U$1315 ( \3448 , RI2b5e785b9d40_327, \2626 );
and \U$1316 ( \3449 , RI2b5e785b93e0_347, \2628 );
and \U$1317 ( \3450 , RI2b5e785b78b0_367, \2630 );
and \U$1318 ( \3451 , RI2b5e785b6f50_387, \2632 );
and \U$1319 ( \3452 , RI2b5e785b57e0_407, \2634 );
and \U$1320 ( \3453 , RI2b5e785b4e80_427, \2636 );
and \U$1321 ( \3454 , RI2b5e785b3ad0_447, \2638 );
and \U$1322 ( \3455 , RI2b5e785b3170_467, \2640 );
and \U$1323 ( \3456 , RI2b5e785b2810_487, \2642 );
and \U$1324 ( \3457 , RI2b5e785b1820_507, \2644 );
and \U$1325 ( \3458 , RI2b5e785b0ec0_527, \2646 );
and \U$1326 ( \3459 , RI2b5e785b0560_547, \2648 );
and \U$1327 ( \3460 , RI2b5e785afc00_567, \2650 );
and \U$1328 ( \3461 , RI2b5e785aefd0_587, \2652 );
or \U$1329 ( \3462 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 );
_DC g1a4f ( \3463_nG1a4f , \3462 , \2671 );
buf \U$1330 ( \3464 , \3463_nG1a4f );
nand \U$1331 ( \3465 , \3464 , \2774 );
xnor \U$1332 ( \3466 , \3465 , 1'b0 );
and \U$1333 ( \3467 , \3443 , \3466 );
and \U$1334 ( \3468 , \3439 , \3466 );
or \U$1335 ( \3469 , \3444 , \3467 , \3468 );
and \U$1336 ( \3470 , \3434 , \3469 );
and \U$1337 ( \3471 , \3418 , \3469 );
or \U$1338 ( \3472 , \3435 , \3470 , \3471 );
xor \U$1339 ( \3473 , \3311 , \3334 );
xor \U$1340 ( \3474 , \3174 , \3218 );
xor \U$1341 ( \3475 , \3474 , \3263 );
and \U$1342 ( \3476 , \3473 , \3475 );
xor \U$1343 ( \3477 , \2997 , \3056 );
xor \U$1344 ( \3478 , \3477 , \3116 );
and \U$1345 ( \3479 , \3475 , \3478 );
and \U$1346 ( \3480 , \3473 , \3478 );
or \U$1347 ( \3481 , \3476 , \3479 , \3480 );
and \U$1348 ( \3482 , \3472 , \3481 );
and \U$1350 ( \3483 , \2880 , \2993 );
and \U$1351 ( \3484 , \2901 , \2990 );
nor \U$1352 ( \3485 , \3483 , \3484 );
xnor \U$1353 ( \3486 , \3485 , \2987 );
xor \U$1354 ( \3487 , 1'b0 , \3486 );
and \U$1355 ( \3488 , \3050 , \3029 );
and \U$1356 ( \3489 , \2924 , \3027 );
nor \U$1357 ( \3490 , \3488 , \3489 );
xnor \U$1358 ( \3491 , \3490 , \3055 );
xor \U$1359 ( \3492 , \3487 , \3491 );
and \U$1360 ( \3493 , \3481 , \3492 );
and \U$1361 ( \3494 , \3472 , \3492 );
or \U$1362 ( \3495 , \3482 , \3493 , \3494 );
xor \U$1364 ( \3496 , 1'b0 , \3351 );
xor \U$1365 ( \3497 , \3496 , \3365 );
xor \U$1366 ( \3498 , \3119 , \3266 );
xor \U$1367 ( \3499 , \3498 , \3335 );
and \U$1368 ( \3500 , \3497 , \3499 );
xor \U$1369 ( \3501 , \3495 , \3500 );
and \U$1371 ( \3502 , \3486 , \3491 );
or \U$1373 ( \3503 , 1'b0 , \3502 , 1'b0 );
and \U$1374 ( \3504 , \3355 , \3359 );
and \U$1375 ( \3505 , \3359 , \3364 );
and \U$1376 ( \3506 , \3355 , \3364 );
or \U$1377 ( \3507 , \3504 , \3505 , \3506 );
xor \U$1378 ( \3508 , \3503 , \3507 );
and \U$1379 ( \3509 , \3342 , \3346 );
and \U$1380 ( \3510 , \3346 , \3350 );
and \U$1381 ( \3511 , \3342 , \3350 );
or \U$1382 ( \3512 , \3509 , \3510 , \3511 );
xor \U$1383 ( \3513 , \3508 , \3512 );
xor \U$1384 ( \3514 , \3501 , \3513 );
xor \U$1385 ( \3515 , \3408 , \3514 );
and \U$1386 ( \3516 , \3017 , \2993 );
and \U$1387 ( \3517 , \3050 , \2990 );
nor \U$1388 ( \3518 , \3516 , \3517 );
xnor \U$1389 ( \3519 , \3518 , \2987 );
and \U$1390 ( \3520 , \3077 , \3029 );
and \U$1391 ( \3521 , \3110 , \3027 );
nor \U$1392 ( \3522 , \3520 , \3521 );
xnor \U$1393 ( \3523 , \3522 , \3055 );
and \U$1394 ( \3524 , \3519 , \3523 );
and \U$1395 ( \3525 , \3139 , \3089 );
and \U$1396 ( \3526 , \3168 , \3087 );
nor \U$1397 ( \3527 , \3525 , \3526 );
xnor \U$1398 ( \3528 , \3527 , \3115 );
and \U$1399 ( \3529 , \3523 , \3528 );
and \U$1400 ( \3530 , \3519 , \3528 );
or \U$1401 ( \3531 , \3524 , \3529 , \3530 );
and \U$1402 ( \3532 , \3194 , \3147 );
and \U$1403 ( \3533 , \3215 , \3145 );
nor \U$1404 ( \3534 , \3532 , \3533 );
xnor \U$1405 ( \3535 , \3534 , \3173 );
and \U$1406 ( \3536 , \3239 , \2848 );
and \U$1407 ( \3537 , \3260 , \2846 );
nor \U$1408 ( \3538 , \3536 , \3537 );
xnor \U$1409 ( \3539 , \3538 , \2853 );
and \U$1410 ( \3540 , \3535 , \3539 );
and \U$1411 ( \3541 , \3287 , \2783 );
and \U$1412 ( \3542 , \3308 , \2781 );
nor \U$1413 ( \3543 , \3541 , \3542 );
xnor \U$1414 ( \3544 , \3543 , \2550 );
and \U$1415 ( \3545 , \3539 , \3544 );
and \U$1416 ( \3546 , \3535 , \3544 );
or \U$1417 ( \3547 , \3540 , \3545 , \3546 );
and \U$1418 ( \3548 , \3531 , \3547 );
xor \U$1419 ( \3549 , \3439 , \3443 );
xor \U$1420 ( \3550 , \3549 , \3466 );
and \U$1421 ( \3551 , \3547 , \3550 );
and \U$1422 ( \3552 , \3531 , \3550 );
or \U$1423 ( \3553 , \3548 , \3551 , \3552 );
xor \U$1424 ( \3554 , \3422 , \3426 );
xor \U$1425 ( \3555 , \3554 , \3431 );
xor \U$1426 ( \3556 , 1'b0 , \3412 );
xor \U$1427 ( \3557 , \3556 , \3416 );
and \U$1428 ( \3558 , \3555 , \3557 );
and \U$1429 ( \3559 , \3553 , \3558 );
xor \U$1430 ( \3560 , \3473 , \3475 );
xor \U$1431 ( \3561 , \3560 , \3478 );
and \U$1432 ( \3562 , \3558 , \3561 );
and \U$1433 ( \3563 , \3553 , \3561 );
or \U$1434 ( \3564 , \3559 , \3562 , \3563 );
xor \U$1435 ( \3565 , \3497 , \3499 );
and \U$1436 ( \3566 , \3564 , \3565 );
xor \U$1437 ( \3567 , \3472 , \3481 );
xor \U$1438 ( \3568 , \3567 , \3492 );
and \U$1439 ( \3569 , \3565 , \3568 );
and \U$1440 ( \3570 , \3564 , \3568 );
or \U$1441 ( \3571 , \3566 , \3569 , \3570 );
nor \U$1442 ( \3572 , \3515 , \3571 );
and \U$1443 ( \3573 , \3495 , \3500 );
and \U$1444 ( \3574 , \3500 , \3513 );
and \U$1445 ( \3575 , \3495 , \3513 );
or \U$1446 ( \3576 , \3573 , \3574 , \3575 );
and \U$1447 ( \3577 , \3338 , \3367 );
and \U$1448 ( \3578 , \3367 , \3407 );
and \U$1449 ( \3579 , \3338 , \3407 );
or \U$1450 ( \3580 , \3577 , \3578 , \3579 );
and \U$1452 ( \3581 , \2769 , \2993 );
and \U$1453 ( \3582 , \2673 , \2990 );
nor \U$1454 ( \3583 , \3581 , \3582 );
xnor \U$1455 ( \3584 , \3583 , \2987 );
xor \U$1456 ( \3585 , 1'b0 , \3584 );
and \U$1457 ( \3586 , \2880 , \3029 );
and \U$1458 ( \3587 , \2901 , \3027 );
nor \U$1459 ( \3588 , \3586 , \3587 );
xnor \U$1460 ( \3589 , \3588 , \3055 );
xor \U$1461 ( \3590 , \3585 , \3589 );
and \U$1463 ( \3591 , \3215 , \2783 );
and \U$1464 ( \3592 , \3139 , \2781 );
nor \U$1465 ( \3593 , \3591 , \3592 );
xnor \U$1466 ( \3594 , \3593 , \2550 );
and \U$1467 ( \3595 , \3260 , \2721 );
and \U$1468 ( \3596 , \3194 , \2719 );
nor \U$1469 ( \3597 , \3595 , \3596 );
xnor \U$1470 ( \3598 , \3597 , \2747 );
xor \U$1471 ( \3599 , \3594 , \3598 );
and \U$1473 ( \3600 , \3239 , \2774 );
nor \U$1474 ( \3601 , 1'b0 , \3600 );
xnor \U$1475 ( \3602 , \3601 , 1'b0 );
xor \U$1476 ( \3603 , \3599 , \3602 );
xor \U$1477 ( \3604 , 1'b0 , \3603 );
xor \U$1478 ( \3605 , \3590 , \3604 );
and \U$1479 ( \3606 , \3396 , \3400 );
and \U$1480 ( \3607 , \3400 , \3405 );
and \U$1481 ( \3608 , \3396 , \3405 );
or \U$1482 ( \3609 , \3606 , \3607 , \3608 );
and \U$1483 ( \3610 , \3381 , \3385 );
and \U$1484 ( \3611 , \3385 , \3390 );
and \U$1485 ( \3612 , \3381 , \3390 );
or \U$1486 ( \3613 , \3610 , \3611 , \3612 );
xor \U$1487 ( \3614 , \3609 , \3613 );
and \U$1488 ( \3615 , \3372 , \3375 );
or \U$1491 ( \3616 , \3615 , 1'b0 , 1'b0 );
xor \U$1492 ( \3617 , \3614 , \3616 );
xor \U$1493 ( \3618 , \3605 , \3617 );
xor \U$1494 ( \3619 , \3580 , \3618 );
and \U$1495 ( \3620 , \3503 , \3507 );
and \U$1496 ( \3621 , \3507 , \3512 );
and \U$1497 ( \3622 , \3503 , \3512 );
or \U$1498 ( \3623 , \3620 , \3621 , \3622 );
and \U$1499 ( \3624 , \3377 , \3391 );
and \U$1500 ( \3625 , \3391 , \3406 );
and \U$1501 ( \3626 , \3377 , \3406 );
or \U$1502 ( \3627 , \3624 , \3625 , \3626 );
xor \U$1503 ( \3628 , \3623 , \3627 );
and \U$1504 ( \3629 , \3050 , \3089 );
and \U$1505 ( \3630 , \2924 , \3087 );
nor \U$1506 ( \3631 , \3629 , \3630 );
xnor \U$1507 ( \3632 , \3631 , \3115 );
and \U$1508 ( \3633 , \3110 , \3147 );
and \U$1509 ( \3634 , \3017 , \3145 );
nor \U$1510 ( \3635 , \3633 , \3634 );
xnor \U$1511 ( \3636 , \3635 , \3173 );
xor \U$1512 ( \3637 , \3632 , \3636 );
and \U$1513 ( \3638 , \3168 , \2848 );
and \U$1514 ( \3639 , \3077 , \2846 );
nor \U$1515 ( \3640 , \3638 , \3639 );
xnor \U$1516 ( \3641 , \3640 , \2853 );
xor \U$1517 ( \3642 , \3637 , \3641 );
xor \U$1518 ( \3643 , \3628 , \3642 );
xor \U$1519 ( \3644 , \3619 , \3643 );
xor \U$1520 ( \3645 , \3576 , \3644 );
and \U$1521 ( \3646 , \3408 , \3514 );
nor \U$1522 ( \3647 , \3645 , \3646 );
nor \U$1523 ( \3648 , \3572 , \3647 );
and \U$1524 ( \3649 , \3580 , \3618 );
and \U$1525 ( \3650 , \3618 , \3643 );
and \U$1526 ( \3651 , \3580 , \3643 );
or \U$1527 ( \3652 , \3649 , \3650 , \3651 );
and \U$1529 ( \3653 , \3584 , \3589 );
or \U$1531 ( \3654 , 1'b0 , \3653 , 1'b0 );
and \U$1532 ( \3655 , \3632 , \3636 );
and \U$1533 ( \3656 , \3636 , \3641 );
and \U$1534 ( \3657 , \3632 , \3641 );
or \U$1535 ( \3658 , \3655 , \3656 , \3657 );
xor \U$1536 ( \3659 , \3654 , \3658 );
and \U$1537 ( \3660 , \3594 , \3598 );
and \U$1538 ( \3661 , \3598 , \3602 );
and \U$1539 ( \3662 , \3594 , \3602 );
or \U$1540 ( \3663 , \3660 , \3661 , \3662 );
xor \U$1541 ( \3664 , \3659 , \3663 );
and \U$1542 ( \3665 , \3609 , \3613 );
and \U$1543 ( \3666 , \3613 , \3616 );
and \U$1544 ( \3667 , \3609 , \3616 );
or \U$1545 ( \3668 , \3665 , \3666 , \3667 );
xor \U$1547 ( \3669 , \3668 , 1'b0 );
and \U$1548 ( \3670 , \2673 , \2993 );
and \U$1549 ( \3671 , \2742 , \2990 );
nor \U$1550 ( \3672 , \3670 , \3671 );
xnor \U$1551 ( \3673 , \3672 , \2987 );
and \U$1552 ( \3674 , \2901 , \3029 );
and \U$1553 ( \3675 , \2769 , \3027 );
nor \U$1554 ( \3676 , \3674 , \3675 );
xnor \U$1555 ( \3677 , \3676 , \3055 );
xor \U$1556 ( \3678 , \3673 , \3677 );
and \U$1557 ( \3679 , \2924 , \3089 );
and \U$1558 ( \3680 , \2880 , \3087 );
nor \U$1559 ( \3681 , \3679 , \3680 );
xnor \U$1560 ( \3682 , \3681 , \3115 );
xor \U$1561 ( \3683 , \3678 , \3682 );
xor \U$1562 ( \3684 , \3669 , \3683 );
xor \U$1563 ( \3685 , \3664 , \3684 );
xor \U$1564 ( \3686 , \3652 , \3685 );
and \U$1565 ( \3687 , \3623 , \3627 );
and \U$1566 ( \3688 , \3627 , \3642 );
and \U$1567 ( \3689 , \3623 , \3642 );
or \U$1568 ( \3690 , \3687 , \3688 , \3689 );
and \U$1569 ( \3691 , \3590 , \3604 );
and \U$1570 ( \3692 , \3604 , \3617 );
and \U$1571 ( \3693 , \3590 , \3617 );
or \U$1572 ( \3694 , \3691 , \3692 , \3693 );
xor \U$1573 ( \3695 , \3690 , \3694 );
and \U$1575 ( \3696 , \3194 , \2721 );
and \U$1576 ( \3697 , \3215 , \2719 );
nor \U$1577 ( \3698 , \3696 , \3697 );
xnor \U$1578 ( \3699 , \3698 , \2747 );
and \U$1580 ( \3700 , \3260 , \2774 );
nor \U$1581 ( \3701 , 1'b0 , \3700 );
xnor \U$1582 ( \3702 , \3701 , 1'b0 );
xor \U$1583 ( \3703 , \3699 , \3702 );
xor \U$1585 ( \3704 , \3703 , 1'b0 );
xor \U$1586 ( \3705 , 1'b0 , \3704 );
and \U$1587 ( \3706 , \3017 , \3147 );
and \U$1588 ( \3707 , \3050 , \3145 );
nor \U$1589 ( \3708 , \3706 , \3707 );
xnor \U$1590 ( \3709 , \3708 , \3173 );
and \U$1591 ( \3710 , \3077 , \2848 );
and \U$1592 ( \3711 , \3110 , \2846 );
nor \U$1593 ( \3712 , \3710 , \3711 );
xnor \U$1594 ( \3713 , \3712 , \2853 );
xor \U$1595 ( \3714 , \3709 , \3713 );
and \U$1596 ( \3715 , \3139 , \2783 );
and \U$1597 ( \3716 , \3168 , \2781 );
nor \U$1598 ( \3717 , \3715 , \3716 );
xnor \U$1599 ( \3718 , \3717 , \2550 );
xor \U$1600 ( \3719 , \3714 , \3718 );
xor \U$1601 ( \3720 , \3705 , \3719 );
xor \U$1602 ( \3721 , \3695 , \3720 );
xor \U$1603 ( \3722 , \3686 , \3721 );
and \U$1604 ( \3723 , \3576 , \3644 );
nor \U$1605 ( \3724 , \3722 , \3723 );
and \U$1606 ( \3725 , \3690 , \3694 );
and \U$1607 ( \3726 , \3694 , \3720 );
and \U$1608 ( \3727 , \3690 , \3720 );
or \U$1609 ( \3728 , \3725 , \3726 , \3727 );
and \U$1610 ( \3729 , \3664 , \3684 );
xor \U$1611 ( \3730 , \3728 , \3729 );
and \U$1614 ( \3731 , \3668 , \3683 );
or \U$1615 ( \3732 , 1'b0 , 1'b0 , \3731 );
and \U$1617 ( \3733 , \3168 , \2783 );
and \U$1618 ( \3734 , \3077 , \2781 );
nor \U$1619 ( \3735 , \3733 , \3734 );
xnor \U$1620 ( \3736 , \3735 , \2550 );
and \U$1621 ( \3737 , \3215 , \2721 );
and \U$1622 ( \3738 , \3139 , \2719 );
nor \U$1623 ( \3739 , \3737 , \3738 );
xnor \U$1624 ( \3740 , \3739 , \2747 );
xor \U$1625 ( \3741 , \3736 , \3740 );
and \U$1627 ( \3742 , \3194 , \2774 );
nor \U$1628 ( \3743 , 1'b0 , \3742 );
xnor \U$1629 ( \3744 , \3743 , 1'b0 );
xor \U$1630 ( \3745 , \3741 , \3744 );
xor \U$1631 ( \3746 , 1'b0 , \3745 );
and \U$1632 ( \3747 , \2880 , \3089 );
and \U$1633 ( \3748 , \2901 , \3087 );
nor \U$1634 ( \3749 , \3747 , \3748 );
xnor \U$1635 ( \3750 , \3749 , \3115 );
and \U$1636 ( \3751 , \3050 , \3147 );
and \U$1637 ( \3752 , \2924 , \3145 );
nor \U$1638 ( \3753 , \3751 , \3752 );
xnor \U$1639 ( \3754 , \3753 , \3173 );
xor \U$1640 ( \3755 , \3750 , \3754 );
and \U$1641 ( \3756 , \3110 , \2848 );
and \U$1642 ( \3757 , \3017 , \2846 );
nor \U$1643 ( \3758 , \3756 , \3757 );
xnor \U$1644 ( \3759 , \3758 , \2853 );
xor \U$1645 ( \3760 , \3755 , \3759 );
xor \U$1646 ( \3761 , \3746 , \3760 );
and \U$1647 ( \3762 , \3673 , \3677 );
and \U$1648 ( \3763 , \3677 , \3682 );
and \U$1649 ( \3764 , \3673 , \3682 );
or \U$1650 ( \3765 , \3762 , \3763 , \3764 );
and \U$1651 ( \3766 , \3709 , \3713 );
and \U$1652 ( \3767 , \3713 , \3718 );
and \U$1653 ( \3768 , \3709 , \3718 );
or \U$1654 ( \3769 , \3766 , \3767 , \3768 );
xor \U$1655 ( \3770 , \3765 , \3769 );
and \U$1656 ( \3771 , \3699 , \3702 );
or \U$1659 ( \3772 , \3771 , 1'b0 , 1'b0 );
xor \U$1660 ( \3773 , \3770 , \3772 );
xor \U$1661 ( \3774 , \3761 , \3773 );
xor \U$1662 ( \3775 , \3732 , \3774 );
and \U$1663 ( \3776 , \3654 , \3658 );
and \U$1664 ( \3777 , \3658 , \3663 );
and \U$1665 ( \3778 , \3654 , \3663 );
or \U$1666 ( \3779 , \3776 , \3777 , \3778 );
and \U$1668 ( \3780 , \3704 , \3719 );
or \U$1670 ( \3781 , 1'b0 , \3780 , 1'b0 );
xor \U$1671 ( \3782 , \3779 , \3781 );
and \U$1673 ( \3783 , \2742 , \2993 );
not \U$1674 ( \3784 , \3783 );
xnor \U$1675 ( \3785 , \3784 , \2987 );
xor \U$1676 ( \3786 , 1'b0 , \3785 );
and \U$1677 ( \3787 , \2769 , \3029 );
and \U$1678 ( \3788 , \2673 , \3027 );
nor \U$1679 ( \3789 , \3787 , \3788 );
xnor \U$1680 ( \3790 , \3789 , \3055 );
xor \U$1681 ( \3791 , \3786 , \3790 );
xor \U$1682 ( \3792 , \3782 , \3791 );
xor \U$1683 ( \3793 , \3775 , \3792 );
xor \U$1684 ( \3794 , \3730 , \3793 );
and \U$1685 ( \3795 , \3652 , \3685 );
and \U$1686 ( \3796 , \3685 , \3721 );
and \U$1687 ( \3797 , \3652 , \3721 );
or \U$1688 ( \3798 , \3795 , \3796 , \3797 );
nor \U$1689 ( \3799 , \3794 , \3798 );
nor \U$1690 ( \3800 , \3724 , \3799 );
nand \U$1691 ( \3801 , \3648 , \3800 );
and \U$1692 ( \3802 , \3732 , \3774 );
and \U$1693 ( \3803 , \3774 , \3792 );
and \U$1694 ( \3804 , \3732 , \3792 );
or \U$1695 ( \3805 , \3802 , \3803 , \3804 );
and \U$1696 ( \3806 , \3765 , \3769 );
and \U$1697 ( \3807 , \3769 , \3772 );
and \U$1698 ( \3808 , \3765 , \3772 );
or \U$1699 ( \3809 , \3806 , \3807 , \3808 );
and \U$1701 ( \3810 , \3745 , \3760 );
or \U$1703 ( \3811 , 1'b0 , \3810 , 1'b0 );
xor \U$1704 ( \3812 , \3809 , \3811 );
and \U$1705 ( \3813 , \2924 , \3147 );
and \U$1706 ( \3814 , \2880 , \3145 );
nor \U$1707 ( \3815 , \3813 , \3814 );
xnor \U$1708 ( \3816 , \3815 , \3173 );
and \U$1709 ( \3817 , \3017 , \2848 );
and \U$1710 ( \3818 , \3050 , \2846 );
nor \U$1711 ( \3819 , \3817 , \3818 );
xnor \U$1712 ( \3820 , \3819 , \2853 );
xor \U$1713 ( \3821 , \3816 , \3820 );
and \U$1714 ( \3822 , \3077 , \2783 );
and \U$1715 ( \3823 , \3110 , \2781 );
nor \U$1716 ( \3824 , \3822 , \3823 );
xnor \U$1717 ( \3825 , \3824 , \2550 );
xor \U$1718 ( \3826 , \3821 , \3825 );
xor \U$1719 ( \3827 , \3812 , \3826 );
xor \U$1720 ( \3828 , \3805 , \3827 );
and \U$1721 ( \3829 , \3779 , \3781 );
and \U$1722 ( \3830 , \3781 , \3791 );
and \U$1723 ( \3831 , \3779 , \3791 );
or \U$1724 ( \3832 , \3829 , \3830 , \3831 );
and \U$1725 ( \3833 , \3761 , \3773 );
xor \U$1726 ( \3834 , \3832 , \3833 );
not \U$1727 ( \3835 , \2987 );
and \U$1728 ( \3836 , \2673 , \3029 );
and \U$1729 ( \3837 , \2742 , \3027 );
nor \U$1730 ( \3838 , \3836 , \3837 );
xnor \U$1731 ( \3839 , \3838 , \3055 );
xor \U$1732 ( \3840 , \3835 , \3839 );
and \U$1733 ( \3841 , \2901 , \3089 );
and \U$1734 ( \3842 , \2769 , \3087 );
nor \U$1735 ( \3843 , \3841 , \3842 );
xnor \U$1736 ( \3844 , \3843 , \3115 );
xor \U$1737 ( \3845 , \3840 , \3844 );
and \U$1739 ( \3846 , \3139 , \2721 );
and \U$1740 ( \3847 , \3168 , \2719 );
nor \U$1741 ( \3848 , \3846 , \3847 );
xnor \U$1742 ( \3849 , \3848 , \2747 );
and \U$1744 ( \3850 , \3215 , \2774 );
nor \U$1745 ( \3851 , 1'b0 , \3850 );
xnor \U$1746 ( \3852 , \3851 , 1'b0 );
xor \U$1747 ( \3853 , \3849 , \3852 );
xor \U$1749 ( \3854 , \3853 , 1'b0 );
xor \U$1750 ( \3855 , 1'b1 , \3854 );
xor \U$1751 ( \3856 , \3845 , \3855 );
and \U$1753 ( \3857 , \3785 , \3790 );
or \U$1755 ( \3858 , 1'b0 , \3857 , 1'b0 );
and \U$1756 ( \3859 , \3750 , \3754 );
and \U$1757 ( \3860 , \3754 , \3759 );
and \U$1758 ( \3861 , \3750 , \3759 );
or \U$1759 ( \3862 , \3859 , \3860 , \3861 );
xor \U$1760 ( \3863 , \3858 , \3862 );
and \U$1761 ( \3864 , \3736 , \3740 );
and \U$1762 ( \3865 , \3740 , \3744 );
and \U$1763 ( \3866 , \3736 , \3744 );
or \U$1764 ( \3867 , \3864 , \3865 , \3866 );
xor \U$1765 ( \3868 , \3863 , \3867 );
xor \U$1766 ( \3869 , \3856 , \3868 );
xor \U$1767 ( \3870 , \3834 , \3869 );
xor \U$1768 ( \3871 , \3828 , \3870 );
and \U$1769 ( \3872 , \3728 , \3729 );
and \U$1770 ( \3873 , \3729 , \3793 );
and \U$1771 ( \3874 , \3728 , \3793 );
or \U$1772 ( \3875 , \3872 , \3873 , \3874 );
nor \U$1773 ( \3876 , \3871 , \3875 );
and \U$1774 ( \3877 , \3832 , \3833 );
and \U$1775 ( \3878 , \3833 , \3869 );
and \U$1776 ( \3879 , \3832 , \3869 );
or \U$1777 ( \3880 , \3877 , \3878 , \3879 );
and \U$1778 ( \3881 , \3835 , \3839 );
and \U$1779 ( \3882 , \3839 , \3844 );
and \U$1780 ( \3883 , \3835 , \3844 );
or \U$1781 ( \3884 , \3881 , \3882 , \3883 );
and \U$1782 ( \3885 , \3816 , \3820 );
and \U$1783 ( \3886 , \3820 , \3825 );
and \U$1784 ( \3887 , \3816 , \3825 );
or \U$1785 ( \3888 , \3885 , \3886 , \3887 );
xor \U$1786 ( \3889 , \3884 , \3888 );
and \U$1787 ( \3890 , \3849 , \3852 );
or \U$1790 ( \3891 , \3890 , 1'b0 , 1'b0 );
xor \U$1791 ( \3892 , \3889 , \3891 );
and \U$1792 ( \3893 , \3858 , \3862 );
and \U$1793 ( \3894 , \3862 , \3867 );
and \U$1794 ( \3895 , \3858 , \3867 );
or \U$1795 ( \3896 , \3893 , \3894 , \3895 );
and \U$1798 ( \3897 , 1'b1 , \3854 );
or \U$1800 ( \3898 , 1'b0 , \3897 , 1'b0 );
xor \U$1801 ( \3899 , \3896 , \3898 );
and \U$1802 ( \3900 , \3168 , \2721 );
and \U$1803 ( \3901 , \3077 , \2719 );
nor \U$1804 ( \3902 , \3900 , \3901 );
xnor \U$1805 ( \3903 , \3902 , \2747 );
and \U$1807 ( \3904 , \3139 , \2774 );
nor \U$1808 ( \3905 , 1'b0 , \3904 );
xnor \U$1809 ( \3906 , \3905 , 1'b0 );
xor \U$1810 ( \3907 , \3903 , \3906 );
xor \U$1812 ( \3908 , \3907 , 1'b0 );
and \U$1813 ( \3909 , \2880 , \3147 );
and \U$1814 ( \3910 , \2901 , \3145 );
nor \U$1815 ( \3911 , \3909 , \3910 );
xnor \U$1816 ( \3912 , \3911 , \3173 );
and \U$1817 ( \3913 , \3050 , \2848 );
and \U$1818 ( \3914 , \2924 , \2846 );
nor \U$1819 ( \3915 , \3913 , \3914 );
xnor \U$1820 ( \3916 , \3915 , \2853 );
xor \U$1821 ( \3917 , \3912 , \3916 );
and \U$1822 ( \3918 , \3110 , \2783 );
and \U$1823 ( \3919 , \3017 , \2781 );
nor \U$1824 ( \3920 , \3918 , \3919 );
xnor \U$1825 ( \3921 , \3920 , \2550 );
xor \U$1826 ( \3922 , \3917 , \3921 );
xor \U$1827 ( \3923 , \3908 , \3922 );
and \U$1829 ( \3924 , \2742 , \3029 );
not \U$1830 ( \3925 , \3924 );
xnor \U$1831 ( \3926 , \3925 , \3055 );
xor \U$1832 ( \3927 , 1'b0 , \3926 );
and \U$1833 ( \3928 , \2769 , \3089 );
and \U$1834 ( \3929 , \2673 , \3087 );
nor \U$1835 ( \3930 , \3928 , \3929 );
xnor \U$1836 ( \3931 , \3930 , \3115 );
xor \U$1837 ( \3932 , \3927 , \3931 );
xor \U$1838 ( \3933 , \3923 , \3932 );
xor \U$1839 ( \3934 , \3899 , \3933 );
xor \U$1840 ( \3935 , \3892 , \3934 );
xor \U$1841 ( \3936 , \3880 , \3935 );
and \U$1842 ( \3937 , \3809 , \3811 );
and \U$1843 ( \3938 , \3811 , \3826 );
and \U$1844 ( \3939 , \3809 , \3826 );
or \U$1845 ( \3940 , \3937 , \3938 , \3939 );
and \U$1846 ( \3941 , \3845 , \3855 );
and \U$1847 ( \3942 , \3855 , \3868 );
and \U$1848 ( \3943 , \3845 , \3868 );
or \U$1849 ( \3944 , \3941 , \3942 , \3943 );
xor \U$1850 ( \3945 , \3940 , \3944 );
xor \U$1852 ( \3946 , \3945 , 1'b1 );
xor \U$1853 ( \3947 , \3936 , \3946 );
and \U$1854 ( \3948 , \3805 , \3827 );
and \U$1855 ( \3949 , \3827 , \3870 );
and \U$1856 ( \3950 , \3805 , \3870 );
or \U$1857 ( \3951 , \3948 , \3949 , \3950 );
nor \U$1858 ( \3952 , \3947 , \3951 );
nor \U$1859 ( \3953 , \3876 , \3952 );
and \U$1860 ( \3954 , \3940 , \3944 );
and \U$1861 ( \3955 , \3944 , 1'b1 );
and \U$1862 ( \3956 , \3940 , 1'b1 );
or \U$1863 ( \3957 , \3954 , \3955 , \3956 );
and \U$1864 ( \3958 , \3892 , \3934 );
xor \U$1865 ( \3959 , \3957 , \3958 );
and \U$1866 ( \3960 , \3896 , \3898 );
and \U$1867 ( \3961 , \3898 , \3933 );
and \U$1868 ( \3962 , \3896 , \3933 );
or \U$1869 ( \3963 , \3960 , \3961 , \3962 );
and \U$1871 ( \3964 , \3168 , \2774 );
nor \U$1872 ( \3965 , 1'b0 , \3964 );
xnor \U$1873 ( \3966 , \3965 , 1'b0 );
xor \U$1875 ( \3967 , \3966 , 1'b0 );
xor \U$1877 ( \3968 , \3967 , 1'b0 );
and \U$1878 ( \3969 , \2924 , \2848 );
and \U$1879 ( \3970 , \2880 , \2846 );
nor \U$1880 ( \3971 , \3969 , \3970 );
xnor \U$1881 ( \3972 , \3971 , \2853 );
and \U$1882 ( \3973 , \3017 , \2783 );
and \U$1883 ( \3974 , \3050 , \2781 );
nor \U$1884 ( \3975 , \3973 , \3974 );
xnor \U$1885 ( \3976 , \3975 , \2550 );
xor \U$1886 ( \3977 , \3972 , \3976 );
and \U$1887 ( \3978 , \3077 , \2721 );
and \U$1888 ( \3979 , \3110 , \2719 );
nor \U$1889 ( \3980 , \3978 , \3979 );
xnor \U$1890 ( \3981 , \3980 , \2747 );
xor \U$1891 ( \3982 , \3977 , \3981 );
xor \U$1892 ( \3983 , \3968 , \3982 );
not \U$1893 ( \3984 , \3055 );
and \U$1894 ( \3985 , \2673 , \3089 );
and \U$1895 ( \3986 , \2742 , \3087 );
nor \U$1896 ( \3987 , \3985 , \3986 );
xnor \U$1897 ( \3988 , \3987 , \3115 );
xor \U$1898 ( \3989 , \3984 , \3988 );
and \U$1899 ( \3990 , \2901 , \3147 );
and \U$1900 ( \3991 , \2769 , \3145 );
nor \U$1901 ( \3992 , \3990 , \3991 );
xnor \U$1902 ( \3993 , \3992 , \3173 );
xor \U$1903 ( \3994 , \3989 , \3993 );
xor \U$1904 ( \3995 , \3983 , \3994 );
xor \U$1906 ( \3996 , \3995 , 1'b0 );
and \U$1908 ( \3997 , \3926 , \3931 );
or \U$1910 ( \3998 , 1'b0 , \3997 , 1'b0 );
and \U$1911 ( \3999 , \3912 , \3916 );
and \U$1912 ( \4000 , \3916 , \3921 );
and \U$1913 ( \4001 , \3912 , \3921 );
or \U$1914 ( \4002 , \3999 , \4000 , \4001 );
xor \U$1915 ( \4003 , \3998 , \4002 );
and \U$1916 ( \4004 , \3903 , \3906 );
or \U$1919 ( \4005 , \4004 , 1'b0 , 1'b0 );
xor \U$1920 ( \4006 , \4003 , \4005 );
xor \U$1921 ( \4007 , \3996 , \4006 );
xor \U$1922 ( \4008 , \3963 , \4007 );
and \U$1923 ( \4009 , \3884 , \3888 );
and \U$1924 ( \4010 , \3888 , \3891 );
and \U$1925 ( \4011 , \3884 , \3891 );
or \U$1926 ( \4012 , \4009 , \4010 , \4011 );
xor \U$1928 ( \4013 , \4012 , 1'b0 );
and \U$1929 ( \4014 , \3908 , \3922 );
and \U$1930 ( \4015 , \3922 , \3932 );
and \U$1931 ( \4016 , \3908 , \3932 );
or \U$1932 ( \4017 , \4014 , \4015 , \4016 );
xor \U$1933 ( \4018 , \4013 , \4017 );
xor \U$1934 ( \4019 , \4008 , \4018 );
xor \U$1935 ( \4020 , \3959 , \4019 );
and \U$1936 ( \4021 , \3880 , \3935 );
and \U$1937 ( \4022 , \3935 , \3946 );
and \U$1938 ( \4023 , \3880 , \3946 );
or \U$1939 ( \4024 , \4021 , \4022 , \4023 );
nor \U$1940 ( \4025 , \4020 , \4024 );
and \U$1941 ( \4026 , \3963 , \4007 );
and \U$1942 ( \4027 , \4007 , \4018 );
and \U$1943 ( \4028 , \3963 , \4018 );
or \U$1944 ( \4029 , \4026 , \4027 , \4028 );
and \U$1945 ( \4030 , \3998 , \4002 );
and \U$1946 ( \4031 , \4002 , \4005 );
and \U$1947 ( \4032 , \3998 , \4005 );
or \U$1948 ( \4033 , \4030 , \4031 , \4032 );
xor \U$1950 ( \4034 , \4033 , 1'b0 );
and \U$1951 ( \4035 , \3968 , \3982 );
and \U$1952 ( \4036 , \3982 , \3994 );
and \U$1953 ( \4037 , \3968 , \3994 );
or \U$1954 ( \4038 , \4035 , \4036 , \4037 );
xor \U$1955 ( \4039 , \4034 , \4038 );
xor \U$1956 ( \4040 , \4029 , \4039 );
and \U$1959 ( \4041 , \4012 , \4017 );
or \U$1960 ( \4042 , 1'b0 , 1'b0 , \4041 );
and \U$1963 ( \4043 , \3995 , \4006 );
or \U$1964 ( \4044 , 1'b0 , 1'b0 , \4043 );
xor \U$1965 ( \4045 , \4042 , \4044 );
and \U$1966 ( \4046 , \2880 , \2848 );
and \U$1967 ( \4047 , \2901 , \2846 );
nor \U$1968 ( \4048 , \4046 , \4047 );
xnor \U$1969 ( \4049 , \4048 , \2853 );
and \U$1970 ( \4050 , \3050 , \2783 );
and \U$1971 ( \4051 , \2924 , \2781 );
nor \U$1972 ( \4052 , \4050 , \4051 );
xnor \U$1973 ( \4053 , \4052 , \2550 );
xor \U$1974 ( \4054 , \4049 , \4053 );
and \U$1975 ( \4055 , \3110 , \2721 );
and \U$1976 ( \4056 , \3017 , \2719 );
nor \U$1977 ( \4057 , \4055 , \4056 );
xnor \U$1978 ( \4058 , \4057 , \2747 );
xor \U$1979 ( \4059 , \4054 , \4058 );
and \U$1981 ( \4060 , \2742 , \3089 );
not \U$1982 ( \4061 , \4060 );
xnor \U$1983 ( \4062 , \4061 , \3115 );
xor \U$1984 ( \4063 , 1'b0 , \4062 );
and \U$1985 ( \4064 , \2769 , \3147 );
and \U$1986 ( \4065 , \2673 , \3145 );
nor \U$1987 ( \4066 , \4064 , \4065 );
xnor \U$1988 ( \4067 , \4066 , \3173 );
xor \U$1989 ( \4068 , \4063 , \4067 );
xor \U$1990 ( \4069 , \4059 , \4068 );
and \U$1993 ( \4070 , \3077 , \2774 );
nor \U$1994 ( \4071 , 1'b0 , \4070 );
xnor \U$1995 ( \4072 , \4071 , 1'b0 );
xor \U$1997 ( \4073 , \4072 , 1'b0 );
xor \U$1999 ( \4074 , \4073 , 1'b0 );
xnor \U$2000 ( \4075 , 1'b0 , \4074 );
xor \U$2001 ( \4076 , \4069 , \4075 );
and \U$2002 ( \4077 , \3984 , \3988 );
and \U$2003 ( \4078 , \3988 , \3993 );
and \U$2004 ( \4079 , \3984 , \3993 );
or \U$2005 ( \4080 , \4077 , \4078 , \4079 );
and \U$2006 ( \4081 , \3972 , \3976 );
and \U$2007 ( \4082 , \3976 , \3981 );
and \U$2008 ( \4083 , \3972 , \3981 );
or \U$2009 ( \4084 , \4081 , \4082 , \4083 );
xor \U$2010 ( \4085 , \4080 , \4084 );
xor \U$2012 ( \4086 , \4085 , 1'b0 );
xor \U$2013 ( \4087 , \4076 , \4086 );
xor \U$2014 ( \4088 , \4045 , \4087 );
xor \U$2015 ( \4089 , \4040 , \4088 );
and \U$2016 ( \4090 , \3957 , \3958 );
and \U$2017 ( \4091 , \3958 , \4019 );
and \U$2018 ( \4092 , \3957 , \4019 );
or \U$2019 ( \4093 , \4090 , \4091 , \4092 );
nor \U$2020 ( \4094 , \4089 , \4093 );
nor \U$2021 ( \4095 , \4025 , \4094 );
nand \U$2022 ( \4096 , \3953 , \4095 );
nor \U$2023 ( \4097 , \3801 , \4096 );
and \U$2024 ( \4098 , \4042 , \4044 );
and \U$2025 ( \4099 , \4044 , \4087 );
and \U$2026 ( \4100 , \4042 , \4087 );
or \U$2027 ( \4101 , \4098 , \4099 , \4100 );
and \U$2028 ( \4102 , \4080 , \4084 );
or \U$2031 ( \4103 , \4102 , 1'b0 , 1'b0 );
or \U$2032 ( \4104 , 1'b0 , \4074 );
xor \U$2033 ( \4105 , \4103 , \4104 );
and \U$2034 ( \4106 , \4059 , \4068 );
xor \U$2035 ( \4107 , \4105 , \4106 );
xor \U$2036 ( \4108 , \4101 , \4107 );
and \U$2039 ( \4109 , \4033 , \4038 );
or \U$2040 ( \4110 , 1'b0 , 1'b0 , \4109 );
and \U$2041 ( \4111 , \4069 , \4075 );
and \U$2042 ( \4112 , \4075 , \4086 );
and \U$2043 ( \4113 , \4069 , \4086 );
or \U$2044 ( \4114 , \4111 , \4112 , \4113 );
xor \U$2045 ( \4115 , \4110 , \4114 );
and \U$2047 ( \4116 , \2924 , \2783 );
and \U$2048 ( \4117 , \2880 , \2781 );
nor \U$2049 ( \4118 , \4116 , \4117 );
xnor \U$2050 ( \4119 , \4118 , \2550 );
and \U$2051 ( \4120 , \3017 , \2721 );
and \U$2052 ( \4121 , \3050 , \2719 );
nor \U$2053 ( \4122 , \4120 , \4121 );
xnor \U$2054 ( \4123 , \4122 , \2747 );
xor \U$2055 ( \4124 , \4119 , \4123 );
and \U$2057 ( \4125 , \3110 , \2774 );
nor \U$2058 ( \4126 , 1'b0 , \4125 );
xnor \U$2059 ( \4127 , \4126 , 1'b0 );
xor \U$2060 ( \4128 , \4124 , \4127 );
xor \U$2061 ( \4129 , 1'b0 , \4128 );
not \U$2062 ( \4130 , \3115 );
and \U$2063 ( \4131 , \2673 , \3147 );
and \U$2064 ( \4132 , \2742 , \3145 );
nor \U$2065 ( \4133 , \4131 , \4132 );
xnor \U$2066 ( \4134 , \4133 , \3173 );
xor \U$2067 ( \4135 , \4130 , \4134 );
and \U$2068 ( \4136 , \2901 , \2848 );
and \U$2069 ( \4137 , \2769 , \2846 );
nor \U$2070 ( \4138 , \4136 , \4137 );
xnor \U$2071 ( \4139 , \4138 , \2853 );
xor \U$2072 ( \4140 , \4135 , \4139 );
xor \U$2073 ( \4141 , \4129 , \4140 );
xor \U$2075 ( \4142 , \4141 , 1'b0 );
and \U$2077 ( \4143 , \4062 , \4067 );
or \U$2079 ( \4144 , 1'b0 , \4143 , 1'b0 );
and \U$2080 ( \4145 , \4049 , \4053 );
and \U$2081 ( \4146 , \4053 , \4058 );
and \U$2082 ( \4147 , \4049 , \4058 );
or \U$2083 ( \4148 , \4145 , \4146 , \4147 );
xor \U$2084 ( \4149 , \4144 , \4148 );
xor \U$2086 ( \4150 , \4149 , 1'b0 );
xor \U$2087 ( \4151 , \4142 , \4150 );
xor \U$2088 ( \4152 , \4115 , \4151 );
xor \U$2089 ( \4153 , \4108 , \4152 );
and \U$2090 ( \4154 , \4029 , \4039 );
and \U$2091 ( \4155 , \4039 , \4088 );
and \U$2092 ( \4156 , \4029 , \4088 );
or \U$2093 ( \4157 , \4154 , \4155 , \4156 );
nor \U$2094 ( \4158 , \4153 , \4157 );
and \U$2095 ( \4159 , \4110 , \4114 );
and \U$2096 ( \4160 , \4114 , \4151 );
and \U$2097 ( \4161 , \4110 , \4151 );
or \U$2098 ( \4162 , \4159 , \4160 , \4161 );
and \U$2099 ( \4163 , \4144 , \4148 );
or \U$2102 ( \4164 , \4163 , 1'b0 , 1'b0 );
xor \U$2104 ( \4165 , \4164 , 1'b0 );
and \U$2106 ( \4166 , \4128 , \4140 );
or \U$2108 ( \4167 , 1'b0 , \4166 , 1'b0 );
xor \U$2109 ( \4168 , \4165 , \4167 );
xor \U$2110 ( \4169 , \4162 , \4168 );
and \U$2111 ( \4170 , \4103 , \4104 );
and \U$2112 ( \4171 , \4104 , \4106 );
and \U$2113 ( \4172 , \4103 , \4106 );
or \U$2114 ( \4173 , \4170 , \4171 , \4172 );
and \U$2117 ( \4174 , \4141 , \4150 );
or \U$2118 ( \4175 , 1'b0 , 1'b0 , \4174 );
xor \U$2119 ( \4176 , \4173 , \4175 );
and \U$2120 ( \4177 , \2880 , \2783 );
and \U$2121 ( \4178 , \2901 , \2781 );
nor \U$2122 ( \4179 , \4177 , \4178 );
xnor \U$2123 ( \4180 , \4179 , \2550 );
and \U$2124 ( \4181 , \3050 , \2721 );
and \U$2125 ( \4182 , \2924 , \2719 );
nor \U$2126 ( \4183 , \4181 , \4182 );
xnor \U$2127 ( \4184 , \4183 , \2747 );
xor \U$2128 ( \4185 , \4180 , \4184 );
and \U$2130 ( \4186 , \3017 , \2774 );
nor \U$2131 ( \4187 , 1'b0 , \4186 );
xnor \U$2132 ( \4188 , \4187 , 1'b0 );
xor \U$2133 ( \4189 , \4185 , \4188 );
and \U$2135 ( \4190 , \2742 , \3147 );
not \U$2136 ( \4191 , \4190 );
xnor \U$2137 ( \4192 , \4191 , \3173 );
xor \U$2138 ( \4193 , 1'b0 , \4192 );
and \U$2139 ( \4194 , \2769 , \2848 );
and \U$2140 ( \4195 , \2673 , \2846 );
nor \U$2141 ( \4196 , \4194 , \4195 );
xnor \U$2142 ( \4197 , \4196 , \2853 );
xor \U$2143 ( \4198 , \4193 , \4197 );
xor \U$2144 ( \4199 , \4189 , \4198 );
xor \U$2146 ( \4200 , \4199 , 1'b1 );
and \U$2147 ( \4201 , \4130 , \4134 );
and \U$2148 ( \4202 , \4134 , \4139 );
and \U$2149 ( \4203 , \4130 , \4139 );
or \U$2150 ( \4204 , \4201 , \4202 , \4203 );
and \U$2151 ( \4205 , \4119 , \4123 );
and \U$2152 ( \4206 , \4123 , \4127 );
and \U$2153 ( \4207 , \4119 , \4127 );
or \U$2154 ( \4208 , \4205 , \4206 , \4207 );
xor \U$2155 ( \4209 , \4204 , \4208 );
xor \U$2157 ( \4210 , \4209 , 1'b0 );
xor \U$2158 ( \4211 , \4200 , \4210 );
xor \U$2159 ( \4212 , \4176 , \4211 );
xor \U$2160 ( \4213 , \4169 , \4212 );
and \U$2161 ( \4214 , \4101 , \4107 );
and \U$2162 ( \4215 , \4107 , \4152 );
and \U$2163 ( \4216 , \4101 , \4152 );
or \U$2164 ( \4217 , \4214 , \4215 , \4216 );
nor \U$2165 ( \4218 , \4213 , \4217 );
nor \U$2166 ( \4219 , \4158 , \4218 );
and \U$2167 ( \4220 , \4173 , \4175 );
and \U$2168 ( \4221 , \4175 , \4211 );
and \U$2169 ( \4222 , \4173 , \4211 );
or \U$2170 ( \4223 , \4220 , \4221 , \4222 );
and \U$2171 ( \4224 , \4204 , \4208 );
or \U$2174 ( \4225 , \4224 , 1'b0 , 1'b0 );
xor \U$2176 ( \4226 , \4225 , 1'b0 );
and \U$2177 ( \4227 , \4189 , \4198 );
xor \U$2178 ( \4228 , \4226 , \4227 );
xor \U$2179 ( \4229 , \4223 , \4228 );
and \U$2182 ( \4230 , \4164 , \4167 );
or \U$2183 ( \4231 , 1'b0 , 1'b0 , \4230 );
and \U$2184 ( \4232 , \4199 , 1'b1 );
and \U$2185 ( \4233 , 1'b1 , \4210 );
and \U$2186 ( \4234 , \4199 , \4210 );
or \U$2187 ( \4235 , \4232 , \4233 , \4234 );
xor \U$2188 ( \4236 , \4231 , \4235 );
and \U$2190 ( \4237 , \2924 , \2721 );
and \U$2191 ( \4238 , \2880 , \2719 );
nor \U$2192 ( \4239 , \4237 , \4238 );
xnor \U$2193 ( \4240 , \4239 , \2747 );
and \U$2195 ( \4241 , \3050 , \2774 );
nor \U$2196 ( \4242 , 1'b0 , \4241 );
xnor \U$2197 ( \4243 , \4242 , 1'b0 );
xor \U$2198 ( \4244 , \4240 , \4243 );
xor \U$2200 ( \4245 , \4244 , 1'b0 );
xor \U$2201 ( \4246 , 1'b0 , \4245 );
not \U$2202 ( \4247 , \3173 );
and \U$2203 ( \4248 , \2673 , \2848 );
and \U$2204 ( \4249 , \2742 , \2846 );
nor \U$2205 ( \4250 , \4248 , \4249 );
xnor \U$2206 ( \4251 , \4250 , \2853 );
xor \U$2207 ( \4252 , \4247 , \4251 );
and \U$2208 ( \4253 , \2901 , \2783 );
and \U$2209 ( \4254 , \2769 , \2781 );
nor \U$2210 ( \4255 , \4253 , \4254 );
xnor \U$2211 ( \4256 , \4255 , \2550 );
xor \U$2212 ( \4257 , \4252 , \4256 );
xor \U$2213 ( \4258 , \4246 , \4257 );
xor \U$2215 ( \4259 , \4258 , 1'b0 );
and \U$2217 ( \4260 , \4192 , \4197 );
or \U$2219 ( \4261 , 1'b0 , \4260 , 1'b0 );
and \U$2220 ( \4262 , \4180 , \4184 );
and \U$2221 ( \4263 , \4184 , \4188 );
and \U$2222 ( \4264 , \4180 , \4188 );
or \U$2223 ( \4265 , \4262 , \4263 , \4264 );
xor \U$2224 ( \4266 , \4261 , \4265 );
xor \U$2226 ( \4267 , \4266 , 1'b0 );
xor \U$2227 ( \4268 , \4259 , \4267 );
xor \U$2228 ( \4269 , \4236 , \4268 );
xor \U$2229 ( \4270 , \4229 , \4269 );
and \U$2230 ( \4271 , \4162 , \4168 );
and \U$2231 ( \4272 , \4168 , \4212 );
and \U$2232 ( \4273 , \4162 , \4212 );
or \U$2233 ( \4274 , \4271 , \4272 , \4273 );
nor \U$2234 ( \4275 , \4270 , \4274 );
and \U$2235 ( \4276 , \4231 , \4235 );
and \U$2236 ( \4277 , \4235 , \4268 );
and \U$2237 ( \4278 , \4231 , \4268 );
or \U$2238 ( \4279 , \4276 , \4277 , \4278 );
and \U$2239 ( \4280 , \4261 , \4265 );
or \U$2242 ( \4281 , \4280 , 1'b0 , 1'b0 );
xor \U$2244 ( \4282 , \4281 , 1'b0 );
and \U$2246 ( \4283 , \4245 , \4257 );
or \U$2248 ( \4284 , 1'b0 , \4283 , 1'b0 );
xor \U$2249 ( \4285 , \4282 , \4284 );
xor \U$2250 ( \4286 , \4279 , \4285 );
and \U$2253 ( \4287 , \4225 , \4227 );
or \U$2254 ( \4288 , 1'b0 , 1'b0 , \4287 );
and \U$2257 ( \4289 , \4258 , \4267 );
or \U$2258 ( \4290 , 1'b0 , 1'b0 , \4289 );
xor \U$2259 ( \4291 , \4288 , \4290 );
xor \U$2260 ( \4292 , \2904 , \2927 );
xor \U$2262 ( \4293 , \4292 , 1'b0 );
xor \U$2264 ( \4294 , 1'b0 , \2854 );
xor \U$2265 ( \4295 , \4294 , \2858 );
xor \U$2266 ( \4296 , \4293 , \4295 );
xor \U$2268 ( \4297 , \4296 , 1'b1 );
and \U$2269 ( \4298 , \4247 , \4251 );
and \U$2270 ( \4299 , \4251 , \4256 );
and \U$2271 ( \4300 , \4247 , \4256 );
or \U$2272 ( \4301 , \4298 , \4299 , \4300 );
and \U$2273 ( \4302 , \4240 , \4243 );
or \U$2276 ( \4303 , \4302 , 1'b0 , 1'b0 );
xor \U$2277 ( \4304 , \4301 , \4303 );
xor \U$2279 ( \4305 , \4304 , 1'b0 );
xor \U$2280 ( \4306 , \4297 , \4305 );
xor \U$2281 ( \4307 , \4291 , \4306 );
xor \U$2282 ( \4308 , \4286 , \4307 );
and \U$2283 ( \4309 , \4223 , \4228 );
and \U$2284 ( \4310 , \4228 , \4269 );
and \U$2285 ( \4311 , \4223 , \4269 );
or \U$2286 ( \4312 , \4309 , \4310 , \4311 );
nor \U$2287 ( \4313 , \4308 , \4312 );
nor \U$2288 ( \4314 , \4275 , \4313 );
nand \U$2289 ( \4315 , \4219 , \4314 );
and \U$2290 ( \4316 , \4288 , \4290 );
and \U$2291 ( \4317 , \4290 , \4306 );
and \U$2292 ( \4318 , \4288 , \4306 );
or \U$2293 ( \4319 , \4316 , \4317 , \4318 );
and \U$2294 ( \4320 , \4301 , \4303 );
or \U$2297 ( \4321 , \4320 , 1'b0 , 1'b0 );
xor \U$2299 ( \4322 , \4321 , 1'b0 );
and \U$2300 ( \4323 , \4293 , \4295 );
xor \U$2301 ( \4324 , \4322 , \4323 );
xor \U$2302 ( \4325 , \4319 , \4324 );
and \U$2305 ( \4326 , \4281 , \4284 );
or \U$2306 ( \4327 , 1'b0 , 1'b0 , \4326 );
and \U$2307 ( \4328 , \4296 , 1'b1 );
and \U$2308 ( \4329 , 1'b1 , \4305 );
and \U$2309 ( \4330 , \4296 , \4305 );
or \U$2310 ( \4331 , \4328 , \4329 , \4330 );
xor \U$2311 ( \4332 , \4327 , \4331 );
xor \U$2313 ( \4333 , 1'b0 , \2936 );
xor \U$2314 ( \4334 , \4333 , \2947 );
xor \U$2316 ( \4335 , \4334 , 1'b0 );
xor \U$2317 ( \4336 , \2860 , \2929 );
xor \U$2319 ( \4337 , \4336 , 1'b0 );
xor \U$2320 ( \4338 , \4335 , \4337 );
xor \U$2321 ( \4339 , \4332 , \4338 );
xor \U$2322 ( \4340 , \4325 , \4339 );
and \U$2323 ( \4341 , \4279 , \4285 );
and \U$2324 ( \4342 , \4285 , \4307 );
and \U$2325 ( \4343 , \4279 , \4307 );
or \U$2326 ( \4344 , \4341 , \4342 , \4343 );
nor \U$2327 ( \4345 , \4340 , \4344 );
and \U$2328 ( \4346 , \4327 , \4331 );
and \U$2329 ( \4347 , \4331 , \4338 );
and \U$2330 ( \4348 , \4327 , \4338 );
or \U$2331 ( \4349 , \4346 , \4347 , \4348 );
xor \U$2333 ( \4350 , \2931 , 1'b0 );
xor \U$2334 ( \4351 , \4350 , \2949 );
xor \U$2335 ( \4352 , \4349 , \4351 );
and \U$2338 ( \4353 , \4321 , \4323 );
or \U$2339 ( \4354 , 1'b0 , 1'b0 , \4353 );
and \U$2342 ( \4355 , \4334 , \4337 );
or \U$2343 ( \4356 , 1'b0 , 1'b0 , \4355 );
xor \U$2344 ( \4357 , \4354 , \4356 );
xor \U$2345 ( \4358 , \2959 , 1'b1 );
xor \U$2346 ( \4359 , \4358 , \2966 );
xor \U$2347 ( \4360 , \4357 , \4359 );
xor \U$2348 ( \4361 , \4352 , \4360 );
and \U$2349 ( \4362 , \4319 , \4324 );
and \U$2350 ( \4363 , \4324 , \4339 );
and \U$2351 ( \4364 , \4319 , \4339 );
or \U$2352 ( \4365 , \4362 , \4363 , \4364 );
nor \U$2353 ( \4366 , \4361 , \4365 );
nor \U$2354 ( \4367 , \4345 , \4366 );
and \U$2355 ( \4368 , \4354 , \4356 );
and \U$2356 ( \4369 , \4356 , \4359 );
and \U$2357 ( \4370 , \4354 , \4359 );
or \U$2358 ( \4371 , \4368 , \4369 , \4370 );
and \U$2360 ( \4372 , \2956 , \2958 );
xor \U$2361 ( \4373 , 1'b0 , \4372 );
xor \U$2362 ( \4374 , \4371 , \4373 );
xor \U$2363 ( \4375 , \2951 , \2969 );
xor \U$2364 ( \4376 , \4375 , \2972 );
xor \U$2365 ( \4377 , \4374 , \4376 );
and \U$2366 ( \4378 , \4349 , \4351 );
and \U$2367 ( \4379 , \4351 , \4360 );
and \U$2368 ( \4380 , \4349 , \4360 );
or \U$2369 ( \4381 , \4378 , \4379 , \4380 );
nor \U$2370 ( \4382 , \4377 , \4381 );
xor \U$2372 ( \4383 , \2975 , 1'b0 );
xor \U$2373 ( \4384 , \4383 , \2977 );
and \U$2374 ( \4385 , \4371 , \4373 );
and \U$2375 ( \4386 , \4373 , \4376 );
and \U$2376 ( \4387 , \4371 , \4376 );
or \U$2377 ( \4388 , \4385 , \4386 , \4387 );
nor \U$2378 ( \4389 , \4384 , \4388 );
nor \U$2379 ( \4390 , \4382 , \4389 );
nand \U$2380 ( \4391 , \4367 , \4390 );
nor \U$2381 ( \4392 , \4315 , \4391 );
nand \U$2382 ( \4393 , \4097 , \4392 );
and \U$2383 ( \4394 , \3194 , \2993 );
and \U$2384 ( \4395 , \3215 , \2990 );
nor \U$2385 ( \4396 , \4394 , \4395 );
xnor \U$2386 ( \4397 , \4396 , \2987 );
and \U$2387 ( \4398 , \3239 , \3029 );
and \U$2388 ( \4399 , \3260 , \3027 );
nor \U$2389 ( \4400 , \4398 , \4399 );
xnor \U$2390 ( \4401 , \4400 , \3055 );
and \U$2391 ( \4402 , \4397 , \4401 );
and \U$2392 ( \4403 , \3287 , \3089 );
and \U$2393 ( \4404 , \3308 , \3087 );
nor \U$2394 ( \4405 , \4403 , \4404 );
xnor \U$2395 ( \4406 , \4405 , \3115 );
and \U$2396 ( \4407 , \4401 , \4406 );
and \U$2397 ( \4408 , \4397 , \4406 );
or \U$2398 ( \4409 , \4402 , \4407 , \4408 );
and \U$2399 ( \4410 , \3308 , \3089 );
and \U$2400 ( \4411 , \3239 , \3087 );
nor \U$2401 ( \4412 , \4410 , \4411 );
xnor \U$2402 ( \4413 , \4412 , \3115 );
and \U$2403 ( \4414 , \3331 , \3147 );
and \U$2404 ( \4415 , \3287 , \3145 );
nor \U$2405 ( \4416 , \4414 , \4415 );
xnor \U$2406 ( \4417 , \4416 , \3173 );
xor \U$2407 ( \4418 , \4413 , \4417 );
nand \U$2408 ( \4419 , \3464 , \2846 );
xnor \U$2409 ( \4420 , \4419 , \2853 );
xor \U$2410 ( \4421 , \4418 , \4420 );
and \U$2411 ( \4422 , \4409 , \4421 );
and \U$2412 ( \4423 , \3215 , \2993 );
and \U$2413 ( \4424 , \3139 , \2990 );
nor \U$2414 ( \4425 , \4423 , \4424 );
xnor \U$2415 ( \4426 , \4425 , \2987 );
xor \U$2416 ( \4427 , \2853 , \4426 );
and \U$2417 ( \4428 , \3260 , \3029 );
and \U$2418 ( \4429 , \3194 , \3027 );
nor \U$2419 ( \4430 , \4428 , \4429 );
xnor \U$2420 ( \4431 , \4430 , \3055 );
xor \U$2421 ( \4432 , \4427 , \4431 );
and \U$2422 ( \4433 , \4421 , \4432 );
and \U$2423 ( \4434 , \4409 , \4432 );
or \U$2424 ( \4435 , \4422 , \4433 , \4434 );
and \U$2425 ( \4436 , \3464 , \2848 );
and \U$2426 ( \4437 , \3331 , \2846 );
nor \U$2427 ( \4438 , \4436 , \4437 );
xnor \U$2428 ( \4439 , \4438 , \2853 );
and \U$2429 ( \4440 , \3139 , \2993 );
and \U$2430 ( \4441 , \3168 , \2990 );
nor \U$2431 ( \4442 , \4440 , \4441 );
xnor \U$2432 ( \4443 , \4442 , \2987 );
and \U$2433 ( \4444 , \3194 , \3029 );
and \U$2434 ( \4445 , \3215 , \3027 );
nor \U$2435 ( \4446 , \4444 , \4445 );
xnor \U$2436 ( \4447 , \4446 , \3055 );
xor \U$2437 ( \4448 , \4443 , \4447 );
and \U$2438 ( \4449 , \3239 , \3089 );
and \U$2439 ( \4450 , \3260 , \3087 );
nor \U$2440 ( \4451 , \4449 , \4450 );
xnor \U$2441 ( \4452 , \4451 , \3115 );
xor \U$2442 ( \4453 , \4448 , \4452 );
xor \U$2443 ( \4454 , \4439 , \4453 );
xor \U$2444 ( \4455 , \4435 , \4454 );
and \U$2445 ( \4456 , \2853 , \4426 );
and \U$2446 ( \4457 , \4426 , \4431 );
and \U$2447 ( \4458 , \2853 , \4431 );
or \U$2448 ( \4459 , \4456 , \4457 , \4458 );
and \U$2449 ( \4460 , \4413 , \4417 );
and \U$2450 ( \4461 , \4417 , \4420 );
and \U$2451 ( \4462 , \4413 , \4420 );
or \U$2452 ( \4463 , \4460 , \4461 , \4462 );
xor \U$2453 ( \4464 , \4459 , \4463 );
and \U$2454 ( \4465 , \3287 , \3147 );
and \U$2455 ( \4466 , \3308 , \3145 );
nor \U$2456 ( \4467 , \4465 , \4466 );
xnor \U$2457 ( \4468 , \4467 , \3173 );
xor \U$2458 ( \4469 , \4464 , \4468 );
xor \U$2459 ( \4470 , \4455 , \4469 );
and \U$2460 ( \4471 , \3260 , \2993 );
and \U$2461 ( \4472 , \3194 , \2990 );
nor \U$2462 ( \4473 , \4471 , \4472 );
xnor \U$2463 ( \4474 , \4473 , \2987 );
and \U$2464 ( \4475 , \3173 , \4474 );
and \U$2465 ( \4476 , \3308 , \3029 );
and \U$2466 ( \4477 , \3239 , \3027 );
nor \U$2467 ( \4478 , \4476 , \4477 );
xnor \U$2468 ( \4479 , \4478 , \3055 );
and \U$2469 ( \4480 , \4474 , \4479 );
and \U$2470 ( \4481 , \3173 , \4479 );
or \U$2471 ( \4482 , \4475 , \4480 , \4481 );
and \U$2472 ( \4483 , \3331 , \3089 );
and \U$2473 ( \4484 , \3287 , \3087 );
nor \U$2474 ( \4485 , \4483 , \4484 );
xnor \U$2475 ( \4486 , \4485 , \3115 );
nand \U$2476 ( \4487 , \3464 , \3145 );
xnor \U$2477 ( \4488 , \4487 , \3173 );
and \U$2478 ( \4489 , \4486 , \4488 );
and \U$2479 ( \4490 , \4482 , \4489 );
and \U$2480 ( \4491 , \3464 , \3147 );
and \U$2481 ( \4492 , \3331 , \3145 );
nor \U$2482 ( \4493 , \4491 , \4492 );
xnor \U$2483 ( \4494 , \4493 , \3173 );
and \U$2484 ( \4495 , \4489 , \4494 );
and \U$2485 ( \4496 , \4482 , \4494 );
or \U$2486 ( \4497 , \4490 , \4495 , \4496 );
xor \U$2487 ( \4498 , \4409 , \4421 );
xor \U$2488 ( \4499 , \4498 , \4432 );
and \U$2489 ( \4500 , \4497 , \4499 );
nor \U$2490 ( \4501 , \4470 , \4500 );
and \U$2491 ( \4502 , \4443 , \4447 );
and \U$2492 ( \4503 , \4447 , \4452 );
and \U$2493 ( \4504 , \4443 , \4452 );
or \U$2494 ( \4505 , \4502 , \4503 , \4504 );
nand \U$2495 ( \4506 , \3464 , \2781 );
xnor \U$2496 ( \4507 , \4506 , \2550 );
xor \U$2497 ( \4508 , \4505 , \4507 );
and \U$2498 ( \4509 , \3260 , \3089 );
and \U$2499 ( \4510 , \3194 , \3087 );
nor \U$2500 ( \4511 , \4509 , \4510 );
xnor \U$2501 ( \4512 , \4511 , \3115 );
and \U$2502 ( \4513 , \3308 , \3147 );
and \U$2503 ( \4514 , \3239 , \3145 );
nor \U$2504 ( \4515 , \4513 , \4514 );
xnor \U$2505 ( \4516 , \4515 , \3173 );
xor \U$2506 ( \4517 , \4512 , \4516 );
and \U$2507 ( \4518 , \3331 , \2848 );
and \U$2508 ( \4519 , \3287 , \2846 );
nor \U$2509 ( \4520 , \4518 , \4519 );
xnor \U$2510 ( \4521 , \4520 , \2853 );
xor \U$2511 ( \4522 , \4517 , \4521 );
xor \U$2512 ( \4523 , \4508 , \4522 );
and \U$2513 ( \4524 , \4459 , \4463 );
and \U$2514 ( \4525 , \4463 , \4468 );
and \U$2515 ( \4526 , \4459 , \4468 );
or \U$2516 ( \4527 , \4524 , \4525 , \4526 );
and \U$2517 ( \4528 , \4439 , \4453 );
xor \U$2518 ( \4529 , \4527 , \4528 );
and \U$2519 ( \4530 , \3168 , \2993 );
and \U$2520 ( \4531 , \3077 , \2990 );
nor \U$2521 ( \4532 , \4530 , \4531 );
xnor \U$2522 ( \4533 , \4532 , \2987 );
xor \U$2523 ( \4534 , \2550 , \4533 );
and \U$2524 ( \4535 , \3215 , \3029 );
and \U$2525 ( \4536 , \3139 , \3027 );
nor \U$2526 ( \4537 , \4535 , \4536 );
xnor \U$2527 ( \4538 , \4537 , \3055 );
xor \U$2528 ( \4539 , \4534 , \4538 );
xor \U$2529 ( \4540 , \4529 , \4539 );
xor \U$2530 ( \4541 , \4523 , \4540 );
and \U$2531 ( \4542 , \4435 , \4454 );
and \U$2532 ( \4543 , \4454 , \4469 );
and \U$2533 ( \4544 , \4435 , \4469 );
or \U$2534 ( \4545 , \4542 , \4543 , \4544 );
nor \U$2535 ( \4546 , \4541 , \4545 );
nor \U$2536 ( \4547 , \4501 , \4546 );
and \U$2537 ( \4548 , \4527 , \4528 );
and \U$2538 ( \4549 , \4528 , \4539 );
and \U$2539 ( \4550 , \4527 , \4539 );
or \U$2540 ( \4551 , \4548 , \4549 , \4550 );
and \U$2541 ( \4552 , \4505 , \4507 );
and \U$2542 ( \4553 , \4507 , \4522 );
and \U$2543 ( \4554 , \4505 , \4522 );
or \U$2544 ( \4555 , \4552 , \4553 , \4554 );
and \U$2545 ( \4556 , \3077 , \2993 );
and \U$2546 ( \4557 , \3110 , \2990 );
nor \U$2547 ( \4558 , \4556 , \4557 );
xnor \U$2548 ( \4559 , \4558 , \2987 );
and \U$2549 ( \4560 , \3139 , \3029 );
and \U$2550 ( \4561 , \3168 , \3027 );
nor \U$2551 ( \4562 , \4560 , \4561 );
xnor \U$2552 ( \4563 , \4562 , \3055 );
xor \U$2553 ( \4564 , \4559 , \4563 );
and \U$2554 ( \4565 , \3194 , \3089 );
and \U$2555 ( \4566 , \3215 , \3087 );
nor \U$2556 ( \4567 , \4565 , \4566 );
xnor \U$2557 ( \4568 , \4567 , \3115 );
xor \U$2558 ( \4569 , \4564 , \4568 );
xor \U$2559 ( \4570 , \4555 , \4569 );
and \U$2560 ( \4571 , \2550 , \4533 );
and \U$2561 ( \4572 , \4533 , \4538 );
and \U$2562 ( \4573 , \2550 , \4538 );
or \U$2563 ( \4574 , \4571 , \4572 , \4573 );
and \U$2564 ( \4575 , \4512 , \4516 );
and \U$2565 ( \4576 , \4516 , \4521 );
and \U$2566 ( \4577 , \4512 , \4521 );
or \U$2567 ( \4578 , \4575 , \4576 , \4577 );
xor \U$2568 ( \4579 , \4574 , \4578 );
and \U$2569 ( \4580 , \3239 , \3147 );
and \U$2570 ( \4581 , \3260 , \3145 );
nor \U$2571 ( \4582 , \4580 , \4581 );
xnor \U$2572 ( \4583 , \4582 , \3173 );
and \U$2573 ( \4584 , \3287 , \2848 );
and \U$2574 ( \4585 , \3308 , \2846 );
nor \U$2575 ( \4586 , \4584 , \4585 );
xnor \U$2576 ( \4587 , \4586 , \2853 );
xor \U$2577 ( \4588 , \4583 , \4587 );
and \U$2578 ( \4589 , \3464 , \2783 );
and \U$2579 ( \4590 , \3331 , \2781 );
nor \U$2580 ( \4591 , \4589 , \4590 );
xnor \U$2581 ( \4592 , \4591 , \2550 );
xor \U$2582 ( \4593 , \4588 , \4592 );
xor \U$2583 ( \4594 , \4579 , \4593 );
xor \U$2584 ( \4595 , \4570 , \4594 );
xor \U$2585 ( \4596 , \4551 , \4595 );
and \U$2586 ( \4597 , \4523 , \4540 );
nor \U$2587 ( \4598 , \4596 , \4597 );
and \U$2588 ( \4599 , \4555 , \4569 );
and \U$2589 ( \4600 , \4569 , \4594 );
and \U$2590 ( \4601 , \4555 , \4594 );
or \U$2591 ( \4602 , \4599 , \4600 , \4601 );
and \U$2592 ( \4603 , \4574 , \4578 );
and \U$2593 ( \4604 , \4578 , \4593 );
and \U$2594 ( \4605 , \4574 , \4593 );
or \U$2595 ( \4606 , \4603 , \4604 , \4605 );
nand \U$2596 ( \4607 , \3464 , \2719 );
xnor \U$2597 ( \4608 , \4607 , \2747 );
and \U$2598 ( \4609 , \3215 , \3089 );
and \U$2599 ( \4610 , \3139 , \3087 );
nor \U$2600 ( \4611 , \4609 , \4610 );
xnor \U$2601 ( \4612 , \4611 , \3115 );
and \U$2602 ( \4613 , \3260 , \3147 );
and \U$2603 ( \4614 , \3194 , \3145 );
nor \U$2604 ( \4615 , \4613 , \4614 );
xnor \U$2605 ( \4616 , \4615 , \3173 );
xor \U$2606 ( \4617 , \4612 , \4616 );
and \U$2607 ( \4618 , \3308 , \2848 );
and \U$2608 ( \4619 , \3239 , \2846 );
nor \U$2609 ( \4620 , \4618 , \4619 );
xnor \U$2610 ( \4621 , \4620 , \2853 );
xor \U$2611 ( \4622 , \4617 , \4621 );
xor \U$2612 ( \4623 , \4608 , \4622 );
and \U$2613 ( \4624 , \3110 , \2993 );
and \U$2614 ( \4625 , \3017 , \2990 );
nor \U$2615 ( \4626 , \4624 , \4625 );
xnor \U$2616 ( \4627 , \4626 , \2987 );
xor \U$2617 ( \4628 , \2747 , \4627 );
and \U$2618 ( \4629 , \3168 , \3029 );
and \U$2619 ( \4630 , \3077 , \3027 );
nor \U$2620 ( \4631 , \4629 , \4630 );
xnor \U$2621 ( \4632 , \4631 , \3055 );
xor \U$2622 ( \4633 , \4628 , \4632 );
xor \U$2623 ( \4634 , \4623 , \4633 );
xor \U$2624 ( \4635 , \4606 , \4634 );
and \U$2625 ( \4636 , \4559 , \4563 );
and \U$2626 ( \4637 , \4563 , \4568 );
and \U$2627 ( \4638 , \4559 , \4568 );
or \U$2628 ( \4639 , \4636 , \4637 , \4638 );
and \U$2629 ( \4640 , \4583 , \4587 );
and \U$2630 ( \4641 , \4587 , \4592 );
and \U$2631 ( \4642 , \4583 , \4592 );
or \U$2632 ( \4643 , \4640 , \4641 , \4642 );
xor \U$2633 ( \4644 , \4639 , \4643 );
and \U$2634 ( \4645 , \3331 , \2783 );
and \U$2635 ( \4646 , \3287 , \2781 );
nor \U$2636 ( \4647 , \4645 , \4646 );
xnor \U$2637 ( \4648 , \4647 , \2550 );
xor \U$2638 ( \4649 , \4644 , \4648 );
xor \U$2639 ( \4650 , \4635 , \4649 );
xor \U$2640 ( \4651 , \4602 , \4650 );
and \U$2641 ( \4652 , \4551 , \4595 );
nor \U$2642 ( \4653 , \4651 , \4652 );
nor \U$2643 ( \4654 , \4598 , \4653 );
nand \U$2644 ( \4655 , \4547 , \4654 );
and \U$2645 ( \4656 , \4606 , \4634 );
and \U$2646 ( \4657 , \4634 , \4649 );
and \U$2647 ( \4658 , \4606 , \4649 );
or \U$2648 ( \4659 , \4656 , \4657 , \4658 );
xor \U$2649 ( \4660 , \3519 , \3523 );
xor \U$2650 ( \4661 , \4660 , \3528 );
and \U$2651 ( \4662 , \2747 , \4627 );
and \U$2652 ( \4663 , \4627 , \4632 );
and \U$2653 ( \4664 , \2747 , \4632 );
or \U$2654 ( \4665 , \4662 , \4663 , \4664 );
and \U$2655 ( \4666 , \4612 , \4616 );
and \U$2656 ( \4667 , \4616 , \4621 );
and \U$2657 ( \4668 , \4612 , \4621 );
or \U$2658 ( \4669 , \4666 , \4667 , \4668 );
xor \U$2659 ( \4670 , \4665 , \4669 );
and \U$2660 ( \4671 , \3464 , \2721 );
and \U$2661 ( \4672 , \3331 , \2719 );
nor \U$2662 ( \4673 , \4671 , \4672 );
xnor \U$2663 ( \4674 , \4673 , \2747 );
xor \U$2664 ( \4675 , \4670 , \4674 );
xor \U$2665 ( \4676 , \4661 , \4675 );
xor \U$2666 ( \4677 , \4659 , \4676 );
and \U$2667 ( \4678 , \4639 , \4643 );
and \U$2668 ( \4679 , \4643 , \4648 );
and \U$2669 ( \4680 , \4639 , \4648 );
or \U$2670 ( \4681 , \4678 , \4679 , \4680 );
and \U$2671 ( \4682 , \4608 , \4622 );
and \U$2672 ( \4683 , \4622 , \4633 );
and \U$2673 ( \4684 , \4608 , \4633 );
or \U$2674 ( \4685 , \4682 , \4683 , \4684 );
xor \U$2675 ( \4686 , \4681 , \4685 );
xor \U$2676 ( \4687 , \3535 , \3539 );
xor \U$2677 ( \4688 , \4687 , \3544 );
xor \U$2678 ( \4689 , \4686 , \4688 );
xor \U$2679 ( \4690 , \4677 , \4689 );
and \U$2680 ( \4691 , \4602 , \4650 );
nor \U$2681 ( \4692 , \4690 , \4691 );
and \U$2682 ( \4693 , \4681 , \4685 );
and \U$2683 ( \4694 , \4685 , \4688 );
and \U$2684 ( \4695 , \4681 , \4688 );
or \U$2685 ( \4696 , \4693 , \4694 , \4695 );
and \U$2686 ( \4697 , \4661 , \4675 );
xor \U$2687 ( \4698 , \4696 , \4697 );
and \U$2688 ( \4699 , \4665 , \4669 );
and \U$2689 ( \4700 , \4669 , \4674 );
and \U$2690 ( \4701 , \4665 , \4674 );
or \U$2691 ( \4702 , \4699 , \4700 , \4701 );
xor \U$2692 ( \4703 , \3555 , \3557 );
xor \U$2693 ( \4704 , \4702 , \4703 );
xor \U$2694 ( \4705 , \3531 , \3547 );
xor \U$2695 ( \4706 , \4705 , \3550 );
xor \U$2696 ( \4707 , \4704 , \4706 );
xor \U$2697 ( \4708 , \4698 , \4707 );
and \U$2698 ( \4709 , \4659 , \4676 );
and \U$2699 ( \4710 , \4676 , \4689 );
and \U$2700 ( \4711 , \4659 , \4689 );
or \U$2701 ( \4712 , \4709 , \4710 , \4711 );
nor \U$2702 ( \4713 , \4708 , \4712 );
nor \U$2703 ( \4714 , \4692 , \4713 );
and \U$2704 ( \4715 , \4702 , \4703 );
and \U$2705 ( \4716 , \4703 , \4706 );
and \U$2706 ( \4717 , \4702 , \4706 );
or \U$2707 ( \4718 , \4715 , \4716 , \4717 );
xor \U$2708 ( \4719 , \3418 , \3434 );
xor \U$2709 ( \4720 , \4719 , \3469 );
xor \U$2710 ( \4721 , \4718 , \4720 );
xor \U$2711 ( \4722 , \3553 , \3558 );
xor \U$2712 ( \4723 , \4722 , \3561 );
xor \U$2713 ( \4724 , \4721 , \4723 );
and \U$2714 ( \4725 , \4696 , \4697 );
and \U$2715 ( \4726 , \4697 , \4707 );
and \U$2716 ( \4727 , \4696 , \4707 );
or \U$2717 ( \4728 , \4725 , \4726 , \4727 );
nor \U$2718 ( \4729 , \4724 , \4728 );
xor \U$2719 ( \4730 , \3564 , \3565 );
xor \U$2720 ( \4731 , \4730 , \3568 );
and \U$2721 ( \4732 , \4718 , \4720 );
and \U$2722 ( \4733 , \4720 , \4723 );
and \U$2723 ( \4734 , \4718 , \4723 );
or \U$2724 ( \4735 , \4732 , \4733 , \4734 );
nor \U$2725 ( \4736 , \4731 , \4735 );
nor \U$2726 ( \4737 , \4729 , \4736 );
nand \U$2727 ( \4738 , \4714 , \4737 );
nor \U$2728 ( \4739 , \4655 , \4738 );
and \U$2729 ( \4740 , \3308 , \2993 );
and \U$2730 ( \4741 , \3239 , \2990 );
nor \U$2731 ( \4742 , \4740 , \4741 );
xnor \U$2732 ( \4743 , \4742 , \2987 );
and \U$2733 ( \4744 , \3115 , \4743 );
and \U$2734 ( \4745 , \3331 , \3029 );
and \U$2735 ( \4746 , \3287 , \3027 );
nor \U$2736 ( \4747 , \4745 , \4746 );
xnor \U$2737 ( \4748 , \4747 , \3055 );
and \U$2738 ( \4749 , \4743 , \4748 );
and \U$2739 ( \4750 , \3115 , \4748 );
or \U$2740 ( \4751 , \4744 , \4749 , \4750 );
and \U$2741 ( \4752 , \3239 , \2993 );
and \U$2742 ( \4753 , \3260 , \2990 );
nor \U$2743 ( \4754 , \4752 , \4753 );
xnor \U$2744 ( \4755 , \4754 , \2987 );
and \U$2745 ( \4756 , \3287 , \3029 );
and \U$2746 ( \4757 , \3308 , \3027 );
nor \U$2747 ( \4758 , \4756 , \4757 );
xnor \U$2748 ( \4759 , \4758 , \3055 );
xor \U$2749 ( \4760 , \4755 , \4759 );
and \U$2750 ( \4761 , \3464 , \3089 );
and \U$2751 ( \4762 , \3331 , \3087 );
nor \U$2752 ( \4763 , \4761 , \4762 );
xnor \U$2753 ( \4764 , \4763 , \3115 );
xor \U$2754 ( \4765 , \4760 , \4764 );
xor \U$2755 ( \4766 , \4751 , \4765 );
nand \U$2756 ( \4767 , \3464 , \3087 );
xnor \U$2757 ( \4768 , \4767 , \3115 );
xor \U$2758 ( \4769 , \3115 , \4743 );
xor \U$2759 ( \4770 , \4769 , \4748 );
and \U$2760 ( \4771 , \4768 , \4770 );
nor \U$2761 ( \4772 , \4766 , \4771 );
and \U$2762 ( \4773 , \4755 , \4759 );
and \U$2763 ( \4774 , \4759 , \4764 );
and \U$2764 ( \4775 , \4755 , \4764 );
or \U$2765 ( \4776 , \4773 , \4774 , \4775 );
xor \U$2766 ( \4777 , \4486 , \4488 );
xor \U$2767 ( \4778 , \4776 , \4777 );
xor \U$2768 ( \4779 , \3173 , \4474 );
xor \U$2769 ( \4780 , \4779 , \4479 );
xor \U$2770 ( \4781 , \4778 , \4780 );
and \U$2771 ( \4782 , \4751 , \4765 );
nor \U$2772 ( \4783 , \4781 , \4782 );
nor \U$2773 ( \4784 , \4772 , \4783 );
xor \U$2774 ( \4785 , \4397 , \4401 );
xor \U$2775 ( \4786 , \4785 , \4406 );
xor \U$2776 ( \4787 , \4482 , \4489 );
xor \U$2777 ( \4788 , \4787 , \4494 );
xor \U$2778 ( \4789 , \4786 , \4788 );
and \U$2779 ( \4790 , \4776 , \4777 );
and \U$2780 ( \4791 , \4777 , \4780 );
and \U$2781 ( \4792 , \4776 , \4780 );
or \U$2782 ( \4793 , \4790 , \4791 , \4792 );
nor \U$2783 ( \4794 , \4789 , \4793 );
xor \U$2784 ( \4795 , \4497 , \4499 );
and \U$2785 ( \4796 , \4786 , \4788 );
nor \U$2786 ( \4797 , \4795 , \4796 );
nor \U$2787 ( \4798 , \4794 , \4797 );
nand \U$2788 ( \4799 , \4784 , \4798 );
and \U$2789 ( \4800 , \3287 , \2993 );
and \U$2790 ( \4801 , \3308 , \2990 );
nor \U$2791 ( \4802 , \4800 , \4801 );
xnor \U$2792 ( \4803 , \4802 , \2987 );
and \U$2793 ( \4804 , \3464 , \3029 );
and \U$2794 ( \4805 , \3331 , \3027 );
nor \U$2795 ( \4806 , \4804 , \4805 );
xnor \U$2796 ( \4807 , \4806 , \3055 );
xor \U$2797 ( \4808 , \4803 , \4807 );
and \U$2798 ( \4809 , \3331 , \2993 );
and \U$2799 ( \4810 , \3287 , \2990 );
nor \U$2800 ( \4811 , \4809 , \4810 );
xnor \U$2801 ( \4812 , \4811 , \2987 );
and \U$2802 ( \4813 , \4812 , \3055 );
nor \U$2803 ( \4814 , \4808 , \4813 );
xor \U$2804 ( \4815 , \4768 , \4770 );
and \U$2805 ( \4816 , \4803 , \4807 );
nor \U$2806 ( \4817 , \4815 , \4816 );
nor \U$2807 ( \4818 , \4814 , \4817 );
xor \U$2808 ( \4819 , \4812 , \3055 );
nand \U$2809 ( \4820 , \3464 , \3027 );
xnor \U$2810 ( \4821 , \4820 , \3055 );
nor \U$2811 ( \4822 , \4819 , \4821 );
and \U$2812 ( \4823 , \3464 , \2993 );
and \U$2813 ( \4824 , \3331 , \2990 );
nor \U$2814 ( \4825 , \4823 , \4824 );
xnor \U$2815 ( \4826 , \4825 , \2987 );
nand \U$2816 ( \4827 , \3464 , \2990 );
xnor \U$2817 ( \4828 , \4827 , \2987 );
and \U$2818 ( \4829 , \4828 , \2987 );
nand \U$2819 ( \4830 , \4826 , \4829 );
or \U$2820 ( \4831 , \4822 , \4830 );
nand \U$2821 ( \4832 , \4819 , \4821 );
nand \U$2822 ( \4833 , \4831 , \4832 );
and \U$2823 ( \4834 , \4818 , \4833 );
nand \U$2824 ( \4835 , \4808 , \4813 );
or \U$2825 ( \4836 , \4817 , \4835 );
nand \U$2826 ( \4837 , \4815 , \4816 );
nand \U$2827 ( \4838 , \4836 , \4837 );
nor \U$2828 ( \4839 , \4834 , \4838 );
or \U$2829 ( \4840 , \4799 , \4839 );
nand \U$2830 ( \4841 , \4766 , \4771 );
or \U$2831 ( \4842 , \4783 , \4841 );
nand \U$2832 ( \4843 , \4781 , \4782 );
nand \U$2833 ( \4844 , \4842 , \4843 );
and \U$2834 ( \4845 , \4798 , \4844 );
nand \U$2835 ( \4846 , \4789 , \4793 );
or \U$2836 ( \4847 , \4797 , \4846 );
nand \U$2837 ( \4848 , \4795 , \4796 );
nand \U$2838 ( \4849 , \4847 , \4848 );
nor \U$2839 ( \4850 , \4845 , \4849 );
nand \U$2840 ( \4851 , \4840 , \4850 );
and \U$2841 ( \4852 , \4739 , \4851 );
nand \U$2842 ( \4853 , \4470 , \4500 );
or \U$2843 ( \4854 , \4546 , \4853 );
nand \U$2844 ( \4855 , \4541 , \4545 );
nand \U$2845 ( \4856 , \4854 , \4855 );
and \U$2846 ( \4857 , \4654 , \4856 );
nand \U$2847 ( \4858 , \4596 , \4597 );
or \U$2848 ( \4859 , \4653 , \4858 );
nand \U$2849 ( \4860 , \4651 , \4652 );
nand \U$2850 ( \4861 , \4859 , \4860 );
nor \U$2851 ( \4862 , \4857 , \4861 );
or \U$2852 ( \4863 , \4738 , \4862 );
nand \U$2853 ( \4864 , \4690 , \4691 );
or \U$2854 ( \4865 , \4713 , \4864 );
nand \U$2855 ( \4866 , \4708 , \4712 );
nand \U$2856 ( \4867 , \4865 , \4866 );
and \U$2857 ( \4868 , \4737 , \4867 );
nand \U$2858 ( \4869 , \4724 , \4728 );
or \U$2859 ( \4870 , \4736 , \4869 );
nand \U$2860 ( \4871 , \4731 , \4735 );
nand \U$2861 ( \4872 , \4870 , \4871 );
nor \U$2862 ( \4873 , \4868 , \4872 );
nand \U$2863 ( \4874 , \4863 , \4873 );
nor \U$2864 ( \4875 , \4852 , \4874 );
or \U$2865 ( \4876 , \4393 , \4875 );
nand \U$2866 ( \4877 , \3515 , \3571 );
or \U$2867 ( \4878 , \3647 , \4877 );
nand \U$2868 ( \4879 , \3645 , \3646 );
nand \U$2869 ( \4880 , \4878 , \4879 );
and \U$2870 ( \4881 , \3800 , \4880 );
nand \U$2871 ( \4882 , \3722 , \3723 );
or \U$2872 ( \4883 , \3799 , \4882 );
nand \U$2873 ( \4884 , \3794 , \3798 );
nand \U$2874 ( \4885 , \4883 , \4884 );
nor \U$2875 ( \4886 , \4881 , \4885 );
or \U$2876 ( \4887 , \4096 , \4886 );
nand \U$2877 ( \4888 , \3871 , \3875 );
or \U$2878 ( \4889 , \3952 , \4888 );
nand \U$2879 ( \4890 , \3947 , \3951 );
nand \U$2880 ( \4891 , \4889 , \4890 );
and \U$2881 ( \4892 , \4095 , \4891 );
nand \U$2882 ( \4893 , \4020 , \4024 );
or \U$2883 ( \4894 , \4094 , \4893 );
nand \U$2884 ( \4895 , \4089 , \4093 );
nand \U$2885 ( \4896 , \4894 , \4895 );
nor \U$2886 ( \4897 , \4892 , \4896 );
nand \U$2887 ( \4898 , \4887 , \4897 );
and \U$2888 ( \4899 , \4392 , \4898 );
nand \U$2889 ( \4900 , \4153 , \4157 );
or \U$2890 ( \4901 , \4218 , \4900 );
nand \U$2891 ( \4902 , \4213 , \4217 );
nand \U$2892 ( \4903 , \4901 , \4902 );
and \U$2893 ( \4904 , \4314 , \4903 );
nand \U$2894 ( \4905 , \4270 , \4274 );
or \U$2895 ( \4906 , \4313 , \4905 );
nand \U$2896 ( \4907 , \4308 , \4312 );
nand \U$2897 ( \4908 , \4906 , \4907 );
nor \U$2898 ( \4909 , \4904 , \4908 );
or \U$2899 ( \4910 , \4391 , \4909 );
nand \U$2900 ( \4911 , \4340 , \4344 );
or \U$2901 ( \4912 , \4366 , \4911 );
nand \U$2902 ( \4913 , \4361 , \4365 );
nand \U$2903 ( \4914 , \4912 , \4913 );
and \U$2904 ( \4915 , \4390 , \4914 );
nand \U$2905 ( \4916 , \4377 , \4381 );
or \U$2906 ( \4917 , \4389 , \4916 );
nand \U$2907 ( \4918 , \4384 , \4388 );
nand \U$2908 ( \4919 , \4917 , \4918 );
nor \U$2909 ( \4920 , \4915 , \4919 );
nand \U$2910 ( \4921 , \4910 , \4920 );
nor \U$2911 ( \4922 , \4899 , \4921 );
nand \U$2912 ( \4923 , \4876 , \4922 );
not \U$2913 ( \4924 , \4923 );
xor \U$2914 ( \4925 , \2983 , \4924 );
buf g3284_GF_PartitionCandidate( \4926_nG3284 , \4925 );
buf \U$2919 ( \4927 , RI2b5e785ebcf0_2);
buf \U$2920 ( \4928 , RI2b5e785ebc78_3);
buf \U$2921 ( \4929 , RI2b5e785ebc00_4);
buf \U$2922 ( \4930 , RI2b5e785ebb88_5);
buf \U$2923 ( \4931 , RI2b5e785ebb10_6);
buf \U$2924 ( \4932 , RI2b5e785eba98_7);
buf \U$2925 ( \4933 , RI2b5e785eba20_8);
buf \U$2926 ( \4934 , RI2b5e785eb9a8_9);
buf \U$2927 ( \4935 , RI2b5e785eb930_10);
buf \U$2928 ( \4936 , RI2b5e785eb8b8_11);
buf \U$2929 ( \4937 , RI2b5e785eb840_12);
and \U$2930 ( \4938 , \4936 , \4937 );
and \U$2931 ( \4939 , \4935 , \4938 );
and \U$2932 ( \4940 , \4934 , \4939 );
and \U$2933 ( \4941 , \4933 , \4940 );
and \U$2934 ( \4942 , \4932 , \4941 );
and \U$2935 ( \4943 , \4931 , \4942 );
and \U$2936 ( \4944 , \4930 , \4943 );
and \U$2937 ( \4945 , \4929 , \4944 );
and \U$2938 ( \4946 , \4928 , \4945 );
xor \U$2939 ( \4947 , \4927 , \4946 );
buf \U$2940 ( \4948 , \4947 );
buf \U$2941 ( \4949 , \4948 );
buf \U$2942 ( \4950 , RI2b5e785ae9b8_600);
buf \U$2943 ( \4951 , RI2b5e785aeb98_596);
buf \U$2944 ( \4952 , RI2b5e785aec10_595);
buf \U$2945 ( \4953 , RI2b5e785aec88_594);
buf \U$2946 ( \4954 , RI2b5e785aed00_593);
buf \U$2947 ( \4955 , RI2b5e785aed78_592);
buf \U$2948 ( \4956 , RI2b5e785aedf0_591);
buf \U$2949 ( \4957 , RI2b5e785aee68_590);
buf \U$2950 ( \4958 , RI2b5e785aeee0_589);
buf \U$2951 ( \4959 , RI2b5e785aef58_588);
buf \U$2952 ( \4960 , RI2b5e785ae9b8_600);
buf \U$2953 ( \4961 , RI2b5e785aea30_599);
buf \U$2954 ( \4962 , RI2b5e785aeaa8_598);
buf \U$2955 ( \4963 , RI2b5e785aeb20_597);
and \U$2956 ( \4964 , \4960 , \4961 , \4962 , \4963 );
nor \U$2957 ( \4965 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4964 );
buf \U$2958 ( \4966 , \4965 );
buf \U$2959 ( \4967 , \4966 );
xor \U$2960 ( \4968 , \4950 , \4967 );
buf \U$2961 ( \4969 , \4968 );
buf \U$2962 ( \4970 , RI2b5e785aea30_599);
and \U$2963 ( \4971 , \4950 , \4967 );
xor \U$2964 ( \4972 , \4970 , \4971 );
buf \U$2965 ( \4973 , \4972 );
buf \U$2966 ( \4974 , RI2b5e785aeaa8_598);
and \U$2967 ( \4975 , \4970 , \4971 );
xor \U$2968 ( \4976 , \4974 , \4975 );
buf \U$2969 ( \4977 , \4976 );
buf \U$2970 ( \4978 , RI2b5e785aeb20_597);
and \U$2971 ( \4979 , \4974 , \4975 );
xor \U$2972 ( \4980 , \4978 , \4979 );
buf \U$2973 ( \4981 , \4980 );
buf \U$2974 ( \4982 , RI2b5e785aeb98_596);
and \U$2975 ( \4983 , \4978 , \4979 );
xor \U$2976 ( \4984 , \4982 , \4983 );
buf \U$2977 ( \4985 , \4984 );
not \U$2978 ( \4986 , \4985 );
buf \U$2979 ( \4987 , RI2b5e785aec10_595);
and \U$2980 ( \4988 , \4982 , \4983 );
xor \U$2981 ( \4989 , \4987 , \4988 );
buf \U$2982 ( \4990 , \4989 );
buf \U$2983 ( \4991 , RI2b5e785aec88_594);
and \U$2984 ( \4992 , \4987 , \4988 );
xor \U$2985 ( \4993 , \4991 , \4992 );
buf \U$2986 ( \4994 , \4993 );
buf \U$2987 ( \4995 , RI2b5e785aed00_593);
and \U$2988 ( \4996 , \4991 , \4992 );
xor \U$2989 ( \4997 , \4995 , \4996 );
buf \U$2990 ( \4998 , \4997 );
buf \U$2991 ( \4999 , RI2b5e785aed78_592);
and \U$2992 ( \5000 , \4995 , \4996 );
xor \U$2993 ( \5001 , \4999 , \5000 );
buf \U$2994 ( \5002 , \5001 );
buf \U$2995 ( \5003 , RI2b5e785aedf0_591);
and \U$2996 ( \5004 , \4999 , \5000 );
xor \U$2997 ( \5005 , \5003 , \5004 );
buf \U$2998 ( \5006 , \5005 );
buf \U$2999 ( \5007 , RI2b5e785aee68_590);
and \U$3000 ( \5008 , \5003 , \5004 );
xor \U$3001 ( \5009 , \5007 , \5008 );
buf \U$3002 ( \5010 , \5009 );
buf \U$3003 ( \5011 , RI2b5e785aeee0_589);
and \U$3004 ( \5012 , \5007 , \5008 );
xor \U$3005 ( \5013 , \5011 , \5012 );
buf \U$3006 ( \5014 , \5013 );
buf \U$3007 ( \5015 , RI2b5e785aef58_588);
and \U$3008 ( \5016 , \5011 , \5012 );
xor \U$3009 ( \5017 , \5015 , \5016 );
buf \U$3010 ( \5018 , \5017 );
nor \U$3011 ( \5019 , \4969 , \4973 , \4977 , \4981 , \4986 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3012 ( \5020 , RI2b5e785daa40_28, \5019 );
not \U$3013 ( \5021 , \4969 );
not \U$3014 ( \5022 , \4973 );
not \U$3015 ( \5023 , \4977 );
not \U$3016 ( \5024 , \4981 );
nor \U$3017 ( \5025 , \5021 , \5022 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3018 ( \5026 , RI2b5e78549540_41, \5025 );
nor \U$3019 ( \5027 , \4969 , \5022 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3020 ( \5028 , RI2b5e785388a8_54, \5027 );
nor \U$3021 ( \5029 , \5021 , \4973 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3022 ( \5030 , RI2b5e784a6330_67, \5029 );
nor \U$3023 ( \5031 , \4969 , \4973 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3024 ( \5032 , RI2b5e78495698_80, \5031 );
nor \U$3025 ( \5033 , \5021 , \5022 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3026 ( \5034 , RI2b5e78495080_93, \5033 );
nor \U$3027 ( \5035 , \4969 , \5022 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3028 ( \5036 , RI2b5e78403b80_106, \5035 );
nor \U$3029 ( \5037 , \5021 , \4973 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3030 ( \5038 , RI2b5e775b1e60_119, \5037 );
nor \U$3031 ( \5039 , \4969 , \4973 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3032 ( \5040 , RI2b5e7750bdf8_132, \5039 );
nor \U$3033 ( \5041 , \5021 , \5022 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3034 ( \5042 , RI2b5e774ff5d0_145, \5041 );
nor \U$3035 ( \5043 , \4969 , \5022 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3036 ( \5044 , RI2b5e774f65e8_158, \5043 );
nor \U$3037 ( \5045 , \5021 , \4973 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3038 ( \5046 , RI2b5e774eabd0_171, \5045 );
nor \U$3039 ( \5047 , \4969 , \4973 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3040 ( \5048 , RI2b5e774de3a8_184, \5047 );
nor \U$3041 ( \5049 , \5021 , \5022 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3042 ( \5050 , RI2b5e774d53c0_197, \5049 );
nor \U$3043 ( \5051 , \4969 , \5022 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3044 ( \5052 , RI2b5e785f4300_210, \5051 );
nor \U$3045 ( \5053 , \5021 , \4973 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3046 ( \5054 , RI2b5e785f3ce8_223, \5053 );
nor \U$3047 ( \5055 , \4969 , \4973 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$3048 ( \5056 , RI2b5e785eb0c0_236, \5055 );
or \U$3049 ( \5057 , \5020 , \5026 , \5028 , \5030 , \5032 , \5034 , \5036 , \5038 , \5040 , \5042 , \5044 , \5046 , \5048 , \5050 , \5052 , \5054 , \5056 );
buf \U$3050 ( \5058 , \4990 );
buf \U$3051 ( \5059 , \4994 );
buf \U$3052 ( \5060 , \4998 );
buf \U$3053 ( \5061 , \5002 );
buf \U$3054 ( \5062 , \5006 );
buf \U$3055 ( \5063 , \5010 );
buf \U$3056 ( \5064 , \5014 );
buf \U$3057 ( \5065 , \5018 );
buf \U$3058 ( \5066 , \4985 );
buf \U$3059 ( \5067 , \4969 );
buf \U$3060 ( \5068 , \4973 );
buf \U$3061 ( \5069 , \4977 );
buf \U$3062 ( \5070 , \4981 );
or \U$3063 ( \5071 , \5067 , \5068 , \5069 , \5070 );
and \U$3064 ( \5072 , \5066 , \5071 );
or \U$3065 ( \5073 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 , \5072 );
buf \U$3066 ( \5074 , \5073 );
_DC g2232 ( \5075_nG2232 , \5057 , \5074 );
buf \U$3067 ( \5076 , \5075_nG2232 );
not \U$3068 ( \5077 , \5076 );
xor \U$3069 ( \5078 , \4949 , \5077 );
xor \U$3070 ( \5079 , \4928 , \4945 );
buf \U$3071 ( \5080 , \5079 );
buf \U$3072 ( \5081 , \5080 );
and \U$3073 ( \5082 , RI2b5e785da9c8_29, \5019 );
and \U$3074 ( \5083 , RI2b5e785494c8_42, \5025 );
and \U$3075 ( \5084 , RI2b5e78538830_55, \5027 );
and \U$3076 ( \5085 , RI2b5e784a62b8_68, \5029 );
and \U$3077 ( \5086 , RI2b5e78495620_81, \5031 );
and \U$3078 ( \5087 , RI2b5e78495008_94, \5033 );
and \U$3079 ( \5088 , RI2b5e78403b08_107, \5035 );
and \U$3080 ( \5089 , RI2b5e775b1de8_120, \5037 );
and \U$3081 ( \5090 , RI2b5e7750bd80_133, \5039 );
and \U$3082 ( \5091 , RI2b5e774ff558_146, \5041 );
and \U$3083 ( \5092 , RI2b5e774f6570_159, \5043 );
and \U$3084 ( \5093 , RI2b5e774eab58_172, \5045 );
and \U$3085 ( \5094 , RI2b5e774de330_185, \5047 );
and \U$3086 ( \5095 , RI2b5e774d5348_198, \5049 );
and \U$3087 ( \5096 , RI2b5e785f4288_211, \5051 );
and \U$3088 ( \5097 , RI2b5e785f3658_224, \5053 );
and \U$3089 ( \5098 , RI2b5e785eb048_237, \5055 );
or \U$3090 ( \5099 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 );
_DC g220e ( \5100_nG220e , \5099 , \5074 );
buf \U$3091 ( \5101 , \5100_nG220e );
not \U$3092 ( \5102 , \5101 );
and \U$3093 ( \5103 , \5081 , \5102 );
xor \U$3094 ( \5104 , \4929 , \4944 );
buf \U$3095 ( \5105 , \5104 );
buf \U$3096 ( \5106 , \5105 );
and \U$3097 ( \5107 , RI2b5e785da950_30, \5019 );
and \U$3098 ( \5108 , RI2b5e78549450_43, \5025 );
and \U$3099 ( \5109 , RI2b5e785387b8_56, \5027 );
and \U$3100 ( \5110 , RI2b5e784a6240_69, \5029 );
and \U$3101 ( \5111 , RI2b5e784955a8_82, \5031 );
and \U$3102 ( \5112 , RI2b5e78494f90_95, \5033 );
and \U$3103 ( \5113 , RI2b5e78403a90_108, \5035 );
and \U$3104 ( \5114 , RI2b5e775b1d70_121, \5037 );
and \U$3105 ( \5115 , RI2b5e7750bd08_134, \5039 );
and \U$3106 ( \5116 , RI2b5e774ff4e0_147, \5041 );
and \U$3107 ( \5117 , RI2b5e774f64f8_160, \5043 );
and \U$3108 ( \5118 , RI2b5e774eaae0_173, \5045 );
and \U$3109 ( \5119 , RI2b5e774de2b8_186, \5047 );
and \U$3110 ( \5120 , RI2b5e774d52d0_199, \5049 );
and \U$3111 ( \5121 , RI2b5e785f4210_212, \5051 );
and \U$3112 ( \5122 , RI2b5e785eb5e8_225, \5053 );
and \U$3113 ( \5123 , RI2b5e785e6c50_238, \5055 );
or \U$3114 ( \5124 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 );
_DC g207b ( \5125_nG207b , \5124 , \5074 );
buf \U$3115 ( \5126 , \5125_nG207b );
not \U$3116 ( \5127 , \5126 );
and \U$3117 ( \5128 , \5106 , \5127 );
xor \U$3118 ( \5129 , \4930 , \4943 );
buf \U$3119 ( \5130 , \5129 );
buf \U$3120 ( \5131 , \5130 );
and \U$3121 ( \5132 , RI2b5e785da8d8_31, \5019 );
and \U$3122 ( \5133 , RI2b5e785493d8_44, \5025 );
and \U$3123 ( \5134 , RI2b5e78538740_57, \5027 );
and \U$3124 ( \5135 , RI2b5e784a61c8_70, \5029 );
and \U$3125 ( \5136 , RI2b5e78495530_83, \5031 );
and \U$3126 ( \5137 , RI2b5e78494f18_96, \5033 );
and \U$3127 ( \5138 , RI2b5e78403a18_109, \5035 );
and \U$3128 ( \5139 , RI2b5e775b1cf8_122, \5037 );
and \U$3129 ( \5140 , RI2b5e7750bc90_135, \5039 );
and \U$3130 ( \5141 , RI2b5e774ff468_148, \5041 );
and \U$3131 ( \5142 , RI2b5e774f6480_161, \5043 );
and \U$3132 ( \5143 , RI2b5e774eaa68_174, \5045 );
and \U$3133 ( \5144 , RI2b5e774de240_187, \5047 );
and \U$3134 ( \5145 , RI2b5e774d5258_200, \5049 );
and \U$3135 ( \5146 , RI2b5e785f4198_213, \5051 );
and \U$3136 ( \5147 , RI2b5e785eb570_226, \5053 );
and \U$3137 ( \5148 , RI2b5e785e6bd8_239, \5055 );
or \U$3138 ( \5149 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 );
_DC g2057 ( \5150_nG2057 , \5149 , \5074 );
buf \U$3139 ( \5151 , \5150_nG2057 );
not \U$3140 ( \5152 , \5151 );
and \U$3141 ( \5153 , \5131 , \5152 );
xor \U$3142 ( \5154 , \4931 , \4942 );
buf \U$3143 ( \5155 , \5154 );
buf \U$3144 ( \5156 , \5155 );
and \U$3145 ( \5157 , RI2b5e785da860_32, \5019 );
and \U$3146 ( \5158 , RI2b5e78549360_45, \5025 );
and \U$3147 ( \5159 , RI2b5e785386c8_58, \5027 );
and \U$3148 ( \5160 , RI2b5e784a6150_71, \5029 );
and \U$3149 ( \5161 , RI2b5e784954b8_84, \5031 );
and \U$3150 ( \5162 , RI2b5e78494ea0_97, \5033 );
and \U$3151 ( \5163 , RI2b5e784039a0_110, \5035 );
and \U$3152 ( \5164 , RI2b5e775b1c80_123, \5037 );
and \U$3153 ( \5165 , RI2b5e7750bc18_136, \5039 );
and \U$3154 ( \5166 , RI2b5e774ff3f0_149, \5041 );
and \U$3155 ( \5167 , RI2b5e774f6408_162, \5043 );
and \U$3156 ( \5168 , RI2b5e774ea9f0_175, \5045 );
and \U$3157 ( \5169 , RI2b5e774de1c8_188, \5047 );
and \U$3158 ( \5170 , RI2b5e774d51e0_201, \5049 );
and \U$3159 ( \5171 , RI2b5e785f4120_214, \5051 );
and \U$3160 ( \5172 , RI2b5e785eb4f8_227, \5053 );
and \U$3161 ( \5173 , RI2b5e785e64d0_240, \5055 );
or \U$3162 ( \5174 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 );
_DC g1ed8 ( \5175_nG1ed8 , \5174 , \5074 );
buf \U$3163 ( \5176 , \5175_nG1ed8 );
not \U$3164 ( \5177 , \5176 );
and \U$3165 ( \5178 , \5156 , \5177 );
xor \U$3166 ( \5179 , \4932 , \4941 );
buf \U$3167 ( \5180 , \5179 );
buf \U$3168 ( \5181 , \5180 );
and \U$3169 ( \5182 , RI2b5e78549900_33, \5019 );
and \U$3170 ( \5183 , RI2b5e78538c68_46, \5025 );
and \U$3171 ( \5184 , RI2b5e78538650_59, \5027 );
and \U$3172 ( \5185 , RI2b5e784a60d8_72, \5029 );
and \U$3173 ( \5186 , RI2b5e78495440_85, \5031 );
and \U$3174 ( \5187 , RI2b5e78494e28_98, \5033 );
and \U$3175 ( \5188 , RI2b5e78403928_111, \5035 );
and \U$3176 ( \5189 , RI2b5e775b1c08_124, \5037 );
and \U$3177 ( \5190 , RI2b5e7750bba0_137, \5039 );
and \U$3178 ( \5191 , RI2b5e774ff378_150, \5041 );
and \U$3179 ( \5192 , RI2b5e774f6390_163, \5043 );
and \U$3180 ( \5193 , RI2b5e774ea978_176, \5045 );
and \U$3181 ( \5194 , RI2b5e774de150_189, \5047 );
and \U$3182 ( \5195 , RI2b5e774d5168_202, \5049 );
and \U$3183 ( \5196 , RI2b5e785f40a8_215, \5051 );
and \U$3184 ( \5197 , RI2b5e785eb480_228, \5053 );
and \U$3185 ( \5198 , RI2b5e785da608_241, \5055 );
or \U$3186 ( \5199 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 );
_DC g1eb4 ( \5200_nG1eb4 , \5199 , \5074 );
buf \U$3187 ( \5201 , \5200_nG1eb4 );
not \U$3188 ( \5202 , \5201 );
and \U$3189 ( \5203 , \5181 , \5202 );
xor \U$3190 ( \5204 , \4933 , \4940 );
buf \U$3191 ( \5205 , \5204 );
buf \U$3192 ( \5206 , \5205 );
and \U$3193 ( \5207 , RI2b5e78549888_34, \5019 );
and \U$3194 ( \5208 , RI2b5e78538bf0_47, \5025 );
and \U$3195 ( \5209 , RI2b5e785385d8_60, \5027 );
and \U$3196 ( \5210 , RI2b5e784a6060_73, \5029 );
and \U$3197 ( \5211 , RI2b5e784953c8_86, \5031 );
and \U$3198 ( \5212 , RI2b5e78403ec8_99, \5033 );
and \U$3199 ( \5213 , RI2b5e775b21a8_112, \5035 );
and \U$3200 ( \5214 , RI2b5e775b1b90_125, \5037 );
and \U$3201 ( \5215 , RI2b5e7750bb28_138, \5039 );
and \U$3202 ( \5216 , RI2b5e774ff300_151, \5041 );
and \U$3203 ( \5217 , RI2b5e774f6318_164, \5043 );
and \U$3204 ( \5218 , RI2b5e774ea900_177, \5045 );
and \U$3205 ( \5219 , RI2b5e774de0d8_190, \5047 );
and \U$3206 ( \5220 , RI2b5e774d50f0_203, \5049 );
and \U$3207 ( \5221 , RI2b5e785f4030_216, \5051 );
and \U$3208 ( \5222 , RI2b5e785eb408_229, \5053 );
and \U$3209 ( \5223 , RI2b5e785da590_242, \5055 );
or \U$3210 ( \5224 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 );
_DC g1d69 ( \5225_nG1d69 , \5224 , \5074 );
buf \U$3211 ( \5226 , \5225_nG1d69 );
not \U$3212 ( \5227 , \5226 );
and \U$3213 ( \5228 , \5206 , \5227 );
xor \U$3214 ( \5229 , \4934 , \4939 );
buf \U$3215 ( \5230 , \5229 );
buf \U$3216 ( \5231 , \5230 );
and \U$3217 ( \5232 , RI2b5e78549810_35, \5019 );
and \U$3218 ( \5233 , RI2b5e78538b78_48, \5025 );
and \U$3219 ( \5234 , RI2b5e78538560_61, \5027 );
and \U$3220 ( \5235 , RI2b5e784a5fe8_74, \5029 );
and \U$3221 ( \5236 , RI2b5e78495350_87, \5031 );
and \U$3222 ( \5237 , RI2b5e78403e50_100, \5033 );
and \U$3223 ( \5238 , RI2b5e775b2130_113, \5035 );
and \U$3224 ( \5239 , RI2b5e775b1b18_126, \5037 );
and \U$3225 ( \5240 , RI2b5e7750bab0_139, \5039 );
and \U$3226 ( \5241 , RI2b5e774ff288_152, \5041 );
and \U$3227 ( \5242 , RI2b5e774f62a0_165, \5043 );
and \U$3228 ( \5243 , RI2b5e774ea888_178, \5045 );
and \U$3229 ( \5244 , RI2b5e774de060_191, \5047 );
and \U$3230 ( \5245 , RI2b5e774d5078_204, \5049 );
and \U$3231 ( \5246 , RI2b5e785f3fb8_217, \5051 );
and \U$3232 ( \5247 , RI2b5e785eb390_230, \5053 );
and \U$3233 ( \5248 , RI2b5e785da518_243, \5055 );
or \U$3234 ( \5249 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 );
_DC g1d45 ( \5250_nG1d45 , \5249 , \5074 );
buf \U$3235 ( \5251 , \5250_nG1d45 );
not \U$3236 ( \5252 , \5251 );
and \U$3237 ( \5253 , \5231 , \5252 );
xor \U$3238 ( \5254 , \4935 , \4938 );
buf \U$3239 ( \5255 , \5254 );
buf \U$3240 ( \5256 , \5255 );
and \U$3241 ( \5257 , RI2b5e78549798_36, \5019 );
and \U$3242 ( \5258 , RI2b5e78538b00_49, \5025 );
and \U$3243 ( \5259 , RI2b5e785384e8_62, \5027 );
and \U$3244 ( \5260 , RI2b5e784a5f70_75, \5029 );
and \U$3245 ( \5261 , RI2b5e784952d8_88, \5031 );
and \U$3246 ( \5262 , RI2b5e78403dd8_101, \5033 );
and \U$3247 ( \5263 , RI2b5e775b20b8_114, \5035 );
and \U$3248 ( \5264 , RI2b5e775b1aa0_127, \5037 );
and \U$3249 ( \5265 , RI2b5e7750ba38_140, \5039 );
and \U$3250 ( \5266 , RI2b5e774ff210_153, \5041 );
and \U$3251 ( \5267 , RI2b5e774f6228_166, \5043 );
and \U$3252 ( \5268 , RI2b5e774ea810_179, \5045 );
and \U$3253 ( \5269 , RI2b5e774ddfe8_192, \5047 );
and \U$3254 ( \5270 , RI2b5e774d5000_205, \5049 );
and \U$3255 ( \5271 , RI2b5e785f3f40_218, \5051 );
and \U$3256 ( \5272 , RI2b5e785eb318_231, \5053 );
and \U$3257 ( \5273 , RI2b5e785da4a0_244, \5055 );
or \U$3258 ( \5274 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 );
_DC g1c2a ( \5275_nG1c2a , \5274 , \5074 );
buf \U$3259 ( \5276 , \5275_nG1c2a );
not \U$3260 ( \5277 , \5276 );
and \U$3261 ( \5278 , \5256 , \5277 );
xor \U$3262 ( \5279 , \4936 , \4937 );
buf \U$3263 ( \5280 , \5279 );
buf \U$3264 ( \5281 , \5280 );
and \U$3265 ( \5282 , RI2b5e78549720_37, \5019 );
and \U$3266 ( \5283 , RI2b5e78538a88_50, \5025 );
and \U$3267 ( \5284 , RI2b5e78538470_63, \5027 );
and \U$3268 ( \5285 , RI2b5e784a5ef8_76, \5029 );
and \U$3269 ( \5286 , RI2b5e78495260_89, \5031 );
and \U$3270 ( \5287 , RI2b5e78403d60_102, \5033 );
and \U$3271 ( \5288 , RI2b5e775b2040_115, \5035 );
and \U$3272 ( \5289 , RI2b5e775b1a28_128, \5037 );
and \U$3273 ( \5290 , RI2b5e7750b9c0_141, \5039 );
and \U$3274 ( \5291 , RI2b5e774ff198_154, \5041 );
and \U$3275 ( \5292 , RI2b5e774f61b0_167, \5043 );
and \U$3276 ( \5293 , RI2b5e774ea798_180, \5045 );
and \U$3277 ( \5294 , RI2b5e774ddf70_193, \5047 );
and \U$3278 ( \5295 , RI2b5e774d4f88_206, \5049 );
and \U$3279 ( \5296 , RI2b5e785f3ec8_219, \5051 );
and \U$3280 ( \5297 , RI2b5e785eb2a0_232, \5053 );
and \U$3281 ( \5298 , RI2b5e785da428_245, \5055 );
or \U$3282 ( \5299 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 );
_DC g1c43 ( \5300_nG1c43 , \5299 , \5074 );
buf \U$3283 ( \5301 , \5300_nG1c43 );
not \U$3284 ( \5302 , \5301 );
and \U$3285 ( \5303 , \5281 , \5302 );
not \U$3286 ( \5304 , \4937 );
buf \U$3287 ( \5305 , \5304 );
buf \U$3288 ( \5306 , \5305 );
and \U$3289 ( \5307 , RI2b5e785496a8_38, \5019 );
and \U$3290 ( \5308 , RI2b5e78538a10_51, \5025 );
and \U$3291 ( \5309 , RI2b5e785383f8_64, \5027 );
and \U$3292 ( \5310 , RI2b5e784a5e80_77, \5029 );
and \U$3293 ( \5311 , RI2b5e784951e8_90, \5031 );
and \U$3294 ( \5312 , RI2b5e78403ce8_103, \5033 );
and \U$3295 ( \5313 , RI2b5e775b1fc8_116, \5035 );
and \U$3296 ( \5314 , RI2b5e775b19b0_129, \5037 );
and \U$3297 ( \5315 , RI2b5e7750b948_142, \5039 );
and \U$3298 ( \5316 , RI2b5e774ff120_155, \5041 );
and \U$3299 ( \5317 , RI2b5e774f6138_168, \5043 );
and \U$3300 ( \5318 , RI2b5e774ea720_181, \5045 );
and \U$3301 ( \5319 , RI2b5e774ddef8_194, \5047 );
and \U$3302 ( \5320 , RI2b5e774d4f10_207, \5049 );
and \U$3303 ( \5321 , RI2b5e785f3e50_220, \5051 );
and \U$3304 ( \5322 , RI2b5e785eb228_233, \5053 );
and \U$3305 ( \5323 , RI2b5e785da3b0_246, \5055 );
or \U$3306 ( \5324 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 );
_DC g1b40 ( \5325_nG1b40 , \5324 , \5074 );
buf \U$3307 ( \5326 , \5325_nG1b40 );
not \U$3308 ( \5327 , \5326 );
and \U$3309 ( \5328 , \5306 , \5327 );
buf \U$3310 ( \5329 , RI2b5e785db148_13);
buf \U$3313 ( \5330 , \5329 );
and \U$3314 ( \5331 , RI2b5e78549630_39, \5019 );
and \U$3315 ( \5332 , RI2b5e78538998_52, \5025 );
and \U$3316 ( \5333 , RI2b5e78538380_65, \5027 );
and \U$3317 ( \5334 , RI2b5e784a5e08_78, \5029 );
and \U$3318 ( \5335 , RI2b5e78495170_91, \5031 );
and \U$3319 ( \5336 , RI2b5e78403c70_104, \5033 );
and \U$3320 ( \5337 , RI2b5e775b1f50_117, \5035 );
and \U$3321 ( \5338 , RI2b5e775b1938_130, \5037 );
and \U$3322 ( \5339 , RI2b5e7750b8d0_143, \5039 );
and \U$3323 ( \5340 , RI2b5e774ff0a8_156, \5041 );
and \U$3324 ( \5341 , RI2b5e774f60c0_169, \5043 );
and \U$3325 ( \5342 , RI2b5e774ea6a8_182, \5045 );
and \U$3326 ( \5343 , RI2b5e774dde80_195, \5047 );
and \U$3327 ( \5344 , RI2b5e774d4e98_208, \5049 );
and \U$3328 ( \5345 , RI2b5e785f3dd8_221, \5051 );
and \U$3329 ( \5346 , RI2b5e785eb1b0_234, \5053 );
and \U$3330 ( \5347 , RI2b5e785da338_247, \5055 );
or \U$3331 ( \5348 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 );
_DC g1b24 ( \5349_nG1b24 , \5348 , \5074 );
buf \U$3332 ( \5350 , \5349_nG1b24 );
not \U$3333 ( \5351 , \5350 );
or \U$3334 ( \5352 , \5330 , \5351 );
and \U$3335 ( \5353 , \5327 , \5352 );
and \U$3336 ( \5354 , \5306 , \5352 );
or \U$3337 ( \5355 , \5328 , \5353 , \5354 );
and \U$3338 ( \5356 , \5302 , \5355 );
and \U$3339 ( \5357 , \5281 , \5355 );
or \U$3340 ( \5358 , \5303 , \5356 , \5357 );
and \U$3341 ( \5359 , \5277 , \5358 );
and \U$3342 ( \5360 , \5256 , \5358 );
or \U$3343 ( \5361 , \5278 , \5359 , \5360 );
and \U$3344 ( \5362 , \5252 , \5361 );
and \U$3345 ( \5363 , \5231 , \5361 );
or \U$3346 ( \5364 , \5253 , \5362 , \5363 );
and \U$3347 ( \5365 , \5227 , \5364 );
and \U$3348 ( \5366 , \5206 , \5364 );
or \U$3349 ( \5367 , \5228 , \5365 , \5366 );
and \U$3350 ( \5368 , \5202 , \5367 );
and \U$3351 ( \5369 , \5181 , \5367 );
or \U$3352 ( \5370 , \5203 , \5368 , \5369 );
and \U$3353 ( \5371 , \5177 , \5370 );
and \U$3354 ( \5372 , \5156 , \5370 );
or \U$3355 ( \5373 , \5178 , \5371 , \5372 );
and \U$3356 ( \5374 , \5152 , \5373 );
and \U$3357 ( \5375 , \5131 , \5373 );
or \U$3358 ( \5376 , \5153 , \5374 , \5375 );
and \U$3359 ( \5377 , \5127 , \5376 );
and \U$3360 ( \5378 , \5106 , \5376 );
or \U$3361 ( \5379 , \5128 , \5377 , \5378 );
and \U$3362 ( \5380 , \5102 , \5379 );
and \U$3363 ( \5381 , \5081 , \5379 );
or \U$3364 ( \5382 , \5103 , \5380 , \5381 );
xor \U$3365 ( \5383 , \5078 , \5382 );
buf g223b_GF_PartitionCandidate( \5384_nG223b , \5383 );
buf \U$3366 ( \5385 , \5384_nG223b );
xor \U$3367 ( \5386 , \5081 , \5102 );
xor \U$3368 ( \5387 , \5386 , \5379 );
buf g2217_GF_PartitionCandidate( \5388_nG2217 , \5387 );
buf \U$3369 ( \5389 , \5388_nG2217 );
xor \U$3370 ( \5390 , \5106 , \5127 );
xor \U$3371 ( \5391 , \5390 , \5376 );
buf g2084_GF_PartitionCandidate( \5392_nG2084 , \5391 );
buf \U$3372 ( \5393 , \5392_nG2084 );
and \U$3373 ( \5394 , \5389 , \5393 );
not \U$3374 ( \5395 , \5394 );
and \U$3375 ( \5396 , \5385 , \5395 );
not \U$3376 ( \5397 , \5396 );
buf \U$3377 ( \5398 , \4969 );
buf \U$3378 ( \5399 , \4990 );
buf \U$3379 ( \5400 , \4994 );
buf \U$3380 ( \5401 , \4998 );
buf \U$3381 ( \5402 , \5002 );
buf \U$3382 ( \5403 , \5006 );
buf \U$3383 ( \5404 , \5010 );
buf \U$3384 ( \5405 , \5014 );
buf \U$3385 ( \5406 , \5018 );
buf \U$3386 ( \5407 , \4985 );
nor \U$3387 ( \5408 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 );
buf \U$3388 ( \5409 , \5408 );
buf \U$3389 ( \5410 , \5409 );
xor \U$3390 ( \5411 , \5398 , \5410 );
buf \U$3391 ( \5412 , \5411 );
buf \U$3392 ( \5413 , \4973 );
and \U$3393 ( \5414 , \5398 , \5410 );
xor \U$3394 ( \5415 , \5413 , \5414 );
buf \U$3395 ( \5416 , \5415 );
buf \U$3396 ( \5417 , \4977 );
and \U$3397 ( \5418 , \5413 , \5414 );
xor \U$3398 ( \5419 , \5417 , \5418 );
buf \U$3399 ( \5420 , \5419 );
buf \U$3400 ( \5421 , \4981 );
and \U$3401 ( \5422 , \5417 , \5418 );
xor \U$3402 ( \5423 , \5421 , \5422 );
buf \U$3403 ( \5424 , \5423 );
buf \U$3404 ( \5425 , \4985 );
and \U$3405 ( \5426 , \5421 , \5422 );
xor \U$3406 ( \5427 , \5425 , \5426 );
buf \U$3407 ( \5428 , \5427 );
not \U$3408 ( \5429 , \5428 );
buf \U$3409 ( \5430 , \4990 );
and \U$3410 ( \5431 , \5425 , \5426 );
xor \U$3411 ( \5432 , \5430 , \5431 );
buf \U$3412 ( \5433 , \5432 );
buf \U$3413 ( \5434 , \4994 );
and \U$3414 ( \5435 , \5430 , \5431 );
xor \U$3415 ( \5436 , \5434 , \5435 );
buf \U$3416 ( \5437 , \5436 );
buf \U$3417 ( \5438 , \4998 );
and \U$3418 ( \5439 , \5434 , \5435 );
xor \U$3419 ( \5440 , \5438 , \5439 );
buf \U$3420 ( \5441 , \5440 );
buf \U$3421 ( \5442 , \5002 );
and \U$3422 ( \5443 , \5438 , \5439 );
xor \U$3423 ( \5444 , \5442 , \5443 );
buf \U$3424 ( \5445 , \5444 );
buf \U$3425 ( \5446 , \5006 );
and \U$3426 ( \5447 , \5442 , \5443 );
xor \U$3427 ( \5448 , \5446 , \5447 );
buf \U$3428 ( \5449 , \5448 );
buf \U$3429 ( \5450 , \5010 );
and \U$3430 ( \5451 , \5446 , \5447 );
xor \U$3431 ( \5452 , \5450 , \5451 );
buf \U$3432 ( \5453 , \5452 );
buf \U$3433 ( \5454 , \5014 );
and \U$3434 ( \5455 , \5450 , \5451 );
xor \U$3435 ( \5456 , \5454 , \5455 );
buf \U$3436 ( \5457 , \5456 );
buf \U$3437 ( \5458 , \5018 );
and \U$3438 ( \5459 , \5454 , \5455 );
xor \U$3439 ( \5460 , \5458 , \5459 );
buf \U$3440 ( \5461 , \5460 );
nor \U$3441 ( \5462 , \5412 , \5416 , \5420 , \5424 , \5429 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3442 ( \5463 , RI2b5e785da248_249, \5462 );
not \U$3443 ( \5464 , \5412 );
not \U$3444 ( \5465 , \5416 );
not \U$3445 ( \5466 , \5420 );
not \U$3446 ( \5467 , \5424 );
nor \U$3447 ( \5468 , \5464 , \5465 , \5466 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3448 ( \5469 , RI2b5e785be750_269, \5468 );
nor \U$3449 ( \5470 , \5412 , \5465 , \5466 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3450 ( \5471 , RI2b5e785bc4a0_289, \5470 );
nor \U$3451 ( \5472 , \5464 , \5416 , \5466 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3452 ( \5473 , RI2b5e785bbb40_309, \5472 );
nor \U$3453 ( \5474 , \5412 , \5416 , \5466 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3454 ( \5475 , RI2b5e785b9c50_329, \5474 );
nor \U$3455 ( \5476 , \5464 , \5465 , \5420 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3456 ( \5477 , RI2b5e785b8120_349, \5476 );
nor \U$3457 ( \5478 , \5412 , \5465 , \5420 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3458 ( \5479 , RI2b5e785b77c0_369, \5478 );
nor \U$3459 ( \5480 , \5464 , \5416 , \5420 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3460 ( \5481 , RI2b5e785b6e60_389, \5480 );
nor \U$3461 ( \5482 , \5412 , \5416 , \5420 , \5467 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3462 ( \5483 , RI2b5e785b56f0_409, \5482 );
nor \U$3463 ( \5484 , \5464 , \5465 , \5466 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3464 ( \5485 , RI2b5e785b4d90_429, \5484 );
nor \U$3465 ( \5486 , \5412 , \5465 , \5466 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3466 ( \5487 , RI2b5e785b39e0_449, \5486 );
nor \U$3467 ( \5488 , \5464 , \5416 , \5466 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3468 ( \5489 , RI2b5e785b3080_469, \5488 );
nor \U$3469 ( \5490 , \5412 , \5416 , \5466 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3470 ( \5491 , RI2b5e785b2720_489, \5490 );
nor \U$3471 ( \5492 , \5464 , \5465 , \5420 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3472 ( \5493 , RI2b5e785b1730_509, \5492 );
nor \U$3473 ( \5494 , \5412 , \5465 , \5420 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3474 ( \5495 , RI2b5e785b0dd0_529, \5494 );
nor \U$3475 ( \5496 , \5464 , \5416 , \5420 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3476 ( \5497 , RI2b5e785b0470_549, \5496 );
nor \U$3477 ( \5498 , \5412 , \5416 , \5420 , \5424 , \5428 , \5433 , \5437 , \5441 , \5445 , \5449 , \5453 , \5457 , \5461 );
and \U$3478 ( \5499 , RI2b5e785af840_569, \5498 );
or \U$3479 ( \5500 , \5463 , \5469 , \5471 , \5473 , \5475 , \5477 , \5479 , \5481 , \5483 , \5485 , \5487 , \5489 , \5491 , \5493 , \5495 , \5497 , \5499 );
buf \U$3480 ( \5501 , \5433 );
buf \U$3481 ( \5502 , \5437 );
buf \U$3482 ( \5503 , \5441 );
buf \U$3483 ( \5504 , \5445 );
buf \U$3484 ( \5505 , \5449 );
buf \U$3485 ( \5506 , \5453 );
buf \U$3486 ( \5507 , \5457 );
buf \U$3487 ( \5508 , \5461 );
buf \U$3488 ( \5509 , \5428 );
buf \U$3489 ( \5510 , \5412 );
buf \U$3490 ( \5511 , \5416 );
buf \U$3491 ( \5512 , \5420 );
buf \U$3492 ( \5513 , \5424 );
or \U$3493 ( \5514 , \5510 , \5511 , \5512 , \5513 );
and \U$3494 ( \5515 , \5509 , \5514 );
or \U$3495 ( \5516 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5515 );
buf \U$3496 ( \5517 , \5516 );
_DC g290c ( \5518_nG290c , \5500 , \5517 );
buf \U$3497 ( \5519 , \5518_nG290c );
buf \U$3498 ( \5520 , RI2b5e785ebd68_1);
and \U$3499 ( \5521 , \4927 , \4946 );
and \U$3500 ( \5522 , \5520 , \5521 );
buf \U$3501 ( \5523 , \5522 );
buf \U$3502 ( \5524 , \5523 );
xor \U$3503 ( \5525 , \5520 , \5521 );
buf \U$3504 ( \5526 , \5525 );
buf \U$3505 ( \5527 , \5526 );
and \U$3506 ( \5528 , RI2b5e785daab8_27, \5019 );
and \U$3507 ( \5529 , RI2b5e785495b8_40, \5025 );
and \U$3508 ( \5530 , RI2b5e78538920_53, \5027 );
and \U$3509 ( \5531 , RI2b5e784a63a8_66, \5029 );
and \U$3510 ( \5532 , RI2b5e78495710_79, \5031 );
and \U$3511 ( \5533 , RI2b5e784950f8_92, \5033 );
and \U$3512 ( \5534 , RI2b5e78403bf8_105, \5035 );
and \U$3513 ( \5535 , RI2b5e775b1ed8_118, \5037 );
and \U$3514 ( \5536 , RI2b5e775b18c0_131, \5039 );
and \U$3515 ( \5537 , RI2b5e7750b858_144, \5041 );
and \U$3516 ( \5538 , RI2b5e774ff030_157, \5043 );
and \U$3517 ( \5539 , RI2b5e774f6048_170, \5045 );
and \U$3518 ( \5540 , RI2b5e774ea630_183, \5047 );
and \U$3519 ( \5541 , RI2b5e774dde08_196, \5049 );
and \U$3520 ( \5542 , RI2b5e774d4e20_209, \5051 );
and \U$3521 ( \5543 , RI2b5e785f3d60_222, \5053 );
and \U$3522 ( \5544 , RI2b5e785eb138_235, \5055 );
or \U$3523 ( \5545 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 );
_DC g23ed ( \5546_nG23ed , \5545 , \5074 );
buf \U$3524 ( \5547 , \5546_nG23ed );
not \U$3525 ( \5548 , \5547 );
and \U$3526 ( \5549 , \5527 , \5548 );
and \U$3527 ( \5550 , \4949 , \5077 );
and \U$3528 ( \5551 , \5077 , \5382 );
and \U$3529 ( \5552 , \4949 , \5382 );
or \U$3530 ( \5553 , \5550 , \5551 , \5552 );
and \U$3531 ( \5554 , \5548 , \5553 );
and \U$3532 ( \5555 , \5527 , \5553 );
or \U$3533 ( \5556 , \5549 , \5554 , \5555 );
xnor \U$3534 ( \5557 , \5524 , \5556 );
buf g2402_GF_PartitionCandidate( \5558_nG2402 , \5557 );
buf \U$3535 ( \5559 , \5558_nG2402 );
xor \U$3536 ( \5560 , \5527 , \5548 );
xor \U$3537 ( \5561 , \5560 , \5553 );
buf g23f6_GF_PartitionCandidate( \5562_nG23f6 , \5561 );
buf \U$3538 ( \5563 , \5562_nG23f6 );
xor \U$3539 ( \5564 , \5559 , \5563 );
xor \U$3540 ( \5565 , \5563 , \5385 );
not \U$3541 ( \5566 , \5565 );
and \U$3542 ( \5567 , \5564 , \5566 );
and \U$3543 ( \5568 , \5519 , \5567 );
and \U$3544 ( \5569 , RI2b5e785da2c0_248, \5462 );
and \U$3545 ( \5570 , RI2b5e785be7c8_268, \5468 );
and \U$3546 ( \5571 , RI2b5e785bc518_288, \5470 );
and \U$3547 ( \5572 , RI2b5e785bbbb8_308, \5472 );
and \U$3548 ( \5573 , RI2b5e785b9cc8_328, \5474 );
and \U$3549 ( \5574 , RI2b5e785b9368_348, \5476 );
and \U$3550 ( \5575 , RI2b5e785b7838_368, \5478 );
and \U$3551 ( \5576 , RI2b5e785b6ed8_388, \5480 );
and \U$3552 ( \5577 , RI2b5e785b5768_408, \5482 );
and \U$3553 ( \5578 , RI2b5e785b4e08_428, \5484 );
and \U$3554 ( \5579 , RI2b5e785b3a58_448, \5486 );
and \U$3555 ( \5580 , RI2b5e785b30f8_468, \5488 );
and \U$3556 ( \5581 , RI2b5e785b2798_488, \5490 );
and \U$3557 ( \5582 , RI2b5e785b17a8_508, \5492 );
and \U$3558 ( \5583 , RI2b5e785b0e48_528, \5494 );
and \U$3559 ( \5584 , RI2b5e785b04e8_548, \5496 );
and \U$3560 ( \5585 , RI2b5e785afb88_568, \5498 );
or \U$3561 ( \5586 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 );
_DC g2a01 ( \5587_nG2a01 , \5586 , \5517 );
buf \U$3562 ( \5588 , \5587_nG2a01 );
and \U$3563 ( \5589 , \5588 , \5565 );
nor \U$3564 ( \5590 , \5568 , \5589 );
and \U$3565 ( \5591 , \5563 , \5385 );
not \U$3566 ( \5592 , \5591 );
and \U$3567 ( \5593 , \5559 , \5592 );
xnor \U$3568 ( \5594 , \5590 , \5593 );
xor \U$3569 ( \5595 , \5397 , \5594 );
and \U$3571 ( \5596 , RI2b5e785da1d0_250, \5462 );
and \U$3572 ( \5597 , RI2b5e785be6d8_270, \5468 );
and \U$3573 ( \5598 , RI2b5e785bc428_290, \5470 );
and \U$3574 ( \5599 , RI2b5e785bbac8_310, \5472 );
and \U$3575 ( \5600 , RI2b5e785b9bd8_330, \5474 );
and \U$3576 ( \5601 , RI2b5e785b80a8_350, \5476 );
and \U$3577 ( \5602 , RI2b5e785b7748_370, \5478 );
and \U$3578 ( \5603 , RI2b5e785b6de8_390, \5480 );
and \U$3579 ( \5604 , RI2b5e785b5678_410, \5482 );
and \U$3580 ( \5605 , RI2b5e785b4d18_430, \5484 );
and \U$3581 ( \5606 , RI2b5e785b3968_450, \5486 );
and \U$3582 ( \5607 , RI2b5e785b3008_470, \5488 );
and \U$3583 ( \5608 , RI2b5e785b26a8_490, \5490 );
and \U$3584 ( \5609 , RI2b5e785b16b8_510, \5492 );
and \U$3585 ( \5610 , RI2b5e785b0d58_530, \5494 );
and \U$3586 ( \5611 , RI2b5e785b03f8_550, \5496 );
and \U$3587 ( \5612 , RI2b5e785af7c8_570, \5498 );
or \U$3588 ( \5613 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 );
_DC g2843 ( \5614_nG2843 , \5613 , \5517 );
buf \U$3589 ( \5615 , \5614_nG2843 );
or \U$3590 ( \5616 , \5524 , \5556 );
not \U$3591 ( \5617 , \5616 );
buf g25dc_GF_PartitionCandidate( \5618_nG25dc , \5617 );
buf \U$3592 ( \5619 , \5618_nG25dc );
xor \U$3593 ( \5620 , \5619 , \5559 );
and \U$3594 ( \5621 , \5615 , \5620 );
nor \U$3595 ( \5622 , 1'b0 , \5621 );
xnor \U$3597 ( \5623 , \5622 , 1'b0 );
xor \U$3598 ( \5624 , \5595 , \5623 );
xor \U$3599 ( \5625 , 1'b0 , \5624 );
xor \U$3601 ( \5626 , \5385 , \5389 );
xor \U$3602 ( \5627 , \5389 , \5393 );
not \U$3603 ( \5628 , \5627 );
and \U$3604 ( \5629 , \5626 , \5628 );
and \U$3605 ( \5630 , \5588 , \5629 );
not \U$3606 ( \5631 , \5630 );
xnor \U$3607 ( \5632 , \5631 , \5396 );
and \U$3608 ( \5633 , \5615 , \5567 );
and \U$3609 ( \5634 , \5519 , \5565 );
nor \U$3610 ( \5635 , \5633 , \5634 );
xnor \U$3611 ( \5636 , \5635 , \5593 );
and \U$3612 ( \5637 , \5632 , \5636 );
or \U$3614 ( \5638 , 1'b0 , \5637 , 1'b0 );
xor \U$3616 ( \5639 , \5638 , 1'b0 );
xor \U$3618 ( \5640 , \5639 , 1'b0 );
and \U$3619 ( \5641 , \5625 , \5640 );
or \U$3620 ( \5642 , 1'b0 , 1'b0 , \5641 );
and \U$3623 ( \5643 , \5588 , \5567 );
not \U$3624 ( \5644 , \5643 );
xnor \U$3625 ( \5645 , \5644 , \5593 );
xor \U$3626 ( \5646 , 1'b0 , \5645 );
and \U$3628 ( \5647 , \5519 , \5620 );
nor \U$3629 ( \5648 , 1'b0 , \5647 );
xnor \U$3630 ( \5649 , \5648 , 1'b0 );
xor \U$3631 ( \5650 , \5646 , \5649 );
xor \U$3632 ( \5651 , 1'b0 , \5650 );
xor \U$3634 ( \5652 , \5651 , 1'b1 );
and \U$3635 ( \5653 , \5397 , \5594 );
and \U$3636 ( \5654 , \5594 , \5623 );
and \U$3637 ( \5655 , \5397 , \5623 );
or \U$3638 ( \5656 , \5653 , \5654 , \5655 );
xor \U$3640 ( \5657 , \5656 , 1'b0 );
xor \U$3642 ( \5658 , \5657 , 1'b0 );
xor \U$3643 ( \5659 , \5652 , \5658 );
and \U$3644 ( \5660 , \5642 , \5659 );
or \U$3646 ( \5661 , 1'b0 , \5660 , 1'b0 );
xor \U$3648 ( \5662 , \5661 , 1'b0 );
and \U$3650 ( \5663 , \5651 , 1'b1 );
and \U$3651 ( \5664 , 1'b1 , \5658 );
and \U$3652 ( \5665 , \5651 , \5658 );
or \U$3653 ( \5666 , \5663 , \5664 , \5665 );
xor \U$3654 ( \5667 , 1'b0 , \5666 );
not \U$3656 ( \5668 , \5593 );
and \U$3658 ( \5669 , \5588 , \5620 );
nor \U$3659 ( \5670 , 1'b0 , \5669 );
xnor \U$3660 ( \5671 , \5670 , 1'b0 );
xor \U$3661 ( \5672 , \5668 , \5671 );
xor \U$3663 ( \5673 , \5672 , 1'b0 );
xor \U$3664 ( \5674 , 1'b0 , \5673 );
xor \U$3666 ( \5675 , \5674 , 1'b0 );
and \U$3668 ( \5676 , \5645 , \5649 );
or \U$3670 ( \5677 , 1'b0 , \5676 , 1'b0 );
xor \U$3672 ( \5678 , \5677 , 1'b0 );
xor \U$3674 ( \5679 , \5678 , 1'b0 );
xor \U$3675 ( \5680 , \5675 , \5679 );
xor \U$3676 ( \5681 , \5667 , \5680 );
xor \U$3677 ( \5682 , \5662 , \5681 );
xor \U$3683 ( \5683 , \5131 , \5152 );
xor \U$3684 ( \5684 , \5683 , \5373 );
buf g2060_GF_PartitionCandidate( \5685_nG2060 , \5684 );
buf \U$3685 ( \5686 , \5685_nG2060 );
xor \U$3686 ( \5687 , \5393 , \5686 );
xor \U$3687 ( \5688 , \5156 , \5177 );
xor \U$3688 ( \5689 , \5688 , \5370 );
buf g1ee1_GF_PartitionCandidate( \5690_nG1ee1 , \5689 );
buf \U$3689 ( \5691 , \5690_nG1ee1 );
xor \U$3690 ( \5692 , \5686 , \5691 );
not \U$3691 ( \5693 , \5692 );
and \U$3692 ( \5694 , \5687 , \5693 );
and \U$3693 ( \5695 , \5588 , \5694 );
not \U$3694 ( \5696 , \5695 );
and \U$3695 ( \5697 , \5686 , \5691 );
not \U$3696 ( \5698 , \5697 );
and \U$3697 ( \5699 , \5393 , \5698 );
xnor \U$3698 ( \5700 , \5696 , \5699 );
and \U$3699 ( \5701 , \5615 , \5629 );
and \U$3700 ( \5702 , \5519 , \5627 );
nor \U$3701 ( \5703 , \5701 , \5702 );
xnor \U$3702 ( \5704 , \5703 , \5396 );
and \U$3703 ( \5705 , \5700 , \5704 );
or \U$3705 ( \5706 , 1'b0 , \5705 , 1'b0 );
and \U$3706 ( \5707 , RI2b5e785da0e0_252, \5462 );
and \U$3707 ( \5708 , RI2b5e785be5e8_272, \5468 );
and \U$3708 ( \5709 , RI2b5e785bc338_292, \5470 );
and \U$3709 ( \5710 , RI2b5e785bb9d8_312, \5472 );
and \U$3710 ( \5711 , RI2b5e785b9ae8_332, \5474 );
and \U$3711 ( \5712 , RI2b5e785b7fb8_352, \5476 );
and \U$3712 ( \5713 , RI2b5e785b7658_372, \5478 );
and \U$3713 ( \5714 , RI2b5e785b5ee8_392, \5480 );
and \U$3714 ( \5715 , RI2b5e785b5588_412, \5482 );
and \U$3715 ( \5716 , RI2b5e785b4c28_432, \5484 );
and \U$3716 ( \5717 , RI2b5e785b3878_452, \5486 );
and \U$3717 ( \5718 , RI2b5e785b2f18_472, \5488 );
and \U$3718 ( \5719 , RI2b5e785b25b8_492, \5490 );
and \U$3719 ( \5720 , RI2b5e785b15c8_512, \5492 );
and \U$3720 ( \5721 , RI2b5e785b0c68_532, \5494 );
and \U$3721 ( \5722 , RI2b5e785b0308_552, \5496 );
and \U$3722 ( \5723 , RI2b5e785af6d8_572, \5498 );
or \U$3723 ( \5724 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 );
_DC g26a4 ( \5725_nG26a4 , \5724 , \5517 );
buf \U$3724 ( \5726 , \5725_nG26a4 );
and \U$3725 ( \5727 , \5726 , \5567 );
and \U$3726 ( \5728 , RI2b5e785da158_251, \5462 );
and \U$3727 ( \5729 , RI2b5e785be660_271, \5468 );
and \U$3728 ( \5730 , RI2b5e785bc3b0_291, \5470 );
and \U$3729 ( \5731 , RI2b5e785bba50_311, \5472 );
and \U$3730 ( \5732 , RI2b5e785b9b60_331, \5474 );
and \U$3731 ( \5733 , RI2b5e785b8030_351, \5476 );
and \U$3732 ( \5734 , RI2b5e785b76d0_371, \5478 );
and \U$3733 ( \5735 , RI2b5e785b6d70_391, \5480 );
and \U$3734 ( \5736 , RI2b5e785b5600_411, \5482 );
and \U$3735 ( \5737 , RI2b5e785b4ca0_431, \5484 );
and \U$3736 ( \5738 , RI2b5e785b38f0_451, \5486 );
and \U$3737 ( \5739 , RI2b5e785b2f90_471, \5488 );
and \U$3738 ( \5740 , RI2b5e785b2630_491, \5490 );
and \U$3739 ( \5741 , RI2b5e785b1640_511, \5492 );
and \U$3740 ( \5742 , RI2b5e785b0ce0_531, \5494 );
and \U$3741 ( \5743 , RI2b5e785b0380_551, \5496 );
and \U$3742 ( \5744 , RI2b5e785af750_571, \5498 );
or \U$3743 ( \5745 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 );
_DC g2782 ( \5746_nG2782 , \5745 , \5517 );
buf \U$3744 ( \5747 , \5746_nG2782 );
and \U$3745 ( \5748 , \5747 , \5565 );
nor \U$3746 ( \5749 , \5727 , \5748 );
xnor \U$3747 ( \5750 , \5749 , \5593 );
and \U$3749 ( \5751 , RI2b5e785da068_253, \5462 );
and \U$3750 ( \5752 , RI2b5e785be570_273, \5468 );
and \U$3751 ( \5753 , RI2b5e785bc2c0_293, \5470 );
and \U$3752 ( \5754 , RI2b5e785bb960_313, \5472 );
and \U$3753 ( \5755 , RI2b5e785b9a70_333, \5474 );
and \U$3754 ( \5756 , RI2b5e785b7f40_353, \5476 );
and \U$3755 ( \5757 , RI2b5e785b75e0_373, \5478 );
and \U$3756 ( \5758 , RI2b5e785b5e70_393, \5480 );
and \U$3757 ( \5759 , RI2b5e785b5510_413, \5482 );
and \U$3758 ( \5760 , RI2b5e785b4bb0_433, \5484 );
and \U$3759 ( \5761 , RI2b5e785b3800_453, \5486 );
and \U$3760 ( \5762 , RI2b5e785b2ea0_473, \5488 );
and \U$3761 ( \5763 , RI2b5e785b2540_493, \5490 );
and \U$3762 ( \5764 , RI2b5e785b1550_513, \5492 );
and \U$3763 ( \5765 , RI2b5e785b0bf0_533, \5494 );
and \U$3764 ( \5766 , RI2b5e785b0290_553, \5496 );
and \U$3765 ( \5767 , RI2b5e785af660_573, \5498 );
or \U$3766 ( \5768 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 );
_DC g25bb ( \5769_nG25bb , \5768 , \5517 );
buf \U$3767 ( \5770 , \5769_nG25bb );
and \U$3768 ( \5771 , \5770 , \5620 );
nor \U$3769 ( \5772 , 1'b0 , \5771 );
xnor \U$3770 ( \5773 , \5772 , 1'b0 );
and \U$3771 ( \5774 , \5750 , \5773 );
or \U$3774 ( \5775 , \5774 , 1'b0 , 1'b0 );
and \U$3775 ( \5776 , \5706 , \5775 );
or \U$3778 ( \5777 , \5776 , 1'b0 , 1'b0 );
and \U$3781 ( \5778 , \5726 , \5620 );
nor \U$3782 ( \5779 , 1'b0 , \5778 );
xnor \U$3783 ( \5780 , \5779 , 1'b0 );
xor \U$3785 ( \5781 , \5780 , 1'b0 );
xor \U$3787 ( \5782 , \5781 , 1'b0 );
not \U$3788 ( \5783 , \5699 );
and \U$3789 ( \5784 , \5519 , \5629 );
and \U$3790 ( \5785 , \5588 , \5627 );
nor \U$3791 ( \5786 , \5784 , \5785 );
xnor \U$3792 ( \5787 , \5786 , \5396 );
xor \U$3793 ( \5788 , \5783 , \5787 );
and \U$3794 ( \5789 , \5747 , \5567 );
and \U$3795 ( \5790 , \5615 , \5565 );
nor \U$3796 ( \5791 , \5789 , \5790 );
xnor \U$3797 ( \5792 , \5791 , \5593 );
xor \U$3798 ( \5793 , \5788 , \5792 );
and \U$3799 ( \5794 , \5782 , \5793 );
or \U$3801 ( \5795 , 1'b0 , \5794 , 1'b0 );
and \U$3802 ( \5796 , \5777 , \5795 );
or \U$3803 ( \5797 , 1'b0 , 1'b0 , \5796 );
and \U$3805 ( \5798 , \5747 , \5620 );
nor \U$3806 ( \5799 , 1'b0 , \5798 );
xnor \U$3807 ( \5800 , \5799 , 1'b0 );
xor \U$3809 ( \5801 , \5800 , 1'b0 );
xor \U$3811 ( \5802 , \5801 , 1'b0 );
xor \U$3813 ( \5803 , 1'b0 , \5632 );
xor \U$3814 ( \5804 , \5803 , \5636 );
xor \U$3815 ( \5805 , \5802 , \5804 );
and \U$3817 ( \5806 , \5805 , 1'b1 );
and \U$3818 ( \5807 , \5783 , \5787 );
and \U$3819 ( \5808 , \5787 , \5792 );
and \U$3820 ( \5809 , \5783 , \5792 );
or \U$3821 ( \5810 , \5807 , \5808 , \5809 );
xor \U$3823 ( \5811 , \5810 , 1'b0 );
xor \U$3825 ( \5812 , \5811 , 1'b0 );
and \U$3826 ( \5813 , 1'b1 , \5812 );
and \U$3827 ( \5814 , \5805 , \5812 );
or \U$3828 ( \5815 , \5806 , \5813 , \5814 );
and \U$3829 ( \5816 , \5797 , \5815 );
xor \U$3831 ( \5817 , \5625 , 1'b0 );
xor \U$3832 ( \5818 , \5817 , \5640 );
and \U$3833 ( \5819 , \5815 , \5818 );
and \U$3834 ( \5820 , \5797 , \5818 );
or \U$3835 ( \5821 , \5816 , \5819 , \5820 );
xor \U$3837 ( \5822 , 1'b0 , \5642 );
xor \U$3838 ( \5823 , \5822 , \5659 );
and \U$3839 ( \5824 , \5821 , \5823 );
or \U$3840 ( \5825 , 1'b0 , 1'b0 , \5824 );
nand \U$3841 ( \5826 , \5682 , \5825 );
nor \U$3842 ( \5827 , \5682 , \5825 );
not \U$3843 ( \5828 , \5827 );
nand \U$3844 ( \5829 , \5826 , \5828 );
xor \U$3845 ( \5830 , \5306 , \5327 );
xor \U$3846 ( \5831 , \5830 , \5352 );
buf g1b47_GF_PartitionCandidate( \5832_nG1b47 , \5831 );
buf \U$3847 ( \5833 , \5832_nG1b47 );
xor \U$3848 ( \5834 , \5330 , \5350 );
buf g1b27_GF_PartitionCandidate( \5835_nG1b27 , \5834 );
buf \U$3849 ( \5836 , \5835_nG1b27 );
xor \U$3850 ( \5837 , \5833 , \5836 );
not \U$3851 ( \5838 , \5836 );
and \U$3852 ( \5839 , \5837 , \5838 );
and \U$3853 ( \5840 , \5770 , \5839 );
and \U$3854 ( \5841 , \5726 , \5836 );
nor \U$3855 ( \5842 , \5840 , \5841 );
xnor \U$3856 ( \5843 , \5842 , \5833 );
and \U$3857 ( \5844 , RI2b5e785c2bc0_255, \5462 );
and \U$3858 ( \5845 , RI2b5e785be480_275, \5468 );
and \U$3859 ( \5846 , RI2b5e785bc1d0_295, \5470 );
and \U$3860 ( \5847 , RI2b5e785ba2e0_315, \5472 );
and \U$3861 ( \5848 , RI2b5e785b9980_335, \5474 );
and \U$3862 ( \5849 , RI2b5e785b7e50_355, \5476 );
and \U$3863 ( \5850 , RI2b5e785b74f0_375, \5478 );
and \U$3864 ( \5851 , RI2b5e785b5d80_395, \5480 );
and \U$3865 ( \5852 , RI2b5e785b5420_415, \5482 );
and \U$3866 ( \5853 , RI2b5e785b4ac0_435, \5484 );
and \U$3867 ( \5854 , RI2b5e785b3710_455, \5486 );
and \U$3868 ( \5855 , RI2b5e785b2db0_475, \5488 );
and \U$3869 ( \5856 , RI2b5e785b2450_495, \5490 );
and \U$3870 ( \5857 , RI2b5e785b1460_515, \5492 );
and \U$3871 ( \5858 , RI2b5e785b0b00_535, \5494 );
and \U$3872 ( \5859 , RI2b5e785b01a0_555, \5496 );
and \U$3873 ( \5860 , RI2b5e785af570_575, \5498 );
or \U$3874 ( \5861 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 );
_DC g242a ( \5862_nG242a , \5861 , \5517 );
buf \U$3875 ( \5863 , \5862_nG242a );
xor \U$3876 ( \5864 , \5256 , \5277 );
xor \U$3877 ( \5865 , \5864 , \5358 );
buf g1c4f_GF_PartitionCandidate( \5866_nG1c4f , \5865 );
buf \U$3878 ( \5867 , \5866_nG1c4f );
xor \U$3879 ( \5868 , \5281 , \5302 );
xor \U$3880 ( \5869 , \5868 , \5355 );
buf g1c53_GF_PartitionCandidate( \5870_nG1c53 , \5869 );
buf \U$3881 ( \5871 , \5870_nG1c53 );
xor \U$3882 ( \5872 , \5867 , \5871 );
xor \U$3883 ( \5873 , \5871 , \5833 );
not \U$3884 ( \5874 , \5873 );
and \U$3885 ( \5875 , \5872 , \5874 );
and \U$3886 ( \5876 , \5863 , \5875 );
and \U$3887 ( \5877 , RI2b5e785c2c38_254, \5462 );
and \U$3888 ( \5878 , RI2b5e785be4f8_274, \5468 );
and \U$3889 ( \5879 , RI2b5e785bc248_294, \5470 );
and \U$3890 ( \5880 , RI2b5e785ba358_314, \5472 );
and \U$3891 ( \5881 , RI2b5e785b99f8_334, \5474 );
and \U$3892 ( \5882 , RI2b5e785b7ec8_354, \5476 );
and \U$3893 ( \5883 , RI2b5e785b7568_374, \5478 );
and \U$3894 ( \5884 , RI2b5e785b5df8_394, \5480 );
and \U$3895 ( \5885 , RI2b5e785b5498_414, \5482 );
and \U$3896 ( \5886 , RI2b5e785b4b38_434, \5484 );
and \U$3897 ( \5887 , RI2b5e785b3788_454, \5486 );
and \U$3898 ( \5888 , RI2b5e785b2e28_474, \5488 );
and \U$3899 ( \5889 , RI2b5e785b24c8_494, \5490 );
and \U$3900 ( \5890 , RI2b5e785b14d8_514, \5492 );
and \U$3901 ( \5891 , RI2b5e785b0b78_534, \5494 );
and \U$3902 ( \5892 , RI2b5e785b0218_554, \5496 );
and \U$3903 ( \5893 , RI2b5e785af5e8_574, \5498 );
or \U$3904 ( \5894 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 );
_DC g24d7 ( \5895_nG24d7 , \5894 , \5517 );
buf \U$3905 ( \5896 , \5895_nG24d7 );
and \U$3906 ( \5897 , \5896 , \5873 );
nor \U$3907 ( \5898 , \5876 , \5897 );
and \U$3908 ( \5899 , \5871 , \5833 );
not \U$3909 ( \5900 , \5899 );
and \U$3910 ( \5901 , \5867 , \5900 );
xnor \U$3911 ( \5902 , \5898 , \5901 );
and \U$3912 ( \5903 , \5843 , \5902 );
and \U$3913 ( \5904 , RI2b5e785c0a00_257, \5462 );
and \U$3914 ( \5905 , RI2b5e785be390_277, \5468 );
and \U$3915 ( \5906 , RI2b5e785bc0e0_297, \5470 );
and \U$3916 ( \5907 , RI2b5e785ba1f0_317, \5472 );
and \U$3917 ( \5908 , RI2b5e785b9890_337, \5474 );
and \U$3918 ( \5909 , RI2b5e785b7d60_357, \5476 );
and \U$3919 ( \5910 , RI2b5e785b7400_377, \5478 );
and \U$3920 ( \5911 , RI2b5e785b5c90_397, \5480 );
and \U$3921 ( \5912 , RI2b5e785b5330_417, \5482 );
and \U$3922 ( \5913 , RI2b5e785b49d0_437, \5484 );
and \U$3923 ( \5914 , RI2b5e785b3620_457, \5486 );
and \U$3924 ( \5915 , RI2b5e785b2cc0_477, \5488 );
and \U$3925 ( \5916 , RI2b5e785b2360_497, \5490 );
and \U$3926 ( \5917 , RI2b5e785b1370_517, \5492 );
and \U$3927 ( \5918 , RI2b5e785b0a10_537, \5494 );
and \U$3928 ( \5919 , RI2b5e785b00b0_557, \5496 );
and \U$3929 ( \5920 , RI2b5e785af480_577, \5498 );
or \U$3930 ( \5921 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 );
_DC g226a ( \5922_nG226a , \5921 , \5517 );
buf \U$3931 ( \5923 , \5922_nG226a );
xor \U$3932 ( \5924 , \5206 , \5227 );
xor \U$3933 ( \5925 , \5924 , \5364 );
buf g1d72_GF_PartitionCandidate( \5926_nG1d72 , \5925 );
buf \U$3934 ( \5927 , \5926_nG1d72 );
xor \U$3935 ( \5928 , \5231 , \5252 );
xor \U$3936 ( \5929 , \5928 , \5361 );
buf g1d4e_GF_PartitionCandidate( \5930_nG1d4e , \5929 );
buf \U$3937 ( \5931 , \5930_nG1d4e );
xor \U$3938 ( \5932 , \5927 , \5931 );
xor \U$3939 ( \5933 , \5931 , \5867 );
not \U$3940 ( \5934 , \5933 );
and \U$3941 ( \5935 , \5932 , \5934 );
and \U$3942 ( \5936 , \5923 , \5935 );
and \U$3943 ( \5937 , RI2b5e785c2b48_256, \5462 );
and \U$3944 ( \5938 , RI2b5e785be408_276, \5468 );
and \U$3945 ( \5939 , RI2b5e785bc158_296, \5470 );
and \U$3946 ( \5940 , RI2b5e785ba268_316, \5472 );
and \U$3947 ( \5941 , RI2b5e785b9908_336, \5474 );
and \U$3948 ( \5942 , RI2b5e785b7dd8_356, \5476 );
and \U$3949 ( \5943 , RI2b5e785b7478_376, \5478 );
and \U$3950 ( \5944 , RI2b5e785b5d08_396, \5480 );
and \U$3951 ( \5945 , RI2b5e785b53a8_416, \5482 );
and \U$3952 ( \5946 , RI2b5e785b4a48_436, \5484 );
and \U$3953 ( \5947 , RI2b5e785b3698_456, \5486 );
and \U$3954 ( \5948 , RI2b5e785b2d38_476, \5488 );
and \U$3955 ( \5949 , RI2b5e785b23d8_496, \5490 );
and \U$3956 ( \5950 , RI2b5e785b13e8_516, \5492 );
and \U$3957 ( \5951 , RI2b5e785b0a88_536, \5494 );
and \U$3958 ( \5952 , RI2b5e785b0128_556, \5496 );
and \U$3959 ( \5953 , RI2b5e785af4f8_576, \5498 );
or \U$3960 ( \5954 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 );
_DC g2302 ( \5955_nG2302 , \5954 , \5517 );
buf \U$3961 ( \5956 , \5955_nG2302 );
and \U$3962 ( \5957 , \5956 , \5933 );
nor \U$3963 ( \5958 , \5936 , \5957 );
and \U$3964 ( \5959 , \5931 , \5867 );
not \U$3965 ( \5960 , \5959 );
and \U$3966 ( \5961 , \5927 , \5960 );
xnor \U$3967 ( \5962 , \5958 , \5961 );
and \U$3968 ( \5963 , \5902 , \5962 );
and \U$3969 ( \5964 , \5843 , \5962 );
or \U$3970 ( \5965 , \5903 , \5963 , \5964 );
and \U$3971 ( \5966 , RI2b5e785c0910_259, \5462 );
and \U$3972 ( \5967 , RI2b5e785be2a0_279, \5468 );
and \U$3973 ( \5968 , RI2b5e785bbff0_299, \5470 );
and \U$3974 ( \5969 , RI2b5e785ba100_319, \5472 );
and \U$3975 ( \5970 , RI2b5e785b97a0_339, \5474 );
and \U$3976 ( \5971 , RI2b5e785b7c70_359, \5476 );
and \U$3977 ( \5972 , RI2b5e785b7310_379, \5478 );
and \U$3978 ( \5973 , RI2b5e785b5ba0_399, \5480 );
and \U$3979 ( \5974 , RI2b5e785b5240_419, \5482 );
and \U$3980 ( \5975 , RI2b5e785b48e0_439, \5484 );
and \U$3981 ( \5976 , RI2b5e785b3530_459, \5486 );
and \U$3982 ( \5977 , RI2b5e785b2bd0_479, \5488 );
and \U$3983 ( \5978 , RI2b5e785b2270_499, \5490 );
and \U$3984 ( \5979 , RI2b5e785b1280_519, \5492 );
and \U$3985 ( \5980 , RI2b5e785b0920_539, \5494 );
and \U$3986 ( \5981 , RI2b5e785affc0_559, \5496 );
and \U$3987 ( \5982 , RI2b5e785af390_579, \5498 );
or \U$3988 ( \5983 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 );
_DC g209f ( \5984_nG209f , \5983 , \5517 );
buf \U$3989 ( \5985 , \5984_nG209f );
xor \U$3990 ( \5986 , \5181 , \5202 );
xor \U$3991 ( \5987 , \5986 , \5367 );
buf g1ebd_GF_PartitionCandidate( \5988_nG1ebd , \5987 );
buf \U$3992 ( \5989 , \5988_nG1ebd );
xor \U$3993 ( \5990 , \5691 , \5989 );
xor \U$3994 ( \5991 , \5989 , \5927 );
not \U$3995 ( \5992 , \5991 );
and \U$3996 ( \5993 , \5990 , \5992 );
and \U$3997 ( \5994 , \5985 , \5993 );
and \U$3998 ( \5995 , RI2b5e785c0988_258, \5462 );
and \U$3999 ( \5996 , RI2b5e785be318_278, \5468 );
and \U$4000 ( \5997 , RI2b5e785bc068_298, \5470 );
and \U$4001 ( \5998 , RI2b5e785ba178_318, \5472 );
and \U$4002 ( \5999 , RI2b5e785b9818_338, \5474 );
and \U$4003 ( \6000 , RI2b5e785b7ce8_358, \5476 );
and \U$4004 ( \6001 , RI2b5e785b7388_378, \5478 );
and \U$4005 ( \6002 , RI2b5e785b5c18_398, \5480 );
and \U$4006 ( \6003 , RI2b5e785b52b8_418, \5482 );
and \U$4007 ( \6004 , RI2b5e785b4958_438, \5484 );
and \U$4008 ( \6005 , RI2b5e785b35a8_458, \5486 );
and \U$4009 ( \6006 , RI2b5e785b2c48_478, \5488 );
and \U$4010 ( \6007 , RI2b5e785b22e8_498, \5490 );
and \U$4011 ( \6008 , RI2b5e785b12f8_518, \5492 );
and \U$4012 ( \6009 , RI2b5e785b0998_538, \5494 );
and \U$4013 ( \6010 , RI2b5e785b0038_558, \5496 );
and \U$4014 ( \6011 , RI2b5e785af408_578, \5498 );
or \U$4015 ( \6012 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 );
_DC g2129 ( \6013_nG2129 , \6012 , \5517 );
buf \U$4016 ( \6014 , \6013_nG2129 );
and \U$4017 ( \6015 , \6014 , \5991 );
nor \U$4018 ( \6016 , \5994 , \6015 );
and \U$4019 ( \6017 , \5989 , \5927 );
not \U$4020 ( \6018 , \6017 );
and \U$4021 ( \6019 , \5691 , \6018 );
xnor \U$4022 ( \6020 , \6016 , \6019 );
and \U$4023 ( \6021 , RI2b5e785c0820_261, \5462 );
and \U$4024 ( \6022 , RI2b5e785be1b0_281, \5468 );
and \U$4025 ( \6023 , RI2b5e785bbf00_301, \5470 );
and \U$4026 ( \6024 , RI2b5e785ba010_321, \5472 );
and \U$4027 ( \6025 , RI2b5e785b96b0_341, \5474 );
and \U$4028 ( \6026 , RI2b5e785b7b80_361, \5476 );
and \U$4029 ( \6027 , RI2b5e785b7220_381, \5478 );
and \U$4030 ( \6028 , RI2b5e785b5ab0_401, \5480 );
and \U$4031 ( \6029 , RI2b5e785b5150_421, \5482 );
and \U$4032 ( \6030 , RI2b5e785b47f0_441, \5484 );
and \U$4033 ( \6031 , RI2b5e785b3440_461, \5486 );
and \U$4034 ( \6032 , RI2b5e785b2ae0_481, \5488 );
and \U$4035 ( \6033 , RI2b5e785b2180_501, \5490 );
and \U$4036 ( \6034 , RI2b5e785b1190_521, \5492 );
and \U$4037 ( \6035 , RI2b5e785b0830_541, \5494 );
and \U$4038 ( \6036 , RI2b5e785afed0_561, \5496 );
and \U$4039 ( \6037 , RI2b5e785af2a0_581, \5498 );
or \U$4040 ( \6038 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 );
_DC g1efc ( \6039_nG1efc , \6038 , \5517 );
buf \U$4041 ( \6040 , \6039_nG1efc );
and \U$4042 ( \6041 , \6040 , \5694 );
and \U$4043 ( \6042 , RI2b5e785c0898_260, \5462 );
and \U$4044 ( \6043 , RI2b5e785be228_280, \5468 );
and \U$4045 ( \6044 , RI2b5e785bbf78_300, \5470 );
and \U$4046 ( \6045 , RI2b5e785ba088_320, \5472 );
and \U$4047 ( \6046 , RI2b5e785b9728_340, \5474 );
and \U$4048 ( \6047 , RI2b5e785b7bf8_360, \5476 );
and \U$4049 ( \6048 , RI2b5e785b7298_380, \5478 );
and \U$4050 ( \6049 , RI2b5e785b5b28_400, \5480 );
and \U$4051 ( \6050 , RI2b5e785b51c8_420, \5482 );
and \U$4052 ( \6051 , RI2b5e785b4868_440, \5484 );
and \U$4053 ( \6052 , RI2b5e785b34b8_460, \5486 );
and \U$4054 ( \6053 , RI2b5e785b2b58_480, \5488 );
and \U$4055 ( \6054 , RI2b5e785b21f8_500, \5490 );
and \U$4056 ( \6055 , RI2b5e785b1208_520, \5492 );
and \U$4057 ( \6056 , RI2b5e785b08a8_540, \5494 );
and \U$4058 ( \6057 , RI2b5e785aff48_560, \5496 );
and \U$4059 ( \6058 , RI2b5e785af318_580, \5498 );
or \U$4060 ( \6059 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 );
_DC g1f70 ( \6060_nG1f70 , \6059 , \5517 );
buf \U$4061 ( \6061 , \6060_nG1f70 );
and \U$4062 ( \6062 , \6061 , \5692 );
nor \U$4063 ( \6063 , \6041 , \6062 );
xnor \U$4064 ( \6064 , \6063 , \5699 );
and \U$4065 ( \6065 , \6020 , \6064 );
and \U$4066 ( \6066 , RI2b5e785c0730_263, \5462 );
and \U$4067 ( \6067 , RI2b5e785be0c0_283, \5468 );
and \U$4068 ( \6068 , RI2b5e785bbe10_303, \5470 );
and \U$4069 ( \6069 , RI2b5e785b9f20_323, \5472 );
and \U$4070 ( \6070 , RI2b5e785b95c0_343, \5474 );
and \U$4071 ( \6071 , RI2b5e785b7a90_363, \5476 );
and \U$4072 ( \6072 , RI2b5e785b7130_383, \5478 );
and \U$4073 ( \6073 , RI2b5e785b59c0_403, \5480 );
and \U$4074 ( \6074 , RI2b5e785b5060_423, \5482 );
and \U$4075 ( \6075 , RI2b5e785b3cb0_443, \5484 );
and \U$4076 ( \6076 , RI2b5e785b3350_463, \5486 );
and \U$4077 ( \6077 , RI2b5e785b29f0_483, \5488 );
and \U$4078 ( \6078 , RI2b5e785b1a00_503, \5490 );
and \U$4079 ( \6079 , RI2b5e785b10a0_523, \5492 );
and \U$4080 ( \6080 , RI2b5e785b0740_543, \5494 );
and \U$4081 ( \6081 , RI2b5e785afde0_563, \5496 );
and \U$4082 ( \6082 , RI2b5e785af1b0_583, \5498 );
or \U$4083 ( \6083 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 );
_DC g1d8b ( \6084_nG1d8b , \6083 , \5517 );
buf \U$4084 ( \6085 , \6084_nG1d8b );
and \U$4085 ( \6086 , \6085 , \5629 );
and \U$4086 ( \6087 , RI2b5e785c07a8_262, \5462 );
and \U$4087 ( \6088 , RI2b5e785be138_282, \5468 );
and \U$4088 ( \6089 , RI2b5e785bbe88_302, \5470 );
and \U$4089 ( \6090 , RI2b5e785b9f98_322, \5472 );
and \U$4090 ( \6091 , RI2b5e785b9638_342, \5474 );
and \U$4091 ( \6092 , RI2b5e785b7b08_362, \5476 );
and \U$4092 ( \6093 , RI2b5e785b71a8_382, \5478 );
and \U$4093 ( \6094 , RI2b5e785b5a38_402, \5480 );
and \U$4094 ( \6095 , RI2b5e785b50d8_422, \5482 );
and \U$4095 ( \6096 , RI2b5e785b4778_442, \5484 );
and \U$4096 ( \6097 , RI2b5e785b33c8_462, \5486 );
and \U$4097 ( \6098 , RI2b5e785b2a68_482, \5488 );
and \U$4098 ( \6099 , RI2b5e785b1a78_502, \5490 );
and \U$4099 ( \6100 , RI2b5e785b1118_522, \5492 );
and \U$4100 ( \6101 , RI2b5e785b07b8_542, \5494 );
and \U$4101 ( \6102 , RI2b5e785afe58_562, \5496 );
and \U$4102 ( \6103 , RI2b5e785af228_582, \5498 );
or \U$4103 ( \6104 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 );
_DC g1df2 ( \6105_nG1df2 , \6104 , \5517 );
buf \U$4104 ( \6106 , \6105_nG1df2 );
and \U$4105 ( \6107 , \6106 , \5627 );
nor \U$4106 ( \6108 , \6086 , \6107 );
xnor \U$4107 ( \6109 , \6108 , \5396 );
and \U$4108 ( \6110 , \6064 , \6109 );
and \U$4109 ( \6111 , \6020 , \6109 );
or \U$4110 ( \6112 , \6065 , \6110 , \6111 );
and \U$4111 ( \6113 , \5965 , \6112 );
and \U$4112 ( \6114 , RI2b5e785c0640_265, \5462 );
and \U$4113 ( \6115 , RI2b5e785bdfd0_285, \5468 );
and \U$4114 ( \6116 , RI2b5e785bbd20_305, \5470 );
and \U$4115 ( \6117 , RI2b5e785b9e30_325, \5472 );
and \U$4116 ( \6118 , RI2b5e785b94d0_345, \5474 );
and \U$4117 ( \6119 , RI2b5e785b79a0_365, \5476 );
and \U$4118 ( \6120 , RI2b5e785b7040_385, \5478 );
and \U$4119 ( \6121 , RI2b5e785b58d0_405, \5480 );
and \U$4120 ( \6122 , RI2b5e785b4f70_425, \5482 );
and \U$4121 ( \6123 , RI2b5e785b3bc0_445, \5484 );
and \U$4122 ( \6124 , RI2b5e785b3260_465, \5486 );
and \U$4123 ( \6125 , RI2b5e785b2900_485, \5488 );
and \U$4124 ( \6126 , RI2b5e785b1910_505, \5490 );
and \U$4125 ( \6127 , RI2b5e785b0fb0_525, \5492 );
and \U$4126 ( \6128 , RI2b5e785b0650_545, \5494 );
and \U$4127 ( \6129 , RI2b5e785afcf0_565, \5496 );
and \U$4128 ( \6130 , RI2b5e785af0c0_585, \5498 );
or \U$4129 ( \6131 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 );
_DC g1c0d ( \6132_nG1c0d , \6131 , \5517 );
buf \U$4130 ( \6133 , \6132_nG1c0d );
and \U$4131 ( \6134 , \6133 , \5567 );
and \U$4132 ( \6135 , RI2b5e785c06b8_264, \5462 );
and \U$4133 ( \6136 , RI2b5e785be048_284, \5468 );
and \U$4134 ( \6137 , RI2b5e785bbd98_304, \5470 );
and \U$4135 ( \6138 , RI2b5e785b9ea8_324, \5472 );
and \U$4136 ( \6139 , RI2b5e785b9548_344, \5474 );
and \U$4137 ( \6140 , RI2b5e785b7a18_364, \5476 );
and \U$4138 ( \6141 , RI2b5e785b70b8_384, \5478 );
and \U$4139 ( \6142 , RI2b5e785b5948_404, \5480 );
and \U$4140 ( \6143 , RI2b5e785b4fe8_424, \5482 );
and \U$4141 ( \6144 , RI2b5e785b3c38_444, \5484 );
and \U$4142 ( \6145 , RI2b5e785b32d8_464, \5486 );
and \U$4143 ( \6146 , RI2b5e785b2978_484, \5488 );
and \U$4144 ( \6147 , RI2b5e785b1988_504, \5490 );
and \U$4145 ( \6148 , RI2b5e785b1028_524, \5492 );
and \U$4146 ( \6149 , RI2b5e785b06c8_544, \5494 );
and \U$4147 ( \6150 , RI2b5e785afd68_564, \5496 );
and \U$4148 ( \6151 , RI2b5e785af138_584, \5498 );
or \U$4149 ( \6152 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 );
_DC g1ca0 ( \6153_nG1ca0 , \6152 , \5517 );
buf \U$4150 ( \6154 , \6153_nG1ca0 );
and \U$4151 ( \6155 , \6154 , \5565 );
nor \U$4152 ( \6156 , \6134 , \6155 );
xnor \U$4153 ( \6157 , \6156 , \5593 );
and \U$4155 ( \6158 , RI2b5e785c05c8_266, \5462 );
and \U$4156 ( \6159 , RI2b5e785bdf58_286, \5468 );
and \U$4157 ( \6160 , RI2b5e785bbca8_306, \5470 );
and \U$4158 ( \6161 , RI2b5e785b9db8_326, \5472 );
and \U$4159 ( \6162 , RI2b5e785b9458_346, \5474 );
and \U$4160 ( \6163 , RI2b5e785b7928_366, \5476 );
and \U$4161 ( \6164 , RI2b5e785b6fc8_386, \5478 );
and \U$4162 ( \6165 , RI2b5e785b5858_406, \5480 );
and \U$4163 ( \6166 , RI2b5e785b4ef8_426, \5482 );
and \U$4164 ( \6167 , RI2b5e785b3b48_446, \5484 );
and \U$4165 ( \6168 , RI2b5e785b31e8_466, \5486 );
and \U$4166 ( \6169 , RI2b5e785b2888_486, \5488 );
and \U$4167 ( \6170 , RI2b5e785b1898_506, \5490 );
and \U$4168 ( \6171 , RI2b5e785b0f38_526, \5492 );
and \U$4169 ( \6172 , RI2b5e785b05d8_546, \5494 );
and \U$4170 ( \6173 , RI2b5e785afc78_566, \5496 );
and \U$4171 ( \6174 , RI2b5e785af048_586, \5498 );
or \U$4172 ( \6175 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 );
_DC g1b85 ( \6176_nG1b85 , \6175 , \5517 );
buf \U$4173 ( \6177 , \6176_nG1b85 );
and \U$4174 ( \6178 , \6177 , \5620 );
nor \U$4175 ( \6179 , 1'b0 , \6178 );
xnor \U$4176 ( \6180 , \6179 , 1'b0 );
and \U$4177 ( \6181 , \6157 , \6180 );
and \U$4178 ( \6182 , \6112 , \6181 );
and \U$4179 ( \6183 , \5965 , \6181 );
or \U$4180 ( \6184 , \6113 , \6182 , \6183 );
and \U$4182 ( \6185 , \6106 , \5629 );
and \U$4183 ( \6186 , \6040 , \5627 );
nor \U$4184 ( \6187 , \6185 , \6186 );
xnor \U$4185 ( \6188 , \6187 , \5396 );
and \U$4186 ( \6189 , \6154 , \5567 );
and \U$4187 ( \6190 , \6085 , \5565 );
nor \U$4188 ( \6191 , \6189 , \6190 );
xnor \U$4189 ( \6192 , \6191 , \5593 );
xor \U$4190 ( \6193 , \6188 , \6192 );
and \U$4192 ( \6194 , \6133 , \5620 );
nor \U$4193 ( \6195 , 1'b0 , \6194 );
xnor \U$4194 ( \6196 , \6195 , 1'b0 );
xor \U$4195 ( \6197 , \6193 , \6196 );
and \U$4196 ( \6198 , \5956 , \5935 );
and \U$4197 ( \6199 , \5863 , \5933 );
nor \U$4198 ( \6200 , \6198 , \6199 );
xnor \U$4199 ( \6201 , \6200 , \5961 );
and \U$4200 ( \6202 , \6014 , \5993 );
and \U$4201 ( \6203 , \5923 , \5991 );
nor \U$4202 ( \6204 , \6202 , \6203 );
xnor \U$4203 ( \6205 , \6204 , \6019 );
xor \U$4204 ( \6206 , \6201 , \6205 );
and \U$4205 ( \6207 , \6061 , \5694 );
and \U$4206 ( \6208 , \5985 , \5692 );
nor \U$4207 ( \6209 , \6207 , \6208 );
xnor \U$4208 ( \6210 , \6209 , \5699 );
xor \U$4209 ( \6211 , \6206 , \6210 );
and \U$4210 ( \6212 , \6197 , \6211 );
or \U$4212 ( \6213 , 1'b0 , \6212 , 1'b0 );
xor \U$4213 ( \6214 , \6184 , \6213 );
and \U$4214 ( \6215 , \6085 , \5567 );
and \U$4215 ( \6216 , \6106 , \5565 );
nor \U$4216 ( \6217 , \6215 , \6216 );
xnor \U$4217 ( \6218 , \6217 , \5593 );
and \U$4219 ( \6219 , \6154 , \5620 );
nor \U$4220 ( \6220 , 1'b0 , \6219 );
xnor \U$4221 ( \6221 , \6220 , 1'b0 );
xor \U$4222 ( \6222 , \6218 , \6221 );
xor \U$4224 ( \6223 , \6222 , 1'b0 );
and \U$4225 ( \6224 , \5923 , \5993 );
and \U$4226 ( \6225 , \5956 , \5991 );
nor \U$4227 ( \6226 , \6224 , \6225 );
xnor \U$4228 ( \6227 , \6226 , \6019 );
and \U$4229 ( \6228 , \5985 , \5694 );
and \U$4230 ( \6229 , \6014 , \5692 );
nor \U$4231 ( \6230 , \6228 , \6229 );
xnor \U$4232 ( \6231 , \6230 , \5699 );
xor \U$4233 ( \6232 , \6227 , \6231 );
and \U$4234 ( \6233 , \6040 , \5629 );
and \U$4235 ( \6234 , \6061 , \5627 );
nor \U$4236 ( \6235 , \6233 , \6234 );
xnor \U$4237 ( \6236 , \6235 , \5396 );
xor \U$4238 ( \6237 , \6232 , \6236 );
xor \U$4239 ( \6238 , \6223 , \6237 );
and \U$4240 ( \6239 , \5747 , \5839 );
and \U$4241 ( \6240 , \5615 , \5836 );
nor \U$4242 ( \6241 , \6239 , \6240 );
xnor \U$4243 ( \6242 , \6241 , \5833 );
and \U$4244 ( \6243 , \5770 , \5875 );
and \U$4245 ( \6244 , \5726 , \5873 );
nor \U$4246 ( \6245 , \6243 , \6244 );
xnor \U$4247 ( \6246 , \6245 , \5901 );
xor \U$4248 ( \6247 , \6242 , \6246 );
and \U$4249 ( \6248 , \5863 , \5935 );
and \U$4250 ( \6249 , \5896 , \5933 );
nor \U$4251 ( \6250 , \6248 , \6249 );
xnor \U$4252 ( \6251 , \6250 , \5961 );
xor \U$4253 ( \6252 , \6247 , \6251 );
xor \U$4254 ( \6253 , \6238 , \6252 );
xor \U$4255 ( \6254 , \6214 , \6253 );
and \U$4257 ( \6255 , \5896 , \5839 );
and \U$4258 ( \6256 , \5770 , \5836 );
nor \U$4259 ( \6257 , \6255 , \6256 );
xnor \U$4260 ( \6258 , \6257 , \5833 );
and \U$4261 ( \6259 , \5956 , \5875 );
and \U$4262 ( \6260 , \5863 , \5873 );
nor \U$4263 ( \6261 , \6259 , \6260 );
xnor \U$4264 ( \6262 , \6261 , \5901 );
and \U$4265 ( \6263 , \6258 , \6262 );
or \U$4267 ( \6264 , 1'b0 , \6263 , 1'b0 );
and \U$4268 ( \6265 , \6014 , \5935 );
and \U$4269 ( \6266 , \5923 , \5933 );
nor \U$4270 ( \6267 , \6265 , \6266 );
xnor \U$4271 ( \6268 , \6267 , \5961 );
and \U$4272 ( \6269 , \6061 , \5993 );
and \U$4273 ( \6270 , \5985 , \5991 );
nor \U$4274 ( \6271 , \6269 , \6270 );
xnor \U$4275 ( \6272 , \6271 , \6019 );
and \U$4276 ( \6273 , \6268 , \6272 );
and \U$4277 ( \6274 , \6106 , \5694 );
and \U$4278 ( \6275 , \6040 , \5692 );
nor \U$4279 ( \6276 , \6274 , \6275 );
xnor \U$4280 ( \6277 , \6276 , \5699 );
and \U$4281 ( \6278 , \6272 , \6277 );
and \U$4282 ( \6279 , \6268 , \6277 );
or \U$4283 ( \6280 , \6273 , \6278 , \6279 );
and \U$4284 ( \6281 , \6264 , \6280 );
and \U$4285 ( \6282 , \6154 , \5629 );
and \U$4286 ( \6283 , \6085 , \5627 );
nor \U$4287 ( \6284 , \6282 , \6283 );
xnor \U$4288 ( \6285 , \6284 , \5396 );
and \U$4289 ( \6286 , \6177 , \5567 );
and \U$4290 ( \6287 , \6133 , \5565 );
nor \U$4291 ( \6288 , \6286 , \6287 );
xnor \U$4292 ( \6289 , \6288 , \5593 );
and \U$4293 ( \6290 , \6285 , \6289 );
and \U$4294 ( \6291 , RI2b5e785c0550_267, \5462 );
and \U$4295 ( \6292 , RI2b5e785bc590_287, \5468 );
and \U$4296 ( \6293 , RI2b5e785bbc30_307, \5470 );
and \U$4297 ( \6294 , RI2b5e785b9d40_327, \5472 );
and \U$4298 ( \6295 , RI2b5e785b93e0_347, \5474 );
and \U$4299 ( \6296 , RI2b5e785b78b0_367, \5476 );
and \U$4300 ( \6297 , RI2b5e785b6f50_387, \5478 );
and \U$4301 ( \6298 , RI2b5e785b57e0_407, \5480 );
and \U$4302 ( \6299 , RI2b5e785b4e80_427, \5482 );
and \U$4303 ( \6300 , RI2b5e785b3ad0_447, \5484 );
and \U$4304 ( \6301 , RI2b5e785b3170_467, \5486 );
and \U$4305 ( \6302 , RI2b5e785b2810_487, \5488 );
and \U$4306 ( \6303 , RI2b5e785b1820_507, \5490 );
and \U$4307 ( \6304 , RI2b5e785b0ec0_527, \5492 );
and \U$4308 ( \6305 , RI2b5e785b0560_547, \5494 );
and \U$4309 ( \6306 , RI2b5e785afc00_567, \5496 );
and \U$4310 ( \6307 , RI2b5e785aefd0_587, \5498 );
or \U$4311 ( \6308 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 );
_DC g1aea ( \6309_nG1aea , \6308 , \5517 );
buf \U$4312 ( \6310 , \6309_nG1aea );
nand \U$4313 ( \6311 , \6310 , \5620 );
xnor \U$4314 ( \6312 , \6311 , 1'b0 );
and \U$4315 ( \6313 , \6289 , \6312 );
and \U$4316 ( \6314 , \6285 , \6312 );
or \U$4317 ( \6315 , \6290 , \6313 , \6314 );
and \U$4318 ( \6316 , \6280 , \6315 );
and \U$4319 ( \6317 , \6264 , \6315 );
or \U$4320 ( \6318 , \6281 , \6316 , \6317 );
xor \U$4321 ( \6319 , \6157 , \6180 );
xor \U$4322 ( \6320 , \6020 , \6064 );
xor \U$4323 ( \6321 , \6320 , \6109 );
and \U$4324 ( \6322 , \6319 , \6321 );
xor \U$4325 ( \6323 , \5843 , \5902 );
xor \U$4326 ( \6324 , \6323 , \5962 );
and \U$4327 ( \6325 , \6321 , \6324 );
and \U$4328 ( \6326 , \6319 , \6324 );
or \U$4329 ( \6327 , \6322 , \6325 , \6326 );
and \U$4330 ( \6328 , \6318 , \6327 );
and \U$4332 ( \6329 , \5726 , \5839 );
and \U$4333 ( \6330 , \5747 , \5836 );
nor \U$4334 ( \6331 , \6329 , \6330 );
xnor \U$4335 ( \6332 , \6331 , \5833 );
xor \U$4336 ( \6333 , 1'b0 , \6332 );
and \U$4337 ( \6334 , \5896 , \5875 );
and \U$4338 ( \6335 , \5770 , \5873 );
nor \U$4339 ( \6336 , \6334 , \6335 );
xnor \U$4340 ( \6337 , \6336 , \5901 );
xor \U$4341 ( \6338 , \6333 , \6337 );
and \U$4342 ( \6339 , \6327 , \6338 );
and \U$4343 ( \6340 , \6318 , \6338 );
or \U$4344 ( \6341 , \6328 , \6339 , \6340 );
xor \U$4346 ( \6342 , 1'b0 , \6197 );
xor \U$4347 ( \6343 , \6342 , \6211 );
xor \U$4348 ( \6344 , \5965 , \6112 );
xor \U$4349 ( \6345 , \6344 , \6181 );
and \U$4350 ( \6346 , \6343 , \6345 );
xor \U$4351 ( \6347 , \6341 , \6346 );
and \U$4353 ( \6348 , \6332 , \6337 );
or \U$4355 ( \6349 , 1'b0 , \6348 , 1'b0 );
and \U$4356 ( \6350 , \6201 , \6205 );
and \U$4357 ( \6351 , \6205 , \6210 );
and \U$4358 ( \6352 , \6201 , \6210 );
or \U$4359 ( \6353 , \6350 , \6351 , \6352 );
xor \U$4360 ( \6354 , \6349 , \6353 );
and \U$4361 ( \6355 , \6188 , \6192 );
and \U$4362 ( \6356 , \6192 , \6196 );
and \U$4363 ( \6357 , \6188 , \6196 );
or \U$4364 ( \6358 , \6355 , \6356 , \6357 );
xor \U$4365 ( \6359 , \6354 , \6358 );
xor \U$4366 ( \6360 , \6347 , \6359 );
xor \U$4367 ( \6361 , \6254 , \6360 );
and \U$4368 ( \6362 , \5863 , \5839 );
and \U$4369 ( \6363 , \5896 , \5836 );
nor \U$4370 ( \6364 , \6362 , \6363 );
xnor \U$4371 ( \6365 , \6364 , \5833 );
and \U$4372 ( \6366 , \5923 , \5875 );
and \U$4373 ( \6367 , \5956 , \5873 );
nor \U$4374 ( \6368 , \6366 , \6367 );
xnor \U$4375 ( \6369 , \6368 , \5901 );
and \U$4376 ( \6370 , \6365 , \6369 );
and \U$4377 ( \6371 , \5985 , \5935 );
and \U$4378 ( \6372 , \6014 , \5933 );
nor \U$4379 ( \6373 , \6371 , \6372 );
xnor \U$4380 ( \6374 , \6373 , \5961 );
and \U$4381 ( \6375 , \6369 , \6374 );
and \U$4382 ( \6376 , \6365 , \6374 );
or \U$4383 ( \6377 , \6370 , \6375 , \6376 );
and \U$4384 ( \6378 , \6040 , \5993 );
and \U$4385 ( \6379 , \6061 , \5991 );
nor \U$4386 ( \6380 , \6378 , \6379 );
xnor \U$4387 ( \6381 , \6380 , \6019 );
and \U$4388 ( \6382 , \6085 , \5694 );
and \U$4389 ( \6383 , \6106 , \5692 );
nor \U$4390 ( \6384 , \6382 , \6383 );
xnor \U$4391 ( \6385 , \6384 , \5699 );
and \U$4392 ( \6386 , \6381 , \6385 );
and \U$4393 ( \6387 , \6133 , \5629 );
and \U$4394 ( \6388 , \6154 , \5627 );
nor \U$4395 ( \6389 , \6387 , \6388 );
xnor \U$4396 ( \6390 , \6389 , \5396 );
and \U$4397 ( \6391 , \6385 , \6390 );
and \U$4398 ( \6392 , \6381 , \6390 );
or \U$4399 ( \6393 , \6386 , \6391 , \6392 );
and \U$4400 ( \6394 , \6377 , \6393 );
xor \U$4401 ( \6395 , \6285 , \6289 );
xor \U$4402 ( \6396 , \6395 , \6312 );
and \U$4403 ( \6397 , \6393 , \6396 );
and \U$4404 ( \6398 , \6377 , \6396 );
or \U$4405 ( \6399 , \6394 , \6397 , \6398 );
xor \U$4406 ( \6400 , \6268 , \6272 );
xor \U$4407 ( \6401 , \6400 , \6277 );
xor \U$4408 ( \6402 , 1'b0 , \6258 );
xor \U$4409 ( \6403 , \6402 , \6262 );
and \U$4410 ( \6404 , \6401 , \6403 );
and \U$4411 ( \6405 , \6399 , \6404 );
xor \U$4412 ( \6406 , \6319 , \6321 );
xor \U$4413 ( \6407 , \6406 , \6324 );
and \U$4414 ( \6408 , \6404 , \6407 );
and \U$4415 ( \6409 , \6399 , \6407 );
or \U$4416 ( \6410 , \6405 , \6408 , \6409 );
xor \U$4417 ( \6411 , \6343 , \6345 );
and \U$4418 ( \6412 , \6410 , \6411 );
xor \U$4419 ( \6413 , \6318 , \6327 );
xor \U$4420 ( \6414 , \6413 , \6338 );
and \U$4421 ( \6415 , \6411 , \6414 );
and \U$4422 ( \6416 , \6410 , \6414 );
or \U$4423 ( \6417 , \6412 , \6415 , \6416 );
nor \U$4424 ( \6418 , \6361 , \6417 );
and \U$4425 ( \6419 , \6341 , \6346 );
and \U$4426 ( \6420 , \6346 , \6359 );
and \U$4427 ( \6421 , \6341 , \6359 );
or \U$4428 ( \6422 , \6419 , \6420 , \6421 );
and \U$4429 ( \6423 , \6184 , \6213 );
and \U$4430 ( \6424 , \6213 , \6253 );
and \U$4431 ( \6425 , \6184 , \6253 );
or \U$4432 ( \6426 , \6423 , \6424 , \6425 );
and \U$4434 ( \6427 , \5615 , \5839 );
and \U$4435 ( \6428 , \5519 , \5836 );
nor \U$4436 ( \6429 , \6427 , \6428 );
xnor \U$4437 ( \6430 , \6429 , \5833 );
xor \U$4438 ( \6431 , 1'b0 , \6430 );
and \U$4439 ( \6432 , \5726 , \5875 );
and \U$4440 ( \6433 , \5747 , \5873 );
nor \U$4441 ( \6434 , \6432 , \6433 );
xnor \U$4442 ( \6435 , \6434 , \5901 );
xor \U$4443 ( \6436 , \6431 , \6435 );
and \U$4445 ( \6437 , \6061 , \5629 );
and \U$4446 ( \6438 , \5985 , \5627 );
nor \U$4447 ( \6439 , \6437 , \6438 );
xnor \U$4448 ( \6440 , \6439 , \5396 );
and \U$4449 ( \6441 , \6106 , \5567 );
and \U$4450 ( \6442 , \6040 , \5565 );
nor \U$4451 ( \6443 , \6441 , \6442 );
xnor \U$4452 ( \6444 , \6443 , \5593 );
xor \U$4453 ( \6445 , \6440 , \6444 );
and \U$4455 ( \6446 , \6085 , \5620 );
nor \U$4456 ( \6447 , 1'b0 , \6446 );
xnor \U$4457 ( \6448 , \6447 , 1'b0 );
xor \U$4458 ( \6449 , \6445 , \6448 );
xor \U$4459 ( \6450 , 1'b0 , \6449 );
xor \U$4460 ( \6451 , \6436 , \6450 );
and \U$4461 ( \6452 , \6242 , \6246 );
and \U$4462 ( \6453 , \6246 , \6251 );
and \U$4463 ( \6454 , \6242 , \6251 );
or \U$4464 ( \6455 , \6452 , \6453 , \6454 );
and \U$4465 ( \6456 , \6227 , \6231 );
and \U$4466 ( \6457 , \6231 , \6236 );
and \U$4467 ( \6458 , \6227 , \6236 );
or \U$4468 ( \6459 , \6456 , \6457 , \6458 );
xor \U$4469 ( \6460 , \6455 , \6459 );
and \U$4470 ( \6461 , \6218 , \6221 );
or \U$4473 ( \6462 , \6461 , 1'b0 , 1'b0 );
xor \U$4474 ( \6463 , \6460 , \6462 );
xor \U$4475 ( \6464 , \6451 , \6463 );
xor \U$4476 ( \6465 , \6426 , \6464 );
and \U$4477 ( \6466 , \6349 , \6353 );
and \U$4478 ( \6467 , \6353 , \6358 );
and \U$4479 ( \6468 , \6349 , \6358 );
or \U$4480 ( \6469 , \6466 , \6467 , \6468 );
and \U$4481 ( \6470 , \6223 , \6237 );
and \U$4482 ( \6471 , \6237 , \6252 );
and \U$4483 ( \6472 , \6223 , \6252 );
or \U$4484 ( \6473 , \6470 , \6471 , \6472 );
xor \U$4485 ( \6474 , \6469 , \6473 );
and \U$4486 ( \6475 , \5896 , \5935 );
and \U$4487 ( \6476 , \5770 , \5933 );
nor \U$4488 ( \6477 , \6475 , \6476 );
xnor \U$4489 ( \6478 , \6477 , \5961 );
and \U$4490 ( \6479 , \5956 , \5993 );
and \U$4491 ( \6480 , \5863 , \5991 );
nor \U$4492 ( \6481 , \6479 , \6480 );
xnor \U$4493 ( \6482 , \6481 , \6019 );
xor \U$4494 ( \6483 , \6478 , \6482 );
and \U$4495 ( \6484 , \6014 , \5694 );
and \U$4496 ( \6485 , \5923 , \5692 );
nor \U$4497 ( \6486 , \6484 , \6485 );
xnor \U$4498 ( \6487 , \6486 , \5699 );
xor \U$4499 ( \6488 , \6483 , \6487 );
xor \U$4500 ( \6489 , \6474 , \6488 );
xor \U$4501 ( \6490 , \6465 , \6489 );
xor \U$4502 ( \6491 , \6422 , \6490 );
and \U$4503 ( \6492 , \6254 , \6360 );
nor \U$4504 ( \6493 , \6491 , \6492 );
nor \U$4505 ( \6494 , \6418 , \6493 );
and \U$4506 ( \6495 , \6426 , \6464 );
and \U$4507 ( \6496 , \6464 , \6489 );
and \U$4508 ( \6497 , \6426 , \6489 );
or \U$4509 ( \6498 , \6495 , \6496 , \6497 );
and \U$4511 ( \6499 , \6430 , \6435 );
or \U$4513 ( \6500 , 1'b0 , \6499 , 1'b0 );
and \U$4514 ( \6501 , \6478 , \6482 );
and \U$4515 ( \6502 , \6482 , \6487 );
and \U$4516 ( \6503 , \6478 , \6487 );
or \U$4517 ( \6504 , \6501 , \6502 , \6503 );
xor \U$4518 ( \6505 , \6500 , \6504 );
and \U$4519 ( \6506 , \6440 , \6444 );
and \U$4520 ( \6507 , \6444 , \6448 );
and \U$4521 ( \6508 , \6440 , \6448 );
or \U$4522 ( \6509 , \6506 , \6507 , \6508 );
xor \U$4523 ( \6510 , \6505 , \6509 );
and \U$4524 ( \6511 , \6455 , \6459 );
and \U$4525 ( \6512 , \6459 , \6462 );
and \U$4526 ( \6513 , \6455 , \6462 );
or \U$4527 ( \6514 , \6511 , \6512 , \6513 );
xor \U$4529 ( \6515 , \6514 , 1'b0 );
and \U$4530 ( \6516 , \5519 , \5839 );
and \U$4531 ( \6517 , \5588 , \5836 );
nor \U$4532 ( \6518 , \6516 , \6517 );
xnor \U$4533 ( \6519 , \6518 , \5833 );
and \U$4534 ( \6520 , \5747 , \5875 );
and \U$4535 ( \6521 , \5615 , \5873 );
nor \U$4536 ( \6522 , \6520 , \6521 );
xnor \U$4537 ( \6523 , \6522 , \5901 );
xor \U$4538 ( \6524 , \6519 , \6523 );
and \U$4539 ( \6525 , \5770 , \5935 );
and \U$4540 ( \6526 , \5726 , \5933 );
nor \U$4541 ( \6527 , \6525 , \6526 );
xnor \U$4542 ( \6528 , \6527 , \5961 );
xor \U$4543 ( \6529 , \6524 , \6528 );
xor \U$4544 ( \6530 , \6515 , \6529 );
xor \U$4545 ( \6531 , \6510 , \6530 );
xor \U$4546 ( \6532 , \6498 , \6531 );
and \U$4547 ( \6533 , \6469 , \6473 );
and \U$4548 ( \6534 , \6473 , \6488 );
and \U$4549 ( \6535 , \6469 , \6488 );
or \U$4550 ( \6536 , \6533 , \6534 , \6535 );
and \U$4551 ( \6537 , \6436 , \6450 );
and \U$4552 ( \6538 , \6450 , \6463 );
and \U$4553 ( \6539 , \6436 , \6463 );
or \U$4554 ( \6540 , \6537 , \6538 , \6539 );
xor \U$4555 ( \6541 , \6536 , \6540 );
and \U$4557 ( \6542 , \6040 , \5567 );
and \U$4558 ( \6543 , \6061 , \5565 );
nor \U$4559 ( \6544 , \6542 , \6543 );
xnor \U$4560 ( \6545 , \6544 , \5593 );
and \U$4562 ( \6546 , \6106 , \5620 );
nor \U$4563 ( \6547 , 1'b0 , \6546 );
xnor \U$4564 ( \6548 , \6547 , 1'b0 );
xor \U$4565 ( \6549 , \6545 , \6548 );
xor \U$4567 ( \6550 , \6549 , 1'b0 );
xor \U$4568 ( \6551 , 1'b0 , \6550 );
and \U$4569 ( \6552 , \5863 , \5993 );
and \U$4570 ( \6553 , \5896 , \5991 );
nor \U$4571 ( \6554 , \6552 , \6553 );
xnor \U$4572 ( \6555 , \6554 , \6019 );
and \U$4573 ( \6556 , \5923 , \5694 );
and \U$4574 ( \6557 , \5956 , \5692 );
nor \U$4575 ( \6558 , \6556 , \6557 );
xnor \U$4576 ( \6559 , \6558 , \5699 );
xor \U$4577 ( \6560 , \6555 , \6559 );
and \U$4578 ( \6561 , \5985 , \5629 );
and \U$4579 ( \6562 , \6014 , \5627 );
nor \U$4580 ( \6563 , \6561 , \6562 );
xnor \U$4581 ( \6564 , \6563 , \5396 );
xor \U$4582 ( \6565 , \6560 , \6564 );
xor \U$4583 ( \6566 , \6551 , \6565 );
xor \U$4584 ( \6567 , \6541 , \6566 );
xor \U$4585 ( \6568 , \6532 , \6567 );
and \U$4586 ( \6569 , \6422 , \6490 );
nor \U$4587 ( \6570 , \6568 , \6569 );
and \U$4588 ( \6571 , \6536 , \6540 );
and \U$4589 ( \6572 , \6540 , \6566 );
and \U$4590 ( \6573 , \6536 , \6566 );
or \U$4591 ( \6574 , \6571 , \6572 , \6573 );
and \U$4592 ( \6575 , \6510 , \6530 );
xor \U$4593 ( \6576 , \6574 , \6575 );
and \U$4596 ( \6577 , \6514 , \6529 );
or \U$4597 ( \6578 , 1'b0 , 1'b0 , \6577 );
and \U$4599 ( \6579 , \6014 , \5629 );
and \U$4600 ( \6580 , \5923 , \5627 );
nor \U$4601 ( \6581 , \6579 , \6580 );
xnor \U$4602 ( \6582 , \6581 , \5396 );
and \U$4603 ( \6583 , \6061 , \5567 );
and \U$4604 ( \6584 , \5985 , \5565 );
nor \U$4605 ( \6585 , \6583 , \6584 );
xnor \U$4606 ( \6586 , \6585 , \5593 );
xor \U$4607 ( \6587 , \6582 , \6586 );
and \U$4609 ( \6588 , \6040 , \5620 );
nor \U$4610 ( \6589 , 1'b0 , \6588 );
xnor \U$4611 ( \6590 , \6589 , 1'b0 );
xor \U$4612 ( \6591 , \6587 , \6590 );
xor \U$4613 ( \6592 , 1'b0 , \6591 );
and \U$4614 ( \6593 , \5726 , \5935 );
and \U$4615 ( \6594 , \5747 , \5933 );
nor \U$4616 ( \6595 , \6593 , \6594 );
xnor \U$4617 ( \6596 , \6595 , \5961 );
and \U$4618 ( \6597 , \5896 , \5993 );
and \U$4619 ( \6598 , \5770 , \5991 );
nor \U$4620 ( \6599 , \6597 , \6598 );
xnor \U$4621 ( \6600 , \6599 , \6019 );
xor \U$4622 ( \6601 , \6596 , \6600 );
and \U$4623 ( \6602 , \5956 , \5694 );
and \U$4624 ( \6603 , \5863 , \5692 );
nor \U$4625 ( \6604 , \6602 , \6603 );
xnor \U$4626 ( \6605 , \6604 , \5699 );
xor \U$4627 ( \6606 , \6601 , \6605 );
xor \U$4628 ( \6607 , \6592 , \6606 );
and \U$4629 ( \6608 , \6519 , \6523 );
and \U$4630 ( \6609 , \6523 , \6528 );
and \U$4631 ( \6610 , \6519 , \6528 );
or \U$4632 ( \6611 , \6608 , \6609 , \6610 );
and \U$4633 ( \6612 , \6555 , \6559 );
and \U$4634 ( \6613 , \6559 , \6564 );
and \U$4635 ( \6614 , \6555 , \6564 );
or \U$4636 ( \6615 , \6612 , \6613 , \6614 );
xor \U$4637 ( \6616 , \6611 , \6615 );
and \U$4638 ( \6617 , \6545 , \6548 );
or \U$4641 ( \6618 , \6617 , 1'b0 , 1'b0 );
xor \U$4642 ( \6619 , \6616 , \6618 );
xor \U$4643 ( \6620 , \6607 , \6619 );
xor \U$4644 ( \6621 , \6578 , \6620 );
and \U$4645 ( \6622 , \6500 , \6504 );
and \U$4646 ( \6623 , \6504 , \6509 );
and \U$4647 ( \6624 , \6500 , \6509 );
or \U$4648 ( \6625 , \6622 , \6623 , \6624 );
and \U$4650 ( \6626 , \6550 , \6565 );
or \U$4652 ( \6627 , 1'b0 , \6626 , 1'b0 );
xor \U$4653 ( \6628 , \6625 , \6627 );
and \U$4655 ( \6629 , \5588 , \5839 );
not \U$4656 ( \6630 , \6629 );
xnor \U$4657 ( \6631 , \6630 , \5833 );
xor \U$4658 ( \6632 , 1'b0 , \6631 );
and \U$4659 ( \6633 , \5615 , \5875 );
and \U$4660 ( \6634 , \5519 , \5873 );
nor \U$4661 ( \6635 , \6633 , \6634 );
xnor \U$4662 ( \6636 , \6635 , \5901 );
xor \U$4663 ( \6637 , \6632 , \6636 );
xor \U$4664 ( \6638 , \6628 , \6637 );
xor \U$4665 ( \6639 , \6621 , \6638 );
xor \U$4666 ( \6640 , \6576 , \6639 );
and \U$4667 ( \6641 , \6498 , \6531 );
and \U$4668 ( \6642 , \6531 , \6567 );
and \U$4669 ( \6643 , \6498 , \6567 );
or \U$4670 ( \6644 , \6641 , \6642 , \6643 );
nor \U$4671 ( \6645 , \6640 , \6644 );
nor \U$4672 ( \6646 , \6570 , \6645 );
nand \U$4673 ( \6647 , \6494 , \6646 );
and \U$4674 ( \6648 , \6578 , \6620 );
and \U$4675 ( \6649 , \6620 , \6638 );
and \U$4676 ( \6650 , \6578 , \6638 );
or \U$4677 ( \6651 , \6648 , \6649 , \6650 );
and \U$4678 ( \6652 , \6611 , \6615 );
and \U$4679 ( \6653 , \6615 , \6618 );
and \U$4680 ( \6654 , \6611 , \6618 );
or \U$4681 ( \6655 , \6652 , \6653 , \6654 );
and \U$4683 ( \6656 , \6591 , \6606 );
or \U$4685 ( \6657 , 1'b0 , \6656 , 1'b0 );
xor \U$4686 ( \6658 , \6655 , \6657 );
and \U$4687 ( \6659 , \5770 , \5993 );
and \U$4688 ( \6660 , \5726 , \5991 );
nor \U$4689 ( \6661 , \6659 , \6660 );
xnor \U$4690 ( \6662 , \6661 , \6019 );
and \U$4691 ( \6663 , \5863 , \5694 );
and \U$4692 ( \6664 , \5896 , \5692 );
nor \U$4693 ( \6665 , \6663 , \6664 );
xnor \U$4694 ( \6666 , \6665 , \5699 );
xor \U$4695 ( \6667 , \6662 , \6666 );
and \U$4696 ( \6668 , \5923 , \5629 );
and \U$4697 ( \6669 , \5956 , \5627 );
nor \U$4698 ( \6670 , \6668 , \6669 );
xnor \U$4699 ( \6671 , \6670 , \5396 );
xor \U$4700 ( \6672 , \6667 , \6671 );
xor \U$4701 ( \6673 , \6658 , \6672 );
xor \U$4702 ( \6674 , \6651 , \6673 );
and \U$4703 ( \6675 , \6625 , \6627 );
and \U$4704 ( \6676 , \6627 , \6637 );
and \U$4705 ( \6677 , \6625 , \6637 );
or \U$4706 ( \6678 , \6675 , \6676 , \6677 );
and \U$4707 ( \6679 , \6607 , \6619 );
xor \U$4708 ( \6680 , \6678 , \6679 );
not \U$4709 ( \6681 , \5833 );
and \U$4710 ( \6682 , \5519 , \5875 );
and \U$4711 ( \6683 , \5588 , \5873 );
nor \U$4712 ( \6684 , \6682 , \6683 );
xnor \U$4713 ( \6685 , \6684 , \5901 );
xor \U$4714 ( \6686 , \6681 , \6685 );
and \U$4715 ( \6687 , \5747 , \5935 );
and \U$4716 ( \6688 , \5615 , \5933 );
nor \U$4717 ( \6689 , \6687 , \6688 );
xnor \U$4718 ( \6690 , \6689 , \5961 );
xor \U$4719 ( \6691 , \6686 , \6690 );
and \U$4721 ( \6692 , \5985 , \5567 );
and \U$4722 ( \6693 , \6014 , \5565 );
nor \U$4723 ( \6694 , \6692 , \6693 );
xnor \U$4724 ( \6695 , \6694 , \5593 );
and \U$4726 ( \6696 , \6061 , \5620 );
nor \U$4727 ( \6697 , 1'b0 , \6696 );
xnor \U$4728 ( \6698 , \6697 , 1'b0 );
xor \U$4729 ( \6699 , \6695 , \6698 );
xor \U$4731 ( \6700 , \6699 , 1'b0 );
xor \U$4732 ( \6701 , 1'b1 , \6700 );
xor \U$4733 ( \6702 , \6691 , \6701 );
and \U$4735 ( \6703 , \6631 , \6636 );
or \U$4737 ( \6704 , 1'b0 , \6703 , 1'b0 );
and \U$4738 ( \6705 , \6596 , \6600 );
and \U$4739 ( \6706 , \6600 , \6605 );
and \U$4740 ( \6707 , \6596 , \6605 );
or \U$4741 ( \6708 , \6705 , \6706 , \6707 );
xor \U$4742 ( \6709 , \6704 , \6708 );
and \U$4743 ( \6710 , \6582 , \6586 );
and \U$4744 ( \6711 , \6586 , \6590 );
and \U$4745 ( \6712 , \6582 , \6590 );
or \U$4746 ( \6713 , \6710 , \6711 , \6712 );
xor \U$4747 ( \6714 , \6709 , \6713 );
xor \U$4748 ( \6715 , \6702 , \6714 );
xor \U$4749 ( \6716 , \6680 , \6715 );
xor \U$4750 ( \6717 , \6674 , \6716 );
and \U$4751 ( \6718 , \6574 , \6575 );
and \U$4752 ( \6719 , \6575 , \6639 );
and \U$4753 ( \6720 , \6574 , \6639 );
or \U$4754 ( \6721 , \6718 , \6719 , \6720 );
nor \U$4755 ( \6722 , \6717 , \6721 );
and \U$4756 ( \6723 , \6678 , \6679 );
and \U$4757 ( \6724 , \6679 , \6715 );
and \U$4758 ( \6725 , \6678 , \6715 );
or \U$4759 ( \6726 , \6723 , \6724 , \6725 );
and \U$4760 ( \6727 , \6681 , \6685 );
and \U$4761 ( \6728 , \6685 , \6690 );
and \U$4762 ( \6729 , \6681 , \6690 );
or \U$4763 ( \6730 , \6727 , \6728 , \6729 );
and \U$4764 ( \6731 , \6662 , \6666 );
and \U$4765 ( \6732 , \6666 , \6671 );
and \U$4766 ( \6733 , \6662 , \6671 );
or \U$4767 ( \6734 , \6731 , \6732 , \6733 );
xor \U$4768 ( \6735 , \6730 , \6734 );
and \U$4769 ( \6736 , \6695 , \6698 );
or \U$4772 ( \6737 , \6736 , 1'b0 , 1'b0 );
xor \U$4773 ( \6738 , \6735 , \6737 );
and \U$4774 ( \6739 , \6704 , \6708 );
and \U$4775 ( \6740 , \6708 , \6713 );
and \U$4776 ( \6741 , \6704 , \6713 );
or \U$4777 ( \6742 , \6739 , \6740 , \6741 );
and \U$4780 ( \6743 , 1'b1 , \6700 );
or \U$4782 ( \6744 , 1'b0 , \6743 , 1'b0 );
xor \U$4783 ( \6745 , \6742 , \6744 );
and \U$4784 ( \6746 , \6014 , \5567 );
and \U$4785 ( \6747 , \5923 , \5565 );
nor \U$4786 ( \6748 , \6746 , \6747 );
xnor \U$4787 ( \6749 , \6748 , \5593 );
and \U$4789 ( \6750 , \5985 , \5620 );
nor \U$4790 ( \6751 , 1'b0 , \6750 );
xnor \U$4791 ( \6752 , \6751 , 1'b0 );
xor \U$4792 ( \6753 , \6749 , \6752 );
xor \U$4794 ( \6754 , \6753 , 1'b0 );
and \U$4795 ( \6755 , \5726 , \5993 );
and \U$4796 ( \6756 , \5747 , \5991 );
nor \U$4797 ( \6757 , \6755 , \6756 );
xnor \U$4798 ( \6758 , \6757 , \6019 );
and \U$4799 ( \6759 , \5896 , \5694 );
and \U$4800 ( \6760 , \5770 , \5692 );
nor \U$4801 ( \6761 , \6759 , \6760 );
xnor \U$4802 ( \6762 , \6761 , \5699 );
xor \U$4803 ( \6763 , \6758 , \6762 );
and \U$4804 ( \6764 , \5956 , \5629 );
and \U$4805 ( \6765 , \5863 , \5627 );
nor \U$4806 ( \6766 , \6764 , \6765 );
xnor \U$4807 ( \6767 , \6766 , \5396 );
xor \U$4808 ( \6768 , \6763 , \6767 );
xor \U$4809 ( \6769 , \6754 , \6768 );
and \U$4811 ( \6770 , \5588 , \5875 );
not \U$4812 ( \6771 , \6770 );
xnor \U$4813 ( \6772 , \6771 , \5901 );
xor \U$4814 ( \6773 , 1'b0 , \6772 );
and \U$4815 ( \6774 , \5615 , \5935 );
and \U$4816 ( \6775 , \5519 , \5933 );
nor \U$4817 ( \6776 , \6774 , \6775 );
xnor \U$4818 ( \6777 , \6776 , \5961 );
xor \U$4819 ( \6778 , \6773 , \6777 );
xor \U$4820 ( \6779 , \6769 , \6778 );
xor \U$4821 ( \6780 , \6745 , \6779 );
xor \U$4822 ( \6781 , \6738 , \6780 );
xor \U$4823 ( \6782 , \6726 , \6781 );
and \U$4824 ( \6783 , \6655 , \6657 );
and \U$4825 ( \6784 , \6657 , \6672 );
and \U$4826 ( \6785 , \6655 , \6672 );
or \U$4827 ( \6786 , \6783 , \6784 , \6785 );
and \U$4828 ( \6787 , \6691 , \6701 );
and \U$4829 ( \6788 , \6701 , \6714 );
and \U$4830 ( \6789 , \6691 , \6714 );
or \U$4831 ( \6790 , \6787 , \6788 , \6789 );
xor \U$4832 ( \6791 , \6786 , \6790 );
xor \U$4834 ( \6792 , \6791 , 1'b1 );
xor \U$4835 ( \6793 , \6782 , \6792 );
and \U$4836 ( \6794 , \6651 , \6673 );
and \U$4837 ( \6795 , \6673 , \6716 );
and \U$4838 ( \6796 , \6651 , \6716 );
or \U$4839 ( \6797 , \6794 , \6795 , \6796 );
nor \U$4840 ( \6798 , \6793 , \6797 );
nor \U$4841 ( \6799 , \6722 , \6798 );
and \U$4842 ( \6800 , \6786 , \6790 );
and \U$4843 ( \6801 , \6790 , 1'b1 );
and \U$4844 ( \6802 , \6786 , 1'b1 );
or \U$4845 ( \6803 , \6800 , \6801 , \6802 );
and \U$4846 ( \6804 , \6738 , \6780 );
xor \U$4847 ( \6805 , \6803 , \6804 );
and \U$4848 ( \6806 , \6742 , \6744 );
and \U$4849 ( \6807 , \6744 , \6779 );
and \U$4850 ( \6808 , \6742 , \6779 );
or \U$4851 ( \6809 , \6806 , \6807 , \6808 );
and \U$4853 ( \6810 , \6014 , \5620 );
nor \U$4854 ( \6811 , 1'b0 , \6810 );
xnor \U$4855 ( \6812 , \6811 , 1'b0 );
xor \U$4857 ( \6813 , \6812 , 1'b0 );
xor \U$4859 ( \6814 , \6813 , 1'b0 );
and \U$4860 ( \6815 , \5770 , \5694 );
and \U$4861 ( \6816 , \5726 , \5692 );
nor \U$4862 ( \6817 , \6815 , \6816 );
xnor \U$4863 ( \6818 , \6817 , \5699 );
and \U$4864 ( \6819 , \5863 , \5629 );
and \U$4865 ( \6820 , \5896 , \5627 );
nor \U$4866 ( \6821 , \6819 , \6820 );
xnor \U$4867 ( \6822 , \6821 , \5396 );
xor \U$4868 ( \6823 , \6818 , \6822 );
and \U$4869 ( \6824 , \5923 , \5567 );
and \U$4870 ( \6825 , \5956 , \5565 );
nor \U$4871 ( \6826 , \6824 , \6825 );
xnor \U$4872 ( \6827 , \6826 , \5593 );
xor \U$4873 ( \6828 , \6823 , \6827 );
xor \U$4874 ( \6829 , \6814 , \6828 );
not \U$4875 ( \6830 , \5901 );
and \U$4876 ( \6831 , \5519 , \5935 );
and \U$4877 ( \6832 , \5588 , \5933 );
nor \U$4878 ( \6833 , \6831 , \6832 );
xnor \U$4879 ( \6834 , \6833 , \5961 );
xor \U$4880 ( \6835 , \6830 , \6834 );
and \U$4881 ( \6836 , \5747 , \5993 );
and \U$4882 ( \6837 , \5615 , \5991 );
nor \U$4883 ( \6838 , \6836 , \6837 );
xnor \U$4884 ( \6839 , \6838 , \6019 );
xor \U$4885 ( \6840 , \6835 , \6839 );
xor \U$4886 ( \6841 , \6829 , \6840 );
xor \U$4888 ( \6842 , \6841 , 1'b0 );
and \U$4890 ( \6843 , \6772 , \6777 );
or \U$4892 ( \6844 , 1'b0 , \6843 , 1'b0 );
and \U$4893 ( \6845 , \6758 , \6762 );
and \U$4894 ( \6846 , \6762 , \6767 );
and \U$4895 ( \6847 , \6758 , \6767 );
or \U$4896 ( \6848 , \6845 , \6846 , \6847 );
xor \U$4897 ( \6849 , \6844 , \6848 );
and \U$4898 ( \6850 , \6749 , \6752 );
or \U$4901 ( \6851 , \6850 , 1'b0 , 1'b0 );
xor \U$4902 ( \6852 , \6849 , \6851 );
xor \U$4903 ( \6853 , \6842 , \6852 );
xor \U$4904 ( \6854 , \6809 , \6853 );
and \U$4905 ( \6855 , \6730 , \6734 );
and \U$4906 ( \6856 , \6734 , \6737 );
and \U$4907 ( \6857 , \6730 , \6737 );
or \U$4908 ( \6858 , \6855 , \6856 , \6857 );
xor \U$4910 ( \6859 , \6858 , 1'b0 );
and \U$4911 ( \6860 , \6754 , \6768 );
and \U$4912 ( \6861 , \6768 , \6778 );
and \U$4913 ( \6862 , \6754 , \6778 );
or \U$4914 ( \6863 , \6860 , \6861 , \6862 );
xor \U$4915 ( \6864 , \6859 , \6863 );
xor \U$4916 ( \6865 , \6854 , \6864 );
xor \U$4917 ( \6866 , \6805 , \6865 );
and \U$4918 ( \6867 , \6726 , \6781 );
and \U$4919 ( \6868 , \6781 , \6792 );
and \U$4920 ( \6869 , \6726 , \6792 );
or \U$4921 ( \6870 , \6867 , \6868 , \6869 );
nor \U$4922 ( \6871 , \6866 , \6870 );
and \U$4923 ( \6872 , \6809 , \6853 );
and \U$4924 ( \6873 , \6853 , \6864 );
and \U$4925 ( \6874 , \6809 , \6864 );
or \U$4926 ( \6875 , \6872 , \6873 , \6874 );
and \U$4927 ( \6876 , \6844 , \6848 );
and \U$4928 ( \6877 , \6848 , \6851 );
and \U$4929 ( \6878 , \6844 , \6851 );
or \U$4930 ( \6879 , \6876 , \6877 , \6878 );
xor \U$4932 ( \6880 , \6879 , 1'b0 );
and \U$4933 ( \6881 , \6814 , \6828 );
and \U$4934 ( \6882 , \6828 , \6840 );
and \U$4935 ( \6883 , \6814 , \6840 );
or \U$4936 ( \6884 , \6881 , \6882 , \6883 );
xor \U$4937 ( \6885 , \6880 , \6884 );
xor \U$4938 ( \6886 , \6875 , \6885 );
and \U$4941 ( \6887 , \6858 , \6863 );
or \U$4942 ( \6888 , 1'b0 , 1'b0 , \6887 );
and \U$4945 ( \6889 , \6841 , \6852 );
or \U$4946 ( \6890 , 1'b0 , 1'b0 , \6889 );
xor \U$4947 ( \6891 , \6888 , \6890 );
and \U$4948 ( \6892 , \5726 , \5694 );
and \U$4949 ( \6893 , \5747 , \5692 );
nor \U$4950 ( \6894 , \6892 , \6893 );
xnor \U$4951 ( \6895 , \6894 , \5699 );
and \U$4952 ( \6896 , \5896 , \5629 );
and \U$4953 ( \6897 , \5770 , \5627 );
nor \U$4954 ( \6898 , \6896 , \6897 );
xnor \U$4955 ( \6899 , \6898 , \5396 );
xor \U$4956 ( \6900 , \6895 , \6899 );
and \U$4957 ( \6901 , \5956 , \5567 );
and \U$4958 ( \6902 , \5863 , \5565 );
nor \U$4959 ( \6903 , \6901 , \6902 );
xnor \U$4960 ( \6904 , \6903 , \5593 );
xor \U$4961 ( \6905 , \6900 , \6904 );
and \U$4963 ( \6906 , \5588 , \5935 );
not \U$4964 ( \6907 , \6906 );
xnor \U$4965 ( \6908 , \6907 , \5961 );
xor \U$4966 ( \6909 , 1'b0 , \6908 );
and \U$4967 ( \6910 , \5615 , \5993 );
and \U$4968 ( \6911 , \5519 , \5991 );
nor \U$4969 ( \6912 , \6910 , \6911 );
xnor \U$4970 ( \6913 , \6912 , \6019 );
xor \U$4971 ( \6914 , \6909 , \6913 );
xor \U$4972 ( \6915 , \6905 , \6914 );
and \U$4975 ( \6916 , \5923 , \5620 );
nor \U$4976 ( \6917 , 1'b0 , \6916 );
xnor \U$4977 ( \6918 , \6917 , 1'b0 );
xor \U$4979 ( \6919 , \6918 , 1'b0 );
xor \U$4981 ( \6920 , \6919 , 1'b0 );
xnor \U$4982 ( \6921 , 1'b0 , \6920 );
xor \U$4983 ( \6922 , \6915 , \6921 );
and \U$4984 ( \6923 , \6830 , \6834 );
and \U$4985 ( \6924 , \6834 , \6839 );
and \U$4986 ( \6925 , \6830 , \6839 );
or \U$4987 ( \6926 , \6923 , \6924 , \6925 );
and \U$4988 ( \6927 , \6818 , \6822 );
and \U$4989 ( \6928 , \6822 , \6827 );
and \U$4990 ( \6929 , \6818 , \6827 );
or \U$4991 ( \6930 , \6927 , \6928 , \6929 );
xor \U$4992 ( \6931 , \6926 , \6930 );
xor \U$4994 ( \6932 , \6931 , 1'b0 );
xor \U$4995 ( \6933 , \6922 , \6932 );
xor \U$4996 ( \6934 , \6891 , \6933 );
xor \U$4997 ( \6935 , \6886 , \6934 );
and \U$4998 ( \6936 , \6803 , \6804 );
and \U$4999 ( \6937 , \6804 , \6865 );
and \U$5000 ( \6938 , \6803 , \6865 );
or \U$5001 ( \6939 , \6936 , \6937 , \6938 );
nor \U$5002 ( \6940 , \6935 , \6939 );
nor \U$5003 ( \6941 , \6871 , \6940 );
nand \U$5004 ( \6942 , \6799 , \6941 );
nor \U$5005 ( \6943 , \6647 , \6942 );
and \U$5006 ( \6944 , \6888 , \6890 );
and \U$5007 ( \6945 , \6890 , \6933 );
and \U$5008 ( \6946 , \6888 , \6933 );
or \U$5009 ( \6947 , \6944 , \6945 , \6946 );
and \U$5010 ( \6948 , \6926 , \6930 );
or \U$5013 ( \6949 , \6948 , 1'b0 , 1'b0 );
or \U$5014 ( \6950 , 1'b0 , \6920 );
xor \U$5015 ( \6951 , \6949 , \6950 );
and \U$5016 ( \6952 , \6905 , \6914 );
xor \U$5017 ( \6953 , \6951 , \6952 );
xor \U$5018 ( \6954 , \6947 , \6953 );
and \U$5021 ( \6955 , \6879 , \6884 );
or \U$5022 ( \6956 , 1'b0 , 1'b0 , \6955 );
and \U$5023 ( \6957 , \6915 , \6921 );
and \U$5024 ( \6958 , \6921 , \6932 );
and \U$5025 ( \6959 , \6915 , \6932 );
or \U$5026 ( \6960 , \6957 , \6958 , \6959 );
xor \U$5027 ( \6961 , \6956 , \6960 );
and \U$5029 ( \6962 , \5770 , \5629 );
and \U$5030 ( \6963 , \5726 , \5627 );
nor \U$5031 ( \6964 , \6962 , \6963 );
xnor \U$5032 ( \6965 , \6964 , \5396 );
and \U$5033 ( \6966 , \5863 , \5567 );
and \U$5034 ( \6967 , \5896 , \5565 );
nor \U$5035 ( \6968 , \6966 , \6967 );
xnor \U$5036 ( \6969 , \6968 , \5593 );
xor \U$5037 ( \6970 , \6965 , \6969 );
and \U$5039 ( \6971 , \5956 , \5620 );
nor \U$5040 ( \6972 , 1'b0 , \6971 );
xnor \U$5041 ( \6973 , \6972 , 1'b0 );
xor \U$5042 ( \6974 , \6970 , \6973 );
xor \U$5043 ( \6975 , 1'b0 , \6974 );
not \U$5044 ( \6976 , \5961 );
and \U$5045 ( \6977 , \5519 , \5993 );
and \U$5046 ( \6978 , \5588 , \5991 );
nor \U$5047 ( \6979 , \6977 , \6978 );
xnor \U$5048 ( \6980 , \6979 , \6019 );
xor \U$5049 ( \6981 , \6976 , \6980 );
and \U$5050 ( \6982 , \5747 , \5694 );
and \U$5051 ( \6983 , \5615 , \5692 );
nor \U$5052 ( \6984 , \6982 , \6983 );
xnor \U$5053 ( \6985 , \6984 , \5699 );
xor \U$5054 ( \6986 , \6981 , \6985 );
xor \U$5055 ( \6987 , \6975 , \6986 );
xor \U$5057 ( \6988 , \6987 , 1'b0 );
and \U$5059 ( \6989 , \6908 , \6913 );
or \U$5061 ( \6990 , 1'b0 , \6989 , 1'b0 );
and \U$5062 ( \6991 , \6895 , \6899 );
and \U$5063 ( \6992 , \6899 , \6904 );
and \U$5064 ( \6993 , \6895 , \6904 );
or \U$5065 ( \6994 , \6991 , \6992 , \6993 );
xor \U$5066 ( \6995 , \6990 , \6994 );
xor \U$5068 ( \6996 , \6995 , 1'b0 );
xor \U$5069 ( \6997 , \6988 , \6996 );
xor \U$5070 ( \6998 , \6961 , \6997 );
xor \U$5071 ( \6999 , \6954 , \6998 );
and \U$5072 ( \7000 , \6875 , \6885 );
and \U$5073 ( \7001 , \6885 , \6934 );
and \U$5074 ( \7002 , \6875 , \6934 );
or \U$5075 ( \7003 , \7000 , \7001 , \7002 );
nor \U$5076 ( \7004 , \6999 , \7003 );
and \U$5077 ( \7005 , \6956 , \6960 );
and \U$5078 ( \7006 , \6960 , \6997 );
and \U$5079 ( \7007 , \6956 , \6997 );
or \U$5080 ( \7008 , \7005 , \7006 , \7007 );
and \U$5081 ( \7009 , \6990 , \6994 );
or \U$5084 ( \7010 , \7009 , 1'b0 , 1'b0 );
xor \U$5086 ( \7011 , \7010 , 1'b0 );
and \U$5088 ( \7012 , \6974 , \6986 );
or \U$5090 ( \7013 , 1'b0 , \7012 , 1'b0 );
xor \U$5091 ( \7014 , \7011 , \7013 );
xor \U$5092 ( \7015 , \7008 , \7014 );
and \U$5093 ( \7016 , \6949 , \6950 );
and \U$5094 ( \7017 , \6950 , \6952 );
and \U$5095 ( \7018 , \6949 , \6952 );
or \U$5096 ( \7019 , \7016 , \7017 , \7018 );
and \U$5099 ( \7020 , \6987 , \6996 );
or \U$5100 ( \7021 , 1'b0 , 1'b0 , \7020 );
xor \U$5101 ( \7022 , \7019 , \7021 );
and \U$5102 ( \7023 , \5726 , \5629 );
and \U$5103 ( \7024 , \5747 , \5627 );
nor \U$5104 ( \7025 , \7023 , \7024 );
xnor \U$5105 ( \7026 , \7025 , \5396 );
and \U$5106 ( \7027 , \5896 , \5567 );
and \U$5107 ( \7028 , \5770 , \5565 );
nor \U$5108 ( \7029 , \7027 , \7028 );
xnor \U$5109 ( \7030 , \7029 , \5593 );
xor \U$5110 ( \7031 , \7026 , \7030 );
and \U$5112 ( \7032 , \5863 , \5620 );
nor \U$5113 ( \7033 , 1'b0 , \7032 );
xnor \U$5114 ( \7034 , \7033 , 1'b0 );
xor \U$5115 ( \7035 , \7031 , \7034 );
and \U$5117 ( \7036 , \5588 , \5993 );
not \U$5118 ( \7037 , \7036 );
xnor \U$5119 ( \7038 , \7037 , \6019 );
xor \U$5120 ( \7039 , 1'b0 , \7038 );
and \U$5121 ( \7040 , \5615 , \5694 );
and \U$5122 ( \7041 , \5519 , \5692 );
nor \U$5123 ( \7042 , \7040 , \7041 );
xnor \U$5124 ( \7043 , \7042 , \5699 );
xor \U$5125 ( \7044 , \7039 , \7043 );
xor \U$5126 ( \7045 , \7035 , \7044 );
xor \U$5128 ( \7046 , \7045 , 1'b1 );
and \U$5129 ( \7047 , \6976 , \6980 );
and \U$5130 ( \7048 , \6980 , \6985 );
and \U$5131 ( \7049 , \6976 , \6985 );
or \U$5132 ( \7050 , \7047 , \7048 , \7049 );
and \U$5133 ( \7051 , \6965 , \6969 );
and \U$5134 ( \7052 , \6969 , \6973 );
and \U$5135 ( \7053 , \6965 , \6973 );
or \U$5136 ( \7054 , \7051 , \7052 , \7053 );
xor \U$5137 ( \7055 , \7050 , \7054 );
xor \U$5139 ( \7056 , \7055 , 1'b0 );
xor \U$5140 ( \7057 , \7046 , \7056 );
xor \U$5141 ( \7058 , \7022 , \7057 );
xor \U$5142 ( \7059 , \7015 , \7058 );
and \U$5143 ( \7060 , \6947 , \6953 );
and \U$5144 ( \7061 , \6953 , \6998 );
and \U$5145 ( \7062 , \6947 , \6998 );
or \U$5146 ( \7063 , \7060 , \7061 , \7062 );
nor \U$5147 ( \7064 , \7059 , \7063 );
nor \U$5148 ( \7065 , \7004 , \7064 );
and \U$5149 ( \7066 , \7019 , \7021 );
and \U$5150 ( \7067 , \7021 , \7057 );
and \U$5151 ( \7068 , \7019 , \7057 );
or \U$5152 ( \7069 , \7066 , \7067 , \7068 );
and \U$5153 ( \7070 , \7050 , \7054 );
or \U$5156 ( \7071 , \7070 , 1'b0 , 1'b0 );
xor \U$5158 ( \7072 , \7071 , 1'b0 );
and \U$5159 ( \7073 , \7035 , \7044 );
xor \U$5160 ( \7074 , \7072 , \7073 );
xor \U$5161 ( \7075 , \7069 , \7074 );
and \U$5164 ( \7076 , \7010 , \7013 );
or \U$5165 ( \7077 , 1'b0 , 1'b0 , \7076 );
and \U$5166 ( \7078 , \7045 , 1'b1 );
and \U$5167 ( \7079 , 1'b1 , \7056 );
and \U$5168 ( \7080 , \7045 , \7056 );
or \U$5169 ( \7081 , \7078 , \7079 , \7080 );
xor \U$5170 ( \7082 , \7077 , \7081 );
and \U$5172 ( \7083 , \5770 , \5567 );
and \U$5173 ( \7084 , \5726 , \5565 );
nor \U$5174 ( \7085 , \7083 , \7084 );
xnor \U$5175 ( \7086 , \7085 , \5593 );
and \U$5177 ( \7087 , \5896 , \5620 );
nor \U$5178 ( \7088 , 1'b0 , \7087 );
xnor \U$5179 ( \7089 , \7088 , 1'b0 );
xor \U$5180 ( \7090 , \7086 , \7089 );
xor \U$5182 ( \7091 , \7090 , 1'b0 );
xor \U$5183 ( \7092 , 1'b0 , \7091 );
not \U$5184 ( \7093 , \6019 );
and \U$5185 ( \7094 , \5519 , \5694 );
and \U$5186 ( \7095 , \5588 , \5692 );
nor \U$5187 ( \7096 , \7094 , \7095 );
xnor \U$5188 ( \7097 , \7096 , \5699 );
xor \U$5189 ( \7098 , \7093 , \7097 );
and \U$5190 ( \7099 , \5747 , \5629 );
and \U$5191 ( \7100 , \5615 , \5627 );
nor \U$5192 ( \7101 , \7099 , \7100 );
xnor \U$5193 ( \7102 , \7101 , \5396 );
xor \U$5194 ( \7103 , \7098 , \7102 );
xor \U$5195 ( \7104 , \7092 , \7103 );
xor \U$5197 ( \7105 , \7104 , 1'b0 );
and \U$5199 ( \7106 , \7038 , \7043 );
or \U$5201 ( \7107 , 1'b0 , \7106 , 1'b0 );
and \U$5202 ( \7108 , \7026 , \7030 );
and \U$5203 ( \7109 , \7030 , \7034 );
and \U$5204 ( \7110 , \7026 , \7034 );
or \U$5205 ( \7111 , \7108 , \7109 , \7110 );
xor \U$5206 ( \7112 , \7107 , \7111 );
xor \U$5208 ( \7113 , \7112 , 1'b0 );
xor \U$5209 ( \7114 , \7105 , \7113 );
xor \U$5210 ( \7115 , \7082 , \7114 );
xor \U$5211 ( \7116 , \7075 , \7115 );
and \U$5212 ( \7117 , \7008 , \7014 );
and \U$5213 ( \7118 , \7014 , \7058 );
and \U$5214 ( \7119 , \7008 , \7058 );
or \U$5215 ( \7120 , \7117 , \7118 , \7119 );
nor \U$5216 ( \7121 , \7116 , \7120 );
and \U$5217 ( \7122 , \7077 , \7081 );
and \U$5218 ( \7123 , \7081 , \7114 );
and \U$5219 ( \7124 , \7077 , \7114 );
or \U$5220 ( \7125 , \7122 , \7123 , \7124 );
and \U$5221 ( \7126 , \7107 , \7111 );
or \U$5224 ( \7127 , \7126 , 1'b0 , 1'b0 );
xor \U$5226 ( \7128 , \7127 , 1'b0 );
and \U$5228 ( \7129 , \7091 , \7103 );
or \U$5230 ( \7130 , 1'b0 , \7129 , 1'b0 );
xor \U$5231 ( \7131 , \7128 , \7130 );
xor \U$5232 ( \7132 , \7125 , \7131 );
and \U$5235 ( \7133 , \7071 , \7073 );
or \U$5236 ( \7134 , 1'b0 , 1'b0 , \7133 );
and \U$5239 ( \7135 , \7104 , \7113 );
or \U$5240 ( \7136 , 1'b0 , 1'b0 , \7135 );
xor \U$5241 ( \7137 , \7134 , \7136 );
xor \U$5242 ( \7138 , \5750 , \5773 );
xor \U$5244 ( \7139 , \7138 , 1'b0 );
xor \U$5246 ( \7140 , 1'b0 , \5700 );
xor \U$5247 ( \7141 , \7140 , \5704 );
xor \U$5248 ( \7142 , \7139 , \7141 );
xor \U$5250 ( \7143 , \7142 , 1'b1 );
and \U$5251 ( \7144 , \7093 , \7097 );
and \U$5252 ( \7145 , \7097 , \7102 );
and \U$5253 ( \7146 , \7093 , \7102 );
or \U$5254 ( \7147 , \7144 , \7145 , \7146 );
and \U$5255 ( \7148 , \7086 , \7089 );
or \U$5258 ( \7149 , \7148 , 1'b0 , 1'b0 );
xor \U$5259 ( \7150 , \7147 , \7149 );
xor \U$5261 ( \7151 , \7150 , 1'b0 );
xor \U$5262 ( \7152 , \7143 , \7151 );
xor \U$5263 ( \7153 , \7137 , \7152 );
xor \U$5264 ( \7154 , \7132 , \7153 );
and \U$5265 ( \7155 , \7069 , \7074 );
and \U$5266 ( \7156 , \7074 , \7115 );
and \U$5267 ( \7157 , \7069 , \7115 );
or \U$5268 ( \7158 , \7155 , \7156 , \7157 );
nor \U$5269 ( \7159 , \7154 , \7158 );
nor \U$5270 ( \7160 , \7121 , \7159 );
nand \U$5271 ( \7161 , \7065 , \7160 );
and \U$5272 ( \7162 , \7134 , \7136 );
and \U$5273 ( \7163 , \7136 , \7152 );
and \U$5274 ( \7164 , \7134 , \7152 );
or \U$5275 ( \7165 , \7162 , \7163 , \7164 );
and \U$5276 ( \7166 , \7147 , \7149 );
or \U$5279 ( \7167 , \7166 , 1'b0 , 1'b0 );
xor \U$5281 ( \7168 , \7167 , 1'b0 );
and \U$5282 ( \7169 , \7139 , \7141 );
xor \U$5283 ( \7170 , \7168 , \7169 );
xor \U$5284 ( \7171 , \7165 , \7170 );
and \U$5287 ( \7172 , \7127 , \7130 );
or \U$5288 ( \7173 , 1'b0 , 1'b0 , \7172 );
and \U$5289 ( \7174 , \7142 , 1'b1 );
and \U$5290 ( \7175 , 1'b1 , \7151 );
and \U$5291 ( \7176 , \7142 , \7151 );
or \U$5292 ( \7177 , \7174 , \7175 , \7176 );
xor \U$5293 ( \7178 , \7173 , \7177 );
xor \U$5295 ( \7179 , 1'b0 , \5782 );
xor \U$5296 ( \7180 , \7179 , \5793 );
xor \U$5298 ( \7181 , \7180 , 1'b0 );
xor \U$5299 ( \7182 , \5706 , \5775 );
xor \U$5301 ( \7183 , \7182 , 1'b0 );
xor \U$5302 ( \7184 , \7181 , \7183 );
xor \U$5303 ( \7185 , \7178 , \7184 );
xor \U$5304 ( \7186 , \7171 , \7185 );
and \U$5305 ( \7187 , \7125 , \7131 );
and \U$5306 ( \7188 , \7131 , \7153 );
and \U$5307 ( \7189 , \7125 , \7153 );
or \U$5308 ( \7190 , \7187 , \7188 , \7189 );
nor \U$5309 ( \7191 , \7186 , \7190 );
and \U$5310 ( \7192 , \7173 , \7177 );
and \U$5311 ( \7193 , \7177 , \7184 );
and \U$5312 ( \7194 , \7173 , \7184 );
or \U$5313 ( \7195 , \7192 , \7193 , \7194 );
xor \U$5315 ( \7196 , \5777 , 1'b0 );
xor \U$5316 ( \7197 , \7196 , \5795 );
xor \U$5317 ( \7198 , \7195 , \7197 );
and \U$5320 ( \7199 , \7167 , \7169 );
or \U$5321 ( \7200 , 1'b0 , 1'b0 , \7199 );
and \U$5324 ( \7201 , \7180 , \7183 );
or \U$5325 ( \7202 , 1'b0 , 1'b0 , \7201 );
xor \U$5326 ( \7203 , \7200 , \7202 );
xor \U$5327 ( \7204 , \5805 , 1'b1 );
xor \U$5328 ( \7205 , \7204 , \5812 );
xor \U$5329 ( \7206 , \7203 , \7205 );
xor \U$5330 ( \7207 , \7198 , \7206 );
and \U$5331 ( \7208 , \7165 , \7170 );
and \U$5332 ( \7209 , \7170 , \7185 );
and \U$5333 ( \7210 , \7165 , \7185 );
or \U$5334 ( \7211 , \7208 , \7209 , \7210 );
nor \U$5335 ( \7212 , \7207 , \7211 );
nor \U$5336 ( \7213 , \7191 , \7212 );
and \U$5337 ( \7214 , \7200 , \7202 );
and \U$5338 ( \7215 , \7202 , \7205 );
and \U$5339 ( \7216 , \7200 , \7205 );
or \U$5340 ( \7217 , \7214 , \7215 , \7216 );
and \U$5342 ( \7218 , \5802 , \5804 );
xor \U$5343 ( \7219 , 1'b0 , \7218 );
xor \U$5344 ( \7220 , \7217 , \7219 );
xor \U$5345 ( \7221 , \5797 , \5815 );
xor \U$5346 ( \7222 , \7221 , \5818 );
xor \U$5347 ( \7223 , \7220 , \7222 );
and \U$5348 ( \7224 , \7195 , \7197 );
and \U$5349 ( \7225 , \7197 , \7206 );
and \U$5350 ( \7226 , \7195 , \7206 );
or \U$5351 ( \7227 , \7224 , \7225 , \7226 );
nor \U$5352 ( \7228 , \7223 , \7227 );
xor \U$5354 ( \7229 , \5821 , 1'b0 );
xor \U$5355 ( \7230 , \7229 , \5823 );
and \U$5356 ( \7231 , \7217 , \7219 );
and \U$5357 ( \7232 , \7219 , \7222 );
and \U$5358 ( \7233 , \7217 , \7222 );
or \U$5359 ( \7234 , \7231 , \7232 , \7233 );
nor \U$5360 ( \7235 , \7230 , \7234 );
nor \U$5361 ( \7236 , \7228 , \7235 );
nand \U$5362 ( \7237 , \7213 , \7236 );
nor \U$5363 ( \7238 , \7161 , \7237 );
nand \U$5364 ( \7239 , \6943 , \7238 );
and \U$5365 ( \7240 , \6040 , \5839 );
and \U$5366 ( \7241 , \6061 , \5836 );
nor \U$5367 ( \7242 , \7240 , \7241 );
xnor \U$5368 ( \7243 , \7242 , \5833 );
and \U$5369 ( \7244 , \6085 , \5875 );
and \U$5370 ( \7245 , \6106 , \5873 );
nor \U$5371 ( \7246 , \7244 , \7245 );
xnor \U$5372 ( \7247 , \7246 , \5901 );
and \U$5373 ( \7248 , \7243 , \7247 );
and \U$5374 ( \7249 , \6133 , \5935 );
and \U$5375 ( \7250 , \6154 , \5933 );
nor \U$5376 ( \7251 , \7249 , \7250 );
xnor \U$5377 ( \7252 , \7251 , \5961 );
and \U$5378 ( \7253 , \7247 , \7252 );
and \U$5379 ( \7254 , \7243 , \7252 );
or \U$5380 ( \7255 , \7248 , \7253 , \7254 );
and \U$5381 ( \7256 , \6154 , \5935 );
and \U$5382 ( \7257 , \6085 , \5933 );
nor \U$5383 ( \7258 , \7256 , \7257 );
xnor \U$5384 ( \7259 , \7258 , \5961 );
and \U$5385 ( \7260 , \6177 , \5993 );
and \U$5386 ( \7261 , \6133 , \5991 );
nor \U$5387 ( \7262 , \7260 , \7261 );
xnor \U$5388 ( \7263 , \7262 , \6019 );
xor \U$5389 ( \7264 , \7259 , \7263 );
nand \U$5390 ( \7265 , \6310 , \5692 );
xnor \U$5391 ( \7266 , \7265 , \5699 );
xor \U$5392 ( \7267 , \7264 , \7266 );
and \U$5393 ( \7268 , \7255 , \7267 );
and \U$5394 ( \7269 , \6061 , \5839 );
and \U$5395 ( \7270 , \5985 , \5836 );
nor \U$5396 ( \7271 , \7269 , \7270 );
xnor \U$5397 ( \7272 , \7271 , \5833 );
xor \U$5398 ( \7273 , \5699 , \7272 );
and \U$5399 ( \7274 , \6106 , \5875 );
and \U$5400 ( \7275 , \6040 , \5873 );
nor \U$5401 ( \7276 , \7274 , \7275 );
xnor \U$5402 ( \7277 , \7276 , \5901 );
xor \U$5403 ( \7278 , \7273 , \7277 );
and \U$5404 ( \7279 , \7267 , \7278 );
and \U$5405 ( \7280 , \7255 , \7278 );
or \U$5406 ( \7281 , \7268 , \7279 , \7280 );
and \U$5407 ( \7282 , \6310 , \5694 );
and \U$5408 ( \7283 , \6177 , \5692 );
nor \U$5409 ( \7284 , \7282 , \7283 );
xnor \U$5410 ( \7285 , \7284 , \5699 );
and \U$5411 ( \7286 , \5985 , \5839 );
and \U$5412 ( \7287 , \6014 , \5836 );
nor \U$5413 ( \7288 , \7286 , \7287 );
xnor \U$5414 ( \7289 , \7288 , \5833 );
and \U$5415 ( \7290 , \6040 , \5875 );
and \U$5416 ( \7291 , \6061 , \5873 );
nor \U$5417 ( \7292 , \7290 , \7291 );
xnor \U$5418 ( \7293 , \7292 , \5901 );
xor \U$5419 ( \7294 , \7289 , \7293 );
and \U$5420 ( \7295 , \6085 , \5935 );
and \U$5421 ( \7296 , \6106 , \5933 );
nor \U$5422 ( \7297 , \7295 , \7296 );
xnor \U$5423 ( \7298 , \7297 , \5961 );
xor \U$5424 ( \7299 , \7294 , \7298 );
xor \U$5425 ( \7300 , \7285 , \7299 );
xor \U$5426 ( \7301 , \7281 , \7300 );
and \U$5427 ( \7302 , \5699 , \7272 );
and \U$5428 ( \7303 , \7272 , \7277 );
and \U$5429 ( \7304 , \5699 , \7277 );
or \U$5430 ( \7305 , \7302 , \7303 , \7304 );
and \U$5431 ( \7306 , \7259 , \7263 );
and \U$5432 ( \7307 , \7263 , \7266 );
and \U$5433 ( \7308 , \7259 , \7266 );
or \U$5434 ( \7309 , \7306 , \7307 , \7308 );
xor \U$5435 ( \7310 , \7305 , \7309 );
and \U$5436 ( \7311 , \6133 , \5993 );
and \U$5437 ( \7312 , \6154 , \5991 );
nor \U$5438 ( \7313 , \7311 , \7312 );
xnor \U$5439 ( \7314 , \7313 , \6019 );
xor \U$5440 ( \7315 , \7310 , \7314 );
xor \U$5441 ( \7316 , \7301 , \7315 );
and \U$5442 ( \7317 , \6106 , \5839 );
and \U$5443 ( \7318 , \6040 , \5836 );
nor \U$5444 ( \7319 , \7317 , \7318 );
xnor \U$5445 ( \7320 , \7319 , \5833 );
and \U$5446 ( \7321 , \6019 , \7320 );
and \U$5447 ( \7322 , \6154 , \5875 );
and \U$5448 ( \7323 , \6085 , \5873 );
nor \U$5449 ( \7324 , \7322 , \7323 );
xnor \U$5450 ( \7325 , \7324 , \5901 );
and \U$5451 ( \7326 , \7320 , \7325 );
and \U$5452 ( \7327 , \6019 , \7325 );
or \U$5453 ( \7328 , \7321 , \7326 , \7327 );
and \U$5454 ( \7329 , \6177 , \5935 );
and \U$5455 ( \7330 , \6133 , \5933 );
nor \U$5456 ( \7331 , \7329 , \7330 );
xnor \U$5457 ( \7332 , \7331 , \5961 );
nand \U$5458 ( \7333 , \6310 , \5991 );
xnor \U$5459 ( \7334 , \7333 , \6019 );
and \U$5460 ( \7335 , \7332 , \7334 );
and \U$5461 ( \7336 , \7328 , \7335 );
and \U$5462 ( \7337 , \6310 , \5993 );
and \U$5463 ( \7338 , \6177 , \5991 );
nor \U$5464 ( \7339 , \7337 , \7338 );
xnor \U$5465 ( \7340 , \7339 , \6019 );
and \U$5466 ( \7341 , \7335 , \7340 );
and \U$5467 ( \7342 , \7328 , \7340 );
or \U$5468 ( \7343 , \7336 , \7341 , \7342 );
xor \U$5469 ( \7344 , \7255 , \7267 );
xor \U$5470 ( \7345 , \7344 , \7278 );
and \U$5471 ( \7346 , \7343 , \7345 );
nor \U$5472 ( \7347 , \7316 , \7346 );
and \U$5473 ( \7348 , \7289 , \7293 );
and \U$5474 ( \7349 , \7293 , \7298 );
and \U$5475 ( \7350 , \7289 , \7298 );
or \U$5476 ( \7351 , \7348 , \7349 , \7350 );
nand \U$5477 ( \7352 , \6310 , \5627 );
xnor \U$5478 ( \7353 , \7352 , \5396 );
xor \U$5479 ( \7354 , \7351 , \7353 );
and \U$5480 ( \7355 , \6106 , \5935 );
and \U$5481 ( \7356 , \6040 , \5933 );
nor \U$5482 ( \7357 , \7355 , \7356 );
xnor \U$5483 ( \7358 , \7357 , \5961 );
and \U$5484 ( \7359 , \6154 , \5993 );
and \U$5485 ( \7360 , \6085 , \5991 );
nor \U$5486 ( \7361 , \7359 , \7360 );
xnor \U$5487 ( \7362 , \7361 , \6019 );
xor \U$5488 ( \7363 , \7358 , \7362 );
and \U$5489 ( \7364 , \6177 , \5694 );
and \U$5490 ( \7365 , \6133 , \5692 );
nor \U$5491 ( \7366 , \7364 , \7365 );
xnor \U$5492 ( \7367 , \7366 , \5699 );
xor \U$5493 ( \7368 , \7363 , \7367 );
xor \U$5494 ( \7369 , \7354 , \7368 );
and \U$5495 ( \7370 , \7305 , \7309 );
and \U$5496 ( \7371 , \7309 , \7314 );
and \U$5497 ( \7372 , \7305 , \7314 );
or \U$5498 ( \7373 , \7370 , \7371 , \7372 );
and \U$5499 ( \7374 , \7285 , \7299 );
xor \U$5500 ( \7375 , \7373 , \7374 );
and \U$5501 ( \7376 , \6014 , \5839 );
and \U$5502 ( \7377 , \5923 , \5836 );
nor \U$5503 ( \7378 , \7376 , \7377 );
xnor \U$5504 ( \7379 , \7378 , \5833 );
xor \U$5505 ( \7380 , \5396 , \7379 );
and \U$5506 ( \7381 , \6061 , \5875 );
and \U$5507 ( \7382 , \5985 , \5873 );
nor \U$5508 ( \7383 , \7381 , \7382 );
xnor \U$5509 ( \7384 , \7383 , \5901 );
xor \U$5510 ( \7385 , \7380 , \7384 );
xor \U$5511 ( \7386 , \7375 , \7385 );
xor \U$5512 ( \7387 , \7369 , \7386 );
and \U$5513 ( \7388 , \7281 , \7300 );
and \U$5514 ( \7389 , \7300 , \7315 );
and \U$5515 ( \7390 , \7281 , \7315 );
or \U$5516 ( \7391 , \7388 , \7389 , \7390 );
nor \U$5517 ( \7392 , \7387 , \7391 );
nor \U$5518 ( \7393 , \7347 , \7392 );
and \U$5519 ( \7394 , \7373 , \7374 );
and \U$5520 ( \7395 , \7374 , \7385 );
and \U$5521 ( \7396 , \7373 , \7385 );
or \U$5522 ( \7397 , \7394 , \7395 , \7396 );
and \U$5523 ( \7398 , \7351 , \7353 );
and \U$5524 ( \7399 , \7353 , \7368 );
and \U$5525 ( \7400 , \7351 , \7368 );
or \U$5526 ( \7401 , \7398 , \7399 , \7400 );
and \U$5527 ( \7402 , \5923 , \5839 );
and \U$5528 ( \7403 , \5956 , \5836 );
nor \U$5529 ( \7404 , \7402 , \7403 );
xnor \U$5530 ( \7405 , \7404 , \5833 );
and \U$5531 ( \7406 , \5985 , \5875 );
and \U$5532 ( \7407 , \6014 , \5873 );
nor \U$5533 ( \7408 , \7406 , \7407 );
xnor \U$5534 ( \7409 , \7408 , \5901 );
xor \U$5535 ( \7410 , \7405 , \7409 );
and \U$5536 ( \7411 , \6040 , \5935 );
and \U$5537 ( \7412 , \6061 , \5933 );
nor \U$5538 ( \7413 , \7411 , \7412 );
xnor \U$5539 ( \7414 , \7413 , \5961 );
xor \U$5540 ( \7415 , \7410 , \7414 );
xor \U$5541 ( \7416 , \7401 , \7415 );
and \U$5542 ( \7417 , \5396 , \7379 );
and \U$5543 ( \7418 , \7379 , \7384 );
and \U$5544 ( \7419 , \5396 , \7384 );
or \U$5545 ( \7420 , \7417 , \7418 , \7419 );
and \U$5546 ( \7421 , \7358 , \7362 );
and \U$5547 ( \7422 , \7362 , \7367 );
and \U$5548 ( \7423 , \7358 , \7367 );
or \U$5549 ( \7424 , \7421 , \7422 , \7423 );
xor \U$5550 ( \7425 , \7420 , \7424 );
and \U$5551 ( \7426 , \6085 , \5993 );
and \U$5552 ( \7427 , \6106 , \5991 );
nor \U$5553 ( \7428 , \7426 , \7427 );
xnor \U$5554 ( \7429 , \7428 , \6019 );
and \U$5555 ( \7430 , \6133 , \5694 );
and \U$5556 ( \7431 , \6154 , \5692 );
nor \U$5557 ( \7432 , \7430 , \7431 );
xnor \U$5558 ( \7433 , \7432 , \5699 );
xor \U$5559 ( \7434 , \7429 , \7433 );
and \U$5560 ( \7435 , \6310 , \5629 );
and \U$5561 ( \7436 , \6177 , \5627 );
nor \U$5562 ( \7437 , \7435 , \7436 );
xnor \U$5563 ( \7438 , \7437 , \5396 );
xor \U$5564 ( \7439 , \7434 , \7438 );
xor \U$5565 ( \7440 , \7425 , \7439 );
xor \U$5566 ( \7441 , \7416 , \7440 );
xor \U$5567 ( \7442 , \7397 , \7441 );
and \U$5568 ( \7443 , \7369 , \7386 );
nor \U$5569 ( \7444 , \7442 , \7443 );
and \U$5570 ( \7445 , \7401 , \7415 );
and \U$5571 ( \7446 , \7415 , \7440 );
and \U$5572 ( \7447 , \7401 , \7440 );
or \U$5573 ( \7448 , \7445 , \7446 , \7447 );
and \U$5574 ( \7449 , \7420 , \7424 );
and \U$5575 ( \7450 , \7424 , \7439 );
and \U$5576 ( \7451 , \7420 , \7439 );
or \U$5577 ( \7452 , \7449 , \7450 , \7451 );
nand \U$5578 ( \7453 , \6310 , \5565 );
xnor \U$5579 ( \7454 , \7453 , \5593 );
and \U$5580 ( \7455 , \6061 , \5935 );
and \U$5581 ( \7456 , \5985 , \5933 );
nor \U$5582 ( \7457 , \7455 , \7456 );
xnor \U$5583 ( \7458 , \7457 , \5961 );
and \U$5584 ( \7459 , \6106 , \5993 );
and \U$5585 ( \7460 , \6040 , \5991 );
nor \U$5586 ( \7461 , \7459 , \7460 );
xnor \U$5587 ( \7462 , \7461 , \6019 );
xor \U$5588 ( \7463 , \7458 , \7462 );
and \U$5589 ( \7464 , \6154 , \5694 );
and \U$5590 ( \7465 , \6085 , \5692 );
nor \U$5591 ( \7466 , \7464 , \7465 );
xnor \U$5592 ( \7467 , \7466 , \5699 );
xor \U$5593 ( \7468 , \7463 , \7467 );
xor \U$5594 ( \7469 , \7454 , \7468 );
and \U$5595 ( \7470 , \5956 , \5839 );
and \U$5596 ( \7471 , \5863 , \5836 );
nor \U$5597 ( \7472 , \7470 , \7471 );
xnor \U$5598 ( \7473 , \7472 , \5833 );
xor \U$5599 ( \7474 , \5593 , \7473 );
and \U$5600 ( \7475 , \6014 , \5875 );
and \U$5601 ( \7476 , \5923 , \5873 );
nor \U$5602 ( \7477 , \7475 , \7476 );
xnor \U$5603 ( \7478 , \7477 , \5901 );
xor \U$5604 ( \7479 , \7474 , \7478 );
xor \U$5605 ( \7480 , \7469 , \7479 );
xor \U$5606 ( \7481 , \7452 , \7480 );
and \U$5607 ( \7482 , \7405 , \7409 );
and \U$5608 ( \7483 , \7409 , \7414 );
and \U$5609 ( \7484 , \7405 , \7414 );
or \U$5610 ( \7485 , \7482 , \7483 , \7484 );
and \U$5611 ( \7486 , \7429 , \7433 );
and \U$5612 ( \7487 , \7433 , \7438 );
and \U$5613 ( \7488 , \7429 , \7438 );
or \U$5614 ( \7489 , \7486 , \7487 , \7488 );
xor \U$5615 ( \7490 , \7485 , \7489 );
and \U$5616 ( \7491 , \6177 , \5629 );
and \U$5617 ( \7492 , \6133 , \5627 );
nor \U$5618 ( \7493 , \7491 , \7492 );
xnor \U$5619 ( \7494 , \7493 , \5396 );
xor \U$5620 ( \7495 , \7490 , \7494 );
xor \U$5621 ( \7496 , \7481 , \7495 );
xor \U$5622 ( \7497 , \7448 , \7496 );
and \U$5623 ( \7498 , \7397 , \7441 );
nor \U$5624 ( \7499 , \7497 , \7498 );
nor \U$5625 ( \7500 , \7444 , \7499 );
nand \U$5626 ( \7501 , \7393 , \7500 );
and \U$5627 ( \7502 , \7452 , \7480 );
and \U$5628 ( \7503 , \7480 , \7495 );
and \U$5629 ( \7504 , \7452 , \7495 );
or \U$5630 ( \7505 , \7502 , \7503 , \7504 );
xor \U$5631 ( \7506 , \6365 , \6369 );
xor \U$5632 ( \7507 , \7506 , \6374 );
and \U$5633 ( \7508 , \5593 , \7473 );
and \U$5634 ( \7509 , \7473 , \7478 );
and \U$5635 ( \7510 , \5593 , \7478 );
or \U$5636 ( \7511 , \7508 , \7509 , \7510 );
and \U$5637 ( \7512 , \7458 , \7462 );
and \U$5638 ( \7513 , \7462 , \7467 );
and \U$5639 ( \7514 , \7458 , \7467 );
or \U$5640 ( \7515 , \7512 , \7513 , \7514 );
xor \U$5641 ( \7516 , \7511 , \7515 );
and \U$5642 ( \7517 , \6310 , \5567 );
and \U$5643 ( \7518 , \6177 , \5565 );
nor \U$5644 ( \7519 , \7517 , \7518 );
xnor \U$5645 ( \7520 , \7519 , \5593 );
xor \U$5646 ( \7521 , \7516 , \7520 );
xor \U$5647 ( \7522 , \7507 , \7521 );
xor \U$5648 ( \7523 , \7505 , \7522 );
and \U$5649 ( \7524 , \7485 , \7489 );
and \U$5650 ( \7525 , \7489 , \7494 );
and \U$5651 ( \7526 , \7485 , \7494 );
or \U$5652 ( \7527 , \7524 , \7525 , \7526 );
and \U$5653 ( \7528 , \7454 , \7468 );
and \U$5654 ( \7529 , \7468 , \7479 );
and \U$5655 ( \7530 , \7454 , \7479 );
or \U$5656 ( \7531 , \7528 , \7529 , \7530 );
xor \U$5657 ( \7532 , \7527 , \7531 );
xor \U$5658 ( \7533 , \6381 , \6385 );
xor \U$5659 ( \7534 , \7533 , \6390 );
xor \U$5660 ( \7535 , \7532 , \7534 );
xor \U$5661 ( \7536 , \7523 , \7535 );
and \U$5662 ( \7537 , \7448 , \7496 );
nor \U$5663 ( \7538 , \7536 , \7537 );
and \U$5664 ( \7539 , \7527 , \7531 );
and \U$5665 ( \7540 , \7531 , \7534 );
and \U$5666 ( \7541 , \7527 , \7534 );
or \U$5667 ( \7542 , \7539 , \7540 , \7541 );
and \U$5668 ( \7543 , \7507 , \7521 );
xor \U$5669 ( \7544 , \7542 , \7543 );
and \U$5670 ( \7545 , \7511 , \7515 );
and \U$5671 ( \7546 , \7515 , \7520 );
and \U$5672 ( \7547 , \7511 , \7520 );
or \U$5673 ( \7548 , \7545 , \7546 , \7547 );
xor \U$5674 ( \7549 , \6401 , \6403 );
xor \U$5675 ( \7550 , \7548 , \7549 );
xor \U$5676 ( \7551 , \6377 , \6393 );
xor \U$5677 ( \7552 , \7551 , \6396 );
xor \U$5678 ( \7553 , \7550 , \7552 );
xor \U$5679 ( \7554 , \7544 , \7553 );
and \U$5680 ( \7555 , \7505 , \7522 );
and \U$5681 ( \7556 , \7522 , \7535 );
and \U$5682 ( \7557 , \7505 , \7535 );
or \U$5683 ( \7558 , \7555 , \7556 , \7557 );
nor \U$5684 ( \7559 , \7554 , \7558 );
nor \U$5685 ( \7560 , \7538 , \7559 );
and \U$5686 ( \7561 , \7548 , \7549 );
and \U$5687 ( \7562 , \7549 , \7552 );
and \U$5688 ( \7563 , \7548 , \7552 );
or \U$5689 ( \7564 , \7561 , \7562 , \7563 );
xor \U$5690 ( \7565 , \6264 , \6280 );
xor \U$5691 ( \7566 , \7565 , \6315 );
xor \U$5692 ( \7567 , \7564 , \7566 );
xor \U$5693 ( \7568 , \6399 , \6404 );
xor \U$5694 ( \7569 , \7568 , \6407 );
xor \U$5695 ( \7570 , \7567 , \7569 );
and \U$5696 ( \7571 , \7542 , \7543 );
and \U$5697 ( \7572 , \7543 , \7553 );
and \U$5698 ( \7573 , \7542 , \7553 );
or \U$5699 ( \7574 , \7571 , \7572 , \7573 );
nor \U$5700 ( \7575 , \7570 , \7574 );
xor \U$5701 ( \7576 , \6410 , \6411 );
xor \U$5702 ( \7577 , \7576 , \6414 );
and \U$5703 ( \7578 , \7564 , \7566 );
and \U$5704 ( \7579 , \7566 , \7569 );
and \U$5705 ( \7580 , \7564 , \7569 );
or \U$5706 ( \7581 , \7578 , \7579 , \7580 );
nor \U$5707 ( \7582 , \7577 , \7581 );
nor \U$5708 ( \7583 , \7575 , \7582 );
nand \U$5709 ( \7584 , \7560 , \7583 );
nor \U$5710 ( \7585 , \7501 , \7584 );
and \U$5711 ( \7586 , \6154 , \5839 );
and \U$5712 ( \7587 , \6085 , \5836 );
nor \U$5713 ( \7588 , \7586 , \7587 );
xnor \U$5714 ( \7589 , \7588 , \5833 );
and \U$5715 ( \7590 , \5961 , \7589 );
and \U$5716 ( \7591 , \6177 , \5875 );
and \U$5717 ( \7592 , \6133 , \5873 );
nor \U$5718 ( \7593 , \7591 , \7592 );
xnor \U$5719 ( \7594 , \7593 , \5901 );
and \U$5720 ( \7595 , \7589 , \7594 );
and \U$5721 ( \7596 , \5961 , \7594 );
or \U$5722 ( \7597 , \7590 , \7595 , \7596 );
and \U$5723 ( \7598 , \6085 , \5839 );
and \U$5724 ( \7599 , \6106 , \5836 );
nor \U$5725 ( \7600 , \7598 , \7599 );
xnor \U$5726 ( \7601 , \7600 , \5833 );
and \U$5727 ( \7602 , \6133 , \5875 );
and \U$5728 ( \7603 , \6154 , \5873 );
nor \U$5729 ( \7604 , \7602 , \7603 );
xnor \U$5730 ( \7605 , \7604 , \5901 );
xor \U$5731 ( \7606 , \7601 , \7605 );
and \U$5732 ( \7607 , \6310 , \5935 );
and \U$5733 ( \7608 , \6177 , \5933 );
nor \U$5734 ( \7609 , \7607 , \7608 );
xnor \U$5735 ( \7610 , \7609 , \5961 );
xor \U$5736 ( \7611 , \7606 , \7610 );
xor \U$5737 ( \7612 , \7597 , \7611 );
nand \U$5738 ( \7613 , \6310 , \5933 );
xnor \U$5739 ( \7614 , \7613 , \5961 );
xor \U$5740 ( \7615 , \5961 , \7589 );
xor \U$5741 ( \7616 , \7615 , \7594 );
and \U$5742 ( \7617 , \7614 , \7616 );
nor \U$5743 ( \7618 , \7612 , \7617 );
and \U$5744 ( \7619 , \7601 , \7605 );
and \U$5745 ( \7620 , \7605 , \7610 );
and \U$5746 ( \7621 , \7601 , \7610 );
or \U$5747 ( \7622 , \7619 , \7620 , \7621 );
xor \U$5748 ( \7623 , \7332 , \7334 );
xor \U$5749 ( \7624 , \7622 , \7623 );
xor \U$5750 ( \7625 , \6019 , \7320 );
xor \U$5751 ( \7626 , \7625 , \7325 );
xor \U$5752 ( \7627 , \7624 , \7626 );
and \U$5753 ( \7628 , \7597 , \7611 );
nor \U$5754 ( \7629 , \7627 , \7628 );
nor \U$5755 ( \7630 , \7618 , \7629 );
xor \U$5756 ( \7631 , \7243 , \7247 );
xor \U$5757 ( \7632 , \7631 , \7252 );
xor \U$5758 ( \7633 , \7328 , \7335 );
xor \U$5759 ( \7634 , \7633 , \7340 );
xor \U$5760 ( \7635 , \7632 , \7634 );
and \U$5761 ( \7636 , \7622 , \7623 );
and \U$5762 ( \7637 , \7623 , \7626 );
and \U$5763 ( \7638 , \7622 , \7626 );
or \U$5764 ( \7639 , \7636 , \7637 , \7638 );
nor \U$5765 ( \7640 , \7635 , \7639 );
xor \U$5766 ( \7641 , \7343 , \7345 );
and \U$5767 ( \7642 , \7632 , \7634 );
nor \U$5768 ( \7643 , \7641 , \7642 );
nor \U$5769 ( \7644 , \7640 , \7643 );
nand \U$5770 ( \7645 , \7630 , \7644 );
and \U$5771 ( \7646 , \6133 , \5839 );
and \U$5772 ( \7647 , \6154 , \5836 );
nor \U$5773 ( \7648 , \7646 , \7647 );
xnor \U$5774 ( \7649 , \7648 , \5833 );
and \U$5775 ( \7650 , \6310 , \5875 );
and \U$5776 ( \7651 , \6177 , \5873 );
nor \U$5777 ( \7652 , \7650 , \7651 );
xnor \U$5778 ( \7653 , \7652 , \5901 );
xor \U$5779 ( \7654 , \7649 , \7653 );
and \U$5780 ( \7655 , \6177 , \5839 );
and \U$5781 ( \7656 , \6133 , \5836 );
nor \U$5782 ( \7657 , \7655 , \7656 );
xnor \U$5783 ( \7658 , \7657 , \5833 );
and \U$5784 ( \7659 , \7658 , \5901 );
nor \U$5785 ( \7660 , \7654 , \7659 );
xor \U$5786 ( \7661 , \7614 , \7616 );
and \U$5787 ( \7662 , \7649 , \7653 );
nor \U$5788 ( \7663 , \7661 , \7662 );
nor \U$5789 ( \7664 , \7660 , \7663 );
xor \U$5790 ( \7665 , \7658 , \5901 );
nand \U$5791 ( \7666 , \6310 , \5873 );
xnor \U$5792 ( \7667 , \7666 , \5901 );
nor \U$5793 ( \7668 , \7665 , \7667 );
and \U$5794 ( \7669 , \6310 , \5839 );
and \U$5795 ( \7670 , \6177 , \5836 );
nor \U$5796 ( \7671 , \7669 , \7670 );
xnor \U$5797 ( \7672 , \7671 , \5833 );
nand \U$5798 ( \7673 , \6310 , \5836 );
xnor \U$5799 ( \7674 , \7673 , \5833 );
and \U$5800 ( \7675 , \7674 , \5833 );
nand \U$5801 ( \7676 , \7672 , \7675 );
or \U$5802 ( \7677 , \7668 , \7676 );
nand \U$5803 ( \7678 , \7665 , \7667 );
nand \U$5804 ( \7679 , \7677 , \7678 );
and \U$5805 ( \7680 , \7664 , \7679 );
nand \U$5806 ( \7681 , \7654 , \7659 );
or \U$5807 ( \7682 , \7663 , \7681 );
nand \U$5808 ( \7683 , \7661 , \7662 );
nand \U$5809 ( \7684 , \7682 , \7683 );
nor \U$5810 ( \7685 , \7680 , \7684 );
or \U$5811 ( \7686 , \7645 , \7685 );
nand \U$5812 ( \7687 , \7612 , \7617 );
or \U$5813 ( \7688 , \7629 , \7687 );
nand \U$5814 ( \7689 , \7627 , \7628 );
nand \U$5815 ( \7690 , \7688 , \7689 );
and \U$5816 ( \7691 , \7644 , \7690 );
nand \U$5817 ( \7692 , \7635 , \7639 );
or \U$5818 ( \7693 , \7643 , \7692 );
nand \U$5819 ( \7694 , \7641 , \7642 );
nand \U$5820 ( \7695 , \7693 , \7694 );
nor \U$5821 ( \7696 , \7691 , \7695 );
nand \U$5822 ( \7697 , \7686 , \7696 );
and \U$5823 ( \7698 , \7585 , \7697 );
nand \U$5824 ( \7699 , \7316 , \7346 );
or \U$5825 ( \7700 , \7392 , \7699 );
nand \U$5826 ( \7701 , \7387 , \7391 );
nand \U$5827 ( \7702 , \7700 , \7701 );
and \U$5828 ( \7703 , \7500 , \7702 );
nand \U$5829 ( \7704 , \7442 , \7443 );
or \U$5830 ( \7705 , \7499 , \7704 );
nand \U$5831 ( \7706 , \7497 , \7498 );
nand \U$5832 ( \7707 , \7705 , \7706 );
nor \U$5833 ( \7708 , \7703 , \7707 );
or \U$5834 ( \7709 , \7584 , \7708 );
nand \U$5835 ( \7710 , \7536 , \7537 );
or \U$5836 ( \7711 , \7559 , \7710 );
nand \U$5837 ( \7712 , \7554 , \7558 );
nand \U$5838 ( \7713 , \7711 , \7712 );
and \U$5839 ( \7714 , \7583 , \7713 );
nand \U$5840 ( \7715 , \7570 , \7574 );
or \U$5841 ( \7716 , \7582 , \7715 );
nand \U$5842 ( \7717 , \7577 , \7581 );
nand \U$5843 ( \7718 , \7716 , \7717 );
nor \U$5844 ( \7719 , \7714 , \7718 );
nand \U$5845 ( \7720 , \7709 , \7719 );
nor \U$5846 ( \7721 , \7698 , \7720 );
or \U$5847 ( \7722 , \7239 , \7721 );
nand \U$5848 ( \7723 , \6361 , \6417 );
or \U$5849 ( \7724 , \6493 , \7723 );
nand \U$5850 ( \7725 , \6491 , \6492 );
nand \U$5851 ( \7726 , \7724 , \7725 );
and \U$5852 ( \7727 , \6646 , \7726 );
nand \U$5853 ( \7728 , \6568 , \6569 );
or \U$5854 ( \7729 , \6645 , \7728 );
nand \U$5855 ( \7730 , \6640 , \6644 );
nand \U$5856 ( \7731 , \7729 , \7730 );
nor \U$5857 ( \7732 , \7727 , \7731 );
or \U$5858 ( \7733 , \6942 , \7732 );
nand \U$5859 ( \7734 , \6717 , \6721 );
or \U$5860 ( \7735 , \6798 , \7734 );
nand \U$5861 ( \7736 , \6793 , \6797 );
nand \U$5862 ( \7737 , \7735 , \7736 );
and \U$5863 ( \7738 , \6941 , \7737 );
nand \U$5864 ( \7739 , \6866 , \6870 );
or \U$5865 ( \7740 , \6940 , \7739 );
nand \U$5866 ( \7741 , \6935 , \6939 );
nand \U$5867 ( \7742 , \7740 , \7741 );
nor \U$5868 ( \7743 , \7738 , \7742 );
nand \U$5869 ( \7744 , \7733 , \7743 );
and \U$5870 ( \7745 , \7238 , \7744 );
nand \U$5871 ( \7746 , \6999 , \7003 );
or \U$5872 ( \7747 , \7064 , \7746 );
nand \U$5873 ( \7748 , \7059 , \7063 );
nand \U$5874 ( \7749 , \7747 , \7748 );
and \U$5875 ( \7750 , \7160 , \7749 );
nand \U$5876 ( \7751 , \7116 , \7120 );
or \U$5877 ( \7752 , \7159 , \7751 );
nand \U$5878 ( \7753 , \7154 , \7158 );
nand \U$5879 ( \7754 , \7752 , \7753 );
nor \U$5880 ( \7755 , \7750 , \7754 );
or \U$5881 ( \7756 , \7237 , \7755 );
nand \U$5882 ( \7757 , \7186 , \7190 );
or \U$5883 ( \7758 , \7212 , \7757 );
nand \U$5884 ( \7759 , \7207 , \7211 );
nand \U$5885 ( \7760 , \7758 , \7759 );
and \U$5886 ( \7761 , \7236 , \7760 );
nand \U$5887 ( \7762 , \7223 , \7227 );
or \U$5888 ( \7763 , \7235 , \7762 );
nand \U$5889 ( \7764 , \7230 , \7234 );
nand \U$5890 ( \7765 , \7763 , \7764 );
nor \U$5891 ( \7766 , \7761 , \7765 );
nand \U$5892 ( \7767 , \7756 , \7766 );
nor \U$5893 ( \7768 , \7745 , \7767 );
nand \U$5894 ( \7769 , \7722 , \7768 );
not \U$5895 ( \7770 , \7769 );
xor \U$5896 ( \7771 , \5829 , \7770 );
buf g32b2_GF_PartitionCandidate( \7772_nG32b2 , \7771 );
buf \U$5897 ( \7773 , RI2b5e785ebd68_1);
buf \U$5898 ( \7774 , RI2b5e785ebcf0_2);
buf \U$5899 ( \7775 , RI2b5e785ebc78_3);
buf \U$5900 ( \7776 , RI2b5e785ebc00_4);
buf \U$5901 ( \7777 , RI2b5e785ebb88_5);
buf \U$5902 ( \7778 , RI2b5e785ebb10_6);
buf \U$5903 ( \7779 , RI2b5e785eba98_7);
buf \U$5904 ( \7780 , RI2b5e785eba20_8);
buf \U$5905 ( \7781 , RI2b5e785eb9a8_9);
buf \U$5906 ( \7782 , RI2b5e785eb930_10);
buf \U$5907 ( \7783 , RI2b5e785eb8b8_11);
buf \U$5908 ( \7784 , RI2b5e785eb840_12);
not \U$5909 ( \7785 , RI2b5e785ae328_614);
buf \U$5910 ( \7786 , \7785 );
and \U$5911 ( \7787 , \7784 , \7786 );
and \U$5912 ( \7788 , \7783 , \7787 );
and \U$5913 ( \7789 , \7782 , \7788 );
and \U$5914 ( \7790 , \7781 , \7789 );
and \U$5915 ( \7791 , \7780 , \7790 );
and \U$5916 ( \7792 , \7779 , \7791 );
and \U$5917 ( \7793 , \7778 , \7792 );
and \U$5918 ( \7794 , \7777 , \7793 );
and \U$5919 ( \7795 , \7776 , \7794 );
and \U$5920 ( \7796 , \7775 , \7795 );
and \U$5921 ( \7797 , \7774 , \7796 );
xor \U$5922 ( \7798 , \7773 , \7797 );
buf \U$5923 ( \7799 , \7798 );
buf \U$5924 ( \7800 , \7799 );
not \U$5925 ( \7801 , \7800 );
nor \U$5926 ( \7802 , \4969 , \4973 , \4977 , \4981 , \4986 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5927 ( \7803 , RI2b5e785daab8_27, \7802 );
nor \U$5928 ( \7804 , \5021 , \5022 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5929 ( \7805 , RI2b5e785495b8_40, \7804 );
nor \U$5930 ( \7806 , \4969 , \5022 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5931 ( \7807 , RI2b5e78538920_53, \7806 );
nor \U$5932 ( \7808 , \5021 , \4973 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5933 ( \7809 , RI2b5e784a63a8_66, \7808 );
nor \U$5934 ( \7810 , \4969 , \4973 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5935 ( \7811 , RI2b5e78495710_79, \7810 );
nor \U$5936 ( \7812 , \5021 , \5022 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5937 ( \7813 , RI2b5e784950f8_92, \7812 );
nor \U$5938 ( \7814 , \4969 , \5022 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5939 ( \7815 , RI2b5e78403bf8_105, \7814 );
nor \U$5940 ( \7816 , \5021 , \4973 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5941 ( \7817 , RI2b5e775b1ed8_118, \7816 );
nor \U$5942 ( \7818 , \4969 , \4973 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5943 ( \7819 , RI2b5e775b18c0_131, \7818 );
nor \U$5944 ( \7820 , \5021 , \5022 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5945 ( \7821 , RI2b5e7750b858_144, \7820 );
nor \U$5946 ( \7822 , \4969 , \5022 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5947 ( \7823 , RI2b5e774ff030_157, \7822 );
nor \U$5948 ( \7824 , \5021 , \4973 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5949 ( \7825 , RI2b5e774f6048_170, \7824 );
nor \U$5950 ( \7826 , \4969 , \4973 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5951 ( \7827 , RI2b5e774ea630_183, \7826 );
nor \U$5952 ( \7828 , \5021 , \5022 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5953 ( \7829 , RI2b5e774dde08_196, \7828 );
nor \U$5954 ( \7830 , \4969 , \5022 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5955 ( \7831 , RI2b5e774d4e20_209, \7830 );
nor \U$5956 ( \7832 , \5021 , \4973 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5957 ( \7833 , RI2b5e785f3d60_222, \7832 );
nor \U$5958 ( \7834 , \4969 , \4973 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$5959 ( \7835 , RI2b5e785eb138_235, \7834 );
or \U$5960 ( \7836 , \7803 , \7805 , \7807 , \7809 , \7811 , \7813 , \7815 , \7817 , \7819 , \7821 , \7823 , \7825 , \7827 , \7829 , \7831 , \7833 , \7835 );
buf \U$5961 ( \7837 , \4990 );
buf \U$5962 ( \7838 , \4994 );
buf \U$5963 ( \7839 , \4998 );
buf \U$5964 ( \7840 , \5002 );
buf \U$5965 ( \7841 , \5006 );
buf \U$5966 ( \7842 , \5010 );
buf \U$5967 ( \7843 , \5014 );
buf \U$5968 ( \7844 , \5018 );
buf \U$5969 ( \7845 , \4985 );
buf \U$5970 ( \7846 , \4969 );
buf \U$5971 ( \7847 , \4973 );
buf \U$5972 ( \7848 , \4977 );
buf \U$5973 ( \7849 , \4981 );
or \U$5974 ( \7850 , \7846 , \7847 , \7848 , \7849 );
and \U$5975 ( \7851 , \7845 , \7850 );
or \U$5976 ( \7852 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7851 );
buf \U$5977 ( \7853 , \7852 );
_DC g1080 ( \7854_nG1080 , \7836 , \7853 );
buf \U$5978 ( \7855 , \7854_nG1080 );
and \U$5979 ( \7856 , \7801 , \7855 );
xor \U$5980 ( \7857 , \7774 , \7796 );
buf \U$5981 ( \7858 , \7857 );
buf \U$5982 ( \7859 , \7858 );
not \U$5983 ( \7860 , \7859 );
and \U$5984 ( \7861 , RI2b5e785daa40_28, \7802 );
and \U$5985 ( \7862 , RI2b5e78549540_41, \7804 );
and \U$5986 ( \7863 , RI2b5e785388a8_54, \7806 );
and \U$5987 ( \7864 , RI2b5e784a6330_67, \7808 );
and \U$5988 ( \7865 , RI2b5e78495698_80, \7810 );
and \U$5989 ( \7866 , RI2b5e78495080_93, \7812 );
and \U$5990 ( \7867 , RI2b5e78403b80_106, \7814 );
and \U$5991 ( \7868 , RI2b5e775b1e60_119, \7816 );
and \U$5992 ( \7869 , RI2b5e7750bdf8_132, \7818 );
and \U$5993 ( \7870 , RI2b5e774ff5d0_145, \7820 );
and \U$5994 ( \7871 , RI2b5e774f65e8_158, \7822 );
and \U$5995 ( \7872 , RI2b5e774eabd0_171, \7824 );
and \U$5996 ( \7873 , RI2b5e774de3a8_184, \7826 );
and \U$5997 ( \7874 , RI2b5e774d53c0_197, \7828 );
and \U$5998 ( \7875 , RI2b5e785f4300_210, \7830 );
and \U$5999 ( \7876 , RI2b5e785f3ce8_223, \7832 );
and \U$6000 ( \7877 , RI2b5e785eb0c0_236, \7834 );
or \U$6001 ( \7878 , \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 );
_DC g1099 ( \7879_nG1099 , \7878 , \7853 );
buf \U$6002 ( \7880 , \7879_nG1099 );
and \U$6003 ( \7881 , \7860 , \7880 );
xor \U$6004 ( \7882 , \7775 , \7795 );
buf \U$6005 ( \7883 , \7882 );
buf \U$6006 ( \7884 , \7883 );
not \U$6007 ( \7885 , \7884 );
and \U$6008 ( \7886 , RI2b5e785da9c8_29, \7802 );
and \U$6009 ( \7887 , RI2b5e785494c8_42, \7804 );
and \U$6010 ( \7888 , RI2b5e78538830_55, \7806 );
and \U$6011 ( \7889 , RI2b5e784a62b8_68, \7808 );
and \U$6012 ( \7890 , RI2b5e78495620_81, \7810 );
and \U$6013 ( \7891 , RI2b5e78495008_94, \7812 );
and \U$6014 ( \7892 , RI2b5e78403b08_107, \7814 );
and \U$6015 ( \7893 , RI2b5e775b1de8_120, \7816 );
and \U$6016 ( \7894 , RI2b5e7750bd80_133, \7818 );
and \U$6017 ( \7895 , RI2b5e774ff558_146, \7820 );
and \U$6018 ( \7896 , RI2b5e774f6570_159, \7822 );
and \U$6019 ( \7897 , RI2b5e774eab58_172, \7824 );
and \U$6020 ( \7898 , RI2b5e774de330_185, \7826 );
and \U$6021 ( \7899 , RI2b5e774d5348_198, \7828 );
and \U$6022 ( \7900 , RI2b5e785f4288_211, \7830 );
and \U$6023 ( \7901 , RI2b5e785f3658_224, \7832 );
and \U$6024 ( \7902 , RI2b5e785eb048_237, \7834 );
or \U$6025 ( \7903 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 );
_DC g10b2 ( \7904_nG10b2 , \7903 , \7853 );
buf \U$6026 ( \7905 , \7904_nG10b2 );
and \U$6027 ( \7906 , \7885 , \7905 );
xor \U$6028 ( \7907 , \7776 , \7794 );
buf \U$6029 ( \7908 , \7907 );
buf \U$6030 ( \7909 , \7908 );
not \U$6031 ( \7910 , \7909 );
and \U$6032 ( \7911 , RI2b5e785da950_30, \7802 );
and \U$6033 ( \7912 , RI2b5e78549450_43, \7804 );
and \U$6034 ( \7913 , RI2b5e785387b8_56, \7806 );
and \U$6035 ( \7914 , RI2b5e784a6240_69, \7808 );
and \U$6036 ( \7915 , RI2b5e784955a8_82, \7810 );
and \U$6037 ( \7916 , RI2b5e78494f90_95, \7812 );
and \U$6038 ( \7917 , RI2b5e78403a90_108, \7814 );
and \U$6039 ( \7918 , RI2b5e775b1d70_121, \7816 );
and \U$6040 ( \7919 , RI2b5e7750bd08_134, \7818 );
and \U$6041 ( \7920 , RI2b5e774ff4e0_147, \7820 );
and \U$6042 ( \7921 , RI2b5e774f64f8_160, \7822 );
and \U$6043 ( \7922 , RI2b5e774eaae0_173, \7824 );
and \U$6044 ( \7923 , RI2b5e774de2b8_186, \7826 );
and \U$6045 ( \7924 , RI2b5e774d52d0_199, \7828 );
and \U$6046 ( \7925 , RI2b5e785f4210_212, \7830 );
and \U$6047 ( \7926 , RI2b5e785eb5e8_225, \7832 );
and \U$6048 ( \7927 , RI2b5e785e6c50_238, \7834 );
or \U$6049 ( \7928 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 );
_DC g10cb ( \7929_nG10cb , \7928 , \7853 );
buf \U$6050 ( \7930 , \7929_nG10cb );
and \U$6051 ( \7931 , \7910 , \7930 );
xor \U$6052 ( \7932 , \7777 , \7793 );
buf \U$6053 ( \7933 , \7932 );
buf \U$6054 ( \7934 , \7933 );
not \U$6055 ( \7935 , \7934 );
and \U$6056 ( \7936 , RI2b5e785da8d8_31, \7802 );
and \U$6057 ( \7937 , RI2b5e785493d8_44, \7804 );
and \U$6058 ( \7938 , RI2b5e78538740_57, \7806 );
and \U$6059 ( \7939 , RI2b5e784a61c8_70, \7808 );
and \U$6060 ( \7940 , RI2b5e78495530_83, \7810 );
and \U$6061 ( \7941 , RI2b5e78494f18_96, \7812 );
and \U$6062 ( \7942 , RI2b5e78403a18_109, \7814 );
and \U$6063 ( \7943 , RI2b5e775b1cf8_122, \7816 );
and \U$6064 ( \7944 , RI2b5e7750bc90_135, \7818 );
and \U$6065 ( \7945 , RI2b5e774ff468_148, \7820 );
and \U$6066 ( \7946 , RI2b5e774f6480_161, \7822 );
and \U$6067 ( \7947 , RI2b5e774eaa68_174, \7824 );
and \U$6068 ( \7948 , RI2b5e774de240_187, \7826 );
and \U$6069 ( \7949 , RI2b5e774d5258_200, \7828 );
and \U$6070 ( \7950 , RI2b5e785f4198_213, \7830 );
and \U$6071 ( \7951 , RI2b5e785eb570_226, \7832 );
and \U$6072 ( \7952 , RI2b5e785e6bd8_239, \7834 );
or \U$6073 ( \7953 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 );
_DC g10e4 ( \7954_nG10e4 , \7953 , \7853 );
buf \U$6074 ( \7955 , \7954_nG10e4 );
and \U$6075 ( \7956 , \7935 , \7955 );
xor \U$6076 ( \7957 , \7778 , \7792 );
buf \U$6077 ( \7958 , \7957 );
buf \U$6078 ( \7959 , \7958 );
not \U$6079 ( \7960 , \7959 );
and \U$6080 ( \7961 , RI2b5e785da860_32, \7802 );
and \U$6081 ( \7962 , RI2b5e78549360_45, \7804 );
and \U$6082 ( \7963 , RI2b5e785386c8_58, \7806 );
and \U$6083 ( \7964 , RI2b5e784a6150_71, \7808 );
and \U$6084 ( \7965 , RI2b5e784954b8_84, \7810 );
and \U$6085 ( \7966 , RI2b5e78494ea0_97, \7812 );
and \U$6086 ( \7967 , RI2b5e784039a0_110, \7814 );
and \U$6087 ( \7968 , RI2b5e775b1c80_123, \7816 );
and \U$6088 ( \7969 , RI2b5e7750bc18_136, \7818 );
and \U$6089 ( \7970 , RI2b5e774ff3f0_149, \7820 );
and \U$6090 ( \7971 , RI2b5e774f6408_162, \7822 );
and \U$6091 ( \7972 , RI2b5e774ea9f0_175, \7824 );
and \U$6092 ( \7973 , RI2b5e774de1c8_188, \7826 );
and \U$6093 ( \7974 , RI2b5e774d51e0_201, \7828 );
and \U$6094 ( \7975 , RI2b5e785f4120_214, \7830 );
and \U$6095 ( \7976 , RI2b5e785eb4f8_227, \7832 );
and \U$6096 ( \7977 , RI2b5e785e64d0_240, \7834 );
or \U$6097 ( \7978 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 );
_DC g10fd ( \7979_nG10fd , \7978 , \7853 );
buf \U$6098 ( \7980 , \7979_nG10fd );
and \U$6099 ( \7981 , \7960 , \7980 );
xor \U$6100 ( \7982 , \7779 , \7791 );
buf \U$6101 ( \7983 , \7982 );
buf \U$6102 ( \7984 , \7983 );
not \U$6103 ( \7985 , \7984 );
and \U$6104 ( \7986 , RI2b5e78549900_33, \7802 );
and \U$6105 ( \7987 , RI2b5e78538c68_46, \7804 );
and \U$6106 ( \7988 , RI2b5e78538650_59, \7806 );
and \U$6107 ( \7989 , RI2b5e784a60d8_72, \7808 );
and \U$6108 ( \7990 , RI2b5e78495440_85, \7810 );
and \U$6109 ( \7991 , RI2b5e78494e28_98, \7812 );
and \U$6110 ( \7992 , RI2b5e78403928_111, \7814 );
and \U$6111 ( \7993 , RI2b5e775b1c08_124, \7816 );
and \U$6112 ( \7994 , RI2b5e7750bba0_137, \7818 );
and \U$6113 ( \7995 , RI2b5e774ff378_150, \7820 );
and \U$6114 ( \7996 , RI2b5e774f6390_163, \7822 );
and \U$6115 ( \7997 , RI2b5e774ea978_176, \7824 );
and \U$6116 ( \7998 , RI2b5e774de150_189, \7826 );
and \U$6117 ( \7999 , RI2b5e774d5168_202, \7828 );
and \U$6118 ( \8000 , RI2b5e785f40a8_215, \7830 );
and \U$6119 ( \8001 , RI2b5e785eb480_228, \7832 );
and \U$6120 ( \8002 , RI2b5e785da608_241, \7834 );
or \U$6121 ( \8003 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 );
_DC g1116 ( \8004_nG1116 , \8003 , \7853 );
buf \U$6122 ( \8005 , \8004_nG1116 );
and \U$6123 ( \8006 , \7985 , \8005 );
xor \U$6124 ( \8007 , \7780 , \7790 );
buf \U$6125 ( \8008 , \8007 );
buf \U$6126 ( \8009 , \8008 );
not \U$6127 ( \8010 , \8009 );
and \U$6128 ( \8011 , RI2b5e78549888_34, \7802 );
and \U$6129 ( \8012 , RI2b5e78538bf0_47, \7804 );
and \U$6130 ( \8013 , RI2b5e785385d8_60, \7806 );
and \U$6131 ( \8014 , RI2b5e784a6060_73, \7808 );
and \U$6132 ( \8015 , RI2b5e784953c8_86, \7810 );
and \U$6133 ( \8016 , RI2b5e78403ec8_99, \7812 );
and \U$6134 ( \8017 , RI2b5e775b21a8_112, \7814 );
and \U$6135 ( \8018 , RI2b5e775b1b90_125, \7816 );
and \U$6136 ( \8019 , RI2b5e7750bb28_138, \7818 );
and \U$6137 ( \8020 , RI2b5e774ff300_151, \7820 );
and \U$6138 ( \8021 , RI2b5e774f6318_164, \7822 );
and \U$6139 ( \8022 , RI2b5e774ea900_177, \7824 );
and \U$6140 ( \8023 , RI2b5e774de0d8_190, \7826 );
and \U$6141 ( \8024 , RI2b5e774d50f0_203, \7828 );
and \U$6142 ( \8025 , RI2b5e785f4030_216, \7830 );
and \U$6143 ( \8026 , RI2b5e785eb408_229, \7832 );
and \U$6144 ( \8027 , RI2b5e785da590_242, \7834 );
or \U$6145 ( \8028 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 );
_DC g112f ( \8029_nG112f , \8028 , \7853 );
buf \U$6146 ( \8030 , \8029_nG112f );
and \U$6147 ( \8031 , \8010 , \8030 );
xor \U$6148 ( \8032 , \7781 , \7789 );
buf \U$6149 ( \8033 , \8032 );
buf \U$6150 ( \8034 , \8033 );
not \U$6151 ( \8035 , \8034 );
and \U$6152 ( \8036 , RI2b5e78549810_35, \7802 );
and \U$6153 ( \8037 , RI2b5e78538b78_48, \7804 );
and \U$6154 ( \8038 , RI2b5e78538560_61, \7806 );
and \U$6155 ( \8039 , RI2b5e784a5fe8_74, \7808 );
and \U$6156 ( \8040 , RI2b5e78495350_87, \7810 );
and \U$6157 ( \8041 , RI2b5e78403e50_100, \7812 );
and \U$6158 ( \8042 , RI2b5e775b2130_113, \7814 );
and \U$6159 ( \8043 , RI2b5e775b1b18_126, \7816 );
and \U$6160 ( \8044 , RI2b5e7750bab0_139, \7818 );
and \U$6161 ( \8045 , RI2b5e774ff288_152, \7820 );
and \U$6162 ( \8046 , RI2b5e774f62a0_165, \7822 );
and \U$6163 ( \8047 , RI2b5e774ea888_178, \7824 );
and \U$6164 ( \8048 , RI2b5e774de060_191, \7826 );
and \U$6165 ( \8049 , RI2b5e774d5078_204, \7828 );
and \U$6166 ( \8050 , RI2b5e785f3fb8_217, \7830 );
and \U$6167 ( \8051 , RI2b5e785eb390_230, \7832 );
and \U$6168 ( \8052 , RI2b5e785da518_243, \7834 );
or \U$6169 ( \8053 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 );
_DC g1148 ( \8054_nG1148 , \8053 , \7853 );
buf \U$6170 ( \8055 , \8054_nG1148 );
and \U$6171 ( \8056 , \8035 , \8055 );
xor \U$6172 ( \8057 , \7782 , \7788 );
buf \U$6173 ( \8058 , \8057 );
buf \U$6174 ( \8059 , \8058 );
not \U$6175 ( \8060 , \8059 );
and \U$6176 ( \8061 , RI2b5e78549798_36, \7802 );
and \U$6177 ( \8062 , RI2b5e78538b00_49, \7804 );
and \U$6178 ( \8063 , RI2b5e785384e8_62, \7806 );
and \U$6179 ( \8064 , RI2b5e784a5f70_75, \7808 );
and \U$6180 ( \8065 , RI2b5e784952d8_88, \7810 );
and \U$6181 ( \8066 , RI2b5e78403dd8_101, \7812 );
and \U$6182 ( \8067 , RI2b5e775b20b8_114, \7814 );
and \U$6183 ( \8068 , RI2b5e775b1aa0_127, \7816 );
and \U$6184 ( \8069 , RI2b5e7750ba38_140, \7818 );
and \U$6185 ( \8070 , RI2b5e774ff210_153, \7820 );
and \U$6186 ( \8071 , RI2b5e774f6228_166, \7822 );
and \U$6187 ( \8072 , RI2b5e774ea810_179, \7824 );
and \U$6188 ( \8073 , RI2b5e774ddfe8_192, \7826 );
and \U$6189 ( \8074 , RI2b5e774d5000_205, \7828 );
and \U$6190 ( \8075 , RI2b5e785f3f40_218, \7830 );
and \U$6191 ( \8076 , RI2b5e785eb318_231, \7832 );
and \U$6192 ( \8077 , RI2b5e785da4a0_244, \7834 );
or \U$6193 ( \8078 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 );
_DC g1161 ( \8079_nG1161 , \8078 , \7853 );
buf \U$6194 ( \8080 , \8079_nG1161 );
and \U$6195 ( \8081 , \8060 , \8080 );
xor \U$6196 ( \8082 , \7783 , \7787 );
buf \U$6197 ( \8083 , \8082 );
buf \U$6198 ( \8084 , \8083 );
not \U$6199 ( \8085 , \8084 );
and \U$6200 ( \8086 , RI2b5e78549720_37, \7802 );
and \U$6201 ( \8087 , RI2b5e78538a88_50, \7804 );
and \U$6202 ( \8088 , RI2b5e78538470_63, \7806 );
and \U$6203 ( \8089 , RI2b5e784a5ef8_76, \7808 );
and \U$6204 ( \8090 , RI2b5e78495260_89, \7810 );
and \U$6205 ( \8091 , RI2b5e78403d60_102, \7812 );
and \U$6206 ( \8092 , RI2b5e775b2040_115, \7814 );
and \U$6207 ( \8093 , RI2b5e775b1a28_128, \7816 );
and \U$6208 ( \8094 , RI2b5e7750b9c0_141, \7818 );
and \U$6209 ( \8095 , RI2b5e774ff198_154, \7820 );
and \U$6210 ( \8096 , RI2b5e774f61b0_167, \7822 );
and \U$6211 ( \8097 , RI2b5e774ea798_180, \7824 );
and \U$6212 ( \8098 , RI2b5e774ddf70_193, \7826 );
and \U$6213 ( \8099 , RI2b5e774d4f88_206, \7828 );
and \U$6214 ( \8100 , RI2b5e785f3ec8_219, \7830 );
and \U$6215 ( \8101 , RI2b5e785eb2a0_232, \7832 );
and \U$6216 ( \8102 , RI2b5e785da428_245, \7834 );
or \U$6217 ( \8103 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 );
_DC g117a ( \8104_nG117a , \8103 , \7853 );
buf \U$6218 ( \8105 , \8104_nG117a );
and \U$6219 ( \8106 , \8085 , \8105 );
xor \U$6220 ( \8107 , \7784 , \7786 );
buf \U$6221 ( \8108 , \8107 );
buf \U$6222 ( \8109 , \8108 );
not \U$6223 ( \8110 , \8109 );
and \U$6224 ( \8111 , RI2b5e785496a8_38, \7802 );
and \U$6225 ( \8112 , RI2b5e78538a10_51, \7804 );
and \U$6226 ( \8113 , RI2b5e785383f8_64, \7806 );
and \U$6227 ( \8114 , RI2b5e784a5e80_77, \7808 );
and \U$6228 ( \8115 , RI2b5e784951e8_90, \7810 );
and \U$6229 ( \8116 , RI2b5e78403ce8_103, \7812 );
and \U$6230 ( \8117 , RI2b5e775b1fc8_116, \7814 );
and \U$6231 ( \8118 , RI2b5e775b19b0_129, \7816 );
and \U$6232 ( \8119 , RI2b5e7750b948_142, \7818 );
and \U$6233 ( \8120 , RI2b5e774ff120_155, \7820 );
and \U$6234 ( \8121 , RI2b5e774f6138_168, \7822 );
and \U$6235 ( \8122 , RI2b5e774ea720_181, \7824 );
and \U$6236 ( \8123 , RI2b5e774ddef8_194, \7826 );
and \U$6237 ( \8124 , RI2b5e774d4f10_207, \7828 );
and \U$6238 ( \8125 , RI2b5e785f3e50_220, \7830 );
and \U$6239 ( \8126 , RI2b5e785eb228_233, \7832 );
and \U$6240 ( \8127 , RI2b5e785da3b0_246, \7834 );
or \U$6241 ( \8128 , \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 );
_DC g1193 ( \8129_nG1193 , \8128 , \7853 );
buf \U$6242 ( \8130 , \8129_nG1193 );
and \U$6243 ( \8131 , \8110 , \8130 );
buf \U$6244 ( \8132 , RI2b5e785db148_13);
buf \U$6247 ( \8133 , \8132 );
not \U$6248 ( \8134 , \8133 );
and \U$6249 ( \8135 , RI2b5e78549630_39, \7802 );
and \U$6250 ( \8136 , RI2b5e78538998_52, \7804 );
and \U$6251 ( \8137 , RI2b5e78538380_65, \7806 );
and \U$6252 ( \8138 , RI2b5e784a5e08_78, \7808 );
and \U$6253 ( \8139 , RI2b5e78495170_91, \7810 );
and \U$6254 ( \8140 , RI2b5e78403c70_104, \7812 );
and \U$6255 ( \8141 , RI2b5e775b1f50_117, \7814 );
and \U$6256 ( \8142 , RI2b5e775b1938_130, \7816 );
and \U$6257 ( \8143 , RI2b5e7750b8d0_143, \7818 );
and \U$6258 ( \8144 , RI2b5e774ff0a8_156, \7820 );
and \U$6259 ( \8145 , RI2b5e774f60c0_169, \7822 );
and \U$6260 ( \8146 , RI2b5e774ea6a8_182, \7824 );
and \U$6261 ( \8147 , RI2b5e774dde80_195, \7826 );
and \U$6262 ( \8148 , RI2b5e774d4e98_208, \7828 );
and \U$6263 ( \8149 , RI2b5e785f3dd8_221, \7830 );
and \U$6264 ( \8150 , RI2b5e785eb1b0_234, \7832 );
and \U$6265 ( \8151 , RI2b5e785da338_247, \7834 );
or \U$6266 ( \8152 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 );
_DC g11ad ( \8153_nG11ad , \8152 , \7853 );
buf \U$6267 ( \8154 , \8153_nG11ad );
and \U$6268 ( \8155 , \8134 , \8154 );
xnor \U$6269 ( \8156 , \8109 , \8130 );
and \U$6270 ( \8157 , \8155 , \8156 );
or \U$6271 ( \8158 , \8131 , \8157 );
xnor \U$6272 ( \8159 , \8084 , \8105 );
and \U$6273 ( \8160 , \8158 , \8159 );
or \U$6274 ( \8161 , \8106 , \8160 );
xnor \U$6275 ( \8162 , \8059 , \8080 );
and \U$6276 ( \8163 , \8161 , \8162 );
or \U$6277 ( \8164 , \8081 , \8163 );
xnor \U$6278 ( \8165 , \8034 , \8055 );
and \U$6279 ( \8166 , \8164 , \8165 );
or \U$6280 ( \8167 , \8056 , \8166 );
xnor \U$6281 ( \8168 , \8009 , \8030 );
and \U$6282 ( \8169 , \8167 , \8168 );
or \U$6283 ( \8170 , \8031 , \8169 );
xnor \U$6284 ( \8171 , \7984 , \8005 );
and \U$6285 ( \8172 , \8170 , \8171 );
or \U$6286 ( \8173 , \8006 , \8172 );
xnor \U$6287 ( \8174 , \7959 , \7980 );
and \U$6288 ( \8175 , \8173 , \8174 );
or \U$6289 ( \8176 , \7981 , \8175 );
xnor \U$6290 ( \8177 , \7934 , \7955 );
and \U$6291 ( \8178 , \8176 , \8177 );
or \U$6292 ( \8179 , \7956 , \8178 );
xnor \U$6293 ( \8180 , \7909 , \7930 );
and \U$6294 ( \8181 , \8179 , \8180 );
or \U$6295 ( \8182 , \7931 , \8181 );
xnor \U$6296 ( \8183 , \7884 , \7905 );
and \U$6297 ( \8184 , \8182 , \8183 );
or \U$6298 ( \8185 , \7906 , \8184 );
xnor \U$6299 ( \8186 , \7859 , \7880 );
and \U$6300 ( \8187 , \8185 , \8186 );
or \U$6301 ( \8188 , \7881 , \8187 );
xnor \U$6302 ( \8189 , \7800 , \7855 );
and \U$6303 ( \8190 , \8188 , \8189 );
or \U$6304 ( \8191 , \7856 , \8190 );
not \U$6305 ( \8192 , \8191 );
buf \U$6306 ( \8193 , \8192 );
buf \U$6307 ( \8194 , RI2b5e785aeb98_596);
buf \U$6308 ( \8195 , RI2b5e785aec10_595);
buf \U$6309 ( \8196 , RI2b5e785aec88_594);
buf \U$6310 ( \8197 , RI2b5e785aed00_593);
buf \U$6311 ( \8198 , RI2b5e785aed78_592);
buf \U$6312 ( \8199 , RI2b5e785aedf0_591);
buf \U$6313 ( \8200 , RI2b5e785aee68_590);
buf \U$6314 ( \8201 , RI2b5e785aeee0_589);
buf \U$6315 ( \8202 , RI2b5e785aef58_588);
buf \U$6316 ( \8203 , RI2b5e785ae9b8_600);
buf \U$6317 ( \8204 , RI2b5e785aea30_599);
buf \U$6318 ( \8205 , RI2b5e785aeaa8_598);
buf \U$6319 ( \8206 , RI2b5e785aeb20_597);
and \U$6320 ( \8207 , \8203 , \8204 , \8205 , \8206 );
nor \U$6321 ( \8208 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8207 );
buf \U$6322 ( \8209 , \8208 );
and \U$6323 ( \8210 , \8193 , \8209 );
nor \U$6324 ( \8211 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 , RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6325 ( \8212 , RI2b5e785daab8_27, \8211 );
nor \U$6326 ( \8213 , \2175 , \2176 , \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6327 ( \8214 , RI2b5e785495b8_40, \8213 );
nor \U$6328 ( \8215 , RI2b5e785ae9b8_600, \2176 , \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6329 ( \8216 , RI2b5e78538920_53, \8215 );
nor \U$6330 ( \8217 , \2175 , RI2b5e785aea30_599, \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6331 ( \8218 , RI2b5e784a63a8_66, \8217 );
nor \U$6332 ( \8219 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2177 , \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6333 ( \8220 , RI2b5e78495710_79, \8219 );
nor \U$6334 ( \8221 , \2175 , \2176 , RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6335 ( \8222 , RI2b5e784950f8_92, \8221 );
nor \U$6336 ( \8223 , RI2b5e785ae9b8_600, \2176 , RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6337 ( \8224 , RI2b5e78403bf8_105, \8223 );
nor \U$6338 ( \8225 , \2175 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6339 ( \8226 , RI2b5e775b1ed8_118, \8225 );
nor \U$6340 ( \8227 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, \2178 , RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6341 ( \8228 , RI2b5e775b18c0_131, \8227 );
nor \U$6342 ( \8229 , \2175 , \2176 , \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6343 ( \8230 , RI2b5e7750b858_144, \8229 );
nor \U$6344 ( \8231 , RI2b5e785ae9b8_600, \2176 , \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6345 ( \8232 , RI2b5e774ff030_157, \8231 );
nor \U$6346 ( \8233 , \2175 , RI2b5e785aea30_599, \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6347 ( \8234 , RI2b5e774f6048_170, \8233 );
nor \U$6348 ( \8235 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2177 , RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6349 ( \8236 , RI2b5e774ea630_183, \8235 );
nor \U$6350 ( \8237 , \2175 , \2176 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6351 ( \8238 , RI2b5e774dde08_196, \8237 );
nor \U$6352 ( \8239 , RI2b5e785ae9b8_600, \2176 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6353 ( \8240 , RI2b5e774d4e20_209, \8239 );
nor \U$6354 ( \8241 , \2175 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6355 ( \8242 , RI2b5e785f3d60_222, \8241 );
nor \U$6356 ( \8243 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596, RI2b5e785aec10_595, RI2b5e785aec88_594, RI2b5e785aed00_593, RI2b5e785aed78_592, RI2b5e785aedf0_591, RI2b5e785aee68_590, RI2b5e785aeee0_589, RI2b5e785aef58_588);
and \U$6357 ( \8244 , RI2b5e785eb138_235, \8243 );
or \U$6358 ( \8245 , \8212 , \8214 , \8216 , \8218 , \8220 , \8222 , \8224 , \8226 , \8228 , \8230 , \8232 , \8234 , \8236 , \8238 , \8240 , \8242 , \8244 );
buf \U$6359 ( \8246 , RI2b5e785aec10_595);
buf \U$6360 ( \8247 , RI2b5e785aec88_594);
buf \U$6361 ( \8248 , RI2b5e785aed00_593);
buf \U$6362 ( \8249 , RI2b5e785aed78_592);
buf \U$6363 ( \8250 , RI2b5e785aedf0_591);
buf \U$6364 ( \8251 , RI2b5e785aee68_590);
buf \U$6365 ( \8252 , RI2b5e785aeee0_589);
buf \U$6366 ( \8253 , RI2b5e785aef58_588);
buf \U$6367 ( \8254 , RI2b5e785aeb98_596);
buf \U$6368 ( \8255 , RI2b5e785ae9b8_600);
buf \U$6369 ( \8256 , RI2b5e785aea30_599);
buf \U$6370 ( \8257 , RI2b5e785aeaa8_598);
buf \U$6371 ( \8258 , RI2b5e785aeb20_597);
or \U$6372 ( \8259 , \8255 , \8256 , \8257 , \8258 );
and \U$6373 ( \8260 , \8254 , \8259 );
or \U$6374 ( \8261 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8260 );
buf \U$6375 ( \8262 , \8261 );
_DC g1220 ( \8263_nG1220 , \8245 , \8262 );
buf \U$6376 ( \8264 , \8263_nG1220 );
not \U$6377 ( \8265 , \8264 );
nor \U$6378 ( \8266 , \4969 , \4973 , \4977 , \4981 , \4986 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6379 ( \8267 , RI2b5e785daab8_27, \8266 );
nor \U$6380 ( \8268 , \5021 , \5022 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6381 ( \8269 , RI2b5e785495b8_40, \8268 );
nor \U$6382 ( \8270 , \4969 , \5022 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6383 ( \8271 , RI2b5e78538920_53, \8270 );
nor \U$6384 ( \8272 , \5021 , \4973 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6385 ( \8273 , RI2b5e784a63a8_66, \8272 );
nor \U$6386 ( \8274 , \4969 , \4973 , \5023 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6387 ( \8275 , RI2b5e78495710_79, \8274 );
nor \U$6388 ( \8276 , \5021 , \5022 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6389 ( \8277 , RI2b5e784950f8_92, \8276 );
nor \U$6390 ( \8278 , \4969 , \5022 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6391 ( \8279 , RI2b5e78403bf8_105, \8278 );
nor \U$6392 ( \8280 , \5021 , \4973 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6393 ( \8281 , RI2b5e775b1ed8_118, \8280 );
nor \U$6394 ( \8282 , \4969 , \4973 , \4977 , \5024 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6395 ( \8283 , RI2b5e775b18c0_131, \8282 );
nor \U$6396 ( \8284 , \5021 , \5022 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6397 ( \8285 , RI2b5e7750b858_144, \8284 );
nor \U$6398 ( \8286 , \4969 , \5022 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6399 ( \8287 , RI2b5e774ff030_157, \8286 );
nor \U$6400 ( \8288 , \5021 , \4973 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6401 ( \8289 , RI2b5e774f6048_170, \8288 );
nor \U$6402 ( \8290 , \4969 , \4973 , \5023 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6403 ( \8291 , RI2b5e774ea630_183, \8290 );
nor \U$6404 ( \8292 , \5021 , \5022 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6405 ( \8293 , RI2b5e774dde08_196, \8292 );
nor \U$6406 ( \8294 , \4969 , \5022 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6407 ( \8295 , RI2b5e774d4e20_209, \8294 );
nor \U$6408 ( \8296 , \5021 , \4973 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6409 ( \8297 , RI2b5e785f3d60_222, \8296 );
nor \U$6410 ( \8298 , \4969 , \4973 , \4977 , \4981 , \4985 , \4990 , \4994 , \4998 , \5002 , \5006 , \5010 , \5014 , \5018 );
and \U$6411 ( \8299 , RI2b5e785eb138_235, \8298 );
or \U$6412 ( \8300 , \8267 , \8269 , \8271 , \8273 , \8275 , \8277 , \8279 , \8281 , \8283 , \8285 , \8287 , \8289 , \8291 , \8293 , \8295 , \8297 , \8299 );
buf \U$6413 ( \8301 , \4990 );
buf \U$6414 ( \8302 , \4994 );
buf \U$6415 ( \8303 , \4998 );
buf \U$6416 ( \8304 , \5002 );
buf \U$6417 ( \8305 , \5006 );
buf \U$6418 ( \8306 , \5010 );
buf \U$6419 ( \8307 , \5014 );
buf \U$6420 ( \8308 , \5018 );
buf \U$6421 ( \8309 , \4985 );
buf \U$6422 ( \8310 , \4969 );
buf \U$6423 ( \8311 , \4973 );
buf \U$6424 ( \8312 , \4977 );
buf \U$6425 ( \8313 , \4981 );
or \U$6426 ( \8314 , \8310 , \8311 , \8312 , \8313 );
and \U$6427 ( \8315 , \8309 , \8314 );
or \U$6428 ( \8316 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8315 );
buf \U$6429 ( \8317 , \8316 );
_DC g1257 ( \8318_nG1257 , \8300 , \8317 );
buf \U$6430 ( \8319 , \8318_nG1257 );
and \U$6431 ( \8320 , \8265 , \8319 );
and \U$6432 ( \8321 , RI2b5e785daa40_28, \8211 );
and \U$6433 ( \8322 , RI2b5e78549540_41, \8213 );
and \U$6434 ( \8323 , RI2b5e785388a8_54, \8215 );
and \U$6435 ( \8324 , RI2b5e784a6330_67, \8217 );
and \U$6436 ( \8325 , RI2b5e78495698_80, \8219 );
and \U$6437 ( \8326 , RI2b5e78495080_93, \8221 );
and \U$6438 ( \8327 , RI2b5e78403b80_106, \8223 );
and \U$6439 ( \8328 , RI2b5e775b1e60_119, \8225 );
and \U$6440 ( \8329 , RI2b5e7750bdf8_132, \8227 );
and \U$6441 ( \8330 , RI2b5e774ff5d0_145, \8229 );
and \U$6442 ( \8331 , RI2b5e774f65e8_158, \8231 );
and \U$6443 ( \8332 , RI2b5e774eabd0_171, \8233 );
and \U$6444 ( \8333 , RI2b5e774de3a8_184, \8235 );
and \U$6445 ( \8334 , RI2b5e774d53c0_197, \8237 );
and \U$6446 ( \8335 , RI2b5e785f4300_210, \8239 );
and \U$6447 ( \8336 , RI2b5e785f3ce8_223, \8241 );
and \U$6448 ( \8337 , RI2b5e785eb0c0_236, \8243 );
or \U$6449 ( \8338 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 );
_DC g126c ( \8339_nG126c , \8338 , \8262 );
buf \U$6450 ( \8340 , \8339_nG126c );
not \U$6451 ( \8341 , \8340 );
and \U$6452 ( \8342 , RI2b5e785daa40_28, \8266 );
and \U$6453 ( \8343 , RI2b5e78549540_41, \8268 );
and \U$6454 ( \8344 , RI2b5e785388a8_54, \8270 );
and \U$6455 ( \8345 , RI2b5e784a6330_67, \8272 );
and \U$6456 ( \8346 , RI2b5e78495698_80, \8274 );
and \U$6457 ( \8347 , RI2b5e78495080_93, \8276 );
and \U$6458 ( \8348 , RI2b5e78403b80_106, \8278 );
and \U$6459 ( \8349 , RI2b5e775b1e60_119, \8280 );
and \U$6460 ( \8350 , RI2b5e7750bdf8_132, \8282 );
and \U$6461 ( \8351 , RI2b5e774ff5d0_145, \8284 );
and \U$6462 ( \8352 , RI2b5e774f65e8_158, \8286 );
and \U$6463 ( \8353 , RI2b5e774eabd0_171, \8288 );
and \U$6464 ( \8354 , RI2b5e774de3a8_184, \8290 );
and \U$6465 ( \8355 , RI2b5e774d53c0_197, \8292 );
and \U$6466 ( \8356 , RI2b5e785f4300_210, \8294 );
and \U$6467 ( \8357 , RI2b5e785f3ce8_223, \8296 );
and \U$6468 ( \8358 , RI2b5e785eb0c0_236, \8298 );
or \U$6469 ( \8359 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 );
_DC g1281 ( \8360_nG1281 , \8359 , \8317 );
buf \U$6470 ( \8361 , \8360_nG1281 );
and \U$6471 ( \8362 , \8341 , \8361 );
and \U$6472 ( \8363 , RI2b5e785da9c8_29, \8211 );
and \U$6473 ( \8364 , RI2b5e785494c8_42, \8213 );
and \U$6474 ( \8365 , RI2b5e78538830_55, \8215 );
and \U$6475 ( \8366 , RI2b5e784a62b8_68, \8217 );
and \U$6476 ( \8367 , RI2b5e78495620_81, \8219 );
and \U$6477 ( \8368 , RI2b5e78495008_94, \8221 );
and \U$6478 ( \8369 , RI2b5e78403b08_107, \8223 );
and \U$6479 ( \8370 , RI2b5e775b1de8_120, \8225 );
and \U$6480 ( \8371 , RI2b5e7750bd80_133, \8227 );
and \U$6481 ( \8372 , RI2b5e774ff558_146, \8229 );
and \U$6482 ( \8373 , RI2b5e774f6570_159, \8231 );
and \U$6483 ( \8374 , RI2b5e774eab58_172, \8233 );
and \U$6484 ( \8375 , RI2b5e774de330_185, \8235 );
and \U$6485 ( \8376 , RI2b5e774d5348_198, \8237 );
and \U$6486 ( \8377 , RI2b5e785f4288_211, \8239 );
and \U$6487 ( \8378 , RI2b5e785f3658_224, \8241 );
and \U$6488 ( \8379 , RI2b5e785eb048_237, \8243 );
or \U$6489 ( \8380 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 );
_DC g1296 ( \8381_nG1296 , \8380 , \8262 );
buf \U$6490 ( \8382 , \8381_nG1296 );
not \U$6491 ( \8383 , \8382 );
and \U$6492 ( \8384 , RI2b5e785da9c8_29, \8266 );
and \U$6493 ( \8385 , RI2b5e785494c8_42, \8268 );
and \U$6494 ( \8386 , RI2b5e78538830_55, \8270 );
and \U$6495 ( \8387 , RI2b5e784a62b8_68, \8272 );
and \U$6496 ( \8388 , RI2b5e78495620_81, \8274 );
and \U$6497 ( \8389 , RI2b5e78495008_94, \8276 );
and \U$6498 ( \8390 , RI2b5e78403b08_107, \8278 );
and \U$6499 ( \8391 , RI2b5e775b1de8_120, \8280 );
and \U$6500 ( \8392 , RI2b5e7750bd80_133, \8282 );
and \U$6501 ( \8393 , RI2b5e774ff558_146, \8284 );
and \U$6502 ( \8394 , RI2b5e774f6570_159, \8286 );
and \U$6503 ( \8395 , RI2b5e774eab58_172, \8288 );
and \U$6504 ( \8396 , RI2b5e774de330_185, \8290 );
and \U$6505 ( \8397 , RI2b5e774d5348_198, \8292 );
and \U$6506 ( \8398 , RI2b5e785f4288_211, \8294 );
and \U$6507 ( \8399 , RI2b5e785f3658_224, \8296 );
and \U$6508 ( \8400 , RI2b5e785eb048_237, \8298 );
or \U$6509 ( \8401 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 );
_DC g12ab ( \8402_nG12ab , \8401 , \8317 );
buf \U$6510 ( \8403 , \8402_nG12ab );
and \U$6511 ( \8404 , \8383 , \8403 );
and \U$6512 ( \8405 , RI2b5e785da950_30, \8211 );
and \U$6513 ( \8406 , RI2b5e78549450_43, \8213 );
and \U$6514 ( \8407 , RI2b5e785387b8_56, \8215 );
and \U$6515 ( \8408 , RI2b5e784a6240_69, \8217 );
and \U$6516 ( \8409 , RI2b5e784955a8_82, \8219 );
and \U$6517 ( \8410 , RI2b5e78494f90_95, \8221 );
and \U$6518 ( \8411 , RI2b5e78403a90_108, \8223 );
and \U$6519 ( \8412 , RI2b5e775b1d70_121, \8225 );
and \U$6520 ( \8413 , RI2b5e7750bd08_134, \8227 );
and \U$6521 ( \8414 , RI2b5e774ff4e0_147, \8229 );
and \U$6522 ( \8415 , RI2b5e774f64f8_160, \8231 );
and \U$6523 ( \8416 , RI2b5e774eaae0_173, \8233 );
and \U$6524 ( \8417 , RI2b5e774de2b8_186, \8235 );
and \U$6525 ( \8418 , RI2b5e774d52d0_199, \8237 );
and \U$6526 ( \8419 , RI2b5e785f4210_212, \8239 );
and \U$6527 ( \8420 , RI2b5e785eb5e8_225, \8241 );
and \U$6528 ( \8421 , RI2b5e785e6c50_238, \8243 );
or \U$6529 ( \8422 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 );
_DC g12c0 ( \8423_nG12c0 , \8422 , \8262 );
buf \U$6530 ( \8424 , \8423_nG12c0 );
not \U$6531 ( \8425 , \8424 );
and \U$6532 ( \8426 , RI2b5e785da950_30, \8266 );
and \U$6533 ( \8427 , RI2b5e78549450_43, \8268 );
and \U$6534 ( \8428 , RI2b5e785387b8_56, \8270 );
and \U$6535 ( \8429 , RI2b5e784a6240_69, \8272 );
and \U$6536 ( \8430 , RI2b5e784955a8_82, \8274 );
and \U$6537 ( \8431 , RI2b5e78494f90_95, \8276 );
and \U$6538 ( \8432 , RI2b5e78403a90_108, \8278 );
and \U$6539 ( \8433 , RI2b5e775b1d70_121, \8280 );
and \U$6540 ( \8434 , RI2b5e7750bd08_134, \8282 );
and \U$6541 ( \8435 , RI2b5e774ff4e0_147, \8284 );
and \U$6542 ( \8436 , RI2b5e774f64f8_160, \8286 );
and \U$6543 ( \8437 , RI2b5e774eaae0_173, \8288 );
and \U$6544 ( \8438 , RI2b5e774de2b8_186, \8290 );
and \U$6545 ( \8439 , RI2b5e774d52d0_199, \8292 );
and \U$6546 ( \8440 , RI2b5e785f4210_212, \8294 );
and \U$6547 ( \8441 , RI2b5e785eb5e8_225, \8296 );
and \U$6548 ( \8442 , RI2b5e785e6c50_238, \8298 );
or \U$6549 ( \8443 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 );
_DC g12d5 ( \8444_nG12d5 , \8443 , \8317 );
buf \U$6550 ( \8445 , \8444_nG12d5 );
and \U$6551 ( \8446 , \8425 , \8445 );
and \U$6552 ( \8447 , RI2b5e785da8d8_31, \8211 );
and \U$6553 ( \8448 , RI2b5e785493d8_44, \8213 );
and \U$6554 ( \8449 , RI2b5e78538740_57, \8215 );
and \U$6555 ( \8450 , RI2b5e784a61c8_70, \8217 );
and \U$6556 ( \8451 , RI2b5e78495530_83, \8219 );
and \U$6557 ( \8452 , RI2b5e78494f18_96, \8221 );
and \U$6558 ( \8453 , RI2b5e78403a18_109, \8223 );
and \U$6559 ( \8454 , RI2b5e775b1cf8_122, \8225 );
and \U$6560 ( \8455 , RI2b5e7750bc90_135, \8227 );
and \U$6561 ( \8456 , RI2b5e774ff468_148, \8229 );
and \U$6562 ( \8457 , RI2b5e774f6480_161, \8231 );
and \U$6563 ( \8458 , RI2b5e774eaa68_174, \8233 );
and \U$6564 ( \8459 , RI2b5e774de240_187, \8235 );
and \U$6565 ( \8460 , RI2b5e774d5258_200, \8237 );
and \U$6566 ( \8461 , RI2b5e785f4198_213, \8239 );
and \U$6567 ( \8462 , RI2b5e785eb570_226, \8241 );
and \U$6568 ( \8463 , RI2b5e785e6bd8_239, \8243 );
or \U$6569 ( \8464 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 );
_DC g12ea ( \8465_nG12ea , \8464 , \8262 );
buf \U$6570 ( \8466 , \8465_nG12ea );
not \U$6571 ( \8467 , \8466 );
and \U$6572 ( \8468 , RI2b5e785da8d8_31, \8266 );
and \U$6573 ( \8469 , RI2b5e785493d8_44, \8268 );
and \U$6574 ( \8470 , RI2b5e78538740_57, \8270 );
and \U$6575 ( \8471 , RI2b5e784a61c8_70, \8272 );
and \U$6576 ( \8472 , RI2b5e78495530_83, \8274 );
and \U$6577 ( \8473 , RI2b5e78494f18_96, \8276 );
and \U$6578 ( \8474 , RI2b5e78403a18_109, \8278 );
and \U$6579 ( \8475 , RI2b5e775b1cf8_122, \8280 );
and \U$6580 ( \8476 , RI2b5e7750bc90_135, \8282 );
and \U$6581 ( \8477 , RI2b5e774ff468_148, \8284 );
and \U$6582 ( \8478 , RI2b5e774f6480_161, \8286 );
and \U$6583 ( \8479 , RI2b5e774eaa68_174, \8288 );
and \U$6584 ( \8480 , RI2b5e774de240_187, \8290 );
and \U$6585 ( \8481 , RI2b5e774d5258_200, \8292 );
and \U$6586 ( \8482 , RI2b5e785f4198_213, \8294 );
and \U$6587 ( \8483 , RI2b5e785eb570_226, \8296 );
and \U$6588 ( \8484 , RI2b5e785e6bd8_239, \8298 );
or \U$6589 ( \8485 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 );
_DC g12ff ( \8486_nG12ff , \8485 , \8317 );
buf \U$6590 ( \8487 , \8486_nG12ff );
and \U$6591 ( \8488 , \8467 , \8487 );
and \U$6592 ( \8489 , RI2b5e785da860_32, \8211 );
and \U$6593 ( \8490 , RI2b5e78549360_45, \8213 );
and \U$6594 ( \8491 , RI2b5e785386c8_58, \8215 );
and \U$6595 ( \8492 , RI2b5e784a6150_71, \8217 );
and \U$6596 ( \8493 , RI2b5e784954b8_84, \8219 );
and \U$6597 ( \8494 , RI2b5e78494ea0_97, \8221 );
and \U$6598 ( \8495 , RI2b5e784039a0_110, \8223 );
and \U$6599 ( \8496 , RI2b5e775b1c80_123, \8225 );
and \U$6600 ( \8497 , RI2b5e7750bc18_136, \8227 );
and \U$6601 ( \8498 , RI2b5e774ff3f0_149, \8229 );
and \U$6602 ( \8499 , RI2b5e774f6408_162, \8231 );
and \U$6603 ( \8500 , RI2b5e774ea9f0_175, \8233 );
and \U$6604 ( \8501 , RI2b5e774de1c8_188, \8235 );
and \U$6605 ( \8502 , RI2b5e774d51e0_201, \8237 );
and \U$6606 ( \8503 , RI2b5e785f4120_214, \8239 );
and \U$6607 ( \8504 , RI2b5e785eb4f8_227, \8241 );
and \U$6608 ( \8505 , RI2b5e785e64d0_240, \8243 );
or \U$6609 ( \8506 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 );
_DC g1314 ( \8507_nG1314 , \8506 , \8262 );
buf \U$6610 ( \8508 , \8507_nG1314 );
not \U$6611 ( \8509 , \8508 );
and \U$6612 ( \8510 , RI2b5e785da860_32, \8266 );
and \U$6613 ( \8511 , RI2b5e78549360_45, \8268 );
and \U$6614 ( \8512 , RI2b5e785386c8_58, \8270 );
and \U$6615 ( \8513 , RI2b5e784a6150_71, \8272 );
and \U$6616 ( \8514 , RI2b5e784954b8_84, \8274 );
and \U$6617 ( \8515 , RI2b5e78494ea0_97, \8276 );
and \U$6618 ( \8516 , RI2b5e784039a0_110, \8278 );
and \U$6619 ( \8517 , RI2b5e775b1c80_123, \8280 );
and \U$6620 ( \8518 , RI2b5e7750bc18_136, \8282 );
and \U$6621 ( \8519 , RI2b5e774ff3f0_149, \8284 );
and \U$6622 ( \8520 , RI2b5e774f6408_162, \8286 );
and \U$6623 ( \8521 , RI2b5e774ea9f0_175, \8288 );
and \U$6624 ( \8522 , RI2b5e774de1c8_188, \8290 );
and \U$6625 ( \8523 , RI2b5e774d51e0_201, \8292 );
and \U$6626 ( \8524 , RI2b5e785f4120_214, \8294 );
and \U$6627 ( \8525 , RI2b5e785eb4f8_227, \8296 );
and \U$6628 ( \8526 , RI2b5e785e64d0_240, \8298 );
or \U$6629 ( \8527 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 );
_DC g1329 ( \8528_nG1329 , \8527 , \8317 );
buf \U$6630 ( \8529 , \8528_nG1329 );
and \U$6631 ( \8530 , \8509 , \8529 );
and \U$6632 ( \8531 , RI2b5e78549900_33, \8211 );
and \U$6633 ( \8532 , RI2b5e78538c68_46, \8213 );
and \U$6634 ( \8533 , RI2b5e78538650_59, \8215 );
and \U$6635 ( \8534 , RI2b5e784a60d8_72, \8217 );
and \U$6636 ( \8535 , RI2b5e78495440_85, \8219 );
and \U$6637 ( \8536 , RI2b5e78494e28_98, \8221 );
and \U$6638 ( \8537 , RI2b5e78403928_111, \8223 );
and \U$6639 ( \8538 , RI2b5e775b1c08_124, \8225 );
and \U$6640 ( \8539 , RI2b5e7750bba0_137, \8227 );
and \U$6641 ( \8540 , RI2b5e774ff378_150, \8229 );
and \U$6642 ( \8541 , RI2b5e774f6390_163, \8231 );
and \U$6643 ( \8542 , RI2b5e774ea978_176, \8233 );
and \U$6644 ( \8543 , RI2b5e774de150_189, \8235 );
and \U$6645 ( \8544 , RI2b5e774d5168_202, \8237 );
and \U$6646 ( \8545 , RI2b5e785f40a8_215, \8239 );
and \U$6647 ( \8546 , RI2b5e785eb480_228, \8241 );
and \U$6648 ( \8547 , RI2b5e785da608_241, \8243 );
or \U$6649 ( \8548 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 );
_DC g133e ( \8549_nG133e , \8548 , \8262 );
buf \U$6650 ( \8550 , \8549_nG133e );
not \U$6651 ( \8551 , \8550 );
and \U$6652 ( \8552 , RI2b5e78549900_33, \8266 );
and \U$6653 ( \8553 , RI2b5e78538c68_46, \8268 );
and \U$6654 ( \8554 , RI2b5e78538650_59, \8270 );
and \U$6655 ( \8555 , RI2b5e784a60d8_72, \8272 );
and \U$6656 ( \8556 , RI2b5e78495440_85, \8274 );
and \U$6657 ( \8557 , RI2b5e78494e28_98, \8276 );
and \U$6658 ( \8558 , RI2b5e78403928_111, \8278 );
and \U$6659 ( \8559 , RI2b5e775b1c08_124, \8280 );
and \U$6660 ( \8560 , RI2b5e7750bba0_137, \8282 );
and \U$6661 ( \8561 , RI2b5e774ff378_150, \8284 );
and \U$6662 ( \8562 , RI2b5e774f6390_163, \8286 );
and \U$6663 ( \8563 , RI2b5e774ea978_176, \8288 );
and \U$6664 ( \8564 , RI2b5e774de150_189, \8290 );
and \U$6665 ( \8565 , RI2b5e774d5168_202, \8292 );
and \U$6666 ( \8566 , RI2b5e785f40a8_215, \8294 );
and \U$6667 ( \8567 , RI2b5e785eb480_228, \8296 );
and \U$6668 ( \8568 , RI2b5e785da608_241, \8298 );
or \U$6669 ( \8569 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 );
_DC g1353 ( \8570_nG1353 , \8569 , \8317 );
buf \U$6670 ( \8571 , \8570_nG1353 );
and \U$6671 ( \8572 , \8551 , \8571 );
and \U$6672 ( \8573 , RI2b5e78549888_34, \8211 );
and \U$6673 ( \8574 , RI2b5e78538bf0_47, \8213 );
and \U$6674 ( \8575 , RI2b5e785385d8_60, \8215 );
and \U$6675 ( \8576 , RI2b5e784a6060_73, \8217 );
and \U$6676 ( \8577 , RI2b5e784953c8_86, \8219 );
and \U$6677 ( \8578 , RI2b5e78403ec8_99, \8221 );
and \U$6678 ( \8579 , RI2b5e775b21a8_112, \8223 );
and \U$6679 ( \8580 , RI2b5e775b1b90_125, \8225 );
and \U$6680 ( \8581 , RI2b5e7750bb28_138, \8227 );
and \U$6681 ( \8582 , RI2b5e774ff300_151, \8229 );
and \U$6682 ( \8583 , RI2b5e774f6318_164, \8231 );
and \U$6683 ( \8584 , RI2b5e774ea900_177, \8233 );
and \U$6684 ( \8585 , RI2b5e774de0d8_190, \8235 );
and \U$6685 ( \8586 , RI2b5e774d50f0_203, \8237 );
and \U$6686 ( \8587 , RI2b5e785f4030_216, \8239 );
and \U$6687 ( \8588 , RI2b5e785eb408_229, \8241 );
and \U$6688 ( \8589 , RI2b5e785da590_242, \8243 );
or \U$6689 ( \8590 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 );
_DC g1368 ( \8591_nG1368 , \8590 , \8262 );
buf \U$6690 ( \8592 , \8591_nG1368 );
not \U$6691 ( \8593 , \8592 );
and \U$6692 ( \8594 , RI2b5e78549888_34, \8266 );
and \U$6693 ( \8595 , RI2b5e78538bf0_47, \8268 );
and \U$6694 ( \8596 , RI2b5e785385d8_60, \8270 );
and \U$6695 ( \8597 , RI2b5e784a6060_73, \8272 );
and \U$6696 ( \8598 , RI2b5e784953c8_86, \8274 );
and \U$6697 ( \8599 , RI2b5e78403ec8_99, \8276 );
and \U$6698 ( \8600 , RI2b5e775b21a8_112, \8278 );
and \U$6699 ( \8601 , RI2b5e775b1b90_125, \8280 );
and \U$6700 ( \8602 , RI2b5e7750bb28_138, \8282 );
and \U$6701 ( \8603 , RI2b5e774ff300_151, \8284 );
and \U$6702 ( \8604 , RI2b5e774f6318_164, \8286 );
and \U$6703 ( \8605 , RI2b5e774ea900_177, \8288 );
and \U$6704 ( \8606 , RI2b5e774de0d8_190, \8290 );
and \U$6705 ( \8607 , RI2b5e774d50f0_203, \8292 );
and \U$6706 ( \8608 , RI2b5e785f4030_216, \8294 );
and \U$6707 ( \8609 , RI2b5e785eb408_229, \8296 );
and \U$6708 ( \8610 , RI2b5e785da590_242, \8298 );
or \U$6709 ( \8611 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 );
_DC g137d ( \8612_nG137d , \8611 , \8317 );
buf \U$6710 ( \8613 , \8612_nG137d );
and \U$6711 ( \8614 , \8593 , \8613 );
and \U$6712 ( \8615 , RI2b5e78549810_35, \8211 );
and \U$6713 ( \8616 , RI2b5e78538b78_48, \8213 );
and \U$6714 ( \8617 , RI2b5e78538560_61, \8215 );
and \U$6715 ( \8618 , RI2b5e784a5fe8_74, \8217 );
and \U$6716 ( \8619 , RI2b5e78495350_87, \8219 );
and \U$6717 ( \8620 , RI2b5e78403e50_100, \8221 );
and \U$6718 ( \8621 , RI2b5e775b2130_113, \8223 );
and \U$6719 ( \8622 , RI2b5e775b1b18_126, \8225 );
and \U$6720 ( \8623 , RI2b5e7750bab0_139, \8227 );
and \U$6721 ( \8624 , RI2b5e774ff288_152, \8229 );
and \U$6722 ( \8625 , RI2b5e774f62a0_165, \8231 );
and \U$6723 ( \8626 , RI2b5e774ea888_178, \8233 );
and \U$6724 ( \8627 , RI2b5e774de060_191, \8235 );
and \U$6725 ( \8628 , RI2b5e774d5078_204, \8237 );
and \U$6726 ( \8629 , RI2b5e785f3fb8_217, \8239 );
and \U$6727 ( \8630 , RI2b5e785eb390_230, \8241 );
and \U$6728 ( \8631 , RI2b5e785da518_243, \8243 );
or \U$6729 ( \8632 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 );
_DC g1392 ( \8633_nG1392 , \8632 , \8262 );
buf \U$6730 ( \8634 , \8633_nG1392 );
not \U$6731 ( \8635 , \8634 );
and \U$6732 ( \8636 , RI2b5e78549810_35, \8266 );
and \U$6733 ( \8637 , RI2b5e78538b78_48, \8268 );
and \U$6734 ( \8638 , RI2b5e78538560_61, \8270 );
and \U$6735 ( \8639 , RI2b5e784a5fe8_74, \8272 );
and \U$6736 ( \8640 , RI2b5e78495350_87, \8274 );
and \U$6737 ( \8641 , RI2b5e78403e50_100, \8276 );
and \U$6738 ( \8642 , RI2b5e775b2130_113, \8278 );
and \U$6739 ( \8643 , RI2b5e775b1b18_126, \8280 );
and \U$6740 ( \8644 , RI2b5e7750bab0_139, \8282 );
and \U$6741 ( \8645 , RI2b5e774ff288_152, \8284 );
and \U$6742 ( \8646 , RI2b5e774f62a0_165, \8286 );
and \U$6743 ( \8647 , RI2b5e774ea888_178, \8288 );
and \U$6744 ( \8648 , RI2b5e774de060_191, \8290 );
and \U$6745 ( \8649 , RI2b5e774d5078_204, \8292 );
and \U$6746 ( \8650 , RI2b5e785f3fb8_217, \8294 );
and \U$6747 ( \8651 , RI2b5e785eb390_230, \8296 );
and \U$6748 ( \8652 , RI2b5e785da518_243, \8298 );
or \U$6749 ( \8653 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 );
_DC g13a7 ( \8654_nG13a7 , \8653 , \8317 );
buf \U$6750 ( \8655 , \8654_nG13a7 );
and \U$6751 ( \8656 , \8635 , \8655 );
and \U$6752 ( \8657 , RI2b5e78549798_36, \8211 );
and \U$6753 ( \8658 , RI2b5e78538b00_49, \8213 );
and \U$6754 ( \8659 , RI2b5e785384e8_62, \8215 );
and \U$6755 ( \8660 , RI2b5e784a5f70_75, \8217 );
and \U$6756 ( \8661 , RI2b5e784952d8_88, \8219 );
and \U$6757 ( \8662 , RI2b5e78403dd8_101, \8221 );
and \U$6758 ( \8663 , RI2b5e775b20b8_114, \8223 );
and \U$6759 ( \8664 , RI2b5e775b1aa0_127, \8225 );
and \U$6760 ( \8665 , RI2b5e7750ba38_140, \8227 );
and \U$6761 ( \8666 , RI2b5e774ff210_153, \8229 );
and \U$6762 ( \8667 , RI2b5e774f6228_166, \8231 );
and \U$6763 ( \8668 , RI2b5e774ea810_179, \8233 );
and \U$6764 ( \8669 , RI2b5e774ddfe8_192, \8235 );
and \U$6765 ( \8670 , RI2b5e774d5000_205, \8237 );
and \U$6766 ( \8671 , RI2b5e785f3f40_218, \8239 );
and \U$6767 ( \8672 , RI2b5e785eb318_231, \8241 );
and \U$6768 ( \8673 , RI2b5e785da4a0_244, \8243 );
or \U$6769 ( \8674 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 );
_DC g13bc ( \8675_nG13bc , \8674 , \8262 );
buf \U$6770 ( \8676 , \8675_nG13bc );
not \U$6771 ( \8677 , \8676 );
and \U$6772 ( \8678 , RI2b5e78549798_36, \8266 );
and \U$6773 ( \8679 , RI2b5e78538b00_49, \8268 );
and \U$6774 ( \8680 , RI2b5e785384e8_62, \8270 );
and \U$6775 ( \8681 , RI2b5e784a5f70_75, \8272 );
and \U$6776 ( \8682 , RI2b5e784952d8_88, \8274 );
and \U$6777 ( \8683 , RI2b5e78403dd8_101, \8276 );
and \U$6778 ( \8684 , RI2b5e775b20b8_114, \8278 );
and \U$6779 ( \8685 , RI2b5e775b1aa0_127, \8280 );
and \U$6780 ( \8686 , RI2b5e7750ba38_140, \8282 );
and \U$6781 ( \8687 , RI2b5e774ff210_153, \8284 );
and \U$6782 ( \8688 , RI2b5e774f6228_166, \8286 );
and \U$6783 ( \8689 , RI2b5e774ea810_179, \8288 );
and \U$6784 ( \8690 , RI2b5e774ddfe8_192, \8290 );
and \U$6785 ( \8691 , RI2b5e774d5000_205, \8292 );
and \U$6786 ( \8692 , RI2b5e785f3f40_218, \8294 );
and \U$6787 ( \8693 , RI2b5e785eb318_231, \8296 );
and \U$6788 ( \8694 , RI2b5e785da4a0_244, \8298 );
or \U$6789 ( \8695 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 );
_DC g13d1 ( \8696_nG13d1 , \8695 , \8317 );
buf \U$6790 ( \8697 , \8696_nG13d1 );
and \U$6791 ( \8698 , \8677 , \8697 );
and \U$6792 ( \8699 , RI2b5e78549720_37, \8211 );
and \U$6793 ( \8700 , RI2b5e78538a88_50, \8213 );
and \U$6794 ( \8701 , RI2b5e78538470_63, \8215 );
and \U$6795 ( \8702 , RI2b5e784a5ef8_76, \8217 );
and \U$6796 ( \8703 , RI2b5e78495260_89, \8219 );
and \U$6797 ( \8704 , RI2b5e78403d60_102, \8221 );
and \U$6798 ( \8705 , RI2b5e775b2040_115, \8223 );
and \U$6799 ( \8706 , RI2b5e775b1a28_128, \8225 );
and \U$6800 ( \8707 , RI2b5e7750b9c0_141, \8227 );
and \U$6801 ( \8708 , RI2b5e774ff198_154, \8229 );
and \U$6802 ( \8709 , RI2b5e774f61b0_167, \8231 );
and \U$6803 ( \8710 , RI2b5e774ea798_180, \8233 );
and \U$6804 ( \8711 , RI2b5e774ddf70_193, \8235 );
and \U$6805 ( \8712 , RI2b5e774d4f88_206, \8237 );
and \U$6806 ( \8713 , RI2b5e785f3ec8_219, \8239 );
and \U$6807 ( \8714 , RI2b5e785eb2a0_232, \8241 );
and \U$6808 ( \8715 , RI2b5e785da428_245, \8243 );
or \U$6809 ( \8716 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 );
_DC g13e6 ( \8717_nG13e6 , \8716 , \8262 );
buf \U$6810 ( \8718 , \8717_nG13e6 );
not \U$6811 ( \8719 , \8718 );
and \U$6812 ( \8720 , RI2b5e78549720_37, \8266 );
and \U$6813 ( \8721 , RI2b5e78538a88_50, \8268 );
and \U$6814 ( \8722 , RI2b5e78538470_63, \8270 );
and \U$6815 ( \8723 , RI2b5e784a5ef8_76, \8272 );
and \U$6816 ( \8724 , RI2b5e78495260_89, \8274 );
and \U$6817 ( \8725 , RI2b5e78403d60_102, \8276 );
and \U$6818 ( \8726 , RI2b5e775b2040_115, \8278 );
and \U$6819 ( \8727 , RI2b5e775b1a28_128, \8280 );
and \U$6820 ( \8728 , RI2b5e7750b9c0_141, \8282 );
and \U$6821 ( \8729 , RI2b5e774ff198_154, \8284 );
and \U$6822 ( \8730 , RI2b5e774f61b0_167, \8286 );
and \U$6823 ( \8731 , RI2b5e774ea798_180, \8288 );
and \U$6824 ( \8732 , RI2b5e774ddf70_193, \8290 );
and \U$6825 ( \8733 , RI2b5e774d4f88_206, \8292 );
and \U$6826 ( \8734 , RI2b5e785f3ec8_219, \8294 );
and \U$6827 ( \8735 , RI2b5e785eb2a0_232, \8296 );
and \U$6828 ( \8736 , RI2b5e785da428_245, \8298 );
or \U$6829 ( \8737 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 );
_DC g13fb ( \8738_nG13fb , \8737 , \8317 );
buf \U$6830 ( \8739 , \8738_nG13fb );
and \U$6831 ( \8740 , \8719 , \8739 );
and \U$6832 ( \8741 , RI2b5e785496a8_38, \8211 );
and \U$6833 ( \8742 , RI2b5e78538a10_51, \8213 );
and \U$6834 ( \8743 , RI2b5e785383f8_64, \8215 );
and \U$6835 ( \8744 , RI2b5e784a5e80_77, \8217 );
and \U$6836 ( \8745 , RI2b5e784951e8_90, \8219 );
and \U$6837 ( \8746 , RI2b5e78403ce8_103, \8221 );
and \U$6838 ( \8747 , RI2b5e775b1fc8_116, \8223 );
and \U$6839 ( \8748 , RI2b5e775b19b0_129, \8225 );
and \U$6840 ( \8749 , RI2b5e7750b948_142, \8227 );
and \U$6841 ( \8750 , RI2b5e774ff120_155, \8229 );
and \U$6842 ( \8751 , RI2b5e774f6138_168, \8231 );
and \U$6843 ( \8752 , RI2b5e774ea720_181, \8233 );
and \U$6844 ( \8753 , RI2b5e774ddef8_194, \8235 );
and \U$6845 ( \8754 , RI2b5e774d4f10_207, \8237 );
and \U$6846 ( \8755 , RI2b5e785f3e50_220, \8239 );
and \U$6847 ( \8756 , RI2b5e785eb228_233, \8241 );
and \U$6848 ( \8757 , RI2b5e785da3b0_246, \8243 );
or \U$6849 ( \8758 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 );
_DC g1410 ( \8759_nG1410 , \8758 , \8262 );
buf \U$6850 ( \8760 , \8759_nG1410 );
not \U$6851 ( \8761 , \8760 );
and \U$6852 ( \8762 , RI2b5e785496a8_38, \8266 );
and \U$6853 ( \8763 , RI2b5e78538a10_51, \8268 );
and \U$6854 ( \8764 , RI2b5e785383f8_64, \8270 );
and \U$6855 ( \8765 , RI2b5e784a5e80_77, \8272 );
and \U$6856 ( \8766 , RI2b5e784951e8_90, \8274 );
and \U$6857 ( \8767 , RI2b5e78403ce8_103, \8276 );
and \U$6858 ( \8768 , RI2b5e775b1fc8_116, \8278 );
and \U$6859 ( \8769 , RI2b5e775b19b0_129, \8280 );
and \U$6860 ( \8770 , RI2b5e7750b948_142, \8282 );
and \U$6861 ( \8771 , RI2b5e774ff120_155, \8284 );
and \U$6862 ( \8772 , RI2b5e774f6138_168, \8286 );
and \U$6863 ( \8773 , RI2b5e774ea720_181, \8288 );
and \U$6864 ( \8774 , RI2b5e774ddef8_194, \8290 );
and \U$6865 ( \8775 , RI2b5e774d4f10_207, \8292 );
and \U$6866 ( \8776 , RI2b5e785f3e50_220, \8294 );
and \U$6867 ( \8777 , RI2b5e785eb228_233, \8296 );
and \U$6868 ( \8778 , RI2b5e785da3b0_246, \8298 );
or \U$6869 ( \8779 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 );
_DC g1425 ( \8780_nG1425 , \8779 , \8317 );
buf \U$6870 ( \8781 , \8780_nG1425 );
and \U$6871 ( \8782 , \8761 , \8781 );
and \U$6872 ( \8783 , RI2b5e78549630_39, \8211 );
and \U$6873 ( \8784 , RI2b5e78538998_52, \8213 );
and \U$6874 ( \8785 , RI2b5e78538380_65, \8215 );
and \U$6875 ( \8786 , RI2b5e784a5e08_78, \8217 );
and \U$6876 ( \8787 , RI2b5e78495170_91, \8219 );
and \U$6877 ( \8788 , RI2b5e78403c70_104, \8221 );
and \U$6878 ( \8789 , RI2b5e775b1f50_117, \8223 );
and \U$6879 ( \8790 , RI2b5e775b1938_130, \8225 );
and \U$6880 ( \8791 , RI2b5e7750b8d0_143, \8227 );
and \U$6881 ( \8792 , RI2b5e774ff0a8_156, \8229 );
and \U$6882 ( \8793 , RI2b5e774f60c0_169, \8231 );
and \U$6883 ( \8794 , RI2b5e774ea6a8_182, \8233 );
and \U$6884 ( \8795 , RI2b5e774dde80_195, \8235 );
and \U$6885 ( \8796 , RI2b5e774d4e98_208, \8237 );
and \U$6886 ( \8797 , RI2b5e785f3dd8_221, \8239 );
and \U$6887 ( \8798 , RI2b5e785eb1b0_234, \8241 );
and \U$6888 ( \8799 , RI2b5e785da338_247, \8243 );
or \U$6889 ( \8800 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 );
_DC g143a ( \8801_nG143a , \8800 , \8262 );
buf \U$6890 ( \8802 , \8801_nG143a );
not \U$6891 ( \8803 , \8802 );
and \U$6892 ( \8804 , RI2b5e78549630_39, \8266 );
and \U$6893 ( \8805 , RI2b5e78538998_52, \8268 );
and \U$6894 ( \8806 , RI2b5e78538380_65, \8270 );
and \U$6895 ( \8807 , RI2b5e784a5e08_78, \8272 );
and \U$6896 ( \8808 , RI2b5e78495170_91, \8274 );
and \U$6897 ( \8809 , RI2b5e78403c70_104, \8276 );
and \U$6898 ( \8810 , RI2b5e775b1f50_117, \8278 );
and \U$6899 ( \8811 , RI2b5e775b1938_130, \8280 );
and \U$6900 ( \8812 , RI2b5e7750b8d0_143, \8282 );
and \U$6901 ( \8813 , RI2b5e774ff0a8_156, \8284 );
and \U$6902 ( \8814 , RI2b5e774f60c0_169, \8286 );
and \U$6903 ( \8815 , RI2b5e774ea6a8_182, \8288 );
and \U$6904 ( \8816 , RI2b5e774dde80_195, \8290 );
and \U$6905 ( \8817 , RI2b5e774d4e98_208, \8292 );
and \U$6906 ( \8818 , RI2b5e785f3dd8_221, \8294 );
and \U$6907 ( \8819 , RI2b5e785eb1b0_234, \8296 );
and \U$6908 ( \8820 , RI2b5e785da338_247, \8298 );
or \U$6909 ( \8821 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 );
_DC g144f ( \8822_nG144f , \8821 , \8317 );
buf \U$6910 ( \8823 , \8822_nG144f );
and \U$6911 ( \8824 , \8803 , \8823 );
xnor \U$6912 ( \8825 , \8781 , \8760 );
and \U$6913 ( \8826 , \8824 , \8825 );
or \U$6914 ( \8827 , \8782 , \8826 );
xnor \U$6915 ( \8828 , \8739 , \8718 );
and \U$6916 ( \8829 , \8827 , \8828 );
or \U$6917 ( \8830 , \8740 , \8829 );
xnor \U$6918 ( \8831 , \8697 , \8676 );
and \U$6919 ( \8832 , \8830 , \8831 );
or \U$6920 ( \8833 , \8698 , \8832 );
xnor \U$6921 ( \8834 , \8655 , \8634 );
and \U$6922 ( \8835 , \8833 , \8834 );
or \U$6923 ( \8836 , \8656 , \8835 );
xnor \U$6924 ( \8837 , \8613 , \8592 );
and \U$6925 ( \8838 , \8836 , \8837 );
or \U$6926 ( \8839 , \8614 , \8838 );
xnor \U$6927 ( \8840 , \8571 , \8550 );
and \U$6928 ( \8841 , \8839 , \8840 );
or \U$6929 ( \8842 , \8572 , \8841 );
xnor \U$6930 ( \8843 , \8529 , \8508 );
and \U$6931 ( \8844 , \8842 , \8843 );
or \U$6932 ( \8845 , \8530 , \8844 );
xnor \U$6933 ( \8846 , \8487 , \8466 );
and \U$6934 ( \8847 , \8845 , \8846 );
or \U$6935 ( \8848 , \8488 , \8847 );
xnor \U$6936 ( \8849 , \8445 , \8424 );
and \U$6937 ( \8850 , \8848 , \8849 );
or \U$6938 ( \8851 , \8446 , \8850 );
xnor \U$6939 ( \8852 , \8403 , \8382 );
and \U$6940 ( \8853 , \8851 , \8852 );
or \U$6941 ( \8854 , \8404 , \8853 );
xnor \U$6942 ( \8855 , \8361 , \8340 );
and \U$6943 ( \8856 , \8854 , \8855 );
or \U$6944 ( \8857 , \8362 , \8856 );
xnor \U$6945 ( \8858 , \8319 , \8264 );
and \U$6946 ( \8859 , \8857 , \8858 );
or \U$6947 ( \8860 , \8320 , \8859 );
buf \U$6948 ( \8861 , \8860 );
and \U$6949 ( \8862 , \8210 , \8861 );
_HMUX g32b3_GF_PartitionCandidate ( \8863_nG32b3 , \4926_nG3284 , \7772_nG32b2 , \8862 );
buf \U$6950 ( \8864 , \8863_nG32b3 );
not \U$6951 ( \8865 , \4389 );
nand \U$6952 ( \8866 , \4918 , \8865 );
nor \U$6953 ( \8867 , \4736 , \3572 );
nor \U$6954 ( \8868 , \3647 , \3724 );
nand \U$6955 ( \8869 , \8867 , \8868 );
nor \U$6956 ( \8870 , \3799 , \3876 );
nor \U$6957 ( \8871 , \3952 , \4025 );
nand \U$6958 ( \8872 , \8870 , \8871 );
nor \U$6959 ( \8873 , \8869 , \8872 );
nor \U$6960 ( \8874 , \4094 , \4158 );
nor \U$6961 ( \8875 , \4218 , \4275 );
nand \U$6962 ( \8876 , \8874 , \8875 );
nor \U$6963 ( \8877 , \4313 , \4345 );
nor \U$6964 ( \8878 , \4366 , \4382 );
nand \U$6965 ( \8879 , \8877 , \8878 );
nor \U$6966 ( \8880 , \8876 , \8879 );
nand \U$6967 ( \8881 , \8873 , \8880 );
nor \U$6968 ( \8882 , \4797 , \4501 );
nor \U$6969 ( \8883 , \4546 , \4598 );
nand \U$6970 ( \8884 , \8882 , \8883 );
nor \U$6971 ( \8885 , \4653 , \4692 );
nor \U$6972 ( \8886 , \4713 , \4729 );
nand \U$6973 ( \8887 , \8885 , \8886 );
nor \U$6974 ( \8888 , \8884 , \8887 );
nor \U$6975 ( \8889 , \4817 , \4772 );
nor \U$6976 ( \8890 , \4783 , \4794 );
nand \U$6977 ( \8891 , \8889 , \8890 );
nor \U$6978 ( \8892 , \4822 , \4814 );
not \U$6979 ( \8893 , \4830 );
and \U$6980 ( \8894 , \8892 , \8893 );
or \U$6981 ( \8895 , \4814 , \4832 );
nand \U$6982 ( \8896 , \8895 , \4835 );
nor \U$6983 ( \8897 , \8894 , \8896 );
or \U$6984 ( \8898 , \8891 , \8897 );
or \U$6985 ( \8899 , \4772 , \4837 );
nand \U$6986 ( \8900 , \8899 , \4841 );
and \U$6987 ( \8901 , \8890 , \8900 );
or \U$6988 ( \8902 , \4794 , \4843 );
nand \U$6989 ( \8903 , \8902 , \4846 );
nor \U$6990 ( \8904 , \8901 , \8903 );
nand \U$6991 ( \8905 , \8898 , \8904 );
and \U$6992 ( \8906 , \8888 , \8905 );
or \U$6993 ( \8907 , \4501 , \4848 );
nand \U$6994 ( \8908 , \8907 , \4853 );
and \U$6995 ( \8909 , \8883 , \8908 );
or \U$6996 ( \8910 , \4598 , \4855 );
nand \U$6997 ( \8911 , \8910 , \4858 );
nor \U$6998 ( \8912 , \8909 , \8911 );
or \U$6999 ( \8913 , \8887 , \8912 );
or \U$7000 ( \8914 , \4692 , \4860 );
nand \U$7001 ( \8915 , \8914 , \4864 );
and \U$7002 ( \8916 , \8886 , \8915 );
or \U$7003 ( \8917 , \4729 , \4866 );
nand \U$7004 ( \8918 , \8917 , \4869 );
nor \U$7005 ( \8919 , \8916 , \8918 );
nand \U$7006 ( \8920 , \8913 , \8919 );
nor \U$7007 ( \8921 , \8906 , \8920 );
or \U$7008 ( \8922 , \8881 , \8921 );
or \U$7009 ( \8923 , \3572 , \4871 );
nand \U$7010 ( \8924 , \8923 , \4877 );
and \U$7011 ( \8925 , \8868 , \8924 );
or \U$7012 ( \8926 , \3724 , \4879 );
nand \U$7013 ( \8927 , \8926 , \4882 );
nor \U$7014 ( \8928 , \8925 , \8927 );
or \U$7015 ( \8929 , \8872 , \8928 );
or \U$7016 ( \8930 , \3876 , \4884 );
nand \U$7017 ( \8931 , \8930 , \4888 );
and \U$7018 ( \8932 , \8871 , \8931 );
or \U$7019 ( \8933 , \4025 , \4890 );
nand \U$7020 ( \8934 , \8933 , \4893 );
nor \U$7021 ( \8935 , \8932 , \8934 );
nand \U$7022 ( \8936 , \8929 , \8935 );
and \U$7023 ( \8937 , \8880 , \8936 );
or \U$7024 ( \8938 , \4158 , \4895 );
nand \U$7025 ( \8939 , \8938 , \4900 );
and \U$7026 ( \8940 , \8875 , \8939 );
or \U$7027 ( \8941 , \4275 , \4902 );
nand \U$7028 ( \8942 , \8941 , \4905 );
nor \U$7029 ( \8943 , \8940 , \8942 );
or \U$7030 ( \8944 , \8879 , \8943 );
or \U$7031 ( \8945 , \4345 , \4907 );
nand \U$7032 ( \8946 , \8945 , \4911 );
and \U$7033 ( \8947 , \8878 , \8946 );
or \U$7034 ( \8948 , \4382 , \4913 );
nand \U$7035 ( \8949 , \8948 , \4916 );
nor \U$7036 ( \8950 , \8947 , \8949 );
nand \U$7037 ( \8951 , \8944 , \8950 );
nor \U$7038 ( \8952 , \8937 , \8951 );
nand \U$7039 ( \8953 , \8922 , \8952 );
not \U$7040 ( \8954 , \8953 );
xor \U$7041 ( \8955 , \8866 , \8954 );
buf g3221_GF_PartitionCandidate( \8956_nG3221 , \8955 );
not \U$7042 ( \8957 , \7235 );
nand \U$7043 ( \8958 , \7764 , \8957 );
nor \U$7044 ( \8959 , \7582 , \6418 );
nor \U$7045 ( \8960 , \6493 , \6570 );
nand \U$7046 ( \8961 , \8959 , \8960 );
nor \U$7047 ( \8962 , \6645 , \6722 );
nor \U$7048 ( \8963 , \6798 , \6871 );
nand \U$7049 ( \8964 , \8962 , \8963 );
nor \U$7050 ( \8965 , \8961 , \8964 );
nor \U$7051 ( \8966 , \6940 , \7004 );
nor \U$7052 ( \8967 , \7064 , \7121 );
nand \U$7053 ( \8968 , \8966 , \8967 );
nor \U$7054 ( \8969 , \7159 , \7191 );
nor \U$7055 ( \8970 , \7212 , \7228 );
nand \U$7056 ( \8971 , \8969 , \8970 );
nor \U$7057 ( \8972 , \8968 , \8971 );
nand \U$7058 ( \8973 , \8965 , \8972 );
nor \U$7059 ( \8974 , \7643 , \7347 );
nor \U$7060 ( \8975 , \7392 , \7444 );
nand \U$7061 ( \8976 , \8974 , \8975 );
nor \U$7062 ( \8977 , \7499 , \7538 );
nor \U$7063 ( \8978 , \7559 , \7575 );
nand \U$7064 ( \8979 , \8977 , \8978 );
nor \U$7065 ( \8980 , \8976 , \8979 );
nor \U$7066 ( \8981 , \7663 , \7618 );
nor \U$7067 ( \8982 , \7629 , \7640 );
nand \U$7068 ( \8983 , \8981 , \8982 );
nor \U$7069 ( \8984 , \7668 , \7660 );
not \U$7070 ( \8985 , \7676 );
and \U$7071 ( \8986 , \8984 , \8985 );
or \U$7072 ( \8987 , \7660 , \7678 );
nand \U$7073 ( \8988 , \8987 , \7681 );
nor \U$7074 ( \8989 , \8986 , \8988 );
or \U$7075 ( \8990 , \8983 , \8989 );
or \U$7076 ( \8991 , \7618 , \7683 );
nand \U$7077 ( \8992 , \8991 , \7687 );
and \U$7078 ( \8993 , \8982 , \8992 );
or \U$7079 ( \8994 , \7640 , \7689 );
nand \U$7080 ( \8995 , \8994 , \7692 );
nor \U$7081 ( \8996 , \8993 , \8995 );
nand \U$7082 ( \8997 , \8990 , \8996 );
and \U$7083 ( \8998 , \8980 , \8997 );
or \U$7084 ( \8999 , \7347 , \7694 );
nand \U$7085 ( \9000 , \8999 , \7699 );
and \U$7086 ( \9001 , \8975 , \9000 );
or \U$7087 ( \9002 , \7444 , \7701 );
nand \U$7088 ( \9003 , \9002 , \7704 );
nor \U$7089 ( \9004 , \9001 , \9003 );
or \U$7090 ( \9005 , \8979 , \9004 );
or \U$7091 ( \9006 , \7538 , \7706 );
nand \U$7092 ( \9007 , \9006 , \7710 );
and \U$7093 ( \9008 , \8978 , \9007 );
or \U$7094 ( \9009 , \7575 , \7712 );
nand \U$7095 ( \9010 , \9009 , \7715 );
nor \U$7096 ( \9011 , \9008 , \9010 );
nand \U$7097 ( \9012 , \9005 , \9011 );
nor \U$7098 ( \9013 , \8998 , \9012 );
or \U$7099 ( \9014 , \8973 , \9013 );
or \U$7100 ( \9015 , \6418 , \7717 );
nand \U$7101 ( \9016 , \9015 , \7723 );
and \U$7102 ( \9017 , \8960 , \9016 );
or \U$7103 ( \9018 , \6570 , \7725 );
nand \U$7104 ( \9019 , \9018 , \7728 );
nor \U$7105 ( \9020 , \9017 , \9019 );
or \U$7106 ( \9021 , \8964 , \9020 );
or \U$7107 ( \9022 , \6722 , \7730 );
nand \U$7108 ( \9023 , \9022 , \7734 );
and \U$7109 ( \9024 , \8963 , \9023 );
or \U$7110 ( \9025 , \6871 , \7736 );
nand \U$7111 ( \9026 , \9025 , \7739 );
nor \U$7112 ( \9027 , \9024 , \9026 );
nand \U$7113 ( \9028 , \9021 , \9027 );
and \U$7114 ( \9029 , \8972 , \9028 );
or \U$7115 ( \9030 , \7004 , \7741 );
nand \U$7116 ( \9031 , \9030 , \7746 );
and \U$7117 ( \9032 , \8967 , \9031 );
or \U$7118 ( \9033 , \7121 , \7748 );
nand \U$7119 ( \9034 , \9033 , \7751 );
nor \U$7120 ( \9035 , \9032 , \9034 );
or \U$7121 ( \9036 , \8971 , \9035 );
or \U$7122 ( \9037 , \7191 , \7753 );
nand \U$7123 ( \9038 , \9037 , \7757 );
and \U$7124 ( \9039 , \8970 , \9038 );
or \U$7125 ( \9040 , \7228 , \7759 );
nand \U$7126 ( \9041 , \9040 , \7762 );
nor \U$7127 ( \9042 , \9039 , \9041 );
nand \U$7128 ( \9043 , \9036 , \9042 );
nor \U$7129 ( \9044 , \9029 , \9043 );
nand \U$7130 ( \9045 , \9014 , \9044 );
not \U$7131 ( \9046 , \9045 );
xor \U$7132 ( \9047 , \8958 , \9046 );
buf g3255_GF_PartitionCandidate( \9048_nG3255 , \9047 );
_HMUX g3256_GF_PartitionCandidate ( \9049_nG3256 , \8956_nG3221 , \9048_nG3255 , \8862 );
buf \U$7133 ( \9050 , \9049_nG3256 );
not \U$7134 ( \9051 , \4382 );
nand \U$7135 ( \9052 , \4916 , \9051 );
nand \U$7136 ( \9053 , \4737 , \3648 );
nand \U$7137 ( \9054 , \3800 , \3953 );
nor \U$7138 ( \9055 , \9053 , \9054 );
nand \U$7139 ( \9056 , \4095 , \4219 );
nand \U$7140 ( \9057 , \4314 , \4367 );
nor \U$7141 ( \9058 , \9056 , \9057 );
nand \U$7142 ( \9059 , \9055 , \9058 );
nand \U$7143 ( \9060 , \4798 , \4547 );
nand \U$7144 ( \9061 , \4654 , \4714 );
nor \U$7145 ( \9062 , \9060 , \9061 );
nand \U$7146 ( \9063 , \4818 , \4784 );
not \U$7147 ( \9064 , \4833 );
or \U$7148 ( \9065 , \9063 , \9064 );
and \U$7149 ( \9066 , \4784 , \4838 );
nor \U$7150 ( \9067 , \9066 , \4844 );
nand \U$7151 ( \9068 , \9065 , \9067 );
and \U$7152 ( \9069 , \9062 , \9068 );
and \U$7153 ( \9070 , \4547 , \4849 );
nor \U$7154 ( \9071 , \9070 , \4856 );
or \U$7155 ( \9072 , \9061 , \9071 );
and \U$7156 ( \9073 , \4714 , \4861 );
nor \U$7157 ( \9074 , \9073 , \4867 );
nand \U$7158 ( \9075 , \9072 , \9074 );
nor \U$7159 ( \9076 , \9069 , \9075 );
or \U$7160 ( \9077 , \9059 , \9076 );
and \U$7161 ( \9078 , \3648 , \4872 );
nor \U$7162 ( \9079 , \9078 , \4880 );
or \U$7163 ( \9080 , \9054 , \9079 );
and \U$7164 ( \9081 , \3953 , \4885 );
nor \U$7165 ( \9082 , \9081 , \4891 );
nand \U$7166 ( \9083 , \9080 , \9082 );
and \U$7167 ( \9084 , \9058 , \9083 );
and \U$7168 ( \9085 , \4219 , \4896 );
nor \U$7169 ( \9086 , \9085 , \4903 );
or \U$7170 ( \9087 , \9057 , \9086 );
and \U$7171 ( \9088 , \4367 , \4908 );
nor \U$7172 ( \9089 , \9088 , \4914 );
nand \U$7173 ( \9090 , \9087 , \9089 );
nor \U$7174 ( \9091 , \9084 , \9090 );
nand \U$7175 ( \9092 , \9077 , \9091 );
not \U$7176 ( \9093 , \9092 );
xor \U$7177 ( \9094 , \9052 , \9093 );
buf g31b2_GF_PartitionCandidate( \9095_nG31b2 , \9094 );
not \U$7178 ( \9096 , \7228 );
nand \U$7179 ( \9097 , \7762 , \9096 );
nand \U$7180 ( \9098 , \7583 , \6494 );
nand \U$7181 ( \9099 , \6646 , \6799 );
nor \U$7182 ( \9100 , \9098 , \9099 );
nand \U$7183 ( \9101 , \6941 , \7065 );
nand \U$7184 ( \9102 , \7160 , \7213 );
nor \U$7185 ( \9103 , \9101 , \9102 );
nand \U$7186 ( \9104 , \9100 , \9103 );
nand \U$7187 ( \9105 , \7644 , \7393 );
nand \U$7188 ( \9106 , \7500 , \7560 );
nor \U$7189 ( \9107 , \9105 , \9106 );
nand \U$7190 ( \9108 , \7664 , \7630 );
not \U$7191 ( \9109 , \7679 );
or \U$7192 ( \9110 , \9108 , \9109 );
and \U$7193 ( \9111 , \7630 , \7684 );
nor \U$7194 ( \9112 , \9111 , \7690 );
nand \U$7195 ( \9113 , \9110 , \9112 );
and \U$7196 ( \9114 , \9107 , \9113 );
and \U$7197 ( \9115 , \7393 , \7695 );
nor \U$7198 ( \9116 , \9115 , \7702 );
or \U$7199 ( \9117 , \9106 , \9116 );
and \U$7200 ( \9118 , \7560 , \7707 );
nor \U$7201 ( \9119 , \9118 , \7713 );
nand \U$7202 ( \9120 , \9117 , \9119 );
nor \U$7203 ( \9121 , \9114 , \9120 );
or \U$7204 ( \9122 , \9104 , \9121 );
and \U$7205 ( \9123 , \6494 , \7718 );
nor \U$7206 ( \9124 , \9123 , \7726 );
or \U$7207 ( \9125 , \9099 , \9124 );
and \U$7208 ( \9126 , \6799 , \7731 );
nor \U$7209 ( \9127 , \9126 , \7737 );
nand \U$7210 ( \9128 , \9125 , \9127 );
and \U$7211 ( \9129 , \9103 , \9128 );
and \U$7212 ( \9130 , \7065 , \7742 );
nor \U$7213 ( \9131 , \9130 , \7749 );
or \U$7214 ( \9132 , \9102 , \9131 );
and \U$7215 ( \9133 , \7213 , \7754 );
nor \U$7216 ( \9134 , \9133 , \7760 );
nand \U$7217 ( \9135 , \9132 , \9134 );
nor \U$7218 ( \9136 , \9129 , \9135 );
nand \U$7219 ( \9137 , \9122 , \9136 );
not \U$7220 ( \9138 , \9137 );
xor \U$7221 ( \9139 , \9097 , \9138 );
buf g31ec_GF_PartitionCandidate( \9140_nG31ec , \9139 );
_HMUX g31ed_GF_PartitionCandidate ( \9141_nG31ed , \9095_nG31b2 , \9140_nG31ec , \8862 );
buf \U$7222 ( \9142 , \9141_nG31ed );
not \U$7223 ( \9143 , \4366 );
nand \U$7224 ( \9144 , \4913 , \9143 );
nand \U$7225 ( \9145 , \8886 , \8867 );
nand \U$7226 ( \9146 , \8868 , \8870 );
nor \U$7227 ( \9147 , \9145 , \9146 );
nand \U$7228 ( \9148 , \8871 , \8874 );
nand \U$7229 ( \9149 , \8875 , \8877 );
nor \U$7230 ( \9150 , \9148 , \9149 );
nand \U$7231 ( \9151 , \9147 , \9150 );
nand \U$7232 ( \9152 , \8890 , \8882 );
nand \U$7233 ( \9153 , \8883 , \8885 );
nor \U$7234 ( \9154 , \9152 , \9153 );
nand \U$7235 ( \9155 , \8892 , \8889 );
or \U$7236 ( \9156 , \9155 , \4830 );
and \U$7237 ( \9157 , \8889 , \8896 );
nor \U$7238 ( \9158 , \9157 , \8900 );
nand \U$7239 ( \9159 , \9156 , \9158 );
and \U$7240 ( \9160 , \9154 , \9159 );
and \U$7241 ( \9161 , \8882 , \8903 );
nor \U$7242 ( \9162 , \9161 , \8908 );
or \U$7243 ( \9163 , \9153 , \9162 );
and \U$7244 ( \9164 , \8885 , \8911 );
nor \U$7245 ( \9165 , \9164 , \8915 );
nand \U$7246 ( \9166 , \9163 , \9165 );
nor \U$7247 ( \9167 , \9160 , \9166 );
or \U$7248 ( \9168 , \9151 , \9167 );
and \U$7249 ( \9169 , \8867 , \8918 );
nor \U$7250 ( \9170 , \9169 , \8924 );
or \U$7251 ( \9171 , \9146 , \9170 );
and \U$7252 ( \9172 , \8870 , \8927 );
nor \U$7253 ( \9173 , \9172 , \8931 );
nand \U$7254 ( \9174 , \9171 , \9173 );
and \U$7255 ( \9175 , \9150 , \9174 );
and \U$7256 ( \9176 , \8874 , \8934 );
nor \U$7257 ( \9177 , \9176 , \8939 );
or \U$7258 ( \9178 , \9149 , \9177 );
and \U$7259 ( \9179 , \8877 , \8942 );
nor \U$7260 ( \9180 , \9179 , \8946 );
nand \U$7261 ( \9181 , \9178 , \9180 );
nor \U$7262 ( \9182 , \9175 , \9181 );
nand \U$7263 ( \9183 , \9168 , \9182 );
not \U$7264 ( \9184 , \9183 );
xor \U$7265 ( \9185 , \9144 , \9184 );
buf g3135_GF_PartitionCandidate( \9186_nG3135 , \9185 );
not \U$7266 ( \9187 , \7212 );
nand \U$7267 ( \9188 , \7759 , \9187 );
nand \U$7268 ( \9189 , \8978 , \8959 );
nand \U$7269 ( \9190 , \8960 , \8962 );
nor \U$7270 ( \9191 , \9189 , \9190 );
nand \U$7271 ( \9192 , \8963 , \8966 );
nand \U$7272 ( \9193 , \8967 , \8969 );
nor \U$7273 ( \9194 , \9192 , \9193 );
nand \U$7274 ( \9195 , \9191 , \9194 );
nand \U$7275 ( \9196 , \8982 , \8974 );
nand \U$7276 ( \9197 , \8975 , \8977 );
nor \U$7277 ( \9198 , \9196 , \9197 );
nand \U$7278 ( \9199 , \8984 , \8981 );
or \U$7279 ( \9200 , \9199 , \7676 );
and \U$7280 ( \9201 , \8981 , \8988 );
nor \U$7281 ( \9202 , \9201 , \8992 );
nand \U$7282 ( \9203 , \9200 , \9202 );
and \U$7283 ( \9204 , \9198 , \9203 );
and \U$7284 ( \9205 , \8974 , \8995 );
nor \U$7285 ( \9206 , \9205 , \9000 );
or \U$7286 ( \9207 , \9197 , \9206 );
and \U$7287 ( \9208 , \8977 , \9003 );
nor \U$7288 ( \9209 , \9208 , \9007 );
nand \U$7289 ( \9210 , \9207 , \9209 );
nor \U$7290 ( \9211 , \9204 , \9210 );
or \U$7291 ( \9212 , \9195 , \9211 );
and \U$7292 ( \9213 , \8959 , \9010 );
nor \U$7293 ( \9214 , \9213 , \9016 );
or \U$7294 ( \9215 , \9190 , \9214 );
and \U$7295 ( \9216 , \8962 , \9019 );
nor \U$7296 ( \9217 , \9216 , \9023 );
nand \U$7297 ( \9218 , \9215 , \9217 );
and \U$7298 ( \9219 , \9194 , \9218 );
and \U$7299 ( \9220 , \8966 , \9026 );
nor \U$7300 ( \9221 , \9220 , \9031 );
or \U$7301 ( \9222 , \9193 , \9221 );
and \U$7302 ( \9223 , \8969 , \9034 );
nor \U$7303 ( \9224 , \9223 , \9038 );
nand \U$7304 ( \9225 , \9222 , \9224 );
nor \U$7305 ( \9226 , \9219 , \9225 );
nand \U$7306 ( \9227 , \9212 , \9226 );
not \U$7307 ( \9228 , \9227 );
xor \U$7308 ( \9229 , \9188 , \9228 );
buf g3177_GF_PartitionCandidate( \9230_nG3177 , \9229 );
_HMUX g3178_GF_PartitionCandidate ( \9231_nG3178 , \9186_nG3135 , \9230_nG3177 , \8862 );
buf \U$7309 ( \9232 , \9231_nG3178 );
not \U$7310 ( \9233 , \4345 );
nand \U$7311 ( \9234 , \4911 , \9233 );
nor \U$7312 ( \9235 , \4738 , \3801 );
nor \U$7313 ( \9236 , \4096 , \4315 );
nand \U$7314 ( \9237 , \9235 , \9236 );
nor \U$7315 ( \9238 , \4799 , \4655 );
not \U$7316 ( \9239 , \4839 );
and \U$7317 ( \9240 , \9238 , \9239 );
or \U$7318 ( \9241 , \4655 , \4850 );
nand \U$7319 ( \9242 , \9241 , \4862 );
nor \U$7320 ( \9243 , \9240 , \9242 );
or \U$7321 ( \9244 , \9237 , \9243 );
or \U$7322 ( \9245 , \3801 , \4873 );
nand \U$7323 ( \9246 , \9245 , \4886 );
and \U$7324 ( \9247 , \9236 , \9246 );
or \U$7325 ( \9248 , \4315 , \4897 );
nand \U$7326 ( \9249 , \9248 , \4909 );
nor \U$7327 ( \9250 , \9247 , \9249 );
nand \U$7328 ( \9251 , \9244 , \9250 );
not \U$7329 ( \9252 , \9251 );
xor \U$7330 ( \9253 , \9234 , \9252 );
buf g30ac_GF_PartitionCandidate( \9254_nG30ac , \9253 );
not \U$7331 ( \9255 , \7191 );
nand \U$7332 ( \9256 , \7757 , \9255 );
nor \U$7333 ( \9257 , \7584 , \6647 );
nor \U$7334 ( \9258 , \6942 , \7161 );
nand \U$7335 ( \9259 , \9257 , \9258 );
nor \U$7336 ( \9260 , \7645 , \7501 );
not \U$7337 ( \9261 , \7685 );
and \U$7338 ( \9262 , \9260 , \9261 );
or \U$7339 ( \9263 , \7501 , \7696 );
nand \U$7340 ( \9264 , \9263 , \7708 );
nor \U$7341 ( \9265 , \9262 , \9264 );
or \U$7342 ( \9266 , \9259 , \9265 );
or \U$7343 ( \9267 , \6647 , \7719 );
nand \U$7344 ( \9268 , \9267 , \7732 );
and \U$7345 ( \9269 , \9258 , \9268 );
or \U$7346 ( \9270 , \7161 , \7743 );
nand \U$7347 ( \9271 , \9270 , \7755 );
nor \U$7348 ( \9272 , \9269 , \9271 );
nand \U$7349 ( \9273 , \9266 , \9272 );
not \U$7350 ( \9274 , \9273 );
xor \U$7351 ( \9275 , \9256 , \9274 );
buf g30f2_GF_PartitionCandidate( \9276_nG30f2 , \9275 );
_HMUX g30f3_GF_PartitionCandidate ( \9277_nG30f3 , \9254_nG30ac , \9276_nG30f2 , \8862 );
buf \U$7352 ( \9278 , \9277_nG30f3 );
not \U$7353 ( \9279 , \4313 );
nand \U$7354 ( \9280 , \4907 , \9279 );
nor \U$7355 ( \9281 , \8887 , \8869 );
nor \U$7356 ( \9282 , \8872 , \8876 );
nand \U$7357 ( \9283 , \9281 , \9282 );
nor \U$7358 ( \9284 , \8891 , \8884 );
not \U$7359 ( \9285 , \8897 );
and \U$7360 ( \9286 , \9284 , \9285 );
or \U$7361 ( \9287 , \8884 , \8904 );
nand \U$7362 ( \9288 , \9287 , \8912 );
nor \U$7363 ( \9289 , \9286 , \9288 );
or \U$7364 ( \9290 , \9283 , \9289 );
or \U$7365 ( \9291 , \8869 , \8919 );
nand \U$7366 ( \9292 , \9291 , \8928 );
and \U$7367 ( \9293 , \9282 , \9292 );
or \U$7368 ( \9294 , \8876 , \8935 );
nand \U$7369 ( \9295 , \9294 , \8943 );
nor \U$7370 ( \9296 , \9293 , \9295 );
nand \U$7371 ( \9297 , \9290 , \9296 );
not \U$7372 ( \9298 , \9297 );
xor \U$7373 ( \9299 , \9280 , \9298 );
buf g301d_GF_PartitionCandidate( \9300_nG301d , \9299 );
not \U$7374 ( \9301 , \7159 );
nand \U$7375 ( \9302 , \7753 , \9301 );
nor \U$7376 ( \9303 , \8979 , \8961 );
nor \U$7377 ( \9304 , \8964 , \8968 );
nand \U$7378 ( \9305 , \9303 , \9304 );
nor \U$7379 ( \9306 , \8983 , \8976 );
not \U$7380 ( \9307 , \8989 );
and \U$7381 ( \9308 , \9306 , \9307 );
or \U$7382 ( \9309 , \8976 , \8996 );
nand \U$7383 ( \9310 , \9309 , \9004 );
nor \U$7384 ( \9311 , \9308 , \9310 );
or \U$7385 ( \9312 , \9305 , \9311 );
or \U$7386 ( \9313 , \8961 , \9011 );
nand \U$7387 ( \9314 , \9313 , \9020 );
and \U$7388 ( \9315 , \9304 , \9314 );
or \U$7389 ( \9316 , \8968 , \9027 );
nand \U$7390 ( \9317 , \9316 , \9035 );
nor \U$7391 ( \9318 , \9315 , \9317 );
nand \U$7392 ( \9319 , \9312 , \9318 );
not \U$7393 ( \9320 , \9319 );
xor \U$7394 ( \9321 , \9302 , \9320 );
buf g3065_GF_PartitionCandidate( \9322_nG3065 , \9321 );
_HMUX g3066_GF_PartitionCandidate ( \9323_nG3066 , \9300_nG301d , \9322_nG3065 , \8862 );
buf \U$7395 ( \9324 , \9323_nG3066 );
not \U$7396 ( \9325 , \4275 );
nand \U$7397 ( \9326 , \4905 , \9325 );
nor \U$7398 ( \9327 , \9061 , \9053 );
nor \U$7399 ( \9328 , \9054 , \9056 );
nand \U$7400 ( \9329 , \9327 , \9328 );
nor \U$7401 ( \9330 , \9063 , \9060 );
and \U$7402 ( \9331 , \9330 , \4833 );
or \U$7403 ( \9332 , \9060 , \9067 );
nand \U$7404 ( \9333 , \9332 , \9071 );
nor \U$7405 ( \9334 , \9331 , \9333 );
or \U$7406 ( \9335 , \9329 , \9334 );
or \U$7407 ( \9336 , \9053 , \9074 );
nand \U$7408 ( \9337 , \9336 , \9079 );
and \U$7409 ( \9338 , \9328 , \9337 );
or \U$7410 ( \9339 , \9056 , \9082 );
nand \U$7411 ( \9340 , \9339 , \9086 );
nor \U$7412 ( \9341 , \9338 , \9340 );
nand \U$7413 ( \9342 , \9335 , \9341 );
not \U$7414 ( \9343 , \9342 );
xor \U$7415 ( \9344 , \9326 , \9343 );
buf g2f88_GF_PartitionCandidate( \9345_nG2f88 , \9344 );
not \U$7416 ( \9346 , \7121 );
nand \U$7417 ( \9347 , \7751 , \9346 );
nor \U$7418 ( \9348 , \9106 , \9098 );
nor \U$7419 ( \9349 , \9099 , \9101 );
nand \U$7420 ( \9350 , \9348 , \9349 );
nor \U$7421 ( \9351 , \9108 , \9105 );
and \U$7422 ( \9352 , \9351 , \7679 );
or \U$7423 ( \9353 , \9105 , \9112 );
nand \U$7424 ( \9354 , \9353 , \9116 );
nor \U$7425 ( \9355 , \9352 , \9354 );
or \U$7426 ( \9356 , \9350 , \9355 );
or \U$7427 ( \9357 , \9098 , \9119 );
nand \U$7428 ( \9358 , \9357 , \9124 );
and \U$7429 ( \9359 , \9349 , \9358 );
or \U$7430 ( \9360 , \9101 , \9127 );
nand \U$7431 ( \9361 , \9360 , \9131 );
nor \U$7432 ( \9362 , \9359 , \9361 );
nand \U$7433 ( \9363 , \9356 , \9362 );
not \U$7434 ( \9364 , \9363 );
xor \U$7435 ( \9365 , \9347 , \9364 );
buf g2fd4_GF_PartitionCandidate( \9366_nG2fd4 , \9365 );
_HMUX g2fd5_GF_PartitionCandidate ( \9367_nG2fd5 , \9345_nG2f88 , \9366_nG2fd4 , \8862 );
buf \U$7436 ( \9368 , \9367_nG2fd5 );
not \U$7437 ( \9369 , \4218 );
nand \U$7438 ( \9370 , \4902 , \9369 );
nor \U$7439 ( \9371 , \9153 , \9145 );
nor \U$7440 ( \9372 , \9146 , \9148 );
nand \U$7441 ( \9373 , \9371 , \9372 );
nor \U$7442 ( \9374 , \9155 , \9152 );
and \U$7443 ( \9375 , \9374 , \8893 );
or \U$7444 ( \9376 , \9152 , \9158 );
nand \U$7445 ( \9377 , \9376 , \9162 );
nor \U$7446 ( \9378 , \9375 , \9377 );
or \U$7447 ( \9379 , \9373 , \9378 );
or \U$7448 ( \9380 , \9145 , \9165 );
nand \U$7449 ( \9381 , \9380 , \9170 );
and \U$7450 ( \9382 , \9372 , \9381 );
or \U$7451 ( \9383 , \9148 , \9173 );
nand \U$7452 ( \9384 , \9383 , \9177 );
nor \U$7453 ( \9385 , \9382 , \9384 );
nand \U$7454 ( \9386 , \9379 , \9385 );
not \U$7455 ( \9387 , \9386 );
xor \U$7456 ( \9388 , \9370 , \9387 );
buf g2eeb_GF_PartitionCandidate( \9389_nG2eeb , \9388 );
not \U$7457 ( \9390 , \7064 );
nand \U$7458 ( \9391 , \7748 , \9390 );
nor \U$7459 ( \9392 , \9197 , \9189 );
nor \U$7460 ( \9393 , \9190 , \9192 );
nand \U$7461 ( \9394 , \9392 , \9393 );
nor \U$7462 ( \9395 , \9199 , \9196 );
and \U$7463 ( \9396 , \9395 , \8985 );
or \U$7464 ( \9397 , \9196 , \9202 );
nand \U$7465 ( \9398 , \9397 , \9206 );
nor \U$7466 ( \9399 , \9396 , \9398 );
or \U$7467 ( \9400 , \9394 , \9399 );
or \U$7468 ( \9401 , \9189 , \9209 );
nand \U$7469 ( \9402 , \9401 , \9214 );
and \U$7470 ( \9403 , \9393 , \9402 );
or \U$7471 ( \9404 , \9192 , \9217 );
nand \U$7472 ( \9405 , \9404 , \9221 );
nor \U$7473 ( \9406 , \9403 , \9405 );
nand \U$7474 ( \9407 , \9400 , \9406 );
not \U$7475 ( \9408 , \9407 );
xor \U$7476 ( \9409 , \9391 , \9408 );
buf g2f3b_GF_PartitionCandidate( \9410_nG2f3b , \9409 );
_HMUX g2f3c_GF_PartitionCandidate ( \9411_nG2f3c , \9389_nG2eeb , \9410_nG2f3b , \8862 );
buf \U$7477 ( \9412 , \9411_nG2f3c );
not \U$7478 ( \9413 , \4158 );
nand \U$7479 ( \9414 , \4900 , \9413 );
nand \U$7480 ( \9415 , \4739 , \4097 );
not \U$7481 ( \9416 , \4851 );
or \U$7482 ( \9417 , \9415 , \9416 );
and \U$7483 ( \9418 , \4097 , \4874 );
nor \U$7484 ( \9419 , \9418 , \4898 );
nand \U$7485 ( \9420 , \9417 , \9419 );
not \U$7486 ( \9421 , \9420 );
xor \U$7487 ( \9422 , \9414 , \9421 );
buf g2e49_GF_PartitionCandidate( \9423_nG2e49 , \9422 );
not \U$7488 ( \9424 , \7004 );
nand \U$7489 ( \9425 , \7746 , \9424 );
nand \U$7490 ( \9426 , \7585 , \6943 );
not \U$7491 ( \9427 , \7697 );
or \U$7492 ( \9428 , \9426 , \9427 );
and \U$7493 ( \9429 , \6943 , \7720 );
nor \U$7494 ( \9430 , \9429 , \7744 );
nand \U$7495 ( \9431 , \9428 , \9430 );
not \U$7496 ( \9432 , \9431 );
xor \U$7497 ( \9433 , \9425 , \9432 );
buf g2e9a_GF_PartitionCandidate( \9434_nG2e9a , \9433 );
_HMUX g2e9b_GF_PartitionCandidate ( \9435_nG2e9b , \9423_nG2e49 , \9434_nG2e9a , \8862 );
buf \U$7498 ( \9436 , \9435_nG2e9b );
not \U$7499 ( \9437 , \4094 );
nand \U$7500 ( \9438 , \4895 , \9437 );
nand \U$7501 ( \9439 , \8888 , \8873 );
not \U$7502 ( \9440 , \8905 );
or \U$7503 ( \9441 , \9439 , \9440 );
and \U$7504 ( \9442 , \8873 , \8920 );
nor \U$7505 ( \9443 , \9442 , \8936 );
nand \U$7506 ( \9444 , \9441 , \9443 );
not \U$7507 ( \9445 , \9444 );
xor \U$7508 ( \9446 , \9438 , \9445 );
buf g2d9e_GF_PartitionCandidate( \9447_nG2d9e , \9446 );
not \U$7509 ( \9448 , \6940 );
nand \U$7510 ( \9449 , \7741 , \9448 );
nand \U$7511 ( \9450 , \8980 , \8965 );
not \U$7512 ( \9451 , \8997 );
or \U$7513 ( \9452 , \9450 , \9451 );
and \U$7514 ( \9453 , \8965 , \9012 );
nor \U$7515 ( \9454 , \9453 , \9028 );
nand \U$7516 ( \9455 , \9452 , \9454 );
not \U$7517 ( \9456 , \9455 );
xor \U$7518 ( \9457 , \9449 , \9456 );
buf g2df7_GF_PartitionCandidate( \9458_nG2df7 , \9457 );
_HMUX g2df8_GF_PartitionCandidate ( \9459_nG2df8 , \9447_nG2d9e , \9458_nG2df7 , \8862 );
buf \U$7519 ( \9460 , \9459_nG2df8 );
not \U$7520 ( \9461 , \4025 );
nand \U$7521 ( \9462 , \4893 , \9461 );
nand \U$7522 ( \9463 , \9062 , \9055 );
not \U$7523 ( \9464 , \9068 );
or \U$7524 ( \9465 , \9463 , \9464 );
and \U$7525 ( \9466 , \9055 , \9075 );
nor \U$7526 ( \9467 , \9466 , \9083 );
nand \U$7527 ( \9468 , \9465 , \9467 );
not \U$7528 ( \9469 , \9468 );
xor \U$7529 ( \9470 , \9462 , \9469 );
buf g2ce8_GF_PartitionCandidate( \9471_nG2ce8 , \9470 );
not \U$7530 ( \9472 , \6871 );
nand \U$7531 ( \9473 , \7739 , \9472 );
nand \U$7532 ( \9474 , \9107 , \9100 );
not \U$7533 ( \9475 , \9113 );
or \U$7534 ( \9476 , \9474 , \9475 );
and \U$7535 ( \9477 , \9100 , \9120 );
nor \U$7536 ( \9478 , \9477 , \9128 );
nand \U$7537 ( \9479 , \9476 , \9478 );
not \U$7538 ( \9480 , \9479 );
xor \U$7539 ( \9481 , \9473 , \9480 );
buf g2d44_GF_PartitionCandidate( \9482_nG2d44 , \9481 );
_HMUX g2d45_GF_PartitionCandidate ( \9483_nG2d45 , \9471_nG2ce8 , \9482_nG2d44 , \8862 );
buf \U$7540 ( \9484 , \9483_nG2d45 );
not \U$7541 ( \9485 , \3952 );
nand \U$7542 ( \9486 , \4890 , \9485 );
nand \U$7543 ( \9487 , \9154 , \9147 );
not \U$7544 ( \9488 , \9159 );
or \U$7545 ( \9489 , \9487 , \9488 );
and \U$7546 ( \9490 , \9147 , \9166 );
nor \U$7547 ( \9491 , \9490 , \9174 );
nand \U$7548 ( \9492 , \9489 , \9491 );
not \U$7549 ( \9493 , \9492 );
xor \U$7550 ( \9494 , \9486 , \9493 );
buf g2c2b_GF_PartitionCandidate( \9495_nG2c2b , \9494 );
not \U$7551 ( \9496 , \6798 );
nand \U$7552 ( \9497 , \7736 , \9496 );
nand \U$7553 ( \9498 , \9198 , \9191 );
not \U$7554 ( \9499 , \9203 );
or \U$7555 ( \9500 , \9498 , \9499 );
and \U$7556 ( \9501 , \9191 , \9210 );
nor \U$7557 ( \9502 , \9501 , \9218 );
nand \U$7558 ( \9503 , \9500 , \9502 );
not \U$7559 ( \9504 , \9503 );
xor \U$7560 ( \9505 , \9497 , \9504 );
buf g2c8b_GF_PartitionCandidate( \9506_nG2c8b , \9505 );
_HMUX g2c8c_GF_PartitionCandidate ( \9507_nG2c8c , \9495_nG2c2b , \9506_nG2c8b , \8862 );
buf \U$7561 ( \9508 , \9507_nG2c8c );
not \U$7562 ( \9509 , \3876 );
nand \U$7563 ( \9510 , \4888 , \9509 );
nand \U$7564 ( \9511 , \9238 , \9235 );
or \U$7565 ( \9512 , \9511 , \4839 );
and \U$7566 ( \9513 , \9235 , \9242 );
nor \U$7567 ( \9514 , \9513 , \9246 );
nand \U$7568 ( \9515 , \9512 , \9514 );
not \U$7569 ( \9516 , \9515 );
xor \U$7570 ( \9517 , \9510 , \9516 );
buf g2b6b_GF_PartitionCandidate( \9518_nG2b6b , \9517 );
not \U$7571 ( \9519 , \6722 );
nand \U$7572 ( \9520 , \7734 , \9519 );
nand \U$7573 ( \9521 , \9260 , \9257 );
or \U$7574 ( \9522 , \9521 , \7685 );
and \U$7575 ( \9523 , \9257 , \9264 );
nor \U$7576 ( \9524 , \9523 , \9268 );
nand \U$7577 ( \9525 , \9522 , \9524 );
not \U$7578 ( \9526 , \9525 );
xor \U$7579 ( \9527 , \9520 , \9526 );
buf g2bca_GF_PartitionCandidate( \9528_nG2bca , \9527 );
_HMUX g2bcb_GF_PartitionCandidate ( \9529_nG2bcb , \9518_nG2b6b , \9528_nG2bca , \8862 );
buf \U$7580 ( \9530 , \9529_nG2bcb );
not \U$7581 ( \9531 , \3799 );
nand \U$7582 ( \9532 , \4884 , \9531 );
nand \U$7583 ( \9533 , \9284 , \9281 );
or \U$7584 ( \9534 , \9533 , \8897 );
and \U$7585 ( \9535 , \9281 , \9288 );
nor \U$7586 ( \9536 , \9535 , \9292 );
nand \U$7587 ( \9537 , \9534 , \9536 );
not \U$7588 ( \9538 , \9537 );
xor \U$7589 ( \9539 , \9532 , \9538 );
buf g2aac_GF_PartitionCandidate( \9540_nG2aac , \9539 );
not \U$7590 ( \9541 , \6645 );
nand \U$7591 ( \9542 , \7730 , \9541 );
nand \U$7592 ( \9543 , \9306 , \9303 );
or \U$7593 ( \9544 , \9543 , \8989 );
and \U$7594 ( \9545 , \9303 , \9310 );
nor \U$7595 ( \9546 , \9545 , \9314 );
nand \U$7596 ( \9547 , \9544 , \9546 );
not \U$7597 ( \9548 , \9547 );
xor \U$7598 ( \9549 , \9542 , \9548 );
buf g2b0b_GF_PartitionCandidate( \9550_nG2b0b , \9549 );
_HMUX g2b0c_GF_PartitionCandidate ( \9551_nG2b0c , \9540_nG2aac , \9550_nG2b0b , \8862 );
buf \U$7599 ( \9552 , \9551_nG2b0c );
not \U$7600 ( \9553 , \3724 );
nand \U$7601 ( \9554 , \4882 , \9553 );
nand \U$7602 ( \9555 , \9330 , \9327 );
or \U$7603 ( \9556 , \9555 , \9064 );
and \U$7604 ( \9557 , \9327 , \9333 );
nor \U$7605 ( \9558 , \9557 , \9337 );
nand \U$7606 ( \9559 , \9556 , \9558 );
not \U$7607 ( \9560 , \9559 );
xor \U$7608 ( \9561 , \9554 , \9560 );
buf g29d8_GF_PartitionCandidate( \9562_nG29d8 , \9561 );
not \U$7609 ( \9563 , \6570 );
nand \U$7610 ( \9564 , \7728 , \9563 );
nand \U$7611 ( \9565 , \9351 , \9348 );
or \U$7612 ( \9566 , \9565 , \9109 );
and \U$7613 ( \9567 , \9348 , \9354 );
nor \U$7614 ( \9568 , \9567 , \9358 );
nand \U$7615 ( \9569 , \9566 , \9568 );
not \U$7616 ( \9570 , \9569 );
xor \U$7617 ( \9571 , \9564 , \9570 );
buf g2a4c_GF_PartitionCandidate( \9572_nG2a4c , \9571 );
_HMUX g2a4d_GF_PartitionCandidate ( \9573_nG2a4d , \9562_nG29d8 , \9572_nG2a4c , \8862 );
buf \U$7618 ( \9574 , \9573_nG2a4d );
not \U$7619 ( \9575 , \3647 );
nand \U$7620 ( \9576 , \4879 , \9575 );
nand \U$7621 ( \9577 , \9374 , \9371 );
or \U$7622 ( \9578 , \9577 , \4830 );
and \U$7623 ( \9579 , \9371 , \9377 );
nor \U$7624 ( \9580 , \9579 , \9381 );
nand \U$7625 ( \9581 , \9578 , \9580 );
not \U$7626 ( \9582 , \9581 );
xor \U$7627 ( \9583 , \9576 , \9582 );
buf g28f0_GF_PartitionCandidate( \9584_nG28f0 , \9583 );
not \U$7628 ( \9585 , \6493 );
nand \U$7629 ( \9586 , \7725 , \9585 );
nand \U$7630 ( \9587 , \9395 , \9392 );
or \U$7631 ( \9588 , \9587 , \7676 );
and \U$7632 ( \9589 , \9392 , \9398 );
nor \U$7633 ( \9590 , \9589 , \9402 );
nand \U$7634 ( \9591 , \9588 , \9590 );
not \U$7635 ( \9592 , \9591 );
xor \U$7636 ( \9593 , \9586 , \9592 );
buf g2963_GF_PartitionCandidate( \9594_nG2963 , \9593 );
_HMUX g2964_GF_PartitionCandidate ( \9595_nG2964 , \9584_nG28f0 , \9594_nG2963 , \8862 );
buf \U$7637 ( \9596 , \9595_nG2964 );
not \U$7638 ( \9597 , \3572 );
nand \U$7639 ( \9598 , \4877 , \9597 );
xor \U$7640 ( \9599 , \9598 , \4875 );
buf g2810_GF_PartitionCandidate( \9600_nG2810 , \9599 );
not \U$7641 ( \9601 , \6418 );
nand \U$7642 ( \9602 , \7723 , \9601 );
xor \U$7643 ( \9603 , \9602 , \7721 );
buf g287c_GF_PartitionCandidate( \9604_nG287c , \9603 );
_HMUX g287d_GF_PartitionCandidate ( \9605_nG287d , \9600_nG2810 , \9604_nG287c , \8862 );
buf \U$7644 ( \9606 , \9605_nG287d );
not \U$7645 ( \9607 , \4736 );
nand \U$7646 ( \9608 , \4871 , \9607 );
xor \U$7647 ( \9609 , \9608 , \8921 );
buf g2737_GF_PartitionCandidate( \9610_nG2737 , \9609 );
not \U$7648 ( \9611 , \7582 );
nand \U$7649 ( \9612 , \7717 , \9611 );
xor \U$7650 ( \9613 , \9612 , \9013 );
buf g27a3_GF_PartitionCandidate( \9614_nG27a3 , \9613 );
_HMUX g27a4_GF_PartitionCandidate ( \9615_nG27a4 , \9610_nG2737 , \9614_nG27a3 , \8862 );
buf \U$7651 ( \9616 , \9615_nG27a4 );
not \U$7652 ( \9617 , \4729 );
nand \U$7653 ( \9618 , \4869 , \9617 );
xor \U$7654 ( \9619 , \9618 , \9076 );
buf g2662_GF_PartitionCandidate( \9620_nG2662 , \9619 );
not \U$7655 ( \9621 , \7575 );
nand \U$7656 ( \9622 , \7715 , \9621 );
xor \U$7657 ( \9623 , \9622 , \9121 );
buf g26ca_GF_PartitionCandidate( \9624_nG26ca , \9623 );
_HMUX g26cb_GF_PartitionCandidate ( \9625_nG26cb , \9620_nG2662 , \9624_nG26ca , \8862 );
buf \U$7658 ( \9626 , \9625_nG26cb );
not \U$7659 ( \9627 , \4713 );
nand \U$7660 ( \9628 , \4866 , \9627 );
xor \U$7661 ( \9629 , \9628 , \9167 );
buf g258f_GF_PartitionCandidate( \9630_nG258f , \9629 );
not \U$7662 ( \9631 , \7559 );
nand \U$7663 ( \9632 , \7712 , \9631 );
xor \U$7664 ( \9633 , \9632 , \9211 );
buf g25f9_GF_PartitionCandidate( \9634_nG25f9 , \9633 );
_HMUX g25fa_GF_PartitionCandidate ( \9635_nG25fa , \9630_nG258f , \9634_nG25f9 , \8862 );
buf \U$7665 ( \9636 , \9635_nG25fa );
not \U$7666 ( \9637 , \4692 );
nand \U$7667 ( \9638 , \4864 , \9637 );
xor \U$7668 ( \9639 , \9638 , \9243 );
buf g24bf_GF_PartitionCandidate( \9640_nG24bf , \9639 );
not \U$7669 ( \9641 , \7538 );
nand \U$7670 ( \9642 , \7710 , \9641 );
xor \U$7671 ( \9643 , \9642 , \9265 );
buf g2524_GF_PartitionCandidate( \9644_nG2524 , \9643 );
_HMUX g2525_GF_PartitionCandidate ( \9645_nG2525 , \9640_nG24bf , \9644_nG2524 , \8862 );
buf \U$7672 ( \9646 , \9645_nG2525 );
not \U$7673 ( \9647 , \4653 );
nand \U$7674 ( \9648 , \4860 , \9647 );
xor \U$7675 ( \9649 , \9648 , \9289 );
buf g23cd_GF_PartitionCandidate( \9650_nG23cd , \9649 );
not \U$7676 ( \9651 , \7499 );
nand \U$7677 ( \9652 , \7706 , \9651 );
xor \U$7678 ( \9653 , \9652 , \9311 );
buf g2459_GF_PartitionCandidate( \9654_nG2459 , \9653 );
_HMUX g245a_GF_PartitionCandidate ( \9655_nG245a , \9650_nG23cd , \9654_nG2459 , \8862 );
buf \U$7679 ( \9656 , \9655_nG245a );
not \U$7680 ( \9657 , \4598 );
nand \U$7681 ( \9658 , \4858 , \9657 );
xor \U$7682 ( \9659 , \9658 , \9334 );
buf g22e6_GF_PartitionCandidate( \9660_nG22e6 , \9659 );
not \U$7683 ( \9661 , \7444 );
nand \U$7684 ( \9662 , \7704 , \9661 );
xor \U$7685 ( \9663 , \9662 , \9355 );
buf g2340_GF_PartitionCandidate( \9664_nG2340 , \9663 );
_HMUX g2341_GF_PartitionCandidate ( \9665_nG2341 , \9660_nG22e6 , \9664_nG2340 , \8862 );
buf \U$7686 ( \9666 , \9665_nG2341 );
not \U$7687 ( \9667 , \4546 );
nand \U$7688 ( \9668 , \4855 , \9667 );
xor \U$7689 ( \9669 , \9668 , \9378 );
buf g21f2_GF_PartitionCandidate( \9670_nG21f2 , \9669 );
not \U$7690 ( \9671 , \7392 );
nand \U$7691 ( \9672 , \7701 , \9671 );
xor \U$7692 ( \9673 , \9672 , \9399 );
buf g228b_GF_PartitionCandidate( \9674_nG228b , \9673 );
_HMUX g228c_GF_PartitionCandidate ( \9675_nG228c , \9670_nG21f2 , \9674_nG228b , \8862 );
buf \U$7693 ( \9676 , \9675_nG228c );
not \U$7694 ( \9677 , \4501 );
nand \U$7695 ( \9678 , \4853 , \9677 );
xor \U$7696 ( \9679 , \9678 , \9416 );
buf g210a_GF_PartitionCandidate( \9680_nG210a , \9679 );
not \U$7697 ( \9681 , \7347 );
nand \U$7698 ( \9682 , \7699 , \9681 );
xor \U$7699 ( \9683 , \9682 , \9427 );
buf g2158_GF_PartitionCandidate( \9684_nG2158 , \9683 );
_HMUX g2159_GF_PartitionCandidate ( \9685_nG2159 , \9680_nG210a , \9684_nG2158 , \8862 );
buf \U$7700 ( \9686 , \9685_nG2159 );
not \U$7701 ( \9687 , \4797 );
nand \U$7702 ( \9688 , \4848 , \9687 );
xor \U$7703 ( \9689 , \9688 , \9440 );
buf g202e_GF_PartitionCandidate( \9690_nG202e , \9689 );
not \U$7704 ( \9691 , \7643 );
nand \U$7705 ( \9692 , \7694 , \9691 );
xor \U$7706 ( \9693 , \9692 , \9451 );
buf g20bb_GF_PartitionCandidate( \9694_nG20bb , \9693 );
_HMUX g20bc_GF_PartitionCandidate ( \9695_nG20bc , \9690_nG202e , \9694_nG20bb , \8862 );
buf \U$7707 ( \9696 , \9695_nG20bc );
not \U$7708 ( \9697 , \4794 );
nand \U$7709 ( \9698 , \4846 , \9697 );
xor \U$7710 ( \9699 , \9698 , \9464 );
buf g1f5c_GF_PartitionCandidate( \9700_nG1f5c , \9699 );
not \U$7711 ( \9701 , \7640 );
nand \U$7712 ( \9702 , \7692 , \9701 );
xor \U$7713 ( \9703 , \9702 , \9475 );
buf g1fa0_GF_PartitionCandidate( \9704_nG1fa0 , \9703 );
_HMUX g1fa1_GF_PartitionCandidate ( \9705_nG1fa1 , \9700_nG1f5c , \9704_nG1fa0 , \8862 );
buf \U$7714 ( \9706 , \9705_nG1fa1 );
not \U$7715 ( \9707 , \4783 );
nand \U$7716 ( \9708 , \4843 , \9707 );
xor \U$7717 ( \9709 , \9708 , \9488 );
buf g1e94_GF_PartitionCandidate( \9710_nG1e94 , \9709 );
not \U$7718 ( \9711 , \7629 );
nand \U$7719 ( \9712 , \7689 , \9711 );
xor \U$7720 ( \9713 , \9712 , \9499 );
buf g1f17_GF_PartitionCandidate( \9714_nG1f17 , \9713 );
_HMUX g1f18_GF_PartitionCandidate ( \9715_nG1f18 , \9710_nG1e94 , \9714_nG1f17 , \8862 );
buf \U$7721 ( \9716 , \9715_nG1f18 );
not \U$7722 ( \9717 , \4772 );
nand \U$7723 ( \9718 , \4841 , \9717 );
xor \U$7724 ( \9719 , \9718 , \4839 );
buf g1dda_GF_PartitionCandidate( \9720_nG1dda , \9719 );
not \U$7725 ( \9721 , \7618 );
nand \U$7726 ( \9722 , \7687 , \9721 );
xor \U$7727 ( \9723 , \9722 , \7685 );
buf g1e10_GF_PartitionCandidate( \9724_nG1e10 , \9723 );
_HMUX g1e11_GF_PartitionCandidate ( \9725_nG1e11 , \9720_nG1dda , \9724_nG1e10 , \8862 );
buf \U$7728 ( \9726 , \9725_nG1e11 );
not \U$7729 ( \9727 , \4817 );
nand \U$7730 ( \9728 , \4837 , \9727 );
xor \U$7731 ( \9729 , \9728 , \8897 );
buf g1d2d_GF_PartitionCandidate( \9730_nG1d2d , \9729 );
not \U$7732 ( \9731 , \7663 );
nand \U$7733 ( \9732 , \7683 , \9731 );
xor \U$7734 ( \9733 , \9732 , \8989 );
buf g1da3_GF_PartitionCandidate( \9734_nG1da3 , \9733 );
_HMUX g1da4_GF_PartitionCandidate ( \9735_nG1da4 , \9730_nG1d2d , \9734_nG1da3 , \8862 );
buf \U$7735 ( \9736 , \9735_nG1da4 );
not \U$7736 ( \9737 , \4814 );
nand \U$7737 ( \9738 , \4835 , \9737 );
xor \U$7738 ( \9739 , \9738 , \9064 );
buf g1c8c_GF_PartitionCandidate( \9740_nG1c8c , \9739 );
not \U$7739 ( \9741 , \7660 );
nand \U$7740 ( \9742 , \7681 , \9741 );
xor \U$7741 ( \9743 , \9742 , \9109 );
buf g1cb6_GF_PartitionCandidate( \9744_nG1cb6 , \9743 );
_HMUX g1cb7_GF_PartitionCandidate ( \9745_nG1cb7 , \9740_nG1c8c , \9744_nG1cb6 , \8862 );
buf \U$7742 ( \9746 , \9745_nG1cb7 );
not \U$7743 ( \9747 , \4822 );
nand \U$7744 ( \9748 , \4832 , \9747 );
xor \U$7745 ( \9749 , \9748 , \4830 );
buf g1bf9_GF_PartitionCandidate( \9750_nG1bf9 , \9749 );
not \U$7746 ( \9751 , \7668 );
nand \U$7747 ( \9752 , \7678 , \9751 );
xor \U$7748 ( \9753 , \9752 , \7676 );
buf g1c61_GF_PartitionCandidate( \9754_nG1c61 , \9753 );
_HMUX g1c62_GF_PartitionCandidate ( \9755_nG1c62 , \9750_nG1bf9 , \9754_nG1c61 , \8862 );
buf \U$7749 ( \9756 , \9755_nG1c62 );
nor \U$7750 ( \9757 , \4826 , \4829 );
not \U$7751 ( \9758 , \9757 );
nand \U$7752 ( \9759 , \4830 , \9758 );
not \U$7753 ( \9760 , \9759 );
buf g1b6e_GF_PartitionCandidate( \9761_nG1b6e , \9760 );
nor \U$7754 ( \9762 , \7672 , \7675 );
not \U$7755 ( \9763 , \9762 );
nand \U$7756 ( \9764 , \7676 , \9763 );
not \U$7757 ( \9765 , \9764 );
buf g1b90_GF_PartitionCandidate( \9766_nG1b90 , \9765 );
_HMUX g1b91_GF_PartitionCandidate ( \9767_nG1b91 , \9761_nG1b6e , \9766_nG1b90 , \8862 );
buf \U$7758 ( \9768 , \9767_nG1b91 );
xor \U$7759 ( \9769 , \4828 , \2987 );
buf g1ab0_GF_PartitionCandidate( \9770_nG1ab0 , \9769 );
xor \U$7760 ( \9771 , \7674 , \5833 );
buf g1b4b_GF_PartitionCandidate( \9772_nG1b4b , \9771 );
_HMUX g1b4c_GF_PartitionCandidate ( \9773_nG1b4c , \9770_nG1ab0 , \9772_nG1b4b , \8862 );
buf \U$7761 ( \9774 , \9773_nG1b4c );
buf \U$7766 ( \9775 , RI2b5e785db058_15);
buf \U$7767 ( \9776 , RI2b5e785dafe0_16);
buf \U$7768 ( \9777 , RI2b5e785daf68_17);
buf \U$7769 ( \9778 , RI2b5e785daef0_18);
buf \U$7770 ( \9779 , RI2b5e785dae78_19);
buf \U$7771 ( \9780 , RI2b5e785dae00_20);
buf \U$7772 ( \9781 , RI2b5e785dad88_21);
buf \U$7773 ( \9782 , RI2b5e785dad10_22);
buf \U$7774 ( \9783 , RI2b5e785dac98_23);
buf \U$7775 ( \9784 , RI2b5e785dac20_24);
buf \U$7776 ( \9785 , RI2b5e785daba8_25);
and \U$7777 ( \9786 , \9784 , \9785 );
and \U$7778 ( \9787 , \9783 , \9786 );
and \U$7779 ( \9788 , \9782 , \9787 );
and \U$7780 ( \9789 , \9781 , \9788 );
and \U$7781 ( \9790 , \9780 , \9789 );
and \U$7782 ( \9791 , \9779 , \9790 );
and \U$7783 ( \9792 , \9778 , \9791 );
and \U$7784 ( \9793 , \9777 , \9792 );
and \U$7785 ( \9794 , \9776 , \9793 );
xor \U$7786 ( \9795 , \9775 , \9794 );
buf \U$7787 ( \9796 , \9795 );
buf \U$7788 ( \9797 , \9796 );
not \U$7789 ( \9798 , RI2b5e785ae580_609);
nor \U$7790 ( \9799 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9798 , RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7791 ( \9800 , RI2b5e785daa40_28, \9799 );
not \U$7792 ( \9801 , RI2b5e785ae3a0_613);
not \U$7793 ( \9802 , RI2b5e785ae418_612);
not \U$7794 ( \9803 , RI2b5e785ae490_611);
not \U$7795 ( \9804 , RI2b5e785ae508_610);
nor \U$7796 ( \9805 , \9801 , \9802 , \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7797 ( \9806 , RI2b5e78549540_41, \9805 );
nor \U$7798 ( \9807 , RI2b5e785ae3a0_613, \9802 , \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7799 ( \9808 , RI2b5e785388a8_54, \9807 );
nor \U$7800 ( \9809 , \9801 , RI2b5e785ae418_612, \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7801 ( \9810 , RI2b5e784a6330_67, \9809 );
nor \U$7802 ( \9811 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7803 ( \9812 , RI2b5e78495698_80, \9811 );
nor \U$7804 ( \9813 , \9801 , \9802 , RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7805 ( \9814 , RI2b5e78495080_93, \9813 );
nor \U$7806 ( \9815 , RI2b5e785ae3a0_613, \9802 , RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7807 ( \9816 , RI2b5e78403b80_106, \9815 );
nor \U$7808 ( \9817 , \9801 , RI2b5e785ae418_612, RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7809 ( \9818 , RI2b5e775b1e60_119, \9817 );
nor \U$7810 ( \9819 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7811 ( \9820 , RI2b5e7750bdf8_132, \9819 );
nor \U$7812 ( \9821 , \9801 , \9802 , \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7813 ( \9822 , RI2b5e774ff5d0_145, \9821 );
nor \U$7814 ( \9823 , RI2b5e785ae3a0_613, \9802 , \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7815 ( \9824 , RI2b5e774f65e8_158, \9823 );
nor \U$7816 ( \9825 , \9801 , RI2b5e785ae418_612, \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7817 ( \9826 , RI2b5e774eabd0_171, \9825 );
nor \U$7818 ( \9827 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7819 ( \9828 , RI2b5e774de3a8_184, \9827 );
nor \U$7820 ( \9829 , \9801 , \9802 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7821 ( \9830 , RI2b5e774d53c0_197, \9829 );
nor \U$7822 ( \9831 , RI2b5e785ae3a0_613, \9802 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7823 ( \9832 , RI2b5e785f4300_210, \9831 );
nor \U$7824 ( \9833 , \9801 , RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7825 ( \9834 , RI2b5e785f3ce8_223, \9833 );
nor \U$7826 ( \9835 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$7827 ( \9836 , RI2b5e785eb0c0_236, \9835 );
or \U$7828 ( \9837 , \9800 , \9806 , \9808 , \9810 , \9812 , \9814 , \9816 , \9818 , \9820 , \9822 , \9824 , \9826 , \9828 , \9830 , \9832 , \9834 , \9836 );
buf \U$7829 ( \9838 , RI2b5e785ae5f8_608);
buf \U$7830 ( \9839 , RI2b5e785ae670_607);
buf \U$7831 ( \9840 , RI2b5e785ae6e8_606);
buf \U$7832 ( \9841 , RI2b5e785ae760_605);
buf \U$7833 ( \9842 , RI2b5e785ae7d8_604);
buf \U$7834 ( \9843 , RI2b5e785ae850_603);
buf \U$7835 ( \9844 , RI2b5e785ae8c8_602);
buf \U$7836 ( \9845 , RI2b5e785ae940_601);
buf \U$7837 ( \9846 , RI2b5e785ae580_609);
buf \U$7838 ( \9847 , RI2b5e785ae3a0_613);
buf \U$7839 ( \9848 , RI2b5e785ae418_612);
buf \U$7840 ( \9849 , RI2b5e785ae490_611);
buf \U$7841 ( \9850 , RI2b5e785ae508_610);
or \U$7842 ( \9851 , \9847 , \9848 , \9849 , \9850 );
and \U$7843 ( \9852 , \9846 , \9851 );
or \U$7844 ( \9853 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9852 );
buf \U$7845 ( \9854 , \9853 );
_DC g3a87 ( \9855_nG3a87 , \9837 , \9854 );
buf \U$7846 ( \9856 , \9855_nG3a87 );
not \U$7847 ( \9857 , \9856 );
xor \U$7848 ( \9858 , \9797 , \9857 );
xor \U$7849 ( \9859 , \9776 , \9793 );
buf \U$7850 ( \9860 , \9859 );
buf \U$7851 ( \9861 , \9860 );
and \U$7852 ( \9862 , RI2b5e785da9c8_29, \9799 );
and \U$7853 ( \9863 , RI2b5e785494c8_42, \9805 );
and \U$7854 ( \9864 , RI2b5e78538830_55, \9807 );
and \U$7855 ( \9865 , RI2b5e784a62b8_68, \9809 );
and \U$7856 ( \9866 , RI2b5e78495620_81, \9811 );
and \U$7857 ( \9867 , RI2b5e78495008_94, \9813 );
and \U$7858 ( \9868 , RI2b5e78403b08_107, \9815 );
and \U$7859 ( \9869 , RI2b5e775b1de8_120, \9817 );
and \U$7860 ( \9870 , RI2b5e7750bd80_133, \9819 );
and \U$7861 ( \9871 , RI2b5e774ff558_146, \9821 );
and \U$7862 ( \9872 , RI2b5e774f6570_159, \9823 );
and \U$7863 ( \9873 , RI2b5e774eab58_172, \9825 );
and \U$7864 ( \9874 , RI2b5e774de330_185, \9827 );
and \U$7865 ( \9875 , RI2b5e774d5348_198, \9829 );
and \U$7866 ( \9876 , RI2b5e785f4288_211, \9831 );
and \U$7867 ( \9877 , RI2b5e785f3658_224, \9833 );
and \U$7868 ( \9878 , RI2b5e785eb048_237, \9835 );
or \U$7869 ( \9879 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 );
_DC g3a63 ( \9880_nG3a63 , \9879 , \9854 );
buf \U$7870 ( \9881 , \9880_nG3a63 );
not \U$7871 ( \9882 , \9881 );
and \U$7872 ( \9883 , \9861 , \9882 );
xor \U$7873 ( \9884 , \9777 , \9792 );
buf \U$7874 ( \9885 , \9884 );
buf \U$7875 ( \9886 , \9885 );
and \U$7876 ( \9887 , RI2b5e785da950_30, \9799 );
and \U$7877 ( \9888 , RI2b5e78549450_43, \9805 );
and \U$7878 ( \9889 , RI2b5e785387b8_56, \9807 );
and \U$7879 ( \9890 , RI2b5e784a6240_69, \9809 );
and \U$7880 ( \9891 , RI2b5e784955a8_82, \9811 );
and \U$7881 ( \9892 , RI2b5e78494f90_95, \9813 );
and \U$7882 ( \9893 , RI2b5e78403a90_108, \9815 );
and \U$7883 ( \9894 , RI2b5e775b1d70_121, \9817 );
and \U$7884 ( \9895 , RI2b5e7750bd08_134, \9819 );
and \U$7885 ( \9896 , RI2b5e774ff4e0_147, \9821 );
and \U$7886 ( \9897 , RI2b5e774f64f8_160, \9823 );
and \U$7887 ( \9898 , RI2b5e774eaae0_173, \9825 );
and \U$7888 ( \9899 , RI2b5e774de2b8_186, \9827 );
and \U$7889 ( \9900 , RI2b5e774d52d0_199, \9829 );
and \U$7890 ( \9901 , RI2b5e785f4210_212, \9831 );
and \U$7891 ( \9902 , RI2b5e785eb5e8_225, \9833 );
and \U$7892 ( \9903 , RI2b5e785e6c50_238, \9835 );
or \U$7893 ( \9904 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 );
_DC g38dc ( \9905_nG38dc , \9904 , \9854 );
buf \U$7894 ( \9906 , \9905_nG38dc );
not \U$7895 ( \9907 , \9906 );
and \U$7896 ( \9908 , \9886 , \9907 );
xor \U$7897 ( \9909 , \9778 , \9791 );
buf \U$7898 ( \9910 , \9909 );
buf \U$7899 ( \9911 , \9910 );
and \U$7900 ( \9912 , RI2b5e785da8d8_31, \9799 );
and \U$7901 ( \9913 , RI2b5e785493d8_44, \9805 );
and \U$7902 ( \9914 , RI2b5e78538740_57, \9807 );
and \U$7903 ( \9915 , RI2b5e784a61c8_70, \9809 );
and \U$7904 ( \9916 , RI2b5e78495530_83, \9811 );
and \U$7905 ( \9917 , RI2b5e78494f18_96, \9813 );
and \U$7906 ( \9918 , RI2b5e78403a18_109, \9815 );
and \U$7907 ( \9919 , RI2b5e775b1cf8_122, \9817 );
and \U$7908 ( \9920 , RI2b5e7750bc90_135, \9819 );
and \U$7909 ( \9921 , RI2b5e774ff468_148, \9821 );
and \U$7910 ( \9922 , RI2b5e774f6480_161, \9823 );
and \U$7911 ( \9923 , RI2b5e774eaa68_174, \9825 );
and \U$7912 ( \9924 , RI2b5e774de240_187, \9827 );
and \U$7913 ( \9925 , RI2b5e774d5258_200, \9829 );
and \U$7914 ( \9926 , RI2b5e785f4198_213, \9831 );
and \U$7915 ( \9927 , RI2b5e785eb570_226, \9833 );
and \U$7916 ( \9928 , RI2b5e785e6bd8_239, \9835 );
or \U$7917 ( \9929 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 );
_DC g38b8 ( \9930_nG38b8 , \9929 , \9854 );
buf \U$7918 ( \9931 , \9930_nG38b8 );
not \U$7919 ( \9932 , \9931 );
and \U$7920 ( \9933 , \9911 , \9932 );
xor \U$7921 ( \9934 , \9779 , \9790 );
buf \U$7922 ( \9935 , \9934 );
buf \U$7923 ( \9936 , \9935 );
and \U$7924 ( \9937 , RI2b5e785da860_32, \9799 );
and \U$7925 ( \9938 , RI2b5e78549360_45, \9805 );
and \U$7926 ( \9939 , RI2b5e785386c8_58, \9807 );
and \U$7927 ( \9940 , RI2b5e784a6150_71, \9809 );
and \U$7928 ( \9941 , RI2b5e784954b8_84, \9811 );
and \U$7929 ( \9942 , RI2b5e78494ea0_97, \9813 );
and \U$7930 ( \9943 , RI2b5e784039a0_110, \9815 );
and \U$7931 ( \9944 , RI2b5e775b1c80_123, \9817 );
and \U$7932 ( \9945 , RI2b5e7750bc18_136, \9819 );
and \U$7933 ( \9946 , RI2b5e774ff3f0_149, \9821 );
and \U$7934 ( \9947 , RI2b5e774f6408_162, \9823 );
and \U$7935 ( \9948 , RI2b5e774ea9f0_175, \9825 );
and \U$7936 ( \9949 , RI2b5e774de1c8_188, \9827 );
and \U$7937 ( \9950 , RI2b5e774d51e0_201, \9829 );
and \U$7938 ( \9951 , RI2b5e785f4120_214, \9831 );
and \U$7939 ( \9952 , RI2b5e785eb4f8_227, \9833 );
and \U$7940 ( \9953 , RI2b5e785e64d0_240, \9835 );
or \U$7941 ( \9954 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 );
_DC g3743 ( \9955_nG3743 , \9954 , \9854 );
buf \U$7942 ( \9956 , \9955_nG3743 );
not \U$7943 ( \9957 , \9956 );
and \U$7944 ( \9958 , \9936 , \9957 );
xor \U$7945 ( \9959 , \9780 , \9789 );
buf \U$7946 ( \9960 , \9959 );
buf \U$7947 ( \9961 , \9960 );
and \U$7948 ( \9962 , RI2b5e78549900_33, \9799 );
and \U$7949 ( \9963 , RI2b5e78538c68_46, \9805 );
and \U$7950 ( \9964 , RI2b5e78538650_59, \9807 );
and \U$7951 ( \9965 , RI2b5e784a60d8_72, \9809 );
and \U$7952 ( \9966 , RI2b5e78495440_85, \9811 );
and \U$7953 ( \9967 , RI2b5e78494e28_98, \9813 );
and \U$7954 ( \9968 , RI2b5e78403928_111, \9815 );
and \U$7955 ( \9969 , RI2b5e775b1c08_124, \9817 );
and \U$7956 ( \9970 , RI2b5e7750bba0_137, \9819 );
and \U$7957 ( \9971 , RI2b5e774ff378_150, \9821 );
and \U$7958 ( \9972 , RI2b5e774f6390_163, \9823 );
and \U$7959 ( \9973 , RI2b5e774ea978_176, \9825 );
and \U$7960 ( \9974 , RI2b5e774de150_189, \9827 );
and \U$7961 ( \9975 , RI2b5e774d5168_202, \9829 );
and \U$7962 ( \9976 , RI2b5e785f40a8_215, \9831 );
and \U$7963 ( \9977 , RI2b5e785eb480_228, \9833 );
and \U$7964 ( \9978 , RI2b5e785da608_241, \9835 );
or \U$7965 ( \9979 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 );
_DC g371f ( \9980_nG371f , \9979 , \9854 );
buf \U$7966 ( \9981 , \9980_nG371f );
not \U$7967 ( \9982 , \9981 );
and \U$7968 ( \9983 , \9961 , \9982 );
xor \U$7969 ( \9984 , \9781 , \9788 );
buf \U$7970 ( \9985 , \9984 );
buf \U$7971 ( \9986 , \9985 );
and \U$7972 ( \9987 , RI2b5e78549888_34, \9799 );
and \U$7973 ( \9988 , RI2b5e78538bf0_47, \9805 );
and \U$7974 ( \9989 , RI2b5e785385d8_60, \9807 );
and \U$7975 ( \9990 , RI2b5e784a6060_73, \9809 );
and \U$7976 ( \9991 , RI2b5e784953c8_86, \9811 );
and \U$7977 ( \9992 , RI2b5e78403ec8_99, \9813 );
and \U$7978 ( \9993 , RI2b5e775b21a8_112, \9815 );
and \U$7979 ( \9994 , RI2b5e775b1b90_125, \9817 );
and \U$7980 ( \9995 , RI2b5e7750bb28_138, \9819 );
and \U$7981 ( \9996 , RI2b5e774ff300_151, \9821 );
and \U$7982 ( \9997 , RI2b5e774f6318_164, \9823 );
and \U$7983 ( \9998 , RI2b5e774ea900_177, \9825 );
and \U$7984 ( \9999 , RI2b5e774de0d8_190, \9827 );
and \U$7985 ( \10000 , RI2b5e774d50f0_203, \9829 );
and \U$7986 ( \10001 , RI2b5e785f4030_216, \9831 );
and \U$7987 ( \10002 , RI2b5e785eb408_229, \9833 );
and \U$7988 ( \10003 , RI2b5e785da590_242, \9835 );
or \U$7989 ( \10004 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 );
_DC g35e1 ( \10005_nG35e1 , \10004 , \9854 );
buf \U$7990 ( \10006 , \10005_nG35e1 );
not \U$7991 ( \10007 , \10006 );
and \U$7992 ( \10008 , \9986 , \10007 );
xor \U$7993 ( \10009 , \9782 , \9787 );
buf \U$7994 ( \10010 , \10009 );
buf \U$7995 ( \10011 , \10010 );
and \U$7996 ( \10012 , RI2b5e78549810_35, \9799 );
and \U$7997 ( \10013 , RI2b5e78538b78_48, \9805 );
and \U$7998 ( \10014 , RI2b5e78538560_61, \9807 );
and \U$7999 ( \10015 , RI2b5e784a5fe8_74, \9809 );
and \U$8000 ( \10016 , RI2b5e78495350_87, \9811 );
and \U$8001 ( \10017 , RI2b5e78403e50_100, \9813 );
and \U$8002 ( \10018 , RI2b5e775b2130_113, \9815 );
and \U$8003 ( \10019 , RI2b5e775b1b18_126, \9817 );
and \U$8004 ( \10020 , RI2b5e7750bab0_139, \9819 );
and \U$8005 ( \10021 , RI2b5e774ff288_152, \9821 );
and \U$8006 ( \10022 , RI2b5e774f62a0_165, \9823 );
and \U$8007 ( \10023 , RI2b5e774ea888_178, \9825 );
and \U$8008 ( \10024 , RI2b5e774de060_191, \9827 );
and \U$8009 ( \10025 , RI2b5e774d5078_204, \9829 );
and \U$8010 ( \10026 , RI2b5e785f3fb8_217, \9831 );
and \U$8011 ( \10027 , RI2b5e785eb390_230, \9833 );
and \U$8012 ( \10028 , RI2b5e785da518_243, \9835 );
or \U$8013 ( \10029 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 );
_DC g35bd ( \10030_nG35bd , \10029 , \9854 );
buf \U$8014 ( \10031 , \10030_nG35bd );
not \U$8015 ( \10032 , \10031 );
and \U$8016 ( \10033 , \10011 , \10032 );
xor \U$8017 ( \10034 , \9783 , \9786 );
buf \U$8018 ( \10035 , \10034 );
buf \U$8019 ( \10036 , \10035 );
and \U$8020 ( \10037 , RI2b5e78549798_36, \9799 );
and \U$8021 ( \10038 , RI2b5e78538b00_49, \9805 );
and \U$8022 ( \10039 , RI2b5e785384e8_62, \9807 );
and \U$8023 ( \10040 , RI2b5e784a5f70_75, \9809 );
and \U$8024 ( \10041 , RI2b5e784952d8_88, \9811 );
and \U$8025 ( \10042 , RI2b5e78403dd8_101, \9813 );
and \U$8026 ( \10043 , RI2b5e775b20b8_114, \9815 );
and \U$8027 ( \10044 , RI2b5e775b1aa0_127, \9817 );
and \U$8028 ( \10045 , RI2b5e7750ba38_140, \9819 );
and \U$8029 ( \10046 , RI2b5e774ff210_153, \9821 );
and \U$8030 ( \10047 , RI2b5e774f6228_166, \9823 );
and \U$8031 ( \10048 , RI2b5e774ea810_179, \9825 );
and \U$8032 ( \10049 , RI2b5e774ddfe8_192, \9827 );
and \U$8033 ( \10050 , RI2b5e774d5000_205, \9829 );
and \U$8034 ( \10051 , RI2b5e785f3f40_218, \9831 );
and \U$8035 ( \10052 , RI2b5e785eb318_231, \9833 );
and \U$8036 ( \10053 , RI2b5e785da4a0_244, \9835 );
or \U$8037 ( \10054 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 );
_DC g34b0 ( \10055_nG34b0 , \10054 , \9854 );
buf \U$8038 ( \10056 , \10055_nG34b0 );
not \U$8039 ( \10057 , \10056 );
and \U$8040 ( \10058 , \10036 , \10057 );
xor \U$8041 ( \10059 , \9784 , \9785 );
buf \U$8042 ( \10060 , \10059 );
buf \U$8043 ( \10061 , \10060 );
and \U$8044 ( \10062 , RI2b5e78549720_37, \9799 );
and \U$8045 ( \10063 , RI2b5e78538a88_50, \9805 );
and \U$8046 ( \10064 , RI2b5e78538470_63, \9807 );
and \U$8047 ( \10065 , RI2b5e784a5ef8_76, \9809 );
and \U$8048 ( \10066 , RI2b5e78495260_89, \9811 );
and \U$8049 ( \10067 , RI2b5e78403d60_102, \9813 );
and \U$8050 ( \10068 , RI2b5e775b2040_115, \9815 );
and \U$8051 ( \10069 , RI2b5e775b1a28_128, \9817 );
and \U$8052 ( \10070 , RI2b5e7750b9c0_141, \9819 );
and \U$8053 ( \10071 , RI2b5e774ff198_154, \9821 );
and \U$8054 ( \10072 , RI2b5e774f61b0_167, \9823 );
and \U$8055 ( \10073 , RI2b5e774ea798_180, \9825 );
and \U$8056 ( \10074 , RI2b5e774ddf70_193, \9827 );
and \U$8057 ( \10075 , RI2b5e774d4f88_206, \9829 );
and \U$8058 ( \10076 , RI2b5e785f3ec8_219, \9831 );
and \U$8059 ( \10077 , RI2b5e785eb2a0_232, \9833 );
and \U$8060 ( \10078 , RI2b5e785da428_245, \9835 );
or \U$8061 ( \10079 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 );
_DC g34c9 ( \10080_nG34c9 , \10079 , \9854 );
buf \U$8062 ( \10081 , \10080_nG34c9 );
not \U$8063 ( \10082 , \10081 );
and \U$8064 ( \10083 , \10061 , \10082 );
not \U$8065 ( \10084 , \9785 );
buf \U$8066 ( \10085 , \10084 );
buf \U$8067 ( \10086 , \10085 );
and \U$8068 ( \10087 , RI2b5e785496a8_38, \9799 );
and \U$8069 ( \10088 , RI2b5e78538a10_51, \9805 );
and \U$8070 ( \10089 , RI2b5e785383f8_64, \9807 );
and \U$8071 ( \10090 , RI2b5e784a5e80_77, \9809 );
and \U$8072 ( \10091 , RI2b5e784951e8_90, \9811 );
and \U$8073 ( \10092 , RI2b5e78403ce8_103, \9813 );
and \U$8074 ( \10093 , RI2b5e775b1fc8_116, \9815 );
and \U$8075 ( \10094 , RI2b5e775b19b0_129, \9817 );
and \U$8076 ( \10095 , RI2b5e7750b948_142, \9819 );
and \U$8077 ( \10096 , RI2b5e774ff120_155, \9821 );
and \U$8078 ( \10097 , RI2b5e774f6138_168, \9823 );
and \U$8079 ( \10098 , RI2b5e774ea720_181, \9825 );
and \U$8080 ( \10099 , RI2b5e774ddef8_194, \9827 );
and \U$8081 ( \10100 , RI2b5e774d4f10_207, \9829 );
and \U$8082 ( \10101 , RI2b5e785f3e50_220, \9831 );
and \U$8083 ( \10102 , RI2b5e785eb228_233, \9833 );
and \U$8084 ( \10103 , RI2b5e785da3b0_246, \9835 );
or \U$8085 ( \10104 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 );
_DC g3393 ( \10105_nG3393 , \10104 , \9854 );
buf \U$8086 ( \10106 , \10105_nG3393 );
not \U$8087 ( \10107 , \10106 );
and \U$8088 ( \10108 , \10086 , \10107 );
buf \U$8089 ( \10109 , RI2b5e785dab30_26);
buf \U$8092 ( \10110 , \10109 );
and \U$8093 ( \10111 , RI2b5e78549630_39, \9799 );
and \U$8094 ( \10112 , RI2b5e78538998_52, \9805 );
and \U$8095 ( \10113 , RI2b5e78538380_65, \9807 );
and \U$8096 ( \10114 , RI2b5e784a5e08_78, \9809 );
and \U$8097 ( \10115 , RI2b5e78495170_91, \9811 );
and \U$8098 ( \10116 , RI2b5e78403c70_104, \9813 );
and \U$8099 ( \10117 , RI2b5e775b1f50_117, \9815 );
and \U$8100 ( \10118 , RI2b5e775b1938_130, \9817 );
and \U$8101 ( \10119 , RI2b5e7750b8d0_143, \9819 );
and \U$8102 ( \10120 , RI2b5e774ff0a8_156, \9821 );
and \U$8103 ( \10121 , RI2b5e774f60c0_169, \9823 );
and \U$8104 ( \10122 , RI2b5e774ea6a8_182, \9825 );
and \U$8105 ( \10123 , RI2b5e774dde80_195, \9827 );
and \U$8106 ( \10124 , RI2b5e774d4e98_208, \9829 );
and \U$8107 ( \10125 , RI2b5e785f3dd8_221, \9831 );
and \U$8108 ( \10126 , RI2b5e785eb1b0_234, \9833 );
and \U$8109 ( \10127 , RI2b5e785da338_247, \9835 );
or \U$8110 ( \10128 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 );
_DC g3377 ( \10129_nG3377 , \10128 , \9854 );
buf \U$8111 ( \10130 , \10129_nG3377 );
not \U$8112 ( \10131 , \10130 );
or \U$8113 ( \10132 , \10110 , \10131 );
and \U$8114 ( \10133 , \10107 , \10132 );
and \U$8115 ( \10134 , \10086 , \10132 );
or \U$8116 ( \10135 , \10108 , \10133 , \10134 );
and \U$8117 ( \10136 , \10082 , \10135 );
and \U$8118 ( \10137 , \10061 , \10135 );
or \U$8119 ( \10138 , \10083 , \10136 , \10137 );
and \U$8120 ( \10139 , \10057 , \10138 );
and \U$8121 ( \10140 , \10036 , \10138 );
or \U$8122 ( \10141 , \10058 , \10139 , \10140 );
and \U$8123 ( \10142 , \10032 , \10141 );
and \U$8124 ( \10143 , \10011 , \10141 );
or \U$8125 ( \10144 , \10033 , \10142 , \10143 );
and \U$8126 ( \10145 , \10007 , \10144 );
and \U$8127 ( \10146 , \9986 , \10144 );
or \U$8128 ( \10147 , \10008 , \10145 , \10146 );
and \U$8129 ( \10148 , \9982 , \10147 );
and \U$8130 ( \10149 , \9961 , \10147 );
or \U$8131 ( \10150 , \9983 , \10148 , \10149 );
and \U$8132 ( \10151 , \9957 , \10150 );
and \U$8133 ( \10152 , \9936 , \10150 );
or \U$8134 ( \10153 , \9958 , \10151 , \10152 );
and \U$8135 ( \10154 , \9932 , \10153 );
and \U$8136 ( \10155 , \9911 , \10153 );
or \U$8137 ( \10156 , \9933 , \10154 , \10155 );
and \U$8138 ( \10157 , \9907 , \10156 );
and \U$8139 ( \10158 , \9886 , \10156 );
or \U$8140 ( \10159 , \9908 , \10157 , \10158 );
and \U$8141 ( \10160 , \9882 , \10159 );
and \U$8142 ( \10161 , \9861 , \10159 );
or \U$8143 ( \10162 , \9883 , \10160 , \10161 );
xor \U$8144 ( \10163 , \9858 , \10162 );
buf g3a90_GF_PartitionCandidate( \10164_nG3a90 , \10163 );
buf \U$8145 ( \10165 , \10164_nG3a90 );
xor \U$8146 ( \10166 , \9861 , \9882 );
xor \U$8147 ( \10167 , \10166 , \10159 );
buf g3a6c_GF_PartitionCandidate( \10168_nG3a6c , \10167 );
buf \U$8148 ( \10169 , \10168_nG3a6c );
xor \U$8149 ( \10170 , \9886 , \9907 );
xor \U$8150 ( \10171 , \10170 , \10156 );
buf g38e5_GF_PartitionCandidate( \10172_nG38e5 , \10171 );
buf \U$8151 ( \10173 , \10172_nG38e5 );
and \U$8152 ( \10174 , \10169 , \10173 );
not \U$8153 ( \10175 , \10174 );
and \U$8154 ( \10176 , \10165 , \10175 );
not \U$8155 ( \10177 , \10176 );
buf \U$8156 ( \10178 , RI2b5e785ae3a0_613);
buf \U$8157 ( \10179 , RI2b5e785ae5f8_608);
buf \U$8158 ( \10180 , RI2b5e785ae670_607);
buf \U$8159 ( \10181 , RI2b5e785ae6e8_606);
buf \U$8160 ( \10182 , RI2b5e785ae760_605);
buf \U$8161 ( \10183 , RI2b5e785ae7d8_604);
buf \U$8162 ( \10184 , RI2b5e785ae850_603);
buf \U$8163 ( \10185 , RI2b5e785ae8c8_602);
buf \U$8164 ( \10186 , RI2b5e785ae940_601);
buf \U$8165 ( \10187 , RI2b5e785ae580_609);
nor \U$8166 ( \10188 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 );
buf \U$8167 ( \10189 , \10188 );
buf \U$8168 ( \10190 , \10189 );
xor \U$8169 ( \10191 , \10178 , \10190 );
buf \U$8170 ( \10192 , \10191 );
buf \U$8171 ( \10193 , RI2b5e785ae418_612);
and \U$8172 ( \10194 , \10178 , \10190 );
xor \U$8173 ( \10195 , \10193 , \10194 );
buf \U$8174 ( \10196 , \10195 );
buf \U$8175 ( \10197 , RI2b5e785ae490_611);
and \U$8176 ( \10198 , \10193 , \10194 );
xor \U$8177 ( \10199 , \10197 , \10198 );
buf \U$8178 ( \10200 , \10199 );
buf \U$8179 ( \10201 , RI2b5e785ae508_610);
and \U$8180 ( \10202 , \10197 , \10198 );
xor \U$8181 ( \10203 , \10201 , \10202 );
buf \U$8182 ( \10204 , \10203 );
buf \U$8183 ( \10205 , RI2b5e785ae580_609);
and \U$8184 ( \10206 , \10201 , \10202 );
xor \U$8185 ( \10207 , \10205 , \10206 );
buf \U$8186 ( \10208 , \10207 );
not \U$8187 ( \10209 , \10208 );
buf \U$8188 ( \10210 , RI2b5e785ae5f8_608);
and \U$8189 ( \10211 , \10205 , \10206 );
xor \U$8190 ( \10212 , \10210 , \10211 );
buf \U$8191 ( \10213 , \10212 );
buf \U$8192 ( \10214 , RI2b5e785ae670_607);
and \U$8193 ( \10215 , \10210 , \10211 );
xor \U$8194 ( \10216 , \10214 , \10215 );
buf \U$8195 ( \10217 , \10216 );
buf \U$8196 ( \10218 , RI2b5e785ae6e8_606);
and \U$8197 ( \10219 , \10214 , \10215 );
xor \U$8198 ( \10220 , \10218 , \10219 );
buf \U$8199 ( \10221 , \10220 );
buf \U$8200 ( \10222 , RI2b5e785ae760_605);
and \U$8201 ( \10223 , \10218 , \10219 );
xor \U$8202 ( \10224 , \10222 , \10223 );
buf \U$8203 ( \10225 , \10224 );
buf \U$8204 ( \10226 , RI2b5e785ae7d8_604);
and \U$8205 ( \10227 , \10222 , \10223 );
xor \U$8206 ( \10228 , \10226 , \10227 );
buf \U$8207 ( \10229 , \10228 );
buf \U$8208 ( \10230 , RI2b5e785ae850_603);
and \U$8209 ( \10231 , \10226 , \10227 );
xor \U$8210 ( \10232 , \10230 , \10231 );
buf \U$8211 ( \10233 , \10232 );
buf \U$8212 ( \10234 , RI2b5e785ae8c8_602);
and \U$8213 ( \10235 , \10230 , \10231 );
xor \U$8214 ( \10236 , \10234 , \10235 );
buf \U$8215 ( \10237 , \10236 );
buf \U$8216 ( \10238 , RI2b5e785ae940_601);
and \U$8217 ( \10239 , \10234 , \10235 );
xor \U$8218 ( \10240 , \10238 , \10239 );
buf \U$8219 ( \10241 , \10240 );
nor \U$8220 ( \10242 , \10192 , \10196 , \10200 , \10204 , \10209 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8221 ( \10243 , RI2b5e785da248_249, \10242 );
not \U$8222 ( \10244 , \10192 );
not \U$8223 ( \10245 , \10196 );
not \U$8224 ( \10246 , \10200 );
not \U$8225 ( \10247 , \10204 );
nor \U$8226 ( \10248 , \10244 , \10245 , \10246 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8227 ( \10249 , RI2b5e785be750_269, \10248 );
nor \U$8228 ( \10250 , \10192 , \10245 , \10246 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8229 ( \10251 , RI2b5e785bc4a0_289, \10250 );
nor \U$8230 ( \10252 , \10244 , \10196 , \10246 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8231 ( \10253 , RI2b5e785bbb40_309, \10252 );
nor \U$8232 ( \10254 , \10192 , \10196 , \10246 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8233 ( \10255 , RI2b5e785b9c50_329, \10254 );
nor \U$8234 ( \10256 , \10244 , \10245 , \10200 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8235 ( \10257 , RI2b5e785b8120_349, \10256 );
nor \U$8236 ( \10258 , \10192 , \10245 , \10200 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8237 ( \10259 , RI2b5e785b77c0_369, \10258 );
nor \U$8238 ( \10260 , \10244 , \10196 , \10200 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8239 ( \10261 , RI2b5e785b6e60_389, \10260 );
nor \U$8240 ( \10262 , \10192 , \10196 , \10200 , \10247 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8241 ( \10263 , RI2b5e785b56f0_409, \10262 );
nor \U$8242 ( \10264 , \10244 , \10245 , \10246 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8243 ( \10265 , RI2b5e785b4d90_429, \10264 );
nor \U$8244 ( \10266 , \10192 , \10245 , \10246 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8245 ( \10267 , RI2b5e785b39e0_449, \10266 );
nor \U$8246 ( \10268 , \10244 , \10196 , \10246 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8247 ( \10269 , RI2b5e785b3080_469, \10268 );
nor \U$8248 ( \10270 , \10192 , \10196 , \10246 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8249 ( \10271 , RI2b5e785b2720_489, \10270 );
nor \U$8250 ( \10272 , \10244 , \10245 , \10200 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8251 ( \10273 , RI2b5e785b1730_509, \10272 );
nor \U$8252 ( \10274 , \10192 , \10245 , \10200 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8253 ( \10275 , RI2b5e785b0dd0_529, \10274 );
nor \U$8254 ( \10276 , \10244 , \10196 , \10200 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8255 ( \10277 , RI2b5e785b0470_549, \10276 );
nor \U$8256 ( \10278 , \10192 , \10196 , \10200 , \10204 , \10208 , \10213 , \10217 , \10221 , \10225 , \10229 , \10233 , \10237 , \10241 );
and \U$8257 ( \10279 , RI2b5e785af840_569, \10278 );
or \U$8258 ( \10280 , \10243 , \10249 , \10251 , \10253 , \10255 , \10257 , \10259 , \10261 , \10263 , \10265 , \10267 , \10269 , \10271 , \10273 , \10275 , \10277 , \10279 );
buf \U$8259 ( \10281 , \10213 );
buf \U$8260 ( \10282 , \10217 );
buf \U$8261 ( \10283 , \10221 );
buf \U$8262 ( \10284 , \10225 );
buf \U$8263 ( \10285 , \10229 );
buf \U$8264 ( \10286 , \10233 );
buf \U$8265 ( \10287 , \10237 );
buf \U$8266 ( \10288 , \10241 );
buf \U$8267 ( \10289 , \10208 );
buf \U$8268 ( \10290 , \10192 );
buf \U$8269 ( \10291 , \10196 );
buf \U$8270 ( \10292 , \10200 );
buf \U$8271 ( \10293 , \10204 );
or \U$8272 ( \10294 , \10290 , \10291 , \10292 , \10293 );
and \U$8273 ( \10295 , \10289 , \10294 );
or \U$8274 ( \10296 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10295 );
buf \U$8275 ( \10297 , \10296 );
_DC g4187 ( \10298_nG4187 , \10280 , \10297 );
buf \U$8276 ( \10299 , \10298_nG4187 );
buf \U$8277 ( \10300 , RI2b5e785db0d0_14);
and \U$8278 ( \10301 , \9775 , \9794 );
and \U$8279 ( \10302 , \10300 , \10301 );
buf \U$8280 ( \10303 , \10302 );
buf \U$8281 ( \10304 , \10303 );
xor \U$8282 ( \10305 , \10300 , \10301 );
buf \U$8283 ( \10306 , \10305 );
buf \U$8284 ( \10307 , \10306 );
and \U$8285 ( \10308 , RI2b5e785daab8_27, \9799 );
and \U$8286 ( \10309 , RI2b5e785495b8_40, \9805 );
and \U$8287 ( \10310 , RI2b5e78538920_53, \9807 );
and \U$8288 ( \10311 , RI2b5e784a63a8_66, \9809 );
and \U$8289 ( \10312 , RI2b5e78495710_79, \9811 );
and \U$8290 ( \10313 , RI2b5e784950f8_92, \9813 );
and \U$8291 ( \10314 , RI2b5e78403bf8_105, \9815 );
and \U$8292 ( \10315 , RI2b5e775b1ed8_118, \9817 );
and \U$8293 ( \10316 , RI2b5e775b18c0_131, \9819 );
and \U$8294 ( \10317 , RI2b5e7750b858_144, \9821 );
and \U$8295 ( \10318 , RI2b5e774ff030_157, \9823 );
and \U$8296 ( \10319 , RI2b5e774f6048_170, \9825 );
and \U$8297 ( \10320 , RI2b5e774ea630_183, \9827 );
and \U$8298 ( \10321 , RI2b5e774dde08_196, \9829 );
and \U$8299 ( \10322 , RI2b5e774d4e20_209, \9831 );
and \U$8300 ( \10323 , RI2b5e785f3d60_222, \9833 );
and \U$8301 ( \10324 , RI2b5e785eb138_235, \9835 );
or \U$8302 ( \10325 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 );
_DC g3c4f ( \10326_nG3c4f , \10325 , \9854 );
buf \U$8303 ( \10327 , \10326_nG3c4f );
not \U$8304 ( \10328 , \10327 );
and \U$8305 ( \10329 , \10307 , \10328 );
and \U$8306 ( \10330 , \9797 , \9857 );
and \U$8307 ( \10331 , \9857 , \10162 );
and \U$8308 ( \10332 , \9797 , \10162 );
or \U$8309 ( \10333 , \10330 , \10331 , \10332 );
and \U$8310 ( \10334 , \10328 , \10333 );
and \U$8311 ( \10335 , \10307 , \10333 );
or \U$8312 ( \10336 , \10329 , \10334 , \10335 );
xnor \U$8313 ( \10337 , \10304 , \10336 );
buf g3c64_GF_PartitionCandidate( \10338_nG3c64 , \10337 );
buf \U$8314 ( \10339 , \10338_nG3c64 );
xor \U$8315 ( \10340 , \10307 , \10328 );
xor \U$8316 ( \10341 , \10340 , \10333 );
buf g3c58_GF_PartitionCandidate( \10342_nG3c58 , \10341 );
buf \U$8317 ( \10343 , \10342_nG3c58 );
xor \U$8318 ( \10344 , \10339 , \10343 );
xor \U$8319 ( \10345 , \10343 , \10165 );
not \U$8320 ( \10346 , \10345 );
and \U$8321 ( \10347 , \10344 , \10346 );
and \U$8322 ( \10348 , \10299 , \10347 );
and \U$8323 ( \10349 , RI2b5e785da2c0_248, \10242 );
and \U$8324 ( \10350 , RI2b5e785be7c8_268, \10248 );
and \U$8325 ( \10351 , RI2b5e785bc518_288, \10250 );
and \U$8326 ( \10352 , RI2b5e785bbbb8_308, \10252 );
and \U$8327 ( \10353 , RI2b5e785b9cc8_328, \10254 );
and \U$8328 ( \10354 , RI2b5e785b9368_348, \10256 );
and \U$8329 ( \10355 , RI2b5e785b7838_368, \10258 );
and \U$8330 ( \10356 , RI2b5e785b6ed8_388, \10260 );
and \U$8331 ( \10357 , RI2b5e785b5768_408, \10262 );
and \U$8332 ( \10358 , RI2b5e785b4e08_428, \10264 );
and \U$8333 ( \10359 , RI2b5e785b3a58_448, \10266 );
and \U$8334 ( \10360 , RI2b5e785b30f8_468, \10268 );
and \U$8335 ( \10361 , RI2b5e785b2798_488, \10270 );
and \U$8336 ( \10362 , RI2b5e785b17a8_508, \10272 );
and \U$8337 ( \10363 , RI2b5e785b0e48_528, \10274 );
and \U$8338 ( \10364 , RI2b5e785b04e8_548, \10276 );
and \U$8339 ( \10365 , RI2b5e785afb88_568, \10278 );
or \U$8340 ( \10366 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 );
_DC g427b ( \10367_nG427b , \10366 , \10297 );
buf \U$8341 ( \10368 , \10367_nG427b );
and \U$8342 ( \10369 , \10368 , \10345 );
nor \U$8343 ( \10370 , \10348 , \10369 );
and \U$8344 ( \10371 , \10343 , \10165 );
not \U$8345 ( \10372 , \10371 );
and \U$8346 ( \10373 , \10339 , \10372 );
xnor \U$8347 ( \10374 , \10370 , \10373 );
xor \U$8348 ( \10375 , \10177 , \10374 );
and \U$8350 ( \10376 , RI2b5e785da1d0_250, \10242 );
and \U$8351 ( \10377 , RI2b5e785be6d8_270, \10248 );
and \U$8352 ( \10378 , RI2b5e785bc428_290, \10250 );
and \U$8353 ( \10379 , RI2b5e785bbac8_310, \10252 );
and \U$8354 ( \10380 , RI2b5e785b9bd8_330, \10254 );
and \U$8355 ( \10381 , RI2b5e785b80a8_350, \10256 );
and \U$8356 ( \10382 , RI2b5e785b7748_370, \10258 );
and \U$8357 ( \10383 , RI2b5e785b6de8_390, \10260 );
and \U$8358 ( \10384 , RI2b5e785b5678_410, \10262 );
and \U$8359 ( \10385 , RI2b5e785b4d18_430, \10264 );
and \U$8360 ( \10386 , RI2b5e785b3968_450, \10266 );
and \U$8361 ( \10387 , RI2b5e785b3008_470, \10268 );
and \U$8362 ( \10388 , RI2b5e785b26a8_490, \10270 );
and \U$8363 ( \10389 , RI2b5e785b16b8_510, \10272 );
and \U$8364 ( \10390 , RI2b5e785b0d58_530, \10274 );
and \U$8365 ( \10391 , RI2b5e785b03f8_550, \10276 );
and \U$8366 ( \10392 , RI2b5e785af7c8_570, \10278 );
or \U$8367 ( \10393 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 );
_DC g40c5 ( \10394_nG40c5 , \10393 , \10297 );
buf \U$8368 ( \10395 , \10394_nG40c5 );
or \U$8369 ( \10396 , \10304 , \10336 );
not \U$8370 ( \10397 , \10396 );
buf g3e60_GF_PartitionCandidate( \10398_nG3e60 , \10397 );
buf \U$8371 ( \10399 , \10398_nG3e60 );
xor \U$8372 ( \10400 , \10399 , \10339 );
and \U$8373 ( \10401 , \10395 , \10400 );
nor \U$8374 ( \10402 , 1'b0 , \10401 );
xnor \U$8376 ( \10403 , \10402 , 1'b0 );
xor \U$8377 ( \10404 , \10375 , \10403 );
xor \U$8378 ( \10405 , 1'b0 , \10404 );
xor \U$8380 ( \10406 , \10165 , \10169 );
xor \U$8381 ( \10407 , \10169 , \10173 );
not \U$8382 ( \10408 , \10407 );
and \U$8383 ( \10409 , \10406 , \10408 );
and \U$8384 ( \10410 , \10368 , \10409 );
not \U$8385 ( \10411 , \10410 );
xnor \U$8386 ( \10412 , \10411 , \10176 );
and \U$8387 ( \10413 , \10395 , \10347 );
and \U$8388 ( \10414 , \10299 , \10345 );
nor \U$8389 ( \10415 , \10413 , \10414 );
xnor \U$8390 ( \10416 , \10415 , \10373 );
and \U$8391 ( \10417 , \10412 , \10416 );
or \U$8393 ( \10418 , 1'b0 , \10417 , 1'b0 );
xor \U$8395 ( \10419 , \10418 , 1'b0 );
xor \U$8397 ( \10420 , \10419 , 1'b0 );
and \U$8398 ( \10421 , \10405 , \10420 );
or \U$8399 ( \10422 , 1'b0 , 1'b0 , \10421 );
and \U$8402 ( \10423 , \10368 , \10347 );
not \U$8403 ( \10424 , \10423 );
xnor \U$8404 ( \10425 , \10424 , \10373 );
xor \U$8405 ( \10426 , 1'b0 , \10425 );
and \U$8407 ( \10427 , \10299 , \10400 );
nor \U$8408 ( \10428 , 1'b0 , \10427 );
xnor \U$8409 ( \10429 , \10428 , 1'b0 );
xor \U$8410 ( \10430 , \10426 , \10429 );
xor \U$8411 ( \10431 , 1'b0 , \10430 );
xor \U$8413 ( \10432 , \10431 , 1'b1 );
and \U$8414 ( \10433 , \10177 , \10374 );
and \U$8415 ( \10434 , \10374 , \10403 );
and \U$8416 ( \10435 , \10177 , \10403 );
or \U$8417 ( \10436 , \10433 , \10434 , \10435 );
xor \U$8419 ( \10437 , \10436 , 1'b0 );
xor \U$8421 ( \10438 , \10437 , 1'b0 );
xor \U$8422 ( \10439 , \10432 , \10438 );
and \U$8423 ( \10440 , \10422 , \10439 );
or \U$8425 ( \10441 , 1'b0 , \10440 , 1'b0 );
xor \U$8427 ( \10442 , \10441 , 1'b0 );
and \U$8429 ( \10443 , \10431 , 1'b1 );
and \U$8430 ( \10444 , 1'b1 , \10438 );
and \U$8431 ( \10445 , \10431 , \10438 );
or \U$8432 ( \10446 , \10443 , \10444 , \10445 );
xor \U$8433 ( \10447 , 1'b0 , \10446 );
not \U$8435 ( \10448 , \10373 );
and \U$8437 ( \10449 , \10368 , \10400 );
nor \U$8438 ( \10450 , 1'b0 , \10449 );
xnor \U$8439 ( \10451 , \10450 , 1'b0 );
xor \U$8440 ( \10452 , \10448 , \10451 );
xor \U$8442 ( \10453 , \10452 , 1'b0 );
xor \U$8443 ( \10454 , 1'b0 , \10453 );
xor \U$8445 ( \10455 , \10454 , 1'b0 );
and \U$8447 ( \10456 , \10425 , \10429 );
or \U$8449 ( \10457 , 1'b0 , \10456 , 1'b0 );
xor \U$8451 ( \10458 , \10457 , 1'b0 );
xor \U$8453 ( \10459 , \10458 , 1'b0 );
xor \U$8454 ( \10460 , \10455 , \10459 );
xor \U$8455 ( \10461 , \10447 , \10460 );
xor \U$8456 ( \10462 , \10442 , \10461 );
xor \U$8462 ( \10463 , \9911 , \9932 );
xor \U$8463 ( \10464 , \10463 , \10153 );
buf g38c1_GF_PartitionCandidate( \10465_nG38c1 , \10464 );
buf \U$8464 ( \10466 , \10465_nG38c1 );
xor \U$8465 ( \10467 , \10173 , \10466 );
xor \U$8466 ( \10468 , \9936 , \9957 );
xor \U$8467 ( \10469 , \10468 , \10150 );
buf g374c_GF_PartitionCandidate( \10470_nG374c , \10469 );
buf \U$8468 ( \10471 , \10470_nG374c );
xor \U$8469 ( \10472 , \10466 , \10471 );
not \U$8470 ( \10473 , \10472 );
and \U$8471 ( \10474 , \10467 , \10473 );
and \U$8472 ( \10475 , \10368 , \10474 );
not \U$8473 ( \10476 , \10475 );
and \U$8474 ( \10477 , \10466 , \10471 );
not \U$8475 ( \10478 , \10477 );
and \U$8476 ( \10479 , \10173 , \10478 );
xnor \U$8477 ( \10480 , \10476 , \10479 );
and \U$8478 ( \10481 , \10395 , \10409 );
and \U$8479 ( \10482 , \10299 , \10407 );
nor \U$8480 ( \10483 , \10481 , \10482 );
xnor \U$8481 ( \10484 , \10483 , \10176 );
and \U$8482 ( \10485 , \10480 , \10484 );
or \U$8484 ( \10486 , 1'b0 , \10485 , 1'b0 );
and \U$8485 ( \10487 , RI2b5e785da0e0_252, \10242 );
and \U$8486 ( \10488 , RI2b5e785be5e8_272, \10248 );
and \U$8487 ( \10489 , RI2b5e785bc338_292, \10250 );
and \U$8488 ( \10490 , RI2b5e785bb9d8_312, \10252 );
and \U$8489 ( \10491 , RI2b5e785b9ae8_332, \10254 );
and \U$8490 ( \10492 , RI2b5e785b7fb8_352, \10256 );
and \U$8491 ( \10493 , RI2b5e785b7658_372, \10258 );
and \U$8492 ( \10494 , RI2b5e785b5ee8_392, \10260 );
and \U$8493 ( \10495 , RI2b5e785b5588_412, \10262 );
and \U$8494 ( \10496 , RI2b5e785b4c28_432, \10264 );
and \U$8495 ( \10497 , RI2b5e785b3878_452, \10266 );
and \U$8496 ( \10498 , RI2b5e785b2f18_472, \10268 );
and \U$8497 ( \10499 , RI2b5e785b25b8_492, \10270 );
and \U$8498 ( \10500 , RI2b5e785b15c8_512, \10272 );
and \U$8499 ( \10501 , RI2b5e785b0c68_532, \10274 );
and \U$8500 ( \10502 , RI2b5e785b0308_552, \10276 );
and \U$8501 ( \10503 , RI2b5e785af6d8_572, \10278 );
or \U$8502 ( \10504 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 );
_DC g3f2a ( \10505_nG3f2a , \10504 , \10297 );
buf \U$8503 ( \10506 , \10505_nG3f2a );
and \U$8504 ( \10507 , \10506 , \10347 );
and \U$8505 ( \10508 , RI2b5e785da158_251, \10242 );
and \U$8506 ( \10509 , RI2b5e785be660_271, \10248 );
and \U$8507 ( \10510 , RI2b5e785bc3b0_291, \10250 );
and \U$8508 ( \10511 , RI2b5e785bba50_311, \10252 );
and \U$8509 ( \10512 , RI2b5e785b9b60_331, \10254 );
and \U$8510 ( \10513 , RI2b5e785b8030_351, \10256 );
and \U$8511 ( \10514 , RI2b5e785b76d0_371, \10258 );
and \U$8512 ( \10515 , RI2b5e785b6d70_391, \10260 );
and \U$8513 ( \10516 , RI2b5e785b5600_411, \10262 );
and \U$8514 ( \10517 , RI2b5e785b4ca0_431, \10264 );
and \U$8515 ( \10518 , RI2b5e785b38f0_451, \10266 );
and \U$8516 ( \10519 , RI2b5e785b2f90_471, \10268 );
and \U$8517 ( \10520 , RI2b5e785b2630_491, \10270 );
and \U$8518 ( \10521 , RI2b5e785b1640_511, \10272 );
and \U$8519 ( \10522 , RI2b5e785b0ce0_531, \10274 );
and \U$8520 ( \10523 , RI2b5e785b0380_551, \10276 );
and \U$8521 ( \10524 , RI2b5e785af750_571, \10278 );
or \U$8522 ( \10525 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 );
_DC g4004 ( \10526_nG4004 , \10525 , \10297 );
buf \U$8523 ( \10527 , \10526_nG4004 );
and \U$8524 ( \10528 , \10527 , \10345 );
nor \U$8525 ( \10529 , \10507 , \10528 );
xnor \U$8526 ( \10530 , \10529 , \10373 );
and \U$8528 ( \10531 , RI2b5e785da068_253, \10242 );
and \U$8529 ( \10532 , RI2b5e785be570_273, \10248 );
and \U$8530 ( \10533 , RI2b5e785bc2c0_293, \10250 );
and \U$8531 ( \10534 , RI2b5e785bb960_313, \10252 );
and \U$8532 ( \10535 , RI2b5e785b9a70_333, \10254 );
and \U$8533 ( \10536 , RI2b5e785b7f40_353, \10256 );
and \U$8534 ( \10537 , RI2b5e785b75e0_373, \10258 );
and \U$8535 ( \10538 , RI2b5e785b5e70_393, \10260 );
and \U$8536 ( \10539 , RI2b5e785b5510_413, \10262 );
and \U$8537 ( \10540 , RI2b5e785b4bb0_433, \10264 );
and \U$8538 ( \10541 , RI2b5e785b3800_453, \10266 );
and \U$8539 ( \10542 , RI2b5e785b2ea0_473, \10268 );
and \U$8540 ( \10543 , RI2b5e785b2540_493, \10270 );
and \U$8541 ( \10544 , RI2b5e785b1550_513, \10272 );
and \U$8542 ( \10545 , RI2b5e785b0bf0_533, \10274 );
and \U$8543 ( \10546 , RI2b5e785b0290_553, \10276 );
and \U$8544 ( \10547 , RI2b5e785af660_573, \10278 );
or \U$8545 ( \10548 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 );
_DC g3e3f ( \10549_nG3e3f , \10548 , \10297 );
buf \U$8546 ( \10550 , \10549_nG3e3f );
and \U$8547 ( \10551 , \10550 , \10400 );
nor \U$8548 ( \10552 , 1'b0 , \10551 );
xnor \U$8549 ( \10553 , \10552 , 1'b0 );
and \U$8550 ( \10554 , \10530 , \10553 );
or \U$8553 ( \10555 , \10554 , 1'b0 , 1'b0 );
and \U$8554 ( \10556 , \10486 , \10555 );
or \U$8557 ( \10557 , \10556 , 1'b0 , 1'b0 );
and \U$8560 ( \10558 , \10506 , \10400 );
nor \U$8561 ( \10559 , 1'b0 , \10558 );
xnor \U$8562 ( \10560 , \10559 , 1'b0 );
xor \U$8564 ( \10561 , \10560 , 1'b0 );
xor \U$8566 ( \10562 , \10561 , 1'b0 );
not \U$8567 ( \10563 , \10479 );
and \U$8568 ( \10564 , \10299 , \10409 );
and \U$8569 ( \10565 , \10368 , \10407 );
nor \U$8570 ( \10566 , \10564 , \10565 );
xnor \U$8571 ( \10567 , \10566 , \10176 );
xor \U$8572 ( \10568 , \10563 , \10567 );
and \U$8573 ( \10569 , \10527 , \10347 );
and \U$8574 ( \10570 , \10395 , \10345 );
nor \U$8575 ( \10571 , \10569 , \10570 );
xnor \U$8576 ( \10572 , \10571 , \10373 );
xor \U$8577 ( \10573 , \10568 , \10572 );
and \U$8578 ( \10574 , \10562 , \10573 );
or \U$8580 ( \10575 , 1'b0 , \10574 , 1'b0 );
and \U$8581 ( \10576 , \10557 , \10575 );
or \U$8582 ( \10577 , 1'b0 , 1'b0 , \10576 );
and \U$8584 ( \10578 , \10527 , \10400 );
nor \U$8585 ( \10579 , 1'b0 , \10578 );
xnor \U$8586 ( \10580 , \10579 , 1'b0 );
xor \U$8588 ( \10581 , \10580 , 1'b0 );
xor \U$8590 ( \10582 , \10581 , 1'b0 );
xor \U$8592 ( \10583 , 1'b0 , \10412 );
xor \U$8593 ( \10584 , \10583 , \10416 );
xor \U$8594 ( \10585 , \10582 , \10584 );
and \U$8596 ( \10586 , \10585 , 1'b1 );
and \U$8597 ( \10587 , \10563 , \10567 );
and \U$8598 ( \10588 , \10567 , \10572 );
and \U$8599 ( \10589 , \10563 , \10572 );
or \U$8600 ( \10590 , \10587 , \10588 , \10589 );
xor \U$8602 ( \10591 , \10590 , 1'b0 );
xor \U$8604 ( \10592 , \10591 , 1'b0 );
and \U$8605 ( \10593 , 1'b1 , \10592 );
and \U$8606 ( \10594 , \10585 , \10592 );
or \U$8607 ( \10595 , \10586 , \10593 , \10594 );
and \U$8608 ( \10596 , \10577 , \10595 );
xor \U$8610 ( \10597 , \10405 , 1'b0 );
xor \U$8611 ( \10598 , \10597 , \10420 );
and \U$8612 ( \10599 , \10595 , \10598 );
and \U$8613 ( \10600 , \10577 , \10598 );
or \U$8614 ( \10601 , \10596 , \10599 , \10600 );
xor \U$8616 ( \10602 , 1'b0 , \10422 );
xor \U$8617 ( \10603 , \10602 , \10439 );
and \U$8618 ( \10604 , \10601 , \10603 );
or \U$8619 ( \10605 , 1'b0 , 1'b0 , \10604 );
nand \U$8620 ( \10606 , \10462 , \10605 );
nor \U$8621 ( \10607 , \10462 , \10605 );
not \U$8622 ( \10608 , \10607 );
nand \U$8623 ( \10609 , \10606 , \10608 );
xor \U$8624 ( \10610 , \10086 , \10107 );
xor \U$8625 ( \10611 , \10610 , \10132 );
buf g339a_GF_PartitionCandidate( \10612_nG339a , \10611 );
buf \U$8626 ( \10613 , \10612_nG339a );
xor \U$8627 ( \10614 , \10110 , \10130 );
buf g337a_GF_PartitionCandidate( \10615_nG337a , \10614 );
buf \U$8628 ( \10616 , \10615_nG337a );
xor \U$8629 ( \10617 , \10613 , \10616 );
not \U$8630 ( \10618 , \10616 );
and \U$8631 ( \10619 , \10617 , \10618 );
and \U$8632 ( \10620 , \10550 , \10619 );
and \U$8633 ( \10621 , \10506 , \10616 );
nor \U$8634 ( \10622 , \10620 , \10621 );
xnor \U$8635 ( \10623 , \10622 , \10613 );
and \U$8636 ( \10624 , RI2b5e785c2bc0_255, \10242 );
and \U$8637 ( \10625 , RI2b5e785be480_275, \10248 );
and \U$8638 ( \10626 , RI2b5e785bc1d0_295, \10250 );
and \U$8639 ( \10627 , RI2b5e785ba2e0_315, \10252 );
and \U$8640 ( \10628 , RI2b5e785b9980_335, \10254 );
and \U$8641 ( \10629 , RI2b5e785b7e50_355, \10256 );
and \U$8642 ( \10630 , RI2b5e785b74f0_375, \10258 );
and \U$8643 ( \10631 , RI2b5e785b5d80_395, \10260 );
and \U$8644 ( \10632 , RI2b5e785b5420_415, \10262 );
and \U$8645 ( \10633 , RI2b5e785b4ac0_435, \10264 );
and \U$8646 ( \10634 , RI2b5e785b3710_455, \10266 );
and \U$8647 ( \10635 , RI2b5e785b2db0_475, \10268 );
and \U$8648 ( \10636 , RI2b5e785b2450_495, \10270 );
and \U$8649 ( \10637 , RI2b5e785b1460_515, \10272 );
and \U$8650 ( \10638 , RI2b5e785b0b00_535, \10274 );
and \U$8651 ( \10639 , RI2b5e785b01a0_555, \10276 );
and \U$8652 ( \10640 , RI2b5e785af570_575, \10278 );
or \U$8653 ( \10641 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 );
_DC g3c8c ( \10642_nG3c8c , \10641 , \10297 );
buf \U$8654 ( \10643 , \10642_nG3c8c );
xor \U$8655 ( \10644 , \10036 , \10057 );
xor \U$8656 ( \10645 , \10644 , \10138 );
buf g34d5_GF_PartitionCandidate( \10646_nG34d5 , \10645 );
buf \U$8657 ( \10647 , \10646_nG34d5 );
xor \U$8658 ( \10648 , \10061 , \10082 );
xor \U$8659 ( \10649 , \10648 , \10135 );
buf g34d9_GF_PartitionCandidate( \10650_nG34d9 , \10649 );
buf \U$8660 ( \10651 , \10650_nG34d9 );
xor \U$8661 ( \10652 , \10647 , \10651 );
xor \U$8662 ( \10653 , \10651 , \10613 );
not \U$8663 ( \10654 , \10653 );
and \U$8664 ( \10655 , \10652 , \10654 );
and \U$8665 ( \10656 , \10643 , \10655 );
and \U$8666 ( \10657 , RI2b5e785c2c38_254, \10242 );
and \U$8667 ( \10658 , RI2b5e785be4f8_274, \10248 );
and \U$8668 ( \10659 , RI2b5e785bc248_294, \10250 );
and \U$8669 ( \10660 , RI2b5e785ba358_314, \10252 );
and \U$8670 ( \10661 , RI2b5e785b99f8_334, \10254 );
and \U$8671 ( \10662 , RI2b5e785b7ec8_354, \10256 );
and \U$8672 ( \10663 , RI2b5e785b7568_374, \10258 );
and \U$8673 ( \10664 , RI2b5e785b5df8_394, \10260 );
and \U$8674 ( \10665 , RI2b5e785b5498_414, \10262 );
and \U$8675 ( \10666 , RI2b5e785b4b38_434, \10264 );
and \U$8676 ( \10667 , RI2b5e785b3788_454, \10266 );
and \U$8677 ( \10668 , RI2b5e785b2e28_474, \10268 );
and \U$8678 ( \10669 , RI2b5e785b24c8_494, \10270 );
and \U$8679 ( \10670 , RI2b5e785b14d8_514, \10272 );
and \U$8680 ( \10671 , RI2b5e785b0b78_534, \10274 );
and \U$8681 ( \10672 , RI2b5e785b0218_554, \10276 );
and \U$8682 ( \10673 , RI2b5e785af5e8_574, \10278 );
or \U$8683 ( \10674 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 );
_DC g3d60 ( \10675_nG3d60 , \10674 , \10297 );
buf \U$8684 ( \10676 , \10675_nG3d60 );
and \U$8685 ( \10677 , \10676 , \10653 );
nor \U$8686 ( \10678 , \10656 , \10677 );
and \U$8687 ( \10679 , \10651 , \10613 );
not \U$8688 ( \10680 , \10679 );
and \U$8689 ( \10681 , \10647 , \10680 );
xnor \U$8690 ( \10682 , \10678 , \10681 );
and \U$8691 ( \10683 , \10623 , \10682 );
and \U$8692 ( \10684 , RI2b5e785c0a00_257, \10242 );
and \U$8693 ( \10685 , RI2b5e785be390_277, \10248 );
and \U$8694 ( \10686 , RI2b5e785bc0e0_297, \10250 );
and \U$8695 ( \10687 , RI2b5e785ba1f0_317, \10252 );
and \U$8696 ( \10688 , RI2b5e785b9890_337, \10254 );
and \U$8697 ( \10689 , RI2b5e785b7d60_357, \10256 );
and \U$8698 ( \10690 , RI2b5e785b7400_377, \10258 );
and \U$8699 ( \10691 , RI2b5e785b5c90_397, \10260 );
and \U$8700 ( \10692 , RI2b5e785b5330_417, \10262 );
and \U$8701 ( \10693 , RI2b5e785b49d0_437, \10264 );
and \U$8702 ( \10694 , RI2b5e785b3620_457, \10266 );
and \U$8703 ( \10695 , RI2b5e785b2cc0_477, \10268 );
and \U$8704 ( \10696 , RI2b5e785b2360_497, \10270 );
and \U$8705 ( \10697 , RI2b5e785b1370_517, \10272 );
and \U$8706 ( \10698 , RI2b5e785b0a10_537, \10274 );
and \U$8707 ( \10699 , RI2b5e785b00b0_557, \10276 );
and \U$8708 ( \10700 , RI2b5e785af480_577, \10278 );
or \U$8709 ( \10701 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 );
_DC g3abf ( \10702_nG3abf , \10701 , \10297 );
buf \U$8710 ( \10703 , \10702_nG3abf );
xor \U$8711 ( \10704 , \9986 , \10007 );
xor \U$8712 ( \10705 , \10704 , \10144 );
buf g35ea_GF_PartitionCandidate( \10706_nG35ea , \10705 );
buf \U$8713 ( \10707 , \10706_nG35ea );
xor \U$8714 ( \10708 , \10011 , \10032 );
xor \U$8715 ( \10709 , \10708 , \10141 );
buf g35c6_GF_PartitionCandidate( \10710_nG35c6 , \10709 );
buf \U$8716 ( \10711 , \10710_nG35c6 );
xor \U$8717 ( \10712 , \10707 , \10711 );
xor \U$8718 ( \10713 , \10711 , \10647 );
not \U$8719 ( \10714 , \10713 );
and \U$8720 ( \10715 , \10712 , \10714 );
and \U$8721 ( \10716 , \10703 , \10715 );
and \U$8722 ( \10717 , RI2b5e785c2b48_256, \10242 );
and \U$8723 ( \10718 , RI2b5e785be408_276, \10248 );
and \U$8724 ( \10719 , RI2b5e785bc158_296, \10250 );
and \U$8725 ( \10720 , RI2b5e785ba268_316, \10252 );
and \U$8726 ( \10721 , RI2b5e785b9908_336, \10254 );
and \U$8727 ( \10722 , RI2b5e785b7dd8_356, \10256 );
and \U$8728 ( \10723 , RI2b5e785b7478_376, \10258 );
and \U$8729 ( \10724 , RI2b5e785b5d08_396, \10260 );
and \U$8730 ( \10725 , RI2b5e785b53a8_416, \10262 );
and \U$8731 ( \10726 , RI2b5e785b4a48_436, \10264 );
and \U$8732 ( \10727 , RI2b5e785b3698_456, \10266 );
and \U$8733 ( \10728 , RI2b5e785b2d38_476, \10268 );
and \U$8734 ( \10729 , RI2b5e785b23d8_496, \10270 );
and \U$8735 ( \10730 , RI2b5e785b13e8_516, \10272 );
and \U$8736 ( \10731 , RI2b5e785b0a88_536, \10274 );
and \U$8737 ( \10732 , RI2b5e785b0128_556, \10276 );
and \U$8738 ( \10733 , RI2b5e785af4f8_576, \10278 );
or \U$8739 ( \10734 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 );
_DC g3b96 ( \10735_nG3b96 , \10734 , \10297 );
buf \U$8740 ( \10736 , \10735_nG3b96 );
and \U$8741 ( \10737 , \10736 , \10713 );
nor \U$8742 ( \10738 , \10716 , \10737 );
and \U$8743 ( \10739 , \10711 , \10647 );
not \U$8744 ( \10740 , \10739 );
and \U$8745 ( \10741 , \10707 , \10740 );
xnor \U$8746 ( \10742 , \10738 , \10741 );
and \U$8747 ( \10743 , \10682 , \10742 );
and \U$8748 ( \10744 , \10623 , \10742 );
or \U$8749 ( \10745 , \10683 , \10743 , \10744 );
and \U$8750 ( \10746 , RI2b5e785c0910_259, \10242 );
and \U$8751 ( \10747 , RI2b5e785be2a0_279, \10248 );
and \U$8752 ( \10748 , RI2b5e785bbff0_299, \10250 );
and \U$8753 ( \10749 , RI2b5e785ba100_319, \10252 );
and \U$8754 ( \10750 , RI2b5e785b97a0_339, \10254 );
and \U$8755 ( \10751 , RI2b5e785b7c70_359, \10256 );
and \U$8756 ( \10752 , RI2b5e785b7310_379, \10258 );
and \U$8757 ( \10753 , RI2b5e785b5ba0_399, \10260 );
and \U$8758 ( \10754 , RI2b5e785b5240_419, \10262 );
and \U$8759 ( \10755 , RI2b5e785b48e0_439, \10264 );
and \U$8760 ( \10756 , RI2b5e785b3530_459, \10266 );
and \U$8761 ( \10757 , RI2b5e785b2bd0_479, \10268 );
and \U$8762 ( \10758 , RI2b5e785b2270_499, \10270 );
and \U$8763 ( \10759 , RI2b5e785b1280_519, \10272 );
and \U$8764 ( \10760 , RI2b5e785b0920_539, \10274 );
and \U$8765 ( \10761 , RI2b5e785affc0_559, \10276 );
and \U$8766 ( \10762 , RI2b5e785af390_579, \10278 );
or \U$8767 ( \10763 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 );
_DC g3900 ( \10764_nG3900 , \10763 , \10297 );
buf \U$8768 ( \10765 , \10764_nG3900 );
xor \U$8769 ( \10766 , \9961 , \9982 );
xor \U$8770 ( \10767 , \10766 , \10147 );
buf g3728_GF_PartitionCandidate( \10768_nG3728 , \10767 );
buf \U$8771 ( \10769 , \10768_nG3728 );
xor \U$8772 ( \10770 , \10471 , \10769 );
xor \U$8773 ( \10771 , \10769 , \10707 );
not \U$8774 ( \10772 , \10771 );
and \U$8775 ( \10773 , \10770 , \10772 );
and \U$8776 ( \10774 , \10765 , \10773 );
and \U$8777 ( \10775 , RI2b5e785c0988_258, \10242 );
and \U$8778 ( \10776 , RI2b5e785be318_278, \10248 );
and \U$8779 ( \10777 , RI2b5e785bc068_298, \10250 );
and \U$8780 ( \10778 , RI2b5e785ba178_318, \10252 );
and \U$8781 ( \10779 , RI2b5e785b9818_338, \10254 );
and \U$8782 ( \10780 , RI2b5e785b7ce8_358, \10256 );
and \U$8783 ( \10781 , RI2b5e785b7388_378, \10258 );
and \U$8784 ( \10782 , RI2b5e785b5c18_398, \10260 );
and \U$8785 ( \10783 , RI2b5e785b52b8_418, \10262 );
and \U$8786 ( \10784 , RI2b5e785b4958_438, \10264 );
and \U$8787 ( \10785 , RI2b5e785b35a8_458, \10266 );
and \U$8788 ( \10786 , RI2b5e785b2c48_478, \10268 );
and \U$8789 ( \10787 , RI2b5e785b22e8_498, \10270 );
and \U$8790 ( \10788 , RI2b5e785b12f8_518, \10272 );
and \U$8791 ( \10789 , RI2b5e785b0998_538, \10274 );
and \U$8792 ( \10790 , RI2b5e785b0038_558, \10276 );
and \U$8793 ( \10791 , RI2b5e785af408_578, \10278 );
or \U$8794 ( \10792 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 );
_DC g39c9 ( \10793_nG39c9 , \10792 , \10297 );
buf \U$8795 ( \10794 , \10793_nG39c9 );
and \U$8796 ( \10795 , \10794 , \10771 );
nor \U$8797 ( \10796 , \10774 , \10795 );
and \U$8798 ( \10797 , \10769 , \10707 );
not \U$8799 ( \10798 , \10797 );
and \U$8800 ( \10799 , \10471 , \10798 );
xnor \U$8801 ( \10800 , \10796 , \10799 );
and \U$8802 ( \10801 , RI2b5e785c0820_261, \10242 );
and \U$8803 ( \10802 , RI2b5e785be1b0_281, \10248 );
and \U$8804 ( \10803 , RI2b5e785bbf00_301, \10250 );
and \U$8805 ( \10804 , RI2b5e785ba010_321, \10252 );
and \U$8806 ( \10805 , RI2b5e785b96b0_341, \10254 );
and \U$8807 ( \10806 , RI2b5e785b7b80_361, \10256 );
and \U$8808 ( \10807 , RI2b5e785b7220_381, \10258 );
and \U$8809 ( \10808 , RI2b5e785b5ab0_401, \10260 );
and \U$8810 ( \10809 , RI2b5e785b5150_421, \10262 );
and \U$8811 ( \10810 , RI2b5e785b47f0_441, \10264 );
and \U$8812 ( \10811 , RI2b5e785b3440_461, \10266 );
and \U$8813 ( \10812 , RI2b5e785b2ae0_481, \10268 );
and \U$8814 ( \10813 , RI2b5e785b2180_501, \10270 );
and \U$8815 ( \10814 , RI2b5e785b1190_521, \10272 );
and \U$8816 ( \10815 , RI2b5e785b0830_541, \10274 );
and \U$8817 ( \10816 , RI2b5e785afed0_561, \10276 );
and \U$8818 ( \10817 , RI2b5e785af2a0_581, \10278 );
or \U$8819 ( \10818 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 );
_DC g3767 ( \10819_nG3767 , \10818 , \10297 );
buf \U$8820 ( \10820 , \10819_nG3767 );
and \U$8821 ( \10821 , \10820 , \10474 );
and \U$8822 ( \10822 , RI2b5e785c0898_260, \10242 );
and \U$8823 ( \10823 , RI2b5e785be228_280, \10248 );
and \U$8824 ( \10824 , RI2b5e785bbf78_300, \10250 );
and \U$8825 ( \10825 , RI2b5e785ba088_320, \10252 );
and \U$8826 ( \10826 , RI2b5e785b9728_340, \10254 );
and \U$8827 ( \10827 , RI2b5e785b7bf8_360, \10256 );
and \U$8828 ( \10828 , RI2b5e785b7298_380, \10258 );
and \U$8829 ( \10829 , RI2b5e785b5b28_400, \10260 );
and \U$8830 ( \10830 , RI2b5e785b51c8_420, \10262 );
and \U$8831 ( \10831 , RI2b5e785b4868_440, \10264 );
and \U$8832 ( \10832 , RI2b5e785b34b8_460, \10266 );
and \U$8833 ( \10833 , RI2b5e785b2b58_480, \10268 );
and \U$8834 ( \10834 , RI2b5e785b21f8_500, \10270 );
and \U$8835 ( \10835 , RI2b5e785b1208_520, \10272 );
and \U$8836 ( \10836 , RI2b5e785b08a8_540, \10274 );
and \U$8837 ( \10837 , RI2b5e785aff48_560, \10276 );
and \U$8838 ( \10838 , RI2b5e785af318_580, \10278 );
or \U$8839 ( \10839 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 );
_DC g381a ( \10840_nG381a , \10839 , \10297 );
buf \U$8840 ( \10841 , \10840_nG381a );
and \U$8841 ( \10842 , \10841 , \10472 );
nor \U$8842 ( \10843 , \10821 , \10842 );
xnor \U$8843 ( \10844 , \10843 , \10479 );
and \U$8844 ( \10845 , \10800 , \10844 );
and \U$8845 ( \10846 , RI2b5e785c0730_263, \10242 );
and \U$8846 ( \10847 , RI2b5e785be0c0_283, \10248 );
and \U$8847 ( \10848 , RI2b5e785bbe10_303, \10250 );
and \U$8848 ( \10849 , RI2b5e785b9f20_323, \10252 );
and \U$8849 ( \10850 , RI2b5e785b95c0_343, \10254 );
and \U$8850 ( \10851 , RI2b5e785b7a90_363, \10256 );
and \U$8851 ( \10852 , RI2b5e785b7130_383, \10258 );
and \U$8852 ( \10853 , RI2b5e785b59c0_403, \10260 );
and \U$8853 ( \10854 , RI2b5e785b5060_423, \10262 );
and \U$8854 ( \10855 , RI2b5e785b3cb0_443, \10264 );
and \U$8855 ( \10856 , RI2b5e785b3350_463, \10266 );
and \U$8856 ( \10857 , RI2b5e785b29f0_483, \10268 );
and \U$8857 ( \10858 , RI2b5e785b1a00_503, \10270 );
and \U$8858 ( \10859 , RI2b5e785b10a0_523, \10272 );
and \U$8859 ( \10860 , RI2b5e785b0740_543, \10274 );
and \U$8860 ( \10861 , RI2b5e785afde0_563, \10276 );
and \U$8861 ( \10862 , RI2b5e785af1b0_583, \10278 );
or \U$8862 ( \10863 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 );
_DC g3603 ( \10864_nG3603 , \10863 , \10297 );
buf \U$8863 ( \10865 , \10864_nG3603 );
and \U$8864 ( \10866 , \10865 , \10409 );
and \U$8865 ( \10867 , RI2b5e785c07a8_262, \10242 );
and \U$8866 ( \10868 , RI2b5e785be138_282, \10248 );
and \U$8867 ( \10869 , RI2b5e785bbe88_302, \10250 );
and \U$8868 ( \10870 , RI2b5e785b9f98_322, \10252 );
and \U$8869 ( \10871 , RI2b5e785b9638_342, \10254 );
and \U$8870 ( \10872 , RI2b5e785b7b08_362, \10256 );
and \U$8871 ( \10873 , RI2b5e785b71a8_382, \10258 );
and \U$8872 ( \10874 , RI2b5e785b5a38_402, \10260 );
and \U$8873 ( \10875 , RI2b5e785b50d8_422, \10262 );
and \U$8874 ( \10876 , RI2b5e785b4778_442, \10264 );
and \U$8875 ( \10877 , RI2b5e785b33c8_462, \10266 );
and \U$8876 ( \10878 , RI2b5e785b2a68_482, \10268 );
and \U$8877 ( \10879 , RI2b5e785b1a78_502, \10270 );
and \U$8878 ( \10880 , RI2b5e785b1118_522, \10272 );
and \U$8879 ( \10881 , RI2b5e785b07b8_542, \10274 );
and \U$8880 ( \10882 , RI2b5e785afe58_562, \10276 );
and \U$8881 ( \10883 , RI2b5e785af228_582, \10278 );
or \U$8882 ( \10884 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 );
_DC g36aa ( \10885_nG36aa , \10884 , \10297 );
buf \U$8883 ( \10886 , \10885_nG36aa );
and \U$8884 ( \10887 , \10886 , \10407 );
nor \U$8885 ( \10888 , \10866 , \10887 );
xnor \U$8886 ( \10889 , \10888 , \10176 );
and \U$8887 ( \10890 , \10844 , \10889 );
and \U$8888 ( \10891 , \10800 , \10889 );
or \U$8889 ( \10892 , \10845 , \10890 , \10891 );
and \U$8890 ( \10893 , \10745 , \10892 );
and \U$8891 ( \10894 , RI2b5e785c0640_265, \10242 );
and \U$8892 ( \10895 , RI2b5e785bdfd0_285, \10248 );
and \U$8893 ( \10896 , RI2b5e785bbd20_305, \10250 );
and \U$8894 ( \10897 , RI2b5e785b9e30_325, \10252 );
and \U$8895 ( \10898 , RI2b5e785b94d0_345, \10254 );
and \U$8896 ( \10899 , RI2b5e785b79a0_365, \10256 );
and \U$8897 ( \10900 , RI2b5e785b7040_385, \10258 );
and \U$8898 ( \10901 , RI2b5e785b58d0_405, \10260 );
and \U$8899 ( \10902 , RI2b5e785b4f70_425, \10262 );
and \U$8900 ( \10903 , RI2b5e785b3bc0_445, \10264 );
and \U$8901 ( \10904 , RI2b5e785b3260_465, \10266 );
and \U$8902 ( \10905 , RI2b5e785b2900_485, \10268 );
and \U$8903 ( \10906 , RI2b5e785b1910_505, \10270 );
and \U$8904 ( \10907 , RI2b5e785b0fb0_525, \10272 );
and \U$8905 ( \10908 , RI2b5e785b0650_545, \10274 );
and \U$8906 ( \10909 , RI2b5e785afcf0_565, \10276 );
and \U$8907 ( \10910 , RI2b5e785af0c0_585, \10278 );
or \U$8908 ( \10911 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 );
_DC g3493 ( \10912_nG3493 , \10911 , \10297 );
buf \U$8909 ( \10913 , \10912_nG3493 );
and \U$8910 ( \10914 , \10913 , \10347 );
and \U$8911 ( \10915 , RI2b5e785c06b8_264, \10242 );
and \U$8912 ( \10916 , RI2b5e785be048_284, \10248 );
and \U$8913 ( \10917 , RI2b5e785bbd98_304, \10250 );
and \U$8914 ( \10918 , RI2b5e785b9ea8_324, \10252 );
and \U$8915 ( \10919 , RI2b5e785b9548_344, \10254 );
and \U$8916 ( \10920 , RI2b5e785b7a18_364, \10256 );
and \U$8917 ( \10921 , RI2b5e785b70b8_384, \10258 );
and \U$8918 ( \10922 , RI2b5e785b5948_404, \10260 );
and \U$8919 ( \10923 , RI2b5e785b4fe8_424, \10262 );
and \U$8920 ( \10924 , RI2b5e785b3c38_444, \10264 );
and \U$8921 ( \10925 , RI2b5e785b32d8_464, \10266 );
and \U$8922 ( \10926 , RI2b5e785b2978_484, \10268 );
and \U$8923 ( \10927 , RI2b5e785b1988_504, \10270 );
and \U$8924 ( \10928 , RI2b5e785b1028_524, \10272 );
and \U$8925 ( \10929 , RI2b5e785b06c8_544, \10274 );
and \U$8926 ( \10930 , RI2b5e785afd68_564, \10276 );
and \U$8927 ( \10931 , RI2b5e785af138_584, \10278 );
or \U$8928 ( \10932 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 );
_DC g3564 ( \10933_nG3564 , \10932 , \10297 );
buf \U$8929 ( \10934 , \10933_nG3564 );
and \U$8930 ( \10935 , \10934 , \10345 );
nor \U$8931 ( \10936 , \10914 , \10935 );
xnor \U$8932 ( \10937 , \10936 , \10373 );
and \U$8934 ( \10938 , RI2b5e785c05c8_266, \10242 );
and \U$8935 ( \10939 , RI2b5e785bdf58_286, \10248 );
and \U$8936 ( \10940 , RI2b5e785bbca8_306, \10250 );
and \U$8937 ( \10941 , RI2b5e785b9db8_326, \10252 );
and \U$8938 ( \10942 , RI2b5e785b9458_346, \10254 );
and \U$8939 ( \10943 , RI2b5e785b7928_366, \10256 );
and \U$8940 ( \10944 , RI2b5e785b6fc8_386, \10258 );
and \U$8941 ( \10945 , RI2b5e785b5858_406, \10260 );
and \U$8942 ( \10946 , RI2b5e785b4ef8_426, \10262 );
and \U$8943 ( \10947 , RI2b5e785b3b48_446, \10264 );
and \U$8944 ( \10948 , RI2b5e785b31e8_466, \10266 );
and \U$8945 ( \10949 , RI2b5e785b2888_486, \10268 );
and \U$8946 ( \10950 , RI2b5e785b1898_506, \10270 );
and \U$8947 ( \10951 , RI2b5e785b0f38_526, \10272 );
and \U$8948 ( \10952 , RI2b5e785b05d8_546, \10274 );
and \U$8949 ( \10953 , RI2b5e785afc78_566, \10276 );
and \U$8950 ( \10954 , RI2b5e785af048_586, \10278 );
or \U$8951 ( \10955 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 );
_DC g3451 ( \10956_nG3451 , \10955 , \10297 );
buf \U$8952 ( \10957 , \10956_nG3451 );
and \U$8953 ( \10958 , \10957 , \10400 );
nor \U$8954 ( \10959 , 1'b0 , \10958 );
xnor \U$8955 ( \10960 , \10959 , 1'b0 );
and \U$8956 ( \10961 , \10937 , \10960 );
and \U$8957 ( \10962 , \10892 , \10961 );
and \U$8958 ( \10963 , \10745 , \10961 );
or \U$8959 ( \10964 , \10893 , \10962 , \10963 );
and \U$8961 ( \10965 , \10886 , \10409 );
and \U$8962 ( \10966 , \10820 , \10407 );
nor \U$8963 ( \10967 , \10965 , \10966 );
xnor \U$8964 ( \10968 , \10967 , \10176 );
and \U$8965 ( \10969 , \10934 , \10347 );
and \U$8966 ( \10970 , \10865 , \10345 );
nor \U$8967 ( \10971 , \10969 , \10970 );
xnor \U$8968 ( \10972 , \10971 , \10373 );
xor \U$8969 ( \10973 , \10968 , \10972 );
and \U$8971 ( \10974 , \10913 , \10400 );
nor \U$8972 ( \10975 , 1'b0 , \10974 );
xnor \U$8973 ( \10976 , \10975 , 1'b0 );
xor \U$8974 ( \10977 , \10973 , \10976 );
and \U$8975 ( \10978 , \10736 , \10715 );
and \U$8976 ( \10979 , \10643 , \10713 );
nor \U$8977 ( \10980 , \10978 , \10979 );
xnor \U$8978 ( \10981 , \10980 , \10741 );
and \U$8979 ( \10982 , \10794 , \10773 );
and \U$8980 ( \10983 , \10703 , \10771 );
nor \U$8981 ( \10984 , \10982 , \10983 );
xnor \U$8982 ( \10985 , \10984 , \10799 );
xor \U$8983 ( \10986 , \10981 , \10985 );
and \U$8984 ( \10987 , \10841 , \10474 );
and \U$8985 ( \10988 , \10765 , \10472 );
nor \U$8986 ( \10989 , \10987 , \10988 );
xnor \U$8987 ( \10990 , \10989 , \10479 );
xor \U$8988 ( \10991 , \10986 , \10990 );
and \U$8989 ( \10992 , \10977 , \10991 );
or \U$8991 ( \10993 , 1'b0 , \10992 , 1'b0 );
xor \U$8992 ( \10994 , \10964 , \10993 );
and \U$8993 ( \10995 , \10865 , \10347 );
and \U$8994 ( \10996 , \10886 , \10345 );
nor \U$8995 ( \10997 , \10995 , \10996 );
xnor \U$8996 ( \10998 , \10997 , \10373 );
and \U$8998 ( \10999 , \10934 , \10400 );
nor \U$8999 ( \11000 , 1'b0 , \10999 );
xnor \U$9000 ( \11001 , \11000 , 1'b0 );
xor \U$9001 ( \11002 , \10998 , \11001 );
xor \U$9003 ( \11003 , \11002 , 1'b0 );
and \U$9004 ( \11004 , \10703 , \10773 );
and \U$9005 ( \11005 , \10736 , \10771 );
nor \U$9006 ( \11006 , \11004 , \11005 );
xnor \U$9007 ( \11007 , \11006 , \10799 );
and \U$9008 ( \11008 , \10765 , \10474 );
and \U$9009 ( \11009 , \10794 , \10472 );
nor \U$9010 ( \11010 , \11008 , \11009 );
xnor \U$9011 ( \11011 , \11010 , \10479 );
xor \U$9012 ( \11012 , \11007 , \11011 );
and \U$9013 ( \11013 , \10820 , \10409 );
and \U$9014 ( \11014 , \10841 , \10407 );
nor \U$9015 ( \11015 , \11013 , \11014 );
xnor \U$9016 ( \11016 , \11015 , \10176 );
xor \U$9017 ( \11017 , \11012 , \11016 );
xor \U$9018 ( \11018 , \11003 , \11017 );
and \U$9019 ( \11019 , \10527 , \10619 );
and \U$9020 ( \11020 , \10395 , \10616 );
nor \U$9021 ( \11021 , \11019 , \11020 );
xnor \U$9022 ( \11022 , \11021 , \10613 );
and \U$9023 ( \11023 , \10550 , \10655 );
and \U$9024 ( \11024 , \10506 , \10653 );
nor \U$9025 ( \11025 , \11023 , \11024 );
xnor \U$9026 ( \11026 , \11025 , \10681 );
xor \U$9027 ( \11027 , \11022 , \11026 );
and \U$9028 ( \11028 , \10643 , \10715 );
and \U$9029 ( \11029 , \10676 , \10713 );
nor \U$9030 ( \11030 , \11028 , \11029 );
xnor \U$9031 ( \11031 , \11030 , \10741 );
xor \U$9032 ( \11032 , \11027 , \11031 );
xor \U$9033 ( \11033 , \11018 , \11032 );
xor \U$9034 ( \11034 , \10994 , \11033 );
and \U$9036 ( \11035 , \10676 , \10619 );
and \U$9037 ( \11036 , \10550 , \10616 );
nor \U$9038 ( \11037 , \11035 , \11036 );
xnor \U$9039 ( \11038 , \11037 , \10613 );
and \U$9040 ( \11039 , \10736 , \10655 );
and \U$9041 ( \11040 , \10643 , \10653 );
nor \U$9042 ( \11041 , \11039 , \11040 );
xnor \U$9043 ( \11042 , \11041 , \10681 );
and \U$9044 ( \11043 , \11038 , \11042 );
or \U$9046 ( \11044 , 1'b0 , \11043 , 1'b0 );
and \U$9047 ( \11045 , \10794 , \10715 );
and \U$9048 ( \11046 , \10703 , \10713 );
nor \U$9049 ( \11047 , \11045 , \11046 );
xnor \U$9050 ( \11048 , \11047 , \10741 );
and \U$9051 ( \11049 , \10841 , \10773 );
and \U$9052 ( \11050 , \10765 , \10771 );
nor \U$9053 ( \11051 , \11049 , \11050 );
xnor \U$9054 ( \11052 , \11051 , \10799 );
and \U$9055 ( \11053 , \11048 , \11052 );
and \U$9056 ( \11054 , \10886 , \10474 );
and \U$9057 ( \11055 , \10820 , \10472 );
nor \U$9058 ( \11056 , \11054 , \11055 );
xnor \U$9059 ( \11057 , \11056 , \10479 );
and \U$9060 ( \11058 , \11052 , \11057 );
and \U$9061 ( \11059 , \11048 , \11057 );
or \U$9062 ( \11060 , \11053 , \11058 , \11059 );
and \U$9063 ( \11061 , \11044 , \11060 );
and \U$9064 ( \11062 , \10934 , \10409 );
and \U$9065 ( \11063 , \10865 , \10407 );
nor \U$9066 ( \11064 , \11062 , \11063 );
xnor \U$9067 ( \11065 , \11064 , \10176 );
and \U$9068 ( \11066 , \10957 , \10347 );
and \U$9069 ( \11067 , \10913 , \10345 );
nor \U$9070 ( \11068 , \11066 , \11067 );
xnor \U$9071 ( \11069 , \11068 , \10373 );
and \U$9072 ( \11070 , \11065 , \11069 );
and \U$9073 ( \11071 , RI2b5e785c0550_267, \10242 );
and \U$9074 ( \11072 , RI2b5e785bc590_287, \10248 );
and \U$9075 ( \11073 , RI2b5e785bbc30_307, \10250 );
and \U$9076 ( \11074 , RI2b5e785b9d40_327, \10252 );
and \U$9077 ( \11075 , RI2b5e785b93e0_347, \10254 );
and \U$9078 ( \11076 , RI2b5e785b78b0_367, \10256 );
and \U$9079 ( \11077 , RI2b5e785b6f50_387, \10258 );
and \U$9080 ( \11078 , RI2b5e785b57e0_407, \10260 );
and \U$9081 ( \11079 , RI2b5e785b4e80_427, \10262 );
and \U$9082 ( \11080 , RI2b5e785b3ad0_447, \10264 );
and \U$9083 ( \11081 , RI2b5e785b3170_467, \10266 );
and \U$9084 ( \11082 , RI2b5e785b2810_487, \10268 );
and \U$9085 ( \11083 , RI2b5e785b1820_507, \10270 );
and \U$9086 ( \11084 , RI2b5e785b0ec0_527, \10272 );
and \U$9087 ( \11085 , RI2b5e785b0560_547, \10274 );
and \U$9088 ( \11086 , RI2b5e785afc00_567, \10276 );
and \U$9089 ( \11087 , RI2b5e785aefd0_587, \10278 );
or \U$9090 ( \11088 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 );
_DC g333d ( \11089_nG333d , \11088 , \10297 );
buf \U$9091 ( \11090 , \11089_nG333d );
nand \U$9092 ( \11091 , \11090 , \10400 );
xnor \U$9093 ( \11092 , \11091 , 1'b0 );
and \U$9094 ( \11093 , \11069 , \11092 );
and \U$9095 ( \11094 , \11065 , \11092 );
or \U$9096 ( \11095 , \11070 , \11093 , \11094 );
and \U$9097 ( \11096 , \11060 , \11095 );
and \U$9098 ( \11097 , \11044 , \11095 );
or \U$9099 ( \11098 , \11061 , \11096 , \11097 );
xor \U$9100 ( \11099 , \10937 , \10960 );
xor \U$9101 ( \11100 , \10800 , \10844 );
xor \U$9102 ( \11101 , \11100 , \10889 );
and \U$9103 ( \11102 , \11099 , \11101 );
xor \U$9104 ( \11103 , \10623 , \10682 );
xor \U$9105 ( \11104 , \11103 , \10742 );
and \U$9106 ( \11105 , \11101 , \11104 );
and \U$9107 ( \11106 , \11099 , \11104 );
or \U$9108 ( \11107 , \11102 , \11105 , \11106 );
and \U$9109 ( \11108 , \11098 , \11107 );
and \U$9111 ( \11109 , \10506 , \10619 );
and \U$9112 ( \11110 , \10527 , \10616 );
nor \U$9113 ( \11111 , \11109 , \11110 );
xnor \U$9114 ( \11112 , \11111 , \10613 );
xor \U$9115 ( \11113 , 1'b0 , \11112 );
and \U$9116 ( \11114 , \10676 , \10655 );
and \U$9117 ( \11115 , \10550 , \10653 );
nor \U$9118 ( \11116 , \11114 , \11115 );
xnor \U$9119 ( \11117 , \11116 , \10681 );
xor \U$9120 ( \11118 , \11113 , \11117 );
and \U$9121 ( \11119 , \11107 , \11118 );
and \U$9122 ( \11120 , \11098 , \11118 );
or \U$9123 ( \11121 , \11108 , \11119 , \11120 );
xor \U$9125 ( \11122 , 1'b0 , \10977 );
xor \U$9126 ( \11123 , \11122 , \10991 );
xor \U$9127 ( \11124 , \10745 , \10892 );
xor \U$9128 ( \11125 , \11124 , \10961 );
and \U$9129 ( \11126 , \11123 , \11125 );
xor \U$9130 ( \11127 , \11121 , \11126 );
and \U$9132 ( \11128 , \11112 , \11117 );
or \U$9134 ( \11129 , 1'b0 , \11128 , 1'b0 );
and \U$9135 ( \11130 , \10981 , \10985 );
and \U$9136 ( \11131 , \10985 , \10990 );
and \U$9137 ( \11132 , \10981 , \10990 );
or \U$9138 ( \11133 , \11130 , \11131 , \11132 );
xor \U$9139 ( \11134 , \11129 , \11133 );
and \U$9140 ( \11135 , \10968 , \10972 );
and \U$9141 ( \11136 , \10972 , \10976 );
and \U$9142 ( \11137 , \10968 , \10976 );
or \U$9143 ( \11138 , \11135 , \11136 , \11137 );
xor \U$9144 ( \11139 , \11134 , \11138 );
xor \U$9145 ( \11140 , \11127 , \11139 );
xor \U$9146 ( \11141 , \11034 , \11140 );
and \U$9147 ( \11142 , \10643 , \10619 );
and \U$9148 ( \11143 , \10676 , \10616 );
nor \U$9149 ( \11144 , \11142 , \11143 );
xnor \U$9150 ( \11145 , \11144 , \10613 );
and \U$9151 ( \11146 , \10703 , \10655 );
and \U$9152 ( \11147 , \10736 , \10653 );
nor \U$9153 ( \11148 , \11146 , \11147 );
xnor \U$9154 ( \11149 , \11148 , \10681 );
and \U$9155 ( \11150 , \11145 , \11149 );
and \U$9156 ( \11151 , \10765 , \10715 );
and \U$9157 ( \11152 , \10794 , \10713 );
nor \U$9158 ( \11153 , \11151 , \11152 );
xnor \U$9159 ( \11154 , \11153 , \10741 );
and \U$9160 ( \11155 , \11149 , \11154 );
and \U$9161 ( \11156 , \11145 , \11154 );
or \U$9162 ( \11157 , \11150 , \11155 , \11156 );
and \U$9163 ( \11158 , \10820 , \10773 );
and \U$9164 ( \11159 , \10841 , \10771 );
nor \U$9165 ( \11160 , \11158 , \11159 );
xnor \U$9166 ( \11161 , \11160 , \10799 );
and \U$9167 ( \11162 , \10865 , \10474 );
and \U$9168 ( \11163 , \10886 , \10472 );
nor \U$9169 ( \11164 , \11162 , \11163 );
xnor \U$9170 ( \11165 , \11164 , \10479 );
and \U$9171 ( \11166 , \11161 , \11165 );
and \U$9172 ( \11167 , \10913 , \10409 );
and \U$9173 ( \11168 , \10934 , \10407 );
nor \U$9174 ( \11169 , \11167 , \11168 );
xnor \U$9175 ( \11170 , \11169 , \10176 );
and \U$9176 ( \11171 , \11165 , \11170 );
and \U$9177 ( \11172 , \11161 , \11170 );
or \U$9178 ( \11173 , \11166 , \11171 , \11172 );
and \U$9179 ( \11174 , \11157 , \11173 );
xor \U$9180 ( \11175 , \11065 , \11069 );
xor \U$9181 ( \11176 , \11175 , \11092 );
and \U$9182 ( \11177 , \11173 , \11176 );
and \U$9183 ( \11178 , \11157 , \11176 );
or \U$9184 ( \11179 , \11174 , \11177 , \11178 );
xor \U$9185 ( \11180 , \11048 , \11052 );
xor \U$9186 ( \11181 , \11180 , \11057 );
xor \U$9187 ( \11182 , 1'b0 , \11038 );
xor \U$9188 ( \11183 , \11182 , \11042 );
and \U$9189 ( \11184 , \11181 , \11183 );
and \U$9190 ( \11185 , \11179 , \11184 );
xor \U$9191 ( \11186 , \11099 , \11101 );
xor \U$9192 ( \11187 , \11186 , \11104 );
and \U$9193 ( \11188 , \11184 , \11187 );
and \U$9194 ( \11189 , \11179 , \11187 );
or \U$9195 ( \11190 , \11185 , \11188 , \11189 );
xor \U$9196 ( \11191 , \11123 , \11125 );
and \U$9197 ( \11192 , \11190 , \11191 );
xor \U$9198 ( \11193 , \11098 , \11107 );
xor \U$9199 ( \11194 , \11193 , \11118 );
and \U$9200 ( \11195 , \11191 , \11194 );
and \U$9201 ( \11196 , \11190 , \11194 );
or \U$9202 ( \11197 , \11192 , \11195 , \11196 );
nor \U$9203 ( \11198 , \11141 , \11197 );
and \U$9204 ( \11199 , \11121 , \11126 );
and \U$9205 ( \11200 , \11126 , \11139 );
and \U$9206 ( \11201 , \11121 , \11139 );
or \U$9207 ( \11202 , \11199 , \11200 , \11201 );
and \U$9208 ( \11203 , \10964 , \10993 );
and \U$9209 ( \11204 , \10993 , \11033 );
and \U$9210 ( \11205 , \10964 , \11033 );
or \U$9211 ( \11206 , \11203 , \11204 , \11205 );
and \U$9213 ( \11207 , \10395 , \10619 );
and \U$9214 ( \11208 , \10299 , \10616 );
nor \U$9215 ( \11209 , \11207 , \11208 );
xnor \U$9216 ( \11210 , \11209 , \10613 );
xor \U$9217 ( \11211 , 1'b0 , \11210 );
and \U$9218 ( \11212 , \10506 , \10655 );
and \U$9219 ( \11213 , \10527 , \10653 );
nor \U$9220 ( \11214 , \11212 , \11213 );
xnor \U$9221 ( \11215 , \11214 , \10681 );
xor \U$9222 ( \11216 , \11211 , \11215 );
and \U$9224 ( \11217 , \10841 , \10409 );
and \U$9225 ( \11218 , \10765 , \10407 );
nor \U$9226 ( \11219 , \11217 , \11218 );
xnor \U$9227 ( \11220 , \11219 , \10176 );
and \U$9228 ( \11221 , \10886 , \10347 );
and \U$9229 ( \11222 , \10820 , \10345 );
nor \U$9230 ( \11223 , \11221 , \11222 );
xnor \U$9231 ( \11224 , \11223 , \10373 );
xor \U$9232 ( \11225 , \11220 , \11224 );
and \U$9234 ( \11226 , \10865 , \10400 );
nor \U$9235 ( \11227 , 1'b0 , \11226 );
xnor \U$9236 ( \11228 , \11227 , 1'b0 );
xor \U$9237 ( \11229 , \11225 , \11228 );
xor \U$9238 ( \11230 , 1'b0 , \11229 );
xor \U$9239 ( \11231 , \11216 , \11230 );
and \U$9240 ( \11232 , \11022 , \11026 );
and \U$9241 ( \11233 , \11026 , \11031 );
and \U$9242 ( \11234 , \11022 , \11031 );
or \U$9243 ( \11235 , \11232 , \11233 , \11234 );
and \U$9244 ( \11236 , \11007 , \11011 );
and \U$9245 ( \11237 , \11011 , \11016 );
and \U$9246 ( \11238 , \11007 , \11016 );
or \U$9247 ( \11239 , \11236 , \11237 , \11238 );
xor \U$9248 ( \11240 , \11235 , \11239 );
and \U$9249 ( \11241 , \10998 , \11001 );
or \U$9252 ( \11242 , \11241 , 1'b0 , 1'b0 );
xor \U$9253 ( \11243 , \11240 , \11242 );
xor \U$9254 ( \11244 , \11231 , \11243 );
xor \U$9255 ( \11245 , \11206 , \11244 );
and \U$9256 ( \11246 , \11129 , \11133 );
and \U$9257 ( \11247 , \11133 , \11138 );
and \U$9258 ( \11248 , \11129 , \11138 );
or \U$9259 ( \11249 , \11246 , \11247 , \11248 );
and \U$9260 ( \11250 , \11003 , \11017 );
and \U$9261 ( \11251 , \11017 , \11032 );
and \U$9262 ( \11252 , \11003 , \11032 );
or \U$9263 ( \11253 , \11250 , \11251 , \11252 );
xor \U$9264 ( \11254 , \11249 , \11253 );
and \U$9265 ( \11255 , \10676 , \10715 );
and \U$9266 ( \11256 , \10550 , \10713 );
nor \U$9267 ( \11257 , \11255 , \11256 );
xnor \U$9268 ( \11258 , \11257 , \10741 );
and \U$9269 ( \11259 , \10736 , \10773 );
and \U$9270 ( \11260 , \10643 , \10771 );
nor \U$9271 ( \11261 , \11259 , \11260 );
xnor \U$9272 ( \11262 , \11261 , \10799 );
xor \U$9273 ( \11263 , \11258 , \11262 );
and \U$9274 ( \11264 , \10794 , \10474 );
and \U$9275 ( \11265 , \10703 , \10472 );
nor \U$9276 ( \11266 , \11264 , \11265 );
xnor \U$9277 ( \11267 , \11266 , \10479 );
xor \U$9278 ( \11268 , \11263 , \11267 );
xor \U$9279 ( \11269 , \11254 , \11268 );
xor \U$9280 ( \11270 , \11245 , \11269 );
xor \U$9281 ( \11271 , \11202 , \11270 );
and \U$9282 ( \11272 , \11034 , \11140 );
nor \U$9283 ( \11273 , \11271 , \11272 );
nor \U$9284 ( \11274 , \11198 , \11273 );
and \U$9285 ( \11275 , \11206 , \11244 );
and \U$9286 ( \11276 , \11244 , \11269 );
and \U$9287 ( \11277 , \11206 , \11269 );
or \U$9288 ( \11278 , \11275 , \11276 , \11277 );
and \U$9290 ( \11279 , \11210 , \11215 );
or \U$9292 ( \11280 , 1'b0 , \11279 , 1'b0 );
and \U$9293 ( \11281 , \11258 , \11262 );
and \U$9294 ( \11282 , \11262 , \11267 );
and \U$9295 ( \11283 , \11258 , \11267 );
or \U$9296 ( \11284 , \11281 , \11282 , \11283 );
xor \U$9297 ( \11285 , \11280 , \11284 );
and \U$9298 ( \11286 , \11220 , \11224 );
and \U$9299 ( \11287 , \11224 , \11228 );
and \U$9300 ( \11288 , \11220 , \11228 );
or \U$9301 ( \11289 , \11286 , \11287 , \11288 );
xor \U$9302 ( \11290 , \11285 , \11289 );
and \U$9303 ( \11291 , \11235 , \11239 );
and \U$9304 ( \11292 , \11239 , \11242 );
and \U$9305 ( \11293 , \11235 , \11242 );
or \U$9306 ( \11294 , \11291 , \11292 , \11293 );
xor \U$9308 ( \11295 , \11294 , 1'b0 );
and \U$9309 ( \11296 , \10299 , \10619 );
and \U$9310 ( \11297 , \10368 , \10616 );
nor \U$9311 ( \11298 , \11296 , \11297 );
xnor \U$9312 ( \11299 , \11298 , \10613 );
and \U$9313 ( \11300 , \10527 , \10655 );
and \U$9314 ( \11301 , \10395 , \10653 );
nor \U$9315 ( \11302 , \11300 , \11301 );
xnor \U$9316 ( \11303 , \11302 , \10681 );
xor \U$9317 ( \11304 , \11299 , \11303 );
and \U$9318 ( \11305 , \10550 , \10715 );
and \U$9319 ( \11306 , \10506 , \10713 );
nor \U$9320 ( \11307 , \11305 , \11306 );
xnor \U$9321 ( \11308 , \11307 , \10741 );
xor \U$9322 ( \11309 , \11304 , \11308 );
xor \U$9323 ( \11310 , \11295 , \11309 );
xor \U$9324 ( \11311 , \11290 , \11310 );
xor \U$9325 ( \11312 , \11278 , \11311 );
and \U$9326 ( \11313 , \11249 , \11253 );
and \U$9327 ( \11314 , \11253 , \11268 );
and \U$9328 ( \11315 , \11249 , \11268 );
or \U$9329 ( \11316 , \11313 , \11314 , \11315 );
and \U$9330 ( \11317 , \11216 , \11230 );
and \U$9331 ( \11318 , \11230 , \11243 );
and \U$9332 ( \11319 , \11216 , \11243 );
or \U$9333 ( \11320 , \11317 , \11318 , \11319 );
xor \U$9334 ( \11321 , \11316 , \11320 );
and \U$9336 ( \11322 , \10820 , \10347 );
and \U$9337 ( \11323 , \10841 , \10345 );
nor \U$9338 ( \11324 , \11322 , \11323 );
xnor \U$9339 ( \11325 , \11324 , \10373 );
and \U$9341 ( \11326 , \10886 , \10400 );
nor \U$9342 ( \11327 , 1'b0 , \11326 );
xnor \U$9343 ( \11328 , \11327 , 1'b0 );
xor \U$9344 ( \11329 , \11325 , \11328 );
xor \U$9346 ( \11330 , \11329 , 1'b0 );
xor \U$9347 ( \11331 , 1'b0 , \11330 );
and \U$9348 ( \11332 , \10643 , \10773 );
and \U$9349 ( \11333 , \10676 , \10771 );
nor \U$9350 ( \11334 , \11332 , \11333 );
xnor \U$9351 ( \11335 , \11334 , \10799 );
and \U$9352 ( \11336 , \10703 , \10474 );
and \U$9353 ( \11337 , \10736 , \10472 );
nor \U$9354 ( \11338 , \11336 , \11337 );
xnor \U$9355 ( \11339 , \11338 , \10479 );
xor \U$9356 ( \11340 , \11335 , \11339 );
and \U$9357 ( \11341 , \10765 , \10409 );
and \U$9358 ( \11342 , \10794 , \10407 );
nor \U$9359 ( \11343 , \11341 , \11342 );
xnor \U$9360 ( \11344 , \11343 , \10176 );
xor \U$9361 ( \11345 , \11340 , \11344 );
xor \U$9362 ( \11346 , \11331 , \11345 );
xor \U$9363 ( \11347 , \11321 , \11346 );
xor \U$9364 ( \11348 , \11312 , \11347 );
and \U$9365 ( \11349 , \11202 , \11270 );
nor \U$9366 ( \11350 , \11348 , \11349 );
and \U$9367 ( \11351 , \11316 , \11320 );
and \U$9368 ( \11352 , \11320 , \11346 );
and \U$9369 ( \11353 , \11316 , \11346 );
or \U$9370 ( \11354 , \11351 , \11352 , \11353 );
and \U$9371 ( \11355 , \11290 , \11310 );
xor \U$9372 ( \11356 , \11354 , \11355 );
and \U$9375 ( \11357 , \11294 , \11309 );
or \U$9376 ( \11358 , 1'b0 , 1'b0 , \11357 );
and \U$9378 ( \11359 , \10794 , \10409 );
and \U$9379 ( \11360 , \10703 , \10407 );
nor \U$9380 ( \11361 , \11359 , \11360 );
xnor \U$9381 ( \11362 , \11361 , \10176 );
and \U$9382 ( \11363 , \10841 , \10347 );
and \U$9383 ( \11364 , \10765 , \10345 );
nor \U$9384 ( \11365 , \11363 , \11364 );
xnor \U$9385 ( \11366 , \11365 , \10373 );
xor \U$9386 ( \11367 , \11362 , \11366 );
and \U$9388 ( \11368 , \10820 , \10400 );
nor \U$9389 ( \11369 , 1'b0 , \11368 );
xnor \U$9390 ( \11370 , \11369 , 1'b0 );
xor \U$9391 ( \11371 , \11367 , \11370 );
xor \U$9392 ( \11372 , 1'b0 , \11371 );
and \U$9393 ( \11373 , \10506 , \10715 );
and \U$9394 ( \11374 , \10527 , \10713 );
nor \U$9395 ( \11375 , \11373 , \11374 );
xnor \U$9396 ( \11376 , \11375 , \10741 );
and \U$9397 ( \11377 , \10676 , \10773 );
and \U$9398 ( \11378 , \10550 , \10771 );
nor \U$9399 ( \11379 , \11377 , \11378 );
xnor \U$9400 ( \11380 , \11379 , \10799 );
xor \U$9401 ( \11381 , \11376 , \11380 );
and \U$9402 ( \11382 , \10736 , \10474 );
and \U$9403 ( \11383 , \10643 , \10472 );
nor \U$9404 ( \11384 , \11382 , \11383 );
xnor \U$9405 ( \11385 , \11384 , \10479 );
xor \U$9406 ( \11386 , \11381 , \11385 );
xor \U$9407 ( \11387 , \11372 , \11386 );
and \U$9408 ( \11388 , \11299 , \11303 );
and \U$9409 ( \11389 , \11303 , \11308 );
and \U$9410 ( \11390 , \11299 , \11308 );
or \U$9411 ( \11391 , \11388 , \11389 , \11390 );
and \U$9412 ( \11392 , \11335 , \11339 );
and \U$9413 ( \11393 , \11339 , \11344 );
and \U$9414 ( \11394 , \11335 , \11344 );
or \U$9415 ( \11395 , \11392 , \11393 , \11394 );
xor \U$9416 ( \11396 , \11391 , \11395 );
and \U$9417 ( \11397 , \11325 , \11328 );
or \U$9420 ( \11398 , \11397 , 1'b0 , 1'b0 );
xor \U$9421 ( \11399 , \11396 , \11398 );
xor \U$9422 ( \11400 , \11387 , \11399 );
xor \U$9423 ( \11401 , \11358 , \11400 );
and \U$9424 ( \11402 , \11280 , \11284 );
and \U$9425 ( \11403 , \11284 , \11289 );
and \U$9426 ( \11404 , \11280 , \11289 );
or \U$9427 ( \11405 , \11402 , \11403 , \11404 );
and \U$9429 ( \11406 , \11330 , \11345 );
or \U$9431 ( \11407 , 1'b0 , \11406 , 1'b0 );
xor \U$9432 ( \11408 , \11405 , \11407 );
and \U$9434 ( \11409 , \10368 , \10619 );
not \U$9435 ( \11410 , \11409 );
xnor \U$9436 ( \11411 , \11410 , \10613 );
xor \U$9437 ( \11412 , 1'b0 , \11411 );
and \U$9438 ( \11413 , \10395 , \10655 );
and \U$9439 ( \11414 , \10299 , \10653 );
nor \U$9440 ( \11415 , \11413 , \11414 );
xnor \U$9441 ( \11416 , \11415 , \10681 );
xor \U$9442 ( \11417 , \11412 , \11416 );
xor \U$9443 ( \11418 , \11408 , \11417 );
xor \U$9444 ( \11419 , \11401 , \11418 );
xor \U$9445 ( \11420 , \11356 , \11419 );
and \U$9446 ( \11421 , \11278 , \11311 );
and \U$9447 ( \11422 , \11311 , \11347 );
and \U$9448 ( \11423 , \11278 , \11347 );
or \U$9449 ( \11424 , \11421 , \11422 , \11423 );
nor \U$9450 ( \11425 , \11420 , \11424 );
nor \U$9451 ( \11426 , \11350 , \11425 );
nand \U$9452 ( \11427 , \11274 , \11426 );
and \U$9453 ( \11428 , \11358 , \11400 );
and \U$9454 ( \11429 , \11400 , \11418 );
and \U$9455 ( \11430 , \11358 , \11418 );
or \U$9456 ( \11431 , \11428 , \11429 , \11430 );
and \U$9457 ( \11432 , \11391 , \11395 );
and \U$9458 ( \11433 , \11395 , \11398 );
and \U$9459 ( \11434 , \11391 , \11398 );
or \U$9460 ( \11435 , \11432 , \11433 , \11434 );
and \U$9462 ( \11436 , \11371 , \11386 );
or \U$9464 ( \11437 , 1'b0 , \11436 , 1'b0 );
xor \U$9465 ( \11438 , \11435 , \11437 );
and \U$9466 ( \11439 , \10550 , \10773 );
and \U$9467 ( \11440 , \10506 , \10771 );
nor \U$9468 ( \11441 , \11439 , \11440 );
xnor \U$9469 ( \11442 , \11441 , \10799 );
and \U$9470 ( \11443 , \10643 , \10474 );
and \U$9471 ( \11444 , \10676 , \10472 );
nor \U$9472 ( \11445 , \11443 , \11444 );
xnor \U$9473 ( \11446 , \11445 , \10479 );
xor \U$9474 ( \11447 , \11442 , \11446 );
and \U$9475 ( \11448 , \10703 , \10409 );
and \U$9476 ( \11449 , \10736 , \10407 );
nor \U$9477 ( \11450 , \11448 , \11449 );
xnor \U$9478 ( \11451 , \11450 , \10176 );
xor \U$9479 ( \11452 , \11447 , \11451 );
xor \U$9480 ( \11453 , \11438 , \11452 );
xor \U$9481 ( \11454 , \11431 , \11453 );
and \U$9482 ( \11455 , \11405 , \11407 );
and \U$9483 ( \11456 , \11407 , \11417 );
and \U$9484 ( \11457 , \11405 , \11417 );
or \U$9485 ( \11458 , \11455 , \11456 , \11457 );
and \U$9486 ( \11459 , \11387 , \11399 );
xor \U$9487 ( \11460 , \11458 , \11459 );
not \U$9488 ( \11461 , \10613 );
and \U$9489 ( \11462 , \10299 , \10655 );
and \U$9490 ( \11463 , \10368 , \10653 );
nor \U$9491 ( \11464 , \11462 , \11463 );
xnor \U$9492 ( \11465 , \11464 , \10681 );
xor \U$9493 ( \11466 , \11461 , \11465 );
and \U$9494 ( \11467 , \10527 , \10715 );
and \U$9495 ( \11468 , \10395 , \10713 );
nor \U$9496 ( \11469 , \11467 , \11468 );
xnor \U$9497 ( \11470 , \11469 , \10741 );
xor \U$9498 ( \11471 , \11466 , \11470 );
and \U$9500 ( \11472 , \10765 , \10347 );
and \U$9501 ( \11473 , \10794 , \10345 );
nor \U$9502 ( \11474 , \11472 , \11473 );
xnor \U$9503 ( \11475 , \11474 , \10373 );
and \U$9505 ( \11476 , \10841 , \10400 );
nor \U$9506 ( \11477 , 1'b0 , \11476 );
xnor \U$9507 ( \11478 , \11477 , 1'b0 );
xor \U$9508 ( \11479 , \11475 , \11478 );
xor \U$9510 ( \11480 , \11479 , 1'b0 );
xor \U$9511 ( \11481 , 1'b1 , \11480 );
xor \U$9512 ( \11482 , \11471 , \11481 );
and \U$9514 ( \11483 , \11411 , \11416 );
or \U$9516 ( \11484 , 1'b0 , \11483 , 1'b0 );
and \U$9517 ( \11485 , \11376 , \11380 );
and \U$9518 ( \11486 , \11380 , \11385 );
and \U$9519 ( \11487 , \11376 , \11385 );
or \U$9520 ( \11488 , \11485 , \11486 , \11487 );
xor \U$9521 ( \11489 , \11484 , \11488 );
and \U$9522 ( \11490 , \11362 , \11366 );
and \U$9523 ( \11491 , \11366 , \11370 );
and \U$9524 ( \11492 , \11362 , \11370 );
or \U$9525 ( \11493 , \11490 , \11491 , \11492 );
xor \U$9526 ( \11494 , \11489 , \11493 );
xor \U$9527 ( \11495 , \11482 , \11494 );
xor \U$9528 ( \11496 , \11460 , \11495 );
xor \U$9529 ( \11497 , \11454 , \11496 );
and \U$9530 ( \11498 , \11354 , \11355 );
and \U$9531 ( \11499 , \11355 , \11419 );
and \U$9532 ( \11500 , \11354 , \11419 );
or \U$9533 ( \11501 , \11498 , \11499 , \11500 );
nor \U$9534 ( \11502 , \11497 , \11501 );
and \U$9535 ( \11503 , \11458 , \11459 );
and \U$9536 ( \11504 , \11459 , \11495 );
and \U$9537 ( \11505 , \11458 , \11495 );
or \U$9538 ( \11506 , \11503 , \11504 , \11505 );
and \U$9539 ( \11507 , \11461 , \11465 );
and \U$9540 ( \11508 , \11465 , \11470 );
and \U$9541 ( \11509 , \11461 , \11470 );
or \U$9542 ( \11510 , \11507 , \11508 , \11509 );
and \U$9543 ( \11511 , \11442 , \11446 );
and \U$9544 ( \11512 , \11446 , \11451 );
and \U$9545 ( \11513 , \11442 , \11451 );
or \U$9546 ( \11514 , \11511 , \11512 , \11513 );
xor \U$9547 ( \11515 , \11510 , \11514 );
and \U$9548 ( \11516 , \11475 , \11478 );
or \U$9551 ( \11517 , \11516 , 1'b0 , 1'b0 );
xor \U$9552 ( \11518 , \11515 , \11517 );
and \U$9553 ( \11519 , \11484 , \11488 );
and \U$9554 ( \11520 , \11488 , \11493 );
and \U$9555 ( \11521 , \11484 , \11493 );
or \U$9556 ( \11522 , \11519 , \11520 , \11521 );
and \U$9559 ( \11523 , 1'b1 , \11480 );
or \U$9561 ( \11524 , 1'b0 , \11523 , 1'b0 );
xor \U$9562 ( \11525 , \11522 , \11524 );
and \U$9563 ( \11526 , \10794 , \10347 );
and \U$9564 ( \11527 , \10703 , \10345 );
nor \U$9565 ( \11528 , \11526 , \11527 );
xnor \U$9566 ( \11529 , \11528 , \10373 );
and \U$9568 ( \11530 , \10765 , \10400 );
nor \U$9569 ( \11531 , 1'b0 , \11530 );
xnor \U$9570 ( \11532 , \11531 , 1'b0 );
xor \U$9571 ( \11533 , \11529 , \11532 );
xor \U$9573 ( \11534 , \11533 , 1'b0 );
and \U$9574 ( \11535 , \10506 , \10773 );
and \U$9575 ( \11536 , \10527 , \10771 );
nor \U$9576 ( \11537 , \11535 , \11536 );
xnor \U$9577 ( \11538 , \11537 , \10799 );
and \U$9578 ( \11539 , \10676 , \10474 );
and \U$9579 ( \11540 , \10550 , \10472 );
nor \U$9580 ( \11541 , \11539 , \11540 );
xnor \U$9581 ( \11542 , \11541 , \10479 );
xor \U$9582 ( \11543 , \11538 , \11542 );
and \U$9583 ( \11544 , \10736 , \10409 );
and \U$9584 ( \11545 , \10643 , \10407 );
nor \U$9585 ( \11546 , \11544 , \11545 );
xnor \U$9586 ( \11547 , \11546 , \10176 );
xor \U$9587 ( \11548 , \11543 , \11547 );
xor \U$9588 ( \11549 , \11534 , \11548 );
and \U$9590 ( \11550 , \10368 , \10655 );
not \U$9591 ( \11551 , \11550 );
xnor \U$9592 ( \11552 , \11551 , \10681 );
xor \U$9593 ( \11553 , 1'b0 , \11552 );
and \U$9594 ( \11554 , \10395 , \10715 );
and \U$9595 ( \11555 , \10299 , \10713 );
nor \U$9596 ( \11556 , \11554 , \11555 );
xnor \U$9597 ( \11557 , \11556 , \10741 );
xor \U$9598 ( \11558 , \11553 , \11557 );
xor \U$9599 ( \11559 , \11549 , \11558 );
xor \U$9600 ( \11560 , \11525 , \11559 );
xor \U$9601 ( \11561 , \11518 , \11560 );
xor \U$9602 ( \11562 , \11506 , \11561 );
and \U$9603 ( \11563 , \11435 , \11437 );
and \U$9604 ( \11564 , \11437 , \11452 );
and \U$9605 ( \11565 , \11435 , \11452 );
or \U$9606 ( \11566 , \11563 , \11564 , \11565 );
and \U$9607 ( \11567 , \11471 , \11481 );
and \U$9608 ( \11568 , \11481 , \11494 );
and \U$9609 ( \11569 , \11471 , \11494 );
or \U$9610 ( \11570 , \11567 , \11568 , \11569 );
xor \U$9611 ( \11571 , \11566 , \11570 );
xor \U$9613 ( \11572 , \11571 , 1'b1 );
xor \U$9614 ( \11573 , \11562 , \11572 );
and \U$9615 ( \11574 , \11431 , \11453 );
and \U$9616 ( \11575 , \11453 , \11496 );
and \U$9617 ( \11576 , \11431 , \11496 );
or \U$9618 ( \11577 , \11574 , \11575 , \11576 );
nor \U$9619 ( \11578 , \11573 , \11577 );
nor \U$9620 ( \11579 , \11502 , \11578 );
and \U$9621 ( \11580 , \11566 , \11570 );
and \U$9622 ( \11581 , \11570 , 1'b1 );
and \U$9623 ( \11582 , \11566 , 1'b1 );
or \U$9624 ( \11583 , \11580 , \11581 , \11582 );
and \U$9625 ( \11584 , \11518 , \11560 );
xor \U$9626 ( \11585 , \11583 , \11584 );
and \U$9627 ( \11586 , \11522 , \11524 );
and \U$9628 ( \11587 , \11524 , \11559 );
and \U$9629 ( \11588 , \11522 , \11559 );
or \U$9630 ( \11589 , \11586 , \11587 , \11588 );
and \U$9632 ( \11590 , \10794 , \10400 );
nor \U$9633 ( \11591 , 1'b0 , \11590 );
xnor \U$9634 ( \11592 , \11591 , 1'b0 );
xor \U$9636 ( \11593 , \11592 , 1'b0 );
xor \U$9638 ( \11594 , \11593 , 1'b0 );
and \U$9639 ( \11595 , \10550 , \10474 );
and \U$9640 ( \11596 , \10506 , \10472 );
nor \U$9641 ( \11597 , \11595 , \11596 );
xnor \U$9642 ( \11598 , \11597 , \10479 );
and \U$9643 ( \11599 , \10643 , \10409 );
and \U$9644 ( \11600 , \10676 , \10407 );
nor \U$9645 ( \11601 , \11599 , \11600 );
xnor \U$9646 ( \11602 , \11601 , \10176 );
xor \U$9647 ( \11603 , \11598 , \11602 );
and \U$9648 ( \11604 , \10703 , \10347 );
and \U$9649 ( \11605 , \10736 , \10345 );
nor \U$9650 ( \11606 , \11604 , \11605 );
xnor \U$9651 ( \11607 , \11606 , \10373 );
xor \U$9652 ( \11608 , \11603 , \11607 );
xor \U$9653 ( \11609 , \11594 , \11608 );
not \U$9654 ( \11610 , \10681 );
and \U$9655 ( \11611 , \10299 , \10715 );
and \U$9656 ( \11612 , \10368 , \10713 );
nor \U$9657 ( \11613 , \11611 , \11612 );
xnor \U$9658 ( \11614 , \11613 , \10741 );
xor \U$9659 ( \11615 , \11610 , \11614 );
and \U$9660 ( \11616 , \10527 , \10773 );
and \U$9661 ( \11617 , \10395 , \10771 );
nor \U$9662 ( \11618 , \11616 , \11617 );
xnor \U$9663 ( \11619 , \11618 , \10799 );
xor \U$9664 ( \11620 , \11615 , \11619 );
xor \U$9665 ( \11621 , \11609 , \11620 );
xor \U$9667 ( \11622 , \11621 , 1'b0 );
and \U$9669 ( \11623 , \11552 , \11557 );
or \U$9671 ( \11624 , 1'b0 , \11623 , 1'b0 );
and \U$9672 ( \11625 , \11538 , \11542 );
and \U$9673 ( \11626 , \11542 , \11547 );
and \U$9674 ( \11627 , \11538 , \11547 );
or \U$9675 ( \11628 , \11625 , \11626 , \11627 );
xor \U$9676 ( \11629 , \11624 , \11628 );
and \U$9677 ( \11630 , \11529 , \11532 );
or \U$9680 ( \11631 , \11630 , 1'b0 , 1'b0 );
xor \U$9681 ( \11632 , \11629 , \11631 );
xor \U$9682 ( \11633 , \11622 , \11632 );
xor \U$9683 ( \11634 , \11589 , \11633 );
and \U$9684 ( \11635 , \11510 , \11514 );
and \U$9685 ( \11636 , \11514 , \11517 );
and \U$9686 ( \11637 , \11510 , \11517 );
or \U$9687 ( \11638 , \11635 , \11636 , \11637 );
xor \U$9689 ( \11639 , \11638 , 1'b0 );
and \U$9690 ( \11640 , \11534 , \11548 );
and \U$9691 ( \11641 , \11548 , \11558 );
and \U$9692 ( \11642 , \11534 , \11558 );
or \U$9693 ( \11643 , \11640 , \11641 , \11642 );
xor \U$9694 ( \11644 , \11639 , \11643 );
xor \U$9695 ( \11645 , \11634 , \11644 );
xor \U$9696 ( \11646 , \11585 , \11645 );
and \U$9697 ( \11647 , \11506 , \11561 );
and \U$9698 ( \11648 , \11561 , \11572 );
and \U$9699 ( \11649 , \11506 , \11572 );
or \U$9700 ( \11650 , \11647 , \11648 , \11649 );
nor \U$9701 ( \11651 , \11646 , \11650 );
and \U$9702 ( \11652 , \11589 , \11633 );
and \U$9703 ( \11653 , \11633 , \11644 );
and \U$9704 ( \11654 , \11589 , \11644 );
or \U$9705 ( \11655 , \11652 , \11653 , \11654 );
and \U$9706 ( \11656 , \11624 , \11628 );
and \U$9707 ( \11657 , \11628 , \11631 );
and \U$9708 ( \11658 , \11624 , \11631 );
or \U$9709 ( \11659 , \11656 , \11657 , \11658 );
xor \U$9711 ( \11660 , \11659 , 1'b0 );
and \U$9712 ( \11661 , \11594 , \11608 );
and \U$9713 ( \11662 , \11608 , \11620 );
and \U$9714 ( \11663 , \11594 , \11620 );
or \U$9715 ( \11664 , \11661 , \11662 , \11663 );
xor \U$9716 ( \11665 , \11660 , \11664 );
xor \U$9717 ( \11666 , \11655 , \11665 );
and \U$9720 ( \11667 , \11638 , \11643 );
or \U$9721 ( \11668 , 1'b0 , 1'b0 , \11667 );
and \U$9724 ( \11669 , \11621 , \11632 );
or \U$9725 ( \11670 , 1'b0 , 1'b0 , \11669 );
xor \U$9726 ( \11671 , \11668 , \11670 );
and \U$9727 ( \11672 , \10506 , \10474 );
and \U$9728 ( \11673 , \10527 , \10472 );
nor \U$9729 ( \11674 , \11672 , \11673 );
xnor \U$9730 ( \11675 , \11674 , \10479 );
and \U$9731 ( \11676 , \10676 , \10409 );
and \U$9732 ( \11677 , \10550 , \10407 );
nor \U$9733 ( \11678 , \11676 , \11677 );
xnor \U$9734 ( \11679 , \11678 , \10176 );
xor \U$9735 ( \11680 , \11675 , \11679 );
and \U$9736 ( \11681 , \10736 , \10347 );
and \U$9737 ( \11682 , \10643 , \10345 );
nor \U$9738 ( \11683 , \11681 , \11682 );
xnor \U$9739 ( \11684 , \11683 , \10373 );
xor \U$9740 ( \11685 , \11680 , \11684 );
and \U$9742 ( \11686 , \10368 , \10715 );
not \U$9743 ( \11687 , \11686 );
xnor \U$9744 ( \11688 , \11687 , \10741 );
xor \U$9745 ( \11689 , 1'b0 , \11688 );
and \U$9746 ( \11690 , \10395 , \10773 );
and \U$9747 ( \11691 , \10299 , \10771 );
nor \U$9748 ( \11692 , \11690 , \11691 );
xnor \U$9749 ( \11693 , \11692 , \10799 );
xor \U$9750 ( \11694 , \11689 , \11693 );
xor \U$9751 ( \11695 , \11685 , \11694 );
and \U$9754 ( \11696 , \10703 , \10400 );
nor \U$9755 ( \11697 , 1'b0 , \11696 );
xnor \U$9756 ( \11698 , \11697 , 1'b0 );
xor \U$9758 ( \11699 , \11698 , 1'b0 );
xor \U$9760 ( \11700 , \11699 , 1'b0 );
xnor \U$9761 ( \11701 , 1'b0 , \11700 );
xor \U$9762 ( \11702 , \11695 , \11701 );
and \U$9763 ( \11703 , \11610 , \11614 );
and \U$9764 ( \11704 , \11614 , \11619 );
and \U$9765 ( \11705 , \11610 , \11619 );
or \U$9766 ( \11706 , \11703 , \11704 , \11705 );
and \U$9767 ( \11707 , \11598 , \11602 );
and \U$9768 ( \11708 , \11602 , \11607 );
and \U$9769 ( \11709 , \11598 , \11607 );
or \U$9770 ( \11710 , \11707 , \11708 , \11709 );
xor \U$9771 ( \11711 , \11706 , \11710 );
xor \U$9773 ( \11712 , \11711 , 1'b0 );
xor \U$9774 ( \11713 , \11702 , \11712 );
xor \U$9775 ( \11714 , \11671 , \11713 );
xor \U$9776 ( \11715 , \11666 , \11714 );
and \U$9777 ( \11716 , \11583 , \11584 );
and \U$9778 ( \11717 , \11584 , \11645 );
and \U$9779 ( \11718 , \11583 , \11645 );
or \U$9780 ( \11719 , \11716 , \11717 , \11718 );
nor \U$9781 ( \11720 , \11715 , \11719 );
nor \U$9782 ( \11721 , \11651 , \11720 );
nand \U$9783 ( \11722 , \11579 , \11721 );
nor \U$9784 ( \11723 , \11427 , \11722 );
and \U$9785 ( \11724 , \11668 , \11670 );
and \U$9786 ( \11725 , \11670 , \11713 );
and \U$9787 ( \11726 , \11668 , \11713 );
or \U$9788 ( \11727 , \11724 , \11725 , \11726 );
and \U$9789 ( \11728 , \11706 , \11710 );
or \U$9792 ( \11729 , \11728 , 1'b0 , 1'b0 );
or \U$9793 ( \11730 , 1'b0 , \11700 );
xor \U$9794 ( \11731 , \11729 , \11730 );
and \U$9795 ( \11732 , \11685 , \11694 );
xor \U$9796 ( \11733 , \11731 , \11732 );
xor \U$9797 ( \11734 , \11727 , \11733 );
and \U$9800 ( \11735 , \11659 , \11664 );
or \U$9801 ( \11736 , 1'b0 , 1'b0 , \11735 );
and \U$9802 ( \11737 , \11695 , \11701 );
and \U$9803 ( \11738 , \11701 , \11712 );
and \U$9804 ( \11739 , \11695 , \11712 );
or \U$9805 ( \11740 , \11737 , \11738 , \11739 );
xor \U$9806 ( \11741 , \11736 , \11740 );
and \U$9808 ( \11742 , \10550 , \10409 );
and \U$9809 ( \11743 , \10506 , \10407 );
nor \U$9810 ( \11744 , \11742 , \11743 );
xnor \U$9811 ( \11745 , \11744 , \10176 );
and \U$9812 ( \11746 , \10643 , \10347 );
and \U$9813 ( \11747 , \10676 , \10345 );
nor \U$9814 ( \11748 , \11746 , \11747 );
xnor \U$9815 ( \11749 , \11748 , \10373 );
xor \U$9816 ( \11750 , \11745 , \11749 );
and \U$9818 ( \11751 , \10736 , \10400 );
nor \U$9819 ( \11752 , 1'b0 , \11751 );
xnor \U$9820 ( \11753 , \11752 , 1'b0 );
xor \U$9821 ( \11754 , \11750 , \11753 );
xor \U$9822 ( \11755 , 1'b0 , \11754 );
not \U$9823 ( \11756 , \10741 );
and \U$9824 ( \11757 , \10299 , \10773 );
and \U$9825 ( \11758 , \10368 , \10771 );
nor \U$9826 ( \11759 , \11757 , \11758 );
xnor \U$9827 ( \11760 , \11759 , \10799 );
xor \U$9828 ( \11761 , \11756 , \11760 );
and \U$9829 ( \11762 , \10527 , \10474 );
and \U$9830 ( \11763 , \10395 , \10472 );
nor \U$9831 ( \11764 , \11762 , \11763 );
xnor \U$9832 ( \11765 , \11764 , \10479 );
xor \U$9833 ( \11766 , \11761 , \11765 );
xor \U$9834 ( \11767 , \11755 , \11766 );
xor \U$9836 ( \11768 , \11767 , 1'b0 );
and \U$9838 ( \11769 , \11688 , \11693 );
or \U$9840 ( \11770 , 1'b0 , \11769 , 1'b0 );
and \U$9841 ( \11771 , \11675 , \11679 );
and \U$9842 ( \11772 , \11679 , \11684 );
and \U$9843 ( \11773 , \11675 , \11684 );
or \U$9844 ( \11774 , \11771 , \11772 , \11773 );
xor \U$9845 ( \11775 , \11770 , \11774 );
xor \U$9847 ( \11776 , \11775 , 1'b0 );
xor \U$9848 ( \11777 , \11768 , \11776 );
xor \U$9849 ( \11778 , \11741 , \11777 );
xor \U$9850 ( \11779 , \11734 , \11778 );
and \U$9851 ( \11780 , \11655 , \11665 );
and \U$9852 ( \11781 , \11665 , \11714 );
and \U$9853 ( \11782 , \11655 , \11714 );
or \U$9854 ( \11783 , \11780 , \11781 , \11782 );
nor \U$9855 ( \11784 , \11779 , \11783 );
and \U$9856 ( \11785 , \11736 , \11740 );
and \U$9857 ( \11786 , \11740 , \11777 );
and \U$9858 ( \11787 , \11736 , \11777 );
or \U$9859 ( \11788 , \11785 , \11786 , \11787 );
and \U$9860 ( \11789 , \11770 , \11774 );
or \U$9863 ( \11790 , \11789 , 1'b0 , 1'b0 );
xor \U$9865 ( \11791 , \11790 , 1'b0 );
and \U$9867 ( \11792 , \11754 , \11766 );
or \U$9869 ( \11793 , 1'b0 , \11792 , 1'b0 );
xor \U$9870 ( \11794 , \11791 , \11793 );
xor \U$9871 ( \11795 , \11788 , \11794 );
and \U$9872 ( \11796 , \11729 , \11730 );
and \U$9873 ( \11797 , \11730 , \11732 );
and \U$9874 ( \11798 , \11729 , \11732 );
or \U$9875 ( \11799 , \11796 , \11797 , \11798 );
and \U$9878 ( \11800 , \11767 , \11776 );
or \U$9879 ( \11801 , 1'b0 , 1'b0 , \11800 );
xor \U$9880 ( \11802 , \11799 , \11801 );
and \U$9881 ( \11803 , \10506 , \10409 );
and \U$9882 ( \11804 , \10527 , \10407 );
nor \U$9883 ( \11805 , \11803 , \11804 );
xnor \U$9884 ( \11806 , \11805 , \10176 );
and \U$9885 ( \11807 , \10676 , \10347 );
and \U$9886 ( \11808 , \10550 , \10345 );
nor \U$9887 ( \11809 , \11807 , \11808 );
xnor \U$9888 ( \11810 , \11809 , \10373 );
xor \U$9889 ( \11811 , \11806 , \11810 );
and \U$9891 ( \11812 , \10643 , \10400 );
nor \U$9892 ( \11813 , 1'b0 , \11812 );
xnor \U$9893 ( \11814 , \11813 , 1'b0 );
xor \U$9894 ( \11815 , \11811 , \11814 );
and \U$9896 ( \11816 , \10368 , \10773 );
not \U$9897 ( \11817 , \11816 );
xnor \U$9898 ( \11818 , \11817 , \10799 );
xor \U$9899 ( \11819 , 1'b0 , \11818 );
and \U$9900 ( \11820 , \10395 , \10474 );
and \U$9901 ( \11821 , \10299 , \10472 );
nor \U$9902 ( \11822 , \11820 , \11821 );
xnor \U$9903 ( \11823 , \11822 , \10479 );
xor \U$9904 ( \11824 , \11819 , \11823 );
xor \U$9905 ( \11825 , \11815 , \11824 );
xor \U$9907 ( \11826 , \11825 , 1'b1 );
and \U$9908 ( \11827 , \11756 , \11760 );
and \U$9909 ( \11828 , \11760 , \11765 );
and \U$9910 ( \11829 , \11756 , \11765 );
or \U$9911 ( \11830 , \11827 , \11828 , \11829 );
and \U$9912 ( \11831 , \11745 , \11749 );
and \U$9913 ( \11832 , \11749 , \11753 );
and \U$9914 ( \11833 , \11745 , \11753 );
or \U$9915 ( \11834 , \11831 , \11832 , \11833 );
xor \U$9916 ( \11835 , \11830 , \11834 );
xor \U$9918 ( \11836 , \11835 , 1'b0 );
xor \U$9919 ( \11837 , \11826 , \11836 );
xor \U$9920 ( \11838 , \11802 , \11837 );
xor \U$9921 ( \11839 , \11795 , \11838 );
and \U$9922 ( \11840 , \11727 , \11733 );
and \U$9923 ( \11841 , \11733 , \11778 );
and \U$9924 ( \11842 , \11727 , \11778 );
or \U$9925 ( \11843 , \11840 , \11841 , \11842 );
nor \U$9926 ( \11844 , \11839 , \11843 );
nor \U$9927 ( \11845 , \11784 , \11844 );
and \U$9928 ( \11846 , \11799 , \11801 );
and \U$9929 ( \11847 , \11801 , \11837 );
and \U$9930 ( \11848 , \11799 , \11837 );
or \U$9931 ( \11849 , \11846 , \11847 , \11848 );
and \U$9932 ( \11850 , \11830 , \11834 );
or \U$9935 ( \11851 , \11850 , 1'b0 , 1'b0 );
xor \U$9937 ( \11852 , \11851 , 1'b0 );
and \U$9938 ( \11853 , \11815 , \11824 );
xor \U$9939 ( \11854 , \11852 , \11853 );
xor \U$9940 ( \11855 , \11849 , \11854 );
and \U$9943 ( \11856 , \11790 , \11793 );
or \U$9944 ( \11857 , 1'b0 , 1'b0 , \11856 );
and \U$9945 ( \11858 , \11825 , 1'b1 );
and \U$9946 ( \11859 , 1'b1 , \11836 );
and \U$9947 ( \11860 , \11825 , \11836 );
or \U$9948 ( \11861 , \11858 , \11859 , \11860 );
xor \U$9949 ( \11862 , \11857 , \11861 );
and \U$9951 ( \11863 , \10550 , \10347 );
and \U$9952 ( \11864 , \10506 , \10345 );
nor \U$9953 ( \11865 , \11863 , \11864 );
xnor \U$9954 ( \11866 , \11865 , \10373 );
and \U$9956 ( \11867 , \10676 , \10400 );
nor \U$9957 ( \11868 , 1'b0 , \11867 );
xnor \U$9958 ( \11869 , \11868 , 1'b0 );
xor \U$9959 ( \11870 , \11866 , \11869 );
xor \U$9961 ( \11871 , \11870 , 1'b0 );
xor \U$9962 ( \11872 , 1'b0 , \11871 );
not \U$9963 ( \11873 , \10799 );
and \U$9964 ( \11874 , \10299 , \10474 );
and \U$9965 ( \11875 , \10368 , \10472 );
nor \U$9966 ( \11876 , \11874 , \11875 );
xnor \U$9967 ( \11877 , \11876 , \10479 );
xor \U$9968 ( \11878 , \11873 , \11877 );
and \U$9969 ( \11879 , \10527 , \10409 );
and \U$9970 ( \11880 , \10395 , \10407 );
nor \U$9971 ( \11881 , \11879 , \11880 );
xnor \U$9972 ( \11882 , \11881 , \10176 );
xor \U$9973 ( \11883 , \11878 , \11882 );
xor \U$9974 ( \11884 , \11872 , \11883 );
xor \U$9976 ( \11885 , \11884 , 1'b0 );
and \U$9978 ( \11886 , \11818 , \11823 );
or \U$9980 ( \11887 , 1'b0 , \11886 , 1'b0 );
and \U$9981 ( \11888 , \11806 , \11810 );
and \U$9982 ( \11889 , \11810 , \11814 );
and \U$9983 ( \11890 , \11806 , \11814 );
or \U$9984 ( \11891 , \11888 , \11889 , \11890 );
xor \U$9985 ( \11892 , \11887 , \11891 );
xor \U$9987 ( \11893 , \11892 , 1'b0 );
xor \U$9988 ( \11894 , \11885 , \11893 );
xor \U$9989 ( \11895 , \11862 , \11894 );
xor \U$9990 ( \11896 , \11855 , \11895 );
and \U$9991 ( \11897 , \11788 , \11794 );
and \U$9992 ( \11898 , \11794 , \11838 );
and \U$9993 ( \11899 , \11788 , \11838 );
or \U$9994 ( \11900 , \11897 , \11898 , \11899 );
nor \U$9995 ( \11901 , \11896 , \11900 );
and \U$9996 ( \11902 , \11857 , \11861 );
and \U$9997 ( \11903 , \11861 , \11894 );
and \U$9998 ( \11904 , \11857 , \11894 );
or \U$9999 ( \11905 , \11902 , \11903 , \11904 );
and \U$10000 ( \11906 , \11887 , \11891 );
or \U$10003 ( \11907 , \11906 , 1'b0 , 1'b0 );
xor \U$10005 ( \11908 , \11907 , 1'b0 );
and \U$10007 ( \11909 , \11871 , \11883 );
or \U$10009 ( \11910 , 1'b0 , \11909 , 1'b0 );
xor \U$10010 ( \11911 , \11908 , \11910 );
xor \U$10011 ( \11912 , \11905 , \11911 );
and \U$10014 ( \11913 , \11851 , \11853 );
or \U$10015 ( \11914 , 1'b0 , 1'b0 , \11913 );
and \U$10018 ( \11915 , \11884 , \11893 );
or \U$10019 ( \11916 , 1'b0 , 1'b0 , \11915 );
xor \U$10020 ( \11917 , \11914 , \11916 );
xor \U$10021 ( \11918 , \10530 , \10553 );
xor \U$10023 ( \11919 , \11918 , 1'b0 );
xor \U$10025 ( \11920 , 1'b0 , \10480 );
xor \U$10026 ( \11921 , \11920 , \10484 );
xor \U$10027 ( \11922 , \11919 , \11921 );
xor \U$10029 ( \11923 , \11922 , 1'b1 );
and \U$10030 ( \11924 , \11873 , \11877 );
and \U$10031 ( \11925 , \11877 , \11882 );
and \U$10032 ( \11926 , \11873 , \11882 );
or \U$10033 ( \11927 , \11924 , \11925 , \11926 );
and \U$10034 ( \11928 , \11866 , \11869 );
or \U$10037 ( \11929 , \11928 , 1'b0 , 1'b0 );
xor \U$10038 ( \11930 , \11927 , \11929 );
xor \U$10040 ( \11931 , \11930 , 1'b0 );
xor \U$10041 ( \11932 , \11923 , \11931 );
xor \U$10042 ( \11933 , \11917 , \11932 );
xor \U$10043 ( \11934 , \11912 , \11933 );
and \U$10044 ( \11935 , \11849 , \11854 );
and \U$10045 ( \11936 , \11854 , \11895 );
and \U$10046 ( \11937 , \11849 , \11895 );
or \U$10047 ( \11938 , \11935 , \11936 , \11937 );
nor \U$10048 ( \11939 , \11934 , \11938 );
nor \U$10049 ( \11940 , \11901 , \11939 );
nand \U$10050 ( \11941 , \11845 , \11940 );
and \U$10051 ( \11942 , \11914 , \11916 );
and \U$10052 ( \11943 , \11916 , \11932 );
and \U$10053 ( \11944 , \11914 , \11932 );
or \U$10054 ( \11945 , \11942 , \11943 , \11944 );
and \U$10055 ( \11946 , \11927 , \11929 );
or \U$10058 ( \11947 , \11946 , 1'b0 , 1'b0 );
xor \U$10060 ( \11948 , \11947 , 1'b0 );
and \U$10061 ( \11949 , \11919 , \11921 );
xor \U$10062 ( \11950 , \11948 , \11949 );
xor \U$10063 ( \11951 , \11945 , \11950 );
and \U$10066 ( \11952 , \11907 , \11910 );
or \U$10067 ( \11953 , 1'b0 , 1'b0 , \11952 );
and \U$10068 ( \11954 , \11922 , 1'b1 );
and \U$10069 ( \11955 , 1'b1 , \11931 );
and \U$10070 ( \11956 , \11922 , \11931 );
or \U$10071 ( \11957 , \11954 , \11955 , \11956 );
xor \U$10072 ( \11958 , \11953 , \11957 );
xor \U$10074 ( \11959 , 1'b0 , \10562 );
xor \U$10075 ( \11960 , \11959 , \10573 );
xor \U$10077 ( \11961 , \11960 , 1'b0 );
xor \U$10078 ( \11962 , \10486 , \10555 );
xor \U$10080 ( \11963 , \11962 , 1'b0 );
xor \U$10081 ( \11964 , \11961 , \11963 );
xor \U$10082 ( \11965 , \11958 , \11964 );
xor \U$10083 ( \11966 , \11951 , \11965 );
and \U$10084 ( \11967 , \11905 , \11911 );
and \U$10085 ( \11968 , \11911 , \11933 );
and \U$10086 ( \11969 , \11905 , \11933 );
or \U$10087 ( \11970 , \11967 , \11968 , \11969 );
nor \U$10088 ( \11971 , \11966 , \11970 );
and \U$10089 ( \11972 , \11953 , \11957 );
and \U$10090 ( \11973 , \11957 , \11964 );
and \U$10091 ( \11974 , \11953 , \11964 );
or \U$10092 ( \11975 , \11972 , \11973 , \11974 );
xor \U$10094 ( \11976 , \10557 , 1'b0 );
xor \U$10095 ( \11977 , \11976 , \10575 );
xor \U$10096 ( \11978 , \11975 , \11977 );
and \U$10099 ( \11979 , \11947 , \11949 );
or \U$10100 ( \11980 , 1'b0 , 1'b0 , \11979 );
and \U$10103 ( \11981 , \11960 , \11963 );
or \U$10104 ( \11982 , 1'b0 , 1'b0 , \11981 );
xor \U$10105 ( \11983 , \11980 , \11982 );
xor \U$10106 ( \11984 , \10585 , 1'b1 );
xor \U$10107 ( \11985 , \11984 , \10592 );
xor \U$10108 ( \11986 , \11983 , \11985 );
xor \U$10109 ( \11987 , \11978 , \11986 );
and \U$10110 ( \11988 , \11945 , \11950 );
and \U$10111 ( \11989 , \11950 , \11965 );
and \U$10112 ( \11990 , \11945 , \11965 );
or \U$10113 ( \11991 , \11988 , \11989 , \11990 );
nor \U$10114 ( \11992 , \11987 , \11991 );
nor \U$10115 ( \11993 , \11971 , \11992 );
and \U$10116 ( \11994 , \11980 , \11982 );
and \U$10117 ( \11995 , \11982 , \11985 );
and \U$10118 ( \11996 , \11980 , \11985 );
or \U$10119 ( \11997 , \11994 , \11995 , \11996 );
and \U$10121 ( \11998 , \10582 , \10584 );
xor \U$10122 ( \11999 , 1'b0 , \11998 );
xor \U$10123 ( \12000 , \11997 , \11999 );
xor \U$10124 ( \12001 , \10577 , \10595 );
xor \U$10125 ( \12002 , \12001 , \10598 );
xor \U$10126 ( \12003 , \12000 , \12002 );
and \U$10127 ( \12004 , \11975 , \11977 );
and \U$10128 ( \12005 , \11977 , \11986 );
and \U$10129 ( \12006 , \11975 , \11986 );
or \U$10130 ( \12007 , \12004 , \12005 , \12006 );
nor \U$10131 ( \12008 , \12003 , \12007 );
xor \U$10133 ( \12009 , \10601 , 1'b0 );
xor \U$10134 ( \12010 , \12009 , \10603 );
and \U$10135 ( \12011 , \11997 , \11999 );
and \U$10136 ( \12012 , \11999 , \12002 );
and \U$10137 ( \12013 , \11997 , \12002 );
or \U$10138 ( \12014 , \12011 , \12012 , \12013 );
nor \U$10139 ( \12015 , \12010 , \12014 );
nor \U$10140 ( \12016 , \12008 , \12015 );
nand \U$10141 ( \12017 , \11993 , \12016 );
nor \U$10142 ( \12018 , \11941 , \12017 );
nand \U$10143 ( \12019 , \11723 , \12018 );
and \U$10144 ( \12020 , \10820 , \10619 );
and \U$10145 ( \12021 , \10841 , \10616 );
nor \U$10146 ( \12022 , \12020 , \12021 );
xnor \U$10147 ( \12023 , \12022 , \10613 );
and \U$10148 ( \12024 , \10865 , \10655 );
and \U$10149 ( \12025 , \10886 , \10653 );
nor \U$10150 ( \12026 , \12024 , \12025 );
xnor \U$10151 ( \12027 , \12026 , \10681 );
and \U$10152 ( \12028 , \12023 , \12027 );
and \U$10153 ( \12029 , \10913 , \10715 );
and \U$10154 ( \12030 , \10934 , \10713 );
nor \U$10155 ( \12031 , \12029 , \12030 );
xnor \U$10156 ( \12032 , \12031 , \10741 );
and \U$10157 ( \12033 , \12027 , \12032 );
and \U$10158 ( \12034 , \12023 , \12032 );
or \U$10159 ( \12035 , \12028 , \12033 , \12034 );
and \U$10160 ( \12036 , \10934 , \10715 );
and \U$10161 ( \12037 , \10865 , \10713 );
nor \U$10162 ( \12038 , \12036 , \12037 );
xnor \U$10163 ( \12039 , \12038 , \10741 );
and \U$10164 ( \12040 , \10957 , \10773 );
and \U$10165 ( \12041 , \10913 , \10771 );
nor \U$10166 ( \12042 , \12040 , \12041 );
xnor \U$10167 ( \12043 , \12042 , \10799 );
xor \U$10168 ( \12044 , \12039 , \12043 );
nand \U$10169 ( \12045 , \11090 , \10472 );
xnor \U$10170 ( \12046 , \12045 , \10479 );
xor \U$10171 ( \12047 , \12044 , \12046 );
and \U$10172 ( \12048 , \12035 , \12047 );
and \U$10173 ( \12049 , \10841 , \10619 );
and \U$10174 ( \12050 , \10765 , \10616 );
nor \U$10175 ( \12051 , \12049 , \12050 );
xnor \U$10176 ( \12052 , \12051 , \10613 );
xor \U$10177 ( \12053 , \10479 , \12052 );
and \U$10178 ( \12054 , \10886 , \10655 );
and \U$10179 ( \12055 , \10820 , \10653 );
nor \U$10180 ( \12056 , \12054 , \12055 );
xnor \U$10181 ( \12057 , \12056 , \10681 );
xor \U$10182 ( \12058 , \12053 , \12057 );
and \U$10183 ( \12059 , \12047 , \12058 );
and \U$10184 ( \12060 , \12035 , \12058 );
or \U$10185 ( \12061 , \12048 , \12059 , \12060 );
and \U$10186 ( \12062 , \11090 , \10474 );
and \U$10187 ( \12063 , \10957 , \10472 );
nor \U$10188 ( \12064 , \12062 , \12063 );
xnor \U$10189 ( \12065 , \12064 , \10479 );
and \U$10190 ( \12066 , \10765 , \10619 );
and \U$10191 ( \12067 , \10794 , \10616 );
nor \U$10192 ( \12068 , \12066 , \12067 );
xnor \U$10193 ( \12069 , \12068 , \10613 );
and \U$10194 ( \12070 , \10820 , \10655 );
and \U$10195 ( \12071 , \10841 , \10653 );
nor \U$10196 ( \12072 , \12070 , \12071 );
xnor \U$10197 ( \12073 , \12072 , \10681 );
xor \U$10198 ( \12074 , \12069 , \12073 );
and \U$10199 ( \12075 , \10865 , \10715 );
and \U$10200 ( \12076 , \10886 , \10713 );
nor \U$10201 ( \12077 , \12075 , \12076 );
xnor \U$10202 ( \12078 , \12077 , \10741 );
xor \U$10203 ( \12079 , \12074 , \12078 );
xor \U$10204 ( \12080 , \12065 , \12079 );
xor \U$10205 ( \12081 , \12061 , \12080 );
and \U$10206 ( \12082 , \10479 , \12052 );
and \U$10207 ( \12083 , \12052 , \12057 );
and \U$10208 ( \12084 , \10479 , \12057 );
or \U$10209 ( \12085 , \12082 , \12083 , \12084 );
and \U$10210 ( \12086 , \12039 , \12043 );
and \U$10211 ( \12087 , \12043 , \12046 );
and \U$10212 ( \12088 , \12039 , \12046 );
or \U$10213 ( \12089 , \12086 , \12087 , \12088 );
xor \U$10214 ( \12090 , \12085 , \12089 );
and \U$10215 ( \12091 , \10913 , \10773 );
and \U$10216 ( \12092 , \10934 , \10771 );
nor \U$10217 ( \12093 , \12091 , \12092 );
xnor \U$10218 ( \12094 , \12093 , \10799 );
xor \U$10219 ( \12095 , \12090 , \12094 );
xor \U$10220 ( \12096 , \12081 , \12095 );
and \U$10221 ( \12097 , \10886 , \10619 );
and \U$10222 ( \12098 , \10820 , \10616 );
nor \U$10223 ( \12099 , \12097 , \12098 );
xnor \U$10224 ( \12100 , \12099 , \10613 );
and \U$10225 ( \12101 , \10799 , \12100 );
and \U$10226 ( \12102 , \10934 , \10655 );
and \U$10227 ( \12103 , \10865 , \10653 );
nor \U$10228 ( \12104 , \12102 , \12103 );
xnor \U$10229 ( \12105 , \12104 , \10681 );
and \U$10230 ( \12106 , \12100 , \12105 );
and \U$10231 ( \12107 , \10799 , \12105 );
or \U$10232 ( \12108 , \12101 , \12106 , \12107 );
and \U$10233 ( \12109 , \10957 , \10715 );
and \U$10234 ( \12110 , \10913 , \10713 );
nor \U$10235 ( \12111 , \12109 , \12110 );
xnor \U$10236 ( \12112 , \12111 , \10741 );
nand \U$10237 ( \12113 , \11090 , \10771 );
xnor \U$10238 ( \12114 , \12113 , \10799 );
and \U$10239 ( \12115 , \12112 , \12114 );
and \U$10240 ( \12116 , \12108 , \12115 );
and \U$10241 ( \12117 , \11090 , \10773 );
and \U$10242 ( \12118 , \10957 , \10771 );
nor \U$10243 ( \12119 , \12117 , \12118 );
xnor \U$10244 ( \12120 , \12119 , \10799 );
and \U$10245 ( \12121 , \12115 , \12120 );
and \U$10246 ( \12122 , \12108 , \12120 );
or \U$10247 ( \12123 , \12116 , \12121 , \12122 );
xor \U$10248 ( \12124 , \12035 , \12047 );
xor \U$10249 ( \12125 , \12124 , \12058 );
and \U$10250 ( \12126 , \12123 , \12125 );
nor \U$10251 ( \12127 , \12096 , \12126 );
and \U$10252 ( \12128 , \12069 , \12073 );
and \U$10253 ( \12129 , \12073 , \12078 );
and \U$10254 ( \12130 , \12069 , \12078 );
or \U$10255 ( \12131 , \12128 , \12129 , \12130 );
nand \U$10256 ( \12132 , \11090 , \10407 );
xnor \U$10257 ( \12133 , \12132 , \10176 );
xor \U$10258 ( \12134 , \12131 , \12133 );
and \U$10259 ( \12135 , \10886 , \10715 );
and \U$10260 ( \12136 , \10820 , \10713 );
nor \U$10261 ( \12137 , \12135 , \12136 );
xnor \U$10262 ( \12138 , \12137 , \10741 );
and \U$10263 ( \12139 , \10934 , \10773 );
and \U$10264 ( \12140 , \10865 , \10771 );
nor \U$10265 ( \12141 , \12139 , \12140 );
xnor \U$10266 ( \12142 , \12141 , \10799 );
xor \U$10267 ( \12143 , \12138 , \12142 );
and \U$10268 ( \12144 , \10957 , \10474 );
and \U$10269 ( \12145 , \10913 , \10472 );
nor \U$10270 ( \12146 , \12144 , \12145 );
xnor \U$10271 ( \12147 , \12146 , \10479 );
xor \U$10272 ( \12148 , \12143 , \12147 );
xor \U$10273 ( \12149 , \12134 , \12148 );
and \U$10274 ( \12150 , \12085 , \12089 );
and \U$10275 ( \12151 , \12089 , \12094 );
and \U$10276 ( \12152 , \12085 , \12094 );
or \U$10277 ( \12153 , \12150 , \12151 , \12152 );
and \U$10278 ( \12154 , \12065 , \12079 );
xor \U$10279 ( \12155 , \12153 , \12154 );
and \U$10280 ( \12156 , \10794 , \10619 );
and \U$10281 ( \12157 , \10703 , \10616 );
nor \U$10282 ( \12158 , \12156 , \12157 );
xnor \U$10283 ( \12159 , \12158 , \10613 );
xor \U$10284 ( \12160 , \10176 , \12159 );
and \U$10285 ( \12161 , \10841 , \10655 );
and \U$10286 ( \12162 , \10765 , \10653 );
nor \U$10287 ( \12163 , \12161 , \12162 );
xnor \U$10288 ( \12164 , \12163 , \10681 );
xor \U$10289 ( \12165 , \12160 , \12164 );
xor \U$10290 ( \12166 , \12155 , \12165 );
xor \U$10291 ( \12167 , \12149 , \12166 );
and \U$10292 ( \12168 , \12061 , \12080 );
and \U$10293 ( \12169 , \12080 , \12095 );
and \U$10294 ( \12170 , \12061 , \12095 );
or \U$10295 ( \12171 , \12168 , \12169 , \12170 );
nor \U$10296 ( \12172 , \12167 , \12171 );
nor \U$10297 ( \12173 , \12127 , \12172 );
and \U$10298 ( \12174 , \12153 , \12154 );
and \U$10299 ( \12175 , \12154 , \12165 );
and \U$10300 ( \12176 , \12153 , \12165 );
or \U$10301 ( \12177 , \12174 , \12175 , \12176 );
and \U$10302 ( \12178 , \12131 , \12133 );
and \U$10303 ( \12179 , \12133 , \12148 );
and \U$10304 ( \12180 , \12131 , \12148 );
or \U$10305 ( \12181 , \12178 , \12179 , \12180 );
and \U$10306 ( \12182 , \10703 , \10619 );
and \U$10307 ( \12183 , \10736 , \10616 );
nor \U$10308 ( \12184 , \12182 , \12183 );
xnor \U$10309 ( \12185 , \12184 , \10613 );
and \U$10310 ( \12186 , \10765 , \10655 );
and \U$10311 ( \12187 , \10794 , \10653 );
nor \U$10312 ( \12188 , \12186 , \12187 );
xnor \U$10313 ( \12189 , \12188 , \10681 );
xor \U$10314 ( \12190 , \12185 , \12189 );
and \U$10315 ( \12191 , \10820 , \10715 );
and \U$10316 ( \12192 , \10841 , \10713 );
nor \U$10317 ( \12193 , \12191 , \12192 );
xnor \U$10318 ( \12194 , \12193 , \10741 );
xor \U$10319 ( \12195 , \12190 , \12194 );
xor \U$10320 ( \12196 , \12181 , \12195 );
and \U$10321 ( \12197 , \10176 , \12159 );
and \U$10322 ( \12198 , \12159 , \12164 );
and \U$10323 ( \12199 , \10176 , \12164 );
or \U$10324 ( \12200 , \12197 , \12198 , \12199 );
and \U$10325 ( \12201 , \12138 , \12142 );
and \U$10326 ( \12202 , \12142 , \12147 );
and \U$10327 ( \12203 , \12138 , \12147 );
or \U$10328 ( \12204 , \12201 , \12202 , \12203 );
xor \U$10329 ( \12205 , \12200 , \12204 );
and \U$10330 ( \12206 , \10865 , \10773 );
and \U$10331 ( \12207 , \10886 , \10771 );
nor \U$10332 ( \12208 , \12206 , \12207 );
xnor \U$10333 ( \12209 , \12208 , \10799 );
and \U$10334 ( \12210 , \10913 , \10474 );
and \U$10335 ( \12211 , \10934 , \10472 );
nor \U$10336 ( \12212 , \12210 , \12211 );
xnor \U$10337 ( \12213 , \12212 , \10479 );
xor \U$10338 ( \12214 , \12209 , \12213 );
and \U$10339 ( \12215 , \11090 , \10409 );
and \U$10340 ( \12216 , \10957 , \10407 );
nor \U$10341 ( \12217 , \12215 , \12216 );
xnor \U$10342 ( \12218 , \12217 , \10176 );
xor \U$10343 ( \12219 , \12214 , \12218 );
xor \U$10344 ( \12220 , \12205 , \12219 );
xor \U$10345 ( \12221 , \12196 , \12220 );
xor \U$10346 ( \12222 , \12177 , \12221 );
and \U$10347 ( \12223 , \12149 , \12166 );
nor \U$10348 ( \12224 , \12222 , \12223 );
and \U$10349 ( \12225 , \12181 , \12195 );
and \U$10350 ( \12226 , \12195 , \12220 );
and \U$10351 ( \12227 , \12181 , \12220 );
or \U$10352 ( \12228 , \12225 , \12226 , \12227 );
and \U$10353 ( \12229 , \12200 , \12204 );
and \U$10354 ( \12230 , \12204 , \12219 );
and \U$10355 ( \12231 , \12200 , \12219 );
or \U$10356 ( \12232 , \12229 , \12230 , \12231 );
nand \U$10357 ( \12233 , \11090 , \10345 );
xnor \U$10358 ( \12234 , \12233 , \10373 );
and \U$10359 ( \12235 , \10841 , \10715 );
and \U$10360 ( \12236 , \10765 , \10713 );
nor \U$10361 ( \12237 , \12235 , \12236 );
xnor \U$10362 ( \12238 , \12237 , \10741 );
and \U$10363 ( \12239 , \10886 , \10773 );
and \U$10364 ( \12240 , \10820 , \10771 );
nor \U$10365 ( \12241 , \12239 , \12240 );
xnor \U$10366 ( \12242 , \12241 , \10799 );
xor \U$10367 ( \12243 , \12238 , \12242 );
and \U$10368 ( \12244 , \10934 , \10474 );
and \U$10369 ( \12245 , \10865 , \10472 );
nor \U$10370 ( \12246 , \12244 , \12245 );
xnor \U$10371 ( \12247 , \12246 , \10479 );
xor \U$10372 ( \12248 , \12243 , \12247 );
xor \U$10373 ( \12249 , \12234 , \12248 );
and \U$10374 ( \12250 , \10736 , \10619 );
and \U$10375 ( \12251 , \10643 , \10616 );
nor \U$10376 ( \12252 , \12250 , \12251 );
xnor \U$10377 ( \12253 , \12252 , \10613 );
xor \U$10378 ( \12254 , \10373 , \12253 );
and \U$10379 ( \12255 , \10794 , \10655 );
and \U$10380 ( \12256 , \10703 , \10653 );
nor \U$10381 ( \12257 , \12255 , \12256 );
xnor \U$10382 ( \12258 , \12257 , \10681 );
xor \U$10383 ( \12259 , \12254 , \12258 );
xor \U$10384 ( \12260 , \12249 , \12259 );
xor \U$10385 ( \12261 , \12232 , \12260 );
and \U$10386 ( \12262 , \12185 , \12189 );
and \U$10387 ( \12263 , \12189 , \12194 );
and \U$10388 ( \12264 , \12185 , \12194 );
or \U$10389 ( \12265 , \12262 , \12263 , \12264 );
and \U$10390 ( \12266 , \12209 , \12213 );
and \U$10391 ( \12267 , \12213 , \12218 );
and \U$10392 ( \12268 , \12209 , \12218 );
or \U$10393 ( \12269 , \12266 , \12267 , \12268 );
xor \U$10394 ( \12270 , \12265 , \12269 );
and \U$10395 ( \12271 , \10957 , \10409 );
and \U$10396 ( \12272 , \10913 , \10407 );
nor \U$10397 ( \12273 , \12271 , \12272 );
xnor \U$10398 ( \12274 , \12273 , \10176 );
xor \U$10399 ( \12275 , \12270 , \12274 );
xor \U$10400 ( \12276 , \12261 , \12275 );
xor \U$10401 ( \12277 , \12228 , \12276 );
and \U$10402 ( \12278 , \12177 , \12221 );
nor \U$10403 ( \12279 , \12277 , \12278 );
nor \U$10404 ( \12280 , \12224 , \12279 );
nand \U$10405 ( \12281 , \12173 , \12280 );
and \U$10406 ( \12282 , \12232 , \12260 );
and \U$10407 ( \12283 , \12260 , \12275 );
and \U$10408 ( \12284 , \12232 , \12275 );
or \U$10409 ( \12285 , \12282 , \12283 , \12284 );
xor \U$10410 ( \12286 , \11145 , \11149 );
xor \U$10411 ( \12287 , \12286 , \11154 );
and \U$10412 ( \12288 , \10373 , \12253 );
and \U$10413 ( \12289 , \12253 , \12258 );
and \U$10414 ( \12290 , \10373 , \12258 );
or \U$10415 ( \12291 , \12288 , \12289 , \12290 );
and \U$10416 ( \12292 , \12238 , \12242 );
and \U$10417 ( \12293 , \12242 , \12247 );
and \U$10418 ( \12294 , \12238 , \12247 );
or \U$10419 ( \12295 , \12292 , \12293 , \12294 );
xor \U$10420 ( \12296 , \12291 , \12295 );
and \U$10421 ( \12297 , \11090 , \10347 );
and \U$10422 ( \12298 , \10957 , \10345 );
nor \U$10423 ( \12299 , \12297 , \12298 );
xnor \U$10424 ( \12300 , \12299 , \10373 );
xor \U$10425 ( \12301 , \12296 , \12300 );
xor \U$10426 ( \12302 , \12287 , \12301 );
xor \U$10427 ( \12303 , \12285 , \12302 );
and \U$10428 ( \12304 , \12265 , \12269 );
and \U$10429 ( \12305 , \12269 , \12274 );
and \U$10430 ( \12306 , \12265 , \12274 );
or \U$10431 ( \12307 , \12304 , \12305 , \12306 );
and \U$10432 ( \12308 , \12234 , \12248 );
and \U$10433 ( \12309 , \12248 , \12259 );
and \U$10434 ( \12310 , \12234 , \12259 );
or \U$10435 ( \12311 , \12308 , \12309 , \12310 );
xor \U$10436 ( \12312 , \12307 , \12311 );
xor \U$10437 ( \12313 , \11161 , \11165 );
xor \U$10438 ( \12314 , \12313 , \11170 );
xor \U$10439 ( \12315 , \12312 , \12314 );
xor \U$10440 ( \12316 , \12303 , \12315 );
and \U$10441 ( \12317 , \12228 , \12276 );
nor \U$10442 ( \12318 , \12316 , \12317 );
and \U$10443 ( \12319 , \12307 , \12311 );
and \U$10444 ( \12320 , \12311 , \12314 );
and \U$10445 ( \12321 , \12307 , \12314 );
or \U$10446 ( \12322 , \12319 , \12320 , \12321 );
and \U$10447 ( \12323 , \12287 , \12301 );
xor \U$10448 ( \12324 , \12322 , \12323 );
and \U$10449 ( \12325 , \12291 , \12295 );
and \U$10450 ( \12326 , \12295 , \12300 );
and \U$10451 ( \12327 , \12291 , \12300 );
or \U$10452 ( \12328 , \12325 , \12326 , \12327 );
xor \U$10453 ( \12329 , \11181 , \11183 );
xor \U$10454 ( \12330 , \12328 , \12329 );
xor \U$10455 ( \12331 , \11157 , \11173 );
xor \U$10456 ( \12332 , \12331 , \11176 );
xor \U$10457 ( \12333 , \12330 , \12332 );
xor \U$10458 ( \12334 , \12324 , \12333 );
and \U$10459 ( \12335 , \12285 , \12302 );
and \U$10460 ( \12336 , \12302 , \12315 );
and \U$10461 ( \12337 , \12285 , \12315 );
or \U$10462 ( \12338 , \12335 , \12336 , \12337 );
nor \U$10463 ( \12339 , \12334 , \12338 );
nor \U$10464 ( \12340 , \12318 , \12339 );
and \U$10465 ( \12341 , \12328 , \12329 );
and \U$10466 ( \12342 , \12329 , \12332 );
and \U$10467 ( \12343 , \12328 , \12332 );
or \U$10468 ( \12344 , \12341 , \12342 , \12343 );
xor \U$10469 ( \12345 , \11044 , \11060 );
xor \U$10470 ( \12346 , \12345 , \11095 );
xor \U$10471 ( \12347 , \12344 , \12346 );
xor \U$10472 ( \12348 , \11179 , \11184 );
xor \U$10473 ( \12349 , \12348 , \11187 );
xor \U$10474 ( \12350 , \12347 , \12349 );
and \U$10475 ( \12351 , \12322 , \12323 );
and \U$10476 ( \12352 , \12323 , \12333 );
and \U$10477 ( \12353 , \12322 , \12333 );
or \U$10478 ( \12354 , \12351 , \12352 , \12353 );
nor \U$10479 ( \12355 , \12350 , \12354 );
xor \U$10480 ( \12356 , \11190 , \11191 );
xor \U$10481 ( \12357 , \12356 , \11194 );
and \U$10482 ( \12358 , \12344 , \12346 );
and \U$10483 ( \12359 , \12346 , \12349 );
and \U$10484 ( \12360 , \12344 , \12349 );
or \U$10485 ( \12361 , \12358 , \12359 , \12360 );
nor \U$10486 ( \12362 , \12357 , \12361 );
nor \U$10487 ( \12363 , \12355 , \12362 );
nand \U$10488 ( \12364 , \12340 , \12363 );
nor \U$10489 ( \12365 , \12281 , \12364 );
and \U$10490 ( \12366 , \10934 , \10619 );
and \U$10491 ( \12367 , \10865 , \10616 );
nor \U$10492 ( \12368 , \12366 , \12367 );
xnor \U$10493 ( \12369 , \12368 , \10613 );
and \U$10494 ( \12370 , \10741 , \12369 );
and \U$10495 ( \12371 , \10957 , \10655 );
and \U$10496 ( \12372 , \10913 , \10653 );
nor \U$10497 ( \12373 , \12371 , \12372 );
xnor \U$10498 ( \12374 , \12373 , \10681 );
and \U$10499 ( \12375 , \12369 , \12374 );
and \U$10500 ( \12376 , \10741 , \12374 );
or \U$10501 ( \12377 , \12370 , \12375 , \12376 );
and \U$10502 ( \12378 , \10865 , \10619 );
and \U$10503 ( \12379 , \10886 , \10616 );
nor \U$10504 ( \12380 , \12378 , \12379 );
xnor \U$10505 ( \12381 , \12380 , \10613 );
and \U$10506 ( \12382 , \10913 , \10655 );
and \U$10507 ( \12383 , \10934 , \10653 );
nor \U$10508 ( \12384 , \12382 , \12383 );
xnor \U$10509 ( \12385 , \12384 , \10681 );
xor \U$10510 ( \12386 , \12381 , \12385 );
and \U$10511 ( \12387 , \11090 , \10715 );
and \U$10512 ( \12388 , \10957 , \10713 );
nor \U$10513 ( \12389 , \12387 , \12388 );
xnor \U$10514 ( \12390 , \12389 , \10741 );
xor \U$10515 ( \12391 , \12386 , \12390 );
xor \U$10516 ( \12392 , \12377 , \12391 );
nand \U$10517 ( \12393 , \11090 , \10713 );
xnor \U$10518 ( \12394 , \12393 , \10741 );
xor \U$10519 ( \12395 , \10741 , \12369 );
xor \U$10520 ( \12396 , \12395 , \12374 );
and \U$10521 ( \12397 , \12394 , \12396 );
nor \U$10522 ( \12398 , \12392 , \12397 );
and \U$10523 ( \12399 , \12381 , \12385 );
and \U$10524 ( \12400 , \12385 , \12390 );
and \U$10525 ( \12401 , \12381 , \12390 );
or \U$10526 ( \12402 , \12399 , \12400 , \12401 );
xor \U$10527 ( \12403 , \12112 , \12114 );
xor \U$10528 ( \12404 , \12402 , \12403 );
xor \U$10529 ( \12405 , \10799 , \12100 );
xor \U$10530 ( \12406 , \12405 , \12105 );
xor \U$10531 ( \12407 , \12404 , \12406 );
and \U$10532 ( \12408 , \12377 , \12391 );
nor \U$10533 ( \12409 , \12407 , \12408 );
nor \U$10534 ( \12410 , \12398 , \12409 );
xor \U$10535 ( \12411 , \12023 , \12027 );
xor \U$10536 ( \12412 , \12411 , \12032 );
xor \U$10537 ( \12413 , \12108 , \12115 );
xor \U$10538 ( \12414 , \12413 , \12120 );
xor \U$10539 ( \12415 , \12412 , \12414 );
and \U$10540 ( \12416 , \12402 , \12403 );
and \U$10541 ( \12417 , \12403 , \12406 );
and \U$10542 ( \12418 , \12402 , \12406 );
or \U$10543 ( \12419 , \12416 , \12417 , \12418 );
nor \U$10544 ( \12420 , \12415 , \12419 );
xor \U$10545 ( \12421 , \12123 , \12125 );
and \U$10546 ( \12422 , \12412 , \12414 );
nor \U$10547 ( \12423 , \12421 , \12422 );
nor \U$10548 ( \12424 , \12420 , \12423 );
nand \U$10549 ( \12425 , \12410 , \12424 );
and \U$10550 ( \12426 , \10913 , \10619 );
and \U$10551 ( \12427 , \10934 , \10616 );
nor \U$10552 ( \12428 , \12426 , \12427 );
xnor \U$10553 ( \12429 , \12428 , \10613 );
and \U$10554 ( \12430 , \11090 , \10655 );
and \U$10555 ( \12431 , \10957 , \10653 );
nor \U$10556 ( \12432 , \12430 , \12431 );
xnor \U$10557 ( \12433 , \12432 , \10681 );
xor \U$10558 ( \12434 , \12429 , \12433 );
and \U$10559 ( \12435 , \10957 , \10619 );
and \U$10560 ( \12436 , \10913 , \10616 );
nor \U$10561 ( \12437 , \12435 , \12436 );
xnor \U$10562 ( \12438 , \12437 , \10613 );
and \U$10563 ( \12439 , \12438 , \10681 );
nor \U$10564 ( \12440 , \12434 , \12439 );
xor \U$10565 ( \12441 , \12394 , \12396 );
and \U$10566 ( \12442 , \12429 , \12433 );
nor \U$10567 ( \12443 , \12441 , \12442 );
nor \U$10568 ( \12444 , \12440 , \12443 );
xor \U$10569 ( \12445 , \12438 , \10681 );
nand \U$10570 ( \12446 , \11090 , \10653 );
xnor \U$10571 ( \12447 , \12446 , \10681 );
nor \U$10572 ( \12448 , \12445 , \12447 );
and \U$10573 ( \12449 , \11090 , \10619 );
and \U$10574 ( \12450 , \10957 , \10616 );
nor \U$10575 ( \12451 , \12449 , \12450 );
xnor \U$10576 ( \12452 , \12451 , \10613 );
nand \U$10577 ( \12453 , \11090 , \10616 );
xnor \U$10578 ( \12454 , \12453 , \10613 );
and \U$10579 ( \12455 , \12454 , \10613 );
nand \U$10580 ( \12456 , \12452 , \12455 );
or \U$10581 ( \12457 , \12448 , \12456 );
nand \U$10582 ( \12458 , \12445 , \12447 );
nand \U$10583 ( \12459 , \12457 , \12458 );
and \U$10584 ( \12460 , \12444 , \12459 );
nand \U$10585 ( \12461 , \12434 , \12439 );
or \U$10586 ( \12462 , \12443 , \12461 );
nand \U$10587 ( \12463 , \12441 , \12442 );
nand \U$10588 ( \12464 , \12462 , \12463 );
nor \U$10589 ( \12465 , \12460 , \12464 );
or \U$10590 ( \12466 , \12425 , \12465 );
nand \U$10591 ( \12467 , \12392 , \12397 );
or \U$10592 ( \12468 , \12409 , \12467 );
nand \U$10593 ( \12469 , \12407 , \12408 );
nand \U$10594 ( \12470 , \12468 , \12469 );
and \U$10595 ( \12471 , \12424 , \12470 );
nand \U$10596 ( \12472 , \12415 , \12419 );
or \U$10597 ( \12473 , \12423 , \12472 );
nand \U$10598 ( \12474 , \12421 , \12422 );
nand \U$10599 ( \12475 , \12473 , \12474 );
nor \U$10600 ( \12476 , \12471 , \12475 );
nand \U$10601 ( \12477 , \12466 , \12476 );
and \U$10602 ( \12478 , \12365 , \12477 );
nand \U$10603 ( \12479 , \12096 , \12126 );
or \U$10604 ( \12480 , \12172 , \12479 );
nand \U$10605 ( \12481 , \12167 , \12171 );
nand \U$10606 ( \12482 , \12480 , \12481 );
and \U$10607 ( \12483 , \12280 , \12482 );
nand \U$10608 ( \12484 , \12222 , \12223 );
or \U$10609 ( \12485 , \12279 , \12484 );
nand \U$10610 ( \12486 , \12277 , \12278 );
nand \U$10611 ( \12487 , \12485 , \12486 );
nor \U$10612 ( \12488 , \12483 , \12487 );
or \U$10613 ( \12489 , \12364 , \12488 );
nand \U$10614 ( \12490 , \12316 , \12317 );
or \U$10615 ( \12491 , \12339 , \12490 );
nand \U$10616 ( \12492 , \12334 , \12338 );
nand \U$10617 ( \12493 , \12491 , \12492 );
and \U$10618 ( \12494 , \12363 , \12493 );
nand \U$10619 ( \12495 , \12350 , \12354 );
or \U$10620 ( \12496 , \12362 , \12495 );
nand \U$10621 ( \12497 , \12357 , \12361 );
nand \U$10622 ( \12498 , \12496 , \12497 );
nor \U$10623 ( \12499 , \12494 , \12498 );
nand \U$10624 ( \12500 , \12489 , \12499 );
nor \U$10625 ( \12501 , \12478 , \12500 );
or \U$10626 ( \12502 , \12019 , \12501 );
nand \U$10627 ( \12503 , \11141 , \11197 );
or \U$10628 ( \12504 , \11273 , \12503 );
nand \U$10629 ( \12505 , \11271 , \11272 );
nand \U$10630 ( \12506 , \12504 , \12505 );
and \U$10631 ( \12507 , \11426 , \12506 );
nand \U$10632 ( \12508 , \11348 , \11349 );
or \U$10633 ( \12509 , \11425 , \12508 );
nand \U$10634 ( \12510 , \11420 , \11424 );
nand \U$10635 ( \12511 , \12509 , \12510 );
nor \U$10636 ( \12512 , \12507 , \12511 );
or \U$10637 ( \12513 , \11722 , \12512 );
nand \U$10638 ( \12514 , \11497 , \11501 );
or \U$10639 ( \12515 , \11578 , \12514 );
nand \U$10640 ( \12516 , \11573 , \11577 );
nand \U$10641 ( \12517 , \12515 , \12516 );
and \U$10642 ( \12518 , \11721 , \12517 );
nand \U$10643 ( \12519 , \11646 , \11650 );
or \U$10644 ( \12520 , \11720 , \12519 );
nand \U$10645 ( \12521 , \11715 , \11719 );
nand \U$10646 ( \12522 , \12520 , \12521 );
nor \U$10647 ( \12523 , \12518 , \12522 );
nand \U$10648 ( \12524 , \12513 , \12523 );
and \U$10649 ( \12525 , \12018 , \12524 );
nand \U$10650 ( \12526 , \11779 , \11783 );
or \U$10651 ( \12527 , \11844 , \12526 );
nand \U$10652 ( \12528 , \11839 , \11843 );
nand \U$10653 ( \12529 , \12527 , \12528 );
and \U$10654 ( \12530 , \11940 , \12529 );
nand \U$10655 ( \12531 , \11896 , \11900 );
or \U$10656 ( \12532 , \11939 , \12531 );
nand \U$10657 ( \12533 , \11934 , \11938 );
nand \U$10658 ( \12534 , \12532 , \12533 );
nor \U$10659 ( \12535 , \12530 , \12534 );
or \U$10660 ( \12536 , \12017 , \12535 );
nand \U$10661 ( \12537 , \11966 , \11970 );
or \U$10662 ( \12538 , \11992 , \12537 );
nand \U$10663 ( \12539 , \11987 , \11991 );
nand \U$10664 ( \12540 , \12538 , \12539 );
and \U$10665 ( \12541 , \12016 , \12540 );
nand \U$10666 ( \12542 , \12003 , \12007 );
or \U$10667 ( \12543 , \12015 , \12542 );
nand \U$10668 ( \12544 , \12010 , \12014 );
nand \U$10669 ( \12545 , \12543 , \12544 );
nor \U$10670 ( \12546 , \12541 , \12545 );
nand \U$10671 ( \12547 , \12536 , \12546 );
nor \U$10672 ( \12548 , \12525 , \12547 );
nand \U$10673 ( \12549 , \12502 , \12548 );
not \U$10674 ( \12550 , \12549 );
xor \U$10675 ( \12551 , \10609 , \12550 );
buf g4b72_GF_PartitionCandidate( \12552_nG4b72 , \12551 );
buf \U$10680 ( \12553 , RI2b5e785db058_15);
buf \U$10681 ( \12554 , RI2b5e785dafe0_16);
buf \U$10682 ( \12555 , RI2b5e785daf68_17);
buf \U$10683 ( \12556 , RI2b5e785daef0_18);
buf \U$10684 ( \12557 , RI2b5e785dae78_19);
buf \U$10685 ( \12558 , RI2b5e785dae00_20);
buf \U$10686 ( \12559 , RI2b5e785dad88_21);
buf \U$10687 ( \12560 , RI2b5e785dad10_22);
buf \U$10688 ( \12561 , RI2b5e785dac98_23);
buf \U$10689 ( \12562 , RI2b5e785dac20_24);
buf \U$10690 ( \12563 , RI2b5e785daba8_25);
and \U$10691 ( \12564 , \12562 , \12563 );
and \U$10692 ( \12565 , \12561 , \12564 );
and \U$10693 ( \12566 , \12560 , \12565 );
and \U$10694 ( \12567 , \12559 , \12566 );
and \U$10695 ( \12568 , \12558 , \12567 );
and \U$10696 ( \12569 , \12557 , \12568 );
and \U$10697 ( \12570 , \12556 , \12569 );
and \U$10698 ( \12571 , \12555 , \12570 );
and \U$10699 ( \12572 , \12554 , \12571 );
xor \U$10700 ( \12573 , \12553 , \12572 );
buf \U$10701 ( \12574 , \12573 );
buf \U$10702 ( \12575 , \12574 );
buf \U$10703 ( \12576 , RI2b5e785ae3a0_613);
buf \U$10704 ( \12577 , RI2b5e785ae580_609);
buf \U$10705 ( \12578 , RI2b5e785ae5f8_608);
buf \U$10706 ( \12579 , RI2b5e785ae670_607);
buf \U$10707 ( \12580 , RI2b5e785ae6e8_606);
buf \U$10708 ( \12581 , RI2b5e785ae760_605);
buf \U$10709 ( \12582 , RI2b5e785ae7d8_604);
buf \U$10710 ( \12583 , RI2b5e785ae850_603);
buf \U$10711 ( \12584 , RI2b5e785ae8c8_602);
buf \U$10712 ( \12585 , RI2b5e785ae940_601);
buf \U$10713 ( \12586 , RI2b5e785ae3a0_613);
buf \U$10714 ( \12587 , RI2b5e785ae418_612);
buf \U$10715 ( \12588 , RI2b5e785ae490_611);
buf \U$10716 ( \12589 , RI2b5e785ae508_610);
and \U$10717 ( \12590 , \12586 , \12587 , \12588 , \12589 );
nor \U$10718 ( \12591 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12590 );
buf \U$10719 ( \12592 , \12591 );
buf \U$10720 ( \12593 , \12592 );
xor \U$10721 ( \12594 , \12576 , \12593 );
buf \U$10722 ( \12595 , \12594 );
buf \U$10723 ( \12596 , RI2b5e785ae418_612);
and \U$10724 ( \12597 , \12576 , \12593 );
xor \U$10725 ( \12598 , \12596 , \12597 );
buf \U$10726 ( \12599 , \12598 );
buf \U$10727 ( \12600 , RI2b5e785ae490_611);
and \U$10728 ( \12601 , \12596 , \12597 );
xor \U$10729 ( \12602 , \12600 , \12601 );
buf \U$10730 ( \12603 , \12602 );
buf \U$10731 ( \12604 , RI2b5e785ae508_610);
and \U$10732 ( \12605 , \12600 , \12601 );
xor \U$10733 ( \12606 , \12604 , \12605 );
buf \U$10734 ( \12607 , \12606 );
buf \U$10735 ( \12608 , RI2b5e785ae580_609);
and \U$10736 ( \12609 , \12604 , \12605 );
xor \U$10737 ( \12610 , \12608 , \12609 );
buf \U$10738 ( \12611 , \12610 );
not \U$10739 ( \12612 , \12611 );
buf \U$10740 ( \12613 , RI2b5e785ae5f8_608);
and \U$10741 ( \12614 , \12608 , \12609 );
xor \U$10742 ( \12615 , \12613 , \12614 );
buf \U$10743 ( \12616 , \12615 );
buf \U$10744 ( \12617 , RI2b5e785ae670_607);
and \U$10745 ( \12618 , \12613 , \12614 );
xor \U$10746 ( \12619 , \12617 , \12618 );
buf \U$10747 ( \12620 , \12619 );
buf \U$10748 ( \12621 , RI2b5e785ae6e8_606);
and \U$10749 ( \12622 , \12617 , \12618 );
xor \U$10750 ( \12623 , \12621 , \12622 );
buf \U$10751 ( \12624 , \12623 );
buf \U$10752 ( \12625 , RI2b5e785ae760_605);
and \U$10753 ( \12626 , \12621 , \12622 );
xor \U$10754 ( \12627 , \12625 , \12626 );
buf \U$10755 ( \12628 , \12627 );
buf \U$10756 ( \12629 , RI2b5e785ae7d8_604);
and \U$10757 ( \12630 , \12625 , \12626 );
xor \U$10758 ( \12631 , \12629 , \12630 );
buf \U$10759 ( \12632 , \12631 );
buf \U$10760 ( \12633 , RI2b5e785ae850_603);
and \U$10761 ( \12634 , \12629 , \12630 );
xor \U$10762 ( \12635 , \12633 , \12634 );
buf \U$10763 ( \12636 , \12635 );
buf \U$10764 ( \12637 , RI2b5e785ae8c8_602);
and \U$10765 ( \12638 , \12633 , \12634 );
xor \U$10766 ( \12639 , \12637 , \12638 );
buf \U$10767 ( \12640 , \12639 );
buf \U$10768 ( \12641 , RI2b5e785ae940_601);
and \U$10769 ( \12642 , \12637 , \12638 );
xor \U$10770 ( \12643 , \12641 , \12642 );
buf \U$10771 ( \12644 , \12643 );
nor \U$10772 ( \12645 , \12595 , \12599 , \12603 , \12607 , \12612 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10773 ( \12646 , RI2b5e785daa40_28, \12645 );
not \U$10774 ( \12647 , \12595 );
not \U$10775 ( \12648 , \12599 );
not \U$10776 ( \12649 , \12603 );
not \U$10777 ( \12650 , \12607 );
nor \U$10778 ( \12651 , \12647 , \12648 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10779 ( \12652 , RI2b5e78549540_41, \12651 );
nor \U$10780 ( \12653 , \12595 , \12648 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10781 ( \12654 , RI2b5e785388a8_54, \12653 );
nor \U$10782 ( \12655 , \12647 , \12599 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10783 ( \12656 , RI2b5e784a6330_67, \12655 );
nor \U$10784 ( \12657 , \12595 , \12599 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10785 ( \12658 , RI2b5e78495698_80, \12657 );
nor \U$10786 ( \12659 , \12647 , \12648 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10787 ( \12660 , RI2b5e78495080_93, \12659 );
nor \U$10788 ( \12661 , \12595 , \12648 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10789 ( \12662 , RI2b5e78403b80_106, \12661 );
nor \U$10790 ( \12663 , \12647 , \12599 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10791 ( \12664 , RI2b5e775b1e60_119, \12663 );
nor \U$10792 ( \12665 , \12595 , \12599 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10793 ( \12666 , RI2b5e7750bdf8_132, \12665 );
nor \U$10794 ( \12667 , \12647 , \12648 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10795 ( \12668 , RI2b5e774ff5d0_145, \12667 );
nor \U$10796 ( \12669 , \12595 , \12648 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10797 ( \12670 , RI2b5e774f65e8_158, \12669 );
nor \U$10798 ( \12671 , \12647 , \12599 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10799 ( \12672 , RI2b5e774eabd0_171, \12671 );
nor \U$10800 ( \12673 , \12595 , \12599 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10801 ( \12674 , RI2b5e774de3a8_184, \12673 );
nor \U$10802 ( \12675 , \12647 , \12648 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10803 ( \12676 , RI2b5e774d53c0_197, \12675 );
nor \U$10804 ( \12677 , \12595 , \12648 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10805 ( \12678 , RI2b5e785f4300_210, \12677 );
nor \U$10806 ( \12679 , \12647 , \12599 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10807 ( \12680 , RI2b5e785f3ce8_223, \12679 );
nor \U$10808 ( \12681 , \12595 , \12599 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$10809 ( \12682 , RI2b5e785eb0c0_236, \12681 );
or \U$10810 ( \12683 , \12646 , \12652 , \12654 , \12656 , \12658 , \12660 , \12662 , \12664 , \12666 , \12668 , \12670 , \12672 , \12674 , \12676 , \12678 , \12680 , \12682 );
buf \U$10811 ( \12684 , \12616 );
buf \U$10812 ( \12685 , \12620 );
buf \U$10813 ( \12686 , \12624 );
buf \U$10814 ( \12687 , \12628 );
buf \U$10815 ( \12688 , \12632 );
buf \U$10816 ( \12689 , \12636 );
buf \U$10817 ( \12690 , \12640 );
buf \U$10818 ( \12691 , \12644 );
buf \U$10819 ( \12692 , \12611 );
buf \U$10820 ( \12693 , \12595 );
buf \U$10821 ( \12694 , \12599 );
buf \U$10822 ( \12695 , \12603 );
buf \U$10823 ( \12696 , \12607 );
or \U$10824 ( \12697 , \12693 , \12694 , \12695 , \12696 );
and \U$10825 ( \12698 , \12692 , \12697 );
or \U$10826 ( \12699 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12698 );
buf \U$10827 ( \12700 , \12699 );
_DC g3b20 ( \12701_nG3b20 , \12683 , \12700 );
buf \U$10828 ( \12702 , \12701_nG3b20 );
not \U$10829 ( \12703 , \12702 );
xor \U$10830 ( \12704 , \12575 , \12703 );
xor \U$10831 ( \12705 , \12554 , \12571 );
buf \U$10832 ( \12706 , \12705 );
buf \U$10833 ( \12707 , \12706 );
and \U$10834 ( \12708 , RI2b5e785da9c8_29, \12645 );
and \U$10835 ( \12709 , RI2b5e785494c8_42, \12651 );
and \U$10836 ( \12710 , RI2b5e78538830_55, \12653 );
and \U$10837 ( \12711 , RI2b5e784a62b8_68, \12655 );
and \U$10838 ( \12712 , RI2b5e78495620_81, \12657 );
and \U$10839 ( \12713 , RI2b5e78495008_94, \12659 );
and \U$10840 ( \12714 , RI2b5e78403b08_107, \12661 );
and \U$10841 ( \12715 , RI2b5e775b1de8_120, \12663 );
and \U$10842 ( \12716 , RI2b5e7750bd80_133, \12665 );
and \U$10843 ( \12717 , RI2b5e774ff558_146, \12667 );
and \U$10844 ( \12718 , RI2b5e774f6570_159, \12669 );
and \U$10845 ( \12719 , RI2b5e774eab58_172, \12671 );
and \U$10846 ( \12720 , RI2b5e774de330_185, \12673 );
and \U$10847 ( \12721 , RI2b5e774d5348_198, \12675 );
and \U$10848 ( \12722 , RI2b5e785f4288_211, \12677 );
and \U$10849 ( \12723 , RI2b5e785f3658_224, \12679 );
and \U$10850 ( \12724 , RI2b5e785eb048_237, \12681 );
or \U$10851 ( \12725 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 );
_DC g3afc ( \12726_nG3afc , \12725 , \12700 );
buf \U$10852 ( \12727 , \12726_nG3afc );
not \U$10853 ( \12728 , \12727 );
and \U$10854 ( \12729 , \12707 , \12728 );
xor \U$10855 ( \12730 , \12555 , \12570 );
buf \U$10856 ( \12731 , \12730 );
buf \U$10857 ( \12732 , \12731 );
and \U$10858 ( \12733 , RI2b5e785da950_30, \12645 );
and \U$10859 ( \12734 , RI2b5e78549450_43, \12651 );
and \U$10860 ( \12735 , RI2b5e785387b8_56, \12653 );
and \U$10861 ( \12736 , RI2b5e784a6240_69, \12655 );
and \U$10862 ( \12737 , RI2b5e784955a8_82, \12657 );
and \U$10863 ( \12738 , RI2b5e78494f90_95, \12659 );
and \U$10864 ( \12739 , RI2b5e78403a90_108, \12661 );
and \U$10865 ( \12740 , RI2b5e775b1d70_121, \12663 );
and \U$10866 ( \12741 , RI2b5e7750bd08_134, \12665 );
and \U$10867 ( \12742 , RI2b5e774ff4e0_147, \12667 );
and \U$10868 ( \12743 , RI2b5e774f64f8_160, \12669 );
and \U$10869 ( \12744 , RI2b5e774eaae0_173, \12671 );
and \U$10870 ( \12745 , RI2b5e774de2b8_186, \12673 );
and \U$10871 ( \12746 , RI2b5e774d52d0_199, \12675 );
and \U$10872 ( \12747 , RI2b5e785f4210_212, \12677 );
and \U$10873 ( \12748 , RI2b5e785eb5e8_225, \12679 );
and \U$10874 ( \12749 , RI2b5e785e6c50_238, \12681 );
or \U$10875 ( \12750 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 );
_DC g3969 ( \12751_nG3969 , \12750 , \12700 );
buf \U$10876 ( \12752 , \12751_nG3969 );
not \U$10877 ( \12753 , \12752 );
and \U$10878 ( \12754 , \12732 , \12753 );
xor \U$10879 ( \12755 , \12556 , \12569 );
buf \U$10880 ( \12756 , \12755 );
buf \U$10881 ( \12757 , \12756 );
and \U$10882 ( \12758 , RI2b5e785da8d8_31, \12645 );
and \U$10883 ( \12759 , RI2b5e785493d8_44, \12651 );
and \U$10884 ( \12760 , RI2b5e78538740_57, \12653 );
and \U$10885 ( \12761 , RI2b5e784a61c8_70, \12655 );
and \U$10886 ( \12762 , RI2b5e78495530_83, \12657 );
and \U$10887 ( \12763 , RI2b5e78494f18_96, \12659 );
and \U$10888 ( \12764 , RI2b5e78403a18_109, \12661 );
and \U$10889 ( \12765 , RI2b5e775b1cf8_122, \12663 );
and \U$10890 ( \12766 , RI2b5e7750bc90_135, \12665 );
and \U$10891 ( \12767 , RI2b5e774ff468_148, \12667 );
and \U$10892 ( \12768 , RI2b5e774f6480_161, \12669 );
and \U$10893 ( \12769 , RI2b5e774eaa68_174, \12671 );
and \U$10894 ( \12770 , RI2b5e774de240_187, \12673 );
and \U$10895 ( \12771 , RI2b5e774d5258_200, \12675 );
and \U$10896 ( \12772 , RI2b5e785f4198_213, \12677 );
and \U$10897 ( \12773 , RI2b5e785eb570_226, \12679 );
and \U$10898 ( \12774 , RI2b5e785e6bd8_239, \12681 );
or \U$10899 ( \12775 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 );
_DC g3945 ( \12776_nG3945 , \12775 , \12700 );
buf \U$10900 ( \12777 , \12776_nG3945 );
not \U$10901 ( \12778 , \12777 );
and \U$10902 ( \12779 , \12757 , \12778 );
xor \U$10903 ( \12780 , \12557 , \12568 );
buf \U$10904 ( \12781 , \12780 );
buf \U$10905 ( \12782 , \12781 );
and \U$10906 ( \12783 , RI2b5e785da860_32, \12645 );
and \U$10907 ( \12784 , RI2b5e78549360_45, \12651 );
and \U$10908 ( \12785 , RI2b5e785386c8_58, \12653 );
and \U$10909 ( \12786 , RI2b5e784a6150_71, \12655 );
and \U$10910 ( \12787 , RI2b5e784954b8_84, \12657 );
and \U$10911 ( \12788 , RI2b5e78494ea0_97, \12659 );
and \U$10912 ( \12789 , RI2b5e784039a0_110, \12661 );
and \U$10913 ( \12790 , RI2b5e775b1c80_123, \12663 );
and \U$10914 ( \12791 , RI2b5e7750bc18_136, \12665 );
and \U$10915 ( \12792 , RI2b5e774ff3f0_149, \12667 );
and \U$10916 ( \12793 , RI2b5e774f6408_162, \12669 );
and \U$10917 ( \12794 , RI2b5e774ea9f0_175, \12671 );
and \U$10918 ( \12795 , RI2b5e774de1c8_188, \12673 );
and \U$10919 ( \12796 , RI2b5e774d51e0_201, \12675 );
and \U$10920 ( \12797 , RI2b5e785f4120_214, \12677 );
and \U$10921 ( \12798 , RI2b5e785eb4f8_227, \12679 );
and \U$10922 ( \12799 , RI2b5e785e64d0_240, \12681 );
or \U$10923 ( \12800 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 );
_DC g37c6 ( \12801_nG37c6 , \12800 , \12700 );
buf \U$10924 ( \12802 , \12801_nG37c6 );
not \U$10925 ( \12803 , \12802 );
and \U$10926 ( \12804 , \12782 , \12803 );
xor \U$10927 ( \12805 , \12558 , \12567 );
buf \U$10928 ( \12806 , \12805 );
buf \U$10929 ( \12807 , \12806 );
and \U$10930 ( \12808 , RI2b5e78549900_33, \12645 );
and \U$10931 ( \12809 , RI2b5e78538c68_46, \12651 );
and \U$10932 ( \12810 , RI2b5e78538650_59, \12653 );
and \U$10933 ( \12811 , RI2b5e784a60d8_72, \12655 );
and \U$10934 ( \12812 , RI2b5e78495440_85, \12657 );
and \U$10935 ( \12813 , RI2b5e78494e28_98, \12659 );
and \U$10936 ( \12814 , RI2b5e78403928_111, \12661 );
and \U$10937 ( \12815 , RI2b5e775b1c08_124, \12663 );
and \U$10938 ( \12816 , RI2b5e7750bba0_137, \12665 );
and \U$10939 ( \12817 , RI2b5e774ff378_150, \12667 );
and \U$10940 ( \12818 , RI2b5e774f6390_163, \12669 );
and \U$10941 ( \12819 , RI2b5e774ea978_176, \12671 );
and \U$10942 ( \12820 , RI2b5e774de150_189, \12673 );
and \U$10943 ( \12821 , RI2b5e774d5168_202, \12675 );
and \U$10944 ( \12822 , RI2b5e785f40a8_215, \12677 );
and \U$10945 ( \12823 , RI2b5e785eb480_228, \12679 );
and \U$10946 ( \12824 , RI2b5e785da608_241, \12681 );
or \U$10947 ( \12825 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 );
_DC g37a2 ( \12826_nG37a2 , \12825 , \12700 );
buf \U$10948 ( \12827 , \12826_nG37a2 );
not \U$10949 ( \12828 , \12827 );
and \U$10950 ( \12829 , \12807 , \12828 );
xor \U$10951 ( \12830 , \12559 , \12566 );
buf \U$10952 ( \12831 , \12830 );
buf \U$10953 ( \12832 , \12831 );
and \U$10954 ( \12833 , RI2b5e78549888_34, \12645 );
and \U$10955 ( \12834 , RI2b5e78538bf0_47, \12651 );
and \U$10956 ( \12835 , RI2b5e785385d8_60, \12653 );
and \U$10957 ( \12836 , RI2b5e784a6060_73, \12655 );
and \U$10958 ( \12837 , RI2b5e784953c8_86, \12657 );
and \U$10959 ( \12838 , RI2b5e78403ec8_99, \12659 );
and \U$10960 ( \12839 , RI2b5e775b21a8_112, \12661 );
and \U$10961 ( \12840 , RI2b5e775b1b90_125, \12663 );
and \U$10962 ( \12841 , RI2b5e7750bb28_138, \12665 );
and \U$10963 ( \12842 , RI2b5e774ff300_151, \12667 );
and \U$10964 ( \12843 , RI2b5e774f6318_164, \12669 );
and \U$10965 ( \12844 , RI2b5e774ea900_177, \12671 );
and \U$10966 ( \12845 , RI2b5e774de0d8_190, \12673 );
and \U$10967 ( \12846 , RI2b5e774d50f0_203, \12675 );
and \U$10968 ( \12847 , RI2b5e785f4030_216, \12677 );
and \U$10969 ( \12848 , RI2b5e785eb408_229, \12679 );
and \U$10970 ( \12849 , RI2b5e785da590_242, \12681 );
or \U$10971 ( \12850 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 );
_DC g3657 ( \12851_nG3657 , \12850 , \12700 );
buf \U$10972 ( \12852 , \12851_nG3657 );
not \U$10973 ( \12853 , \12852 );
and \U$10974 ( \12854 , \12832 , \12853 );
xor \U$10975 ( \12855 , \12560 , \12565 );
buf \U$10976 ( \12856 , \12855 );
buf \U$10977 ( \12857 , \12856 );
and \U$10978 ( \12858 , RI2b5e78549810_35, \12645 );
and \U$10979 ( \12859 , RI2b5e78538b78_48, \12651 );
and \U$10980 ( \12860 , RI2b5e78538560_61, \12653 );
and \U$10981 ( \12861 , RI2b5e784a5fe8_74, \12655 );
and \U$10982 ( \12862 , RI2b5e78495350_87, \12657 );
and \U$10983 ( \12863 , RI2b5e78403e50_100, \12659 );
and \U$10984 ( \12864 , RI2b5e775b2130_113, \12661 );
and \U$10985 ( \12865 , RI2b5e775b1b18_126, \12663 );
and \U$10986 ( \12866 , RI2b5e7750bab0_139, \12665 );
and \U$10987 ( \12867 , RI2b5e774ff288_152, \12667 );
and \U$10988 ( \12868 , RI2b5e774f62a0_165, \12669 );
and \U$10989 ( \12869 , RI2b5e774ea888_178, \12671 );
and \U$10990 ( \12870 , RI2b5e774de060_191, \12673 );
and \U$10991 ( \12871 , RI2b5e774d5078_204, \12675 );
and \U$10992 ( \12872 , RI2b5e785f3fb8_217, \12677 );
and \U$10993 ( \12873 , RI2b5e785eb390_230, \12679 );
and \U$10994 ( \12874 , RI2b5e785da518_243, \12681 );
or \U$10995 ( \12875 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 );
_DC g3633 ( \12876_nG3633 , \12875 , \12700 );
buf \U$10996 ( \12877 , \12876_nG3633 );
not \U$10997 ( \12878 , \12877 );
and \U$10998 ( \12879 , \12857 , \12878 );
xor \U$10999 ( \12880 , \12561 , \12564 );
buf \U$11000 ( \12881 , \12880 );
buf \U$11001 ( \12882 , \12881 );
and \U$11002 ( \12883 , RI2b5e78549798_36, \12645 );
and \U$11003 ( \12884 , RI2b5e78538b00_49, \12651 );
and \U$11004 ( \12885 , RI2b5e785384e8_62, \12653 );
and \U$11005 ( \12886 , RI2b5e784a5f70_75, \12655 );
and \U$11006 ( \12887 , RI2b5e784952d8_88, \12657 );
and \U$11007 ( \12888 , RI2b5e78403dd8_101, \12659 );
and \U$11008 ( \12889 , RI2b5e775b20b8_114, \12661 );
and \U$11009 ( \12890 , RI2b5e775b1aa0_127, \12663 );
and \U$11010 ( \12891 , RI2b5e7750ba38_140, \12665 );
and \U$11011 ( \12892 , RI2b5e774ff210_153, \12667 );
and \U$11012 ( \12893 , RI2b5e774f6228_166, \12669 );
and \U$11013 ( \12894 , RI2b5e774ea810_179, \12671 );
and \U$11014 ( \12895 , RI2b5e774ddfe8_192, \12673 );
and \U$11015 ( \12896 , RI2b5e774d5000_205, \12675 );
and \U$11016 ( \12897 , RI2b5e785f3f40_218, \12677 );
and \U$11017 ( \12898 , RI2b5e785eb318_231, \12679 );
and \U$11018 ( \12899 , RI2b5e785da4a0_244, \12681 );
or \U$11019 ( \12900 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 );
_DC g3518 ( \12901_nG3518 , \12900 , \12700 );
buf \U$11020 ( \12902 , \12901_nG3518 );
not \U$11021 ( \12903 , \12902 );
and \U$11022 ( \12904 , \12882 , \12903 );
xor \U$11023 ( \12905 , \12562 , \12563 );
buf \U$11024 ( \12906 , \12905 );
buf \U$11025 ( \12907 , \12906 );
and \U$11026 ( \12908 , RI2b5e78549720_37, \12645 );
and \U$11027 ( \12909 , RI2b5e78538a88_50, \12651 );
and \U$11028 ( \12910 , RI2b5e78538470_63, \12653 );
and \U$11029 ( \12911 , RI2b5e784a5ef8_76, \12655 );
and \U$11030 ( \12912 , RI2b5e78495260_89, \12657 );
and \U$11031 ( \12913 , RI2b5e78403d60_102, \12659 );
and \U$11032 ( \12914 , RI2b5e775b2040_115, \12661 );
and \U$11033 ( \12915 , RI2b5e775b1a28_128, \12663 );
and \U$11034 ( \12916 , RI2b5e7750b9c0_141, \12665 );
and \U$11035 ( \12917 , RI2b5e774ff198_154, \12667 );
and \U$11036 ( \12918 , RI2b5e774f61b0_167, \12669 );
and \U$11037 ( \12919 , RI2b5e774ea798_180, \12671 );
and \U$11038 ( \12920 , RI2b5e774ddf70_193, \12673 );
and \U$11039 ( \12921 , RI2b5e774d4f88_206, \12675 );
and \U$11040 ( \12922 , RI2b5e785f3ec8_219, \12677 );
and \U$11041 ( \12923 , RI2b5e785eb2a0_232, \12679 );
and \U$11042 ( \12924 , RI2b5e785da428_245, \12681 );
or \U$11043 ( \12925 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 );
_DC g3531 ( \12926_nG3531 , \12925 , \12700 );
buf \U$11044 ( \12927 , \12926_nG3531 );
not \U$11045 ( \12928 , \12927 );
and \U$11046 ( \12929 , \12907 , \12928 );
not \U$11047 ( \12930 , \12563 );
buf \U$11048 ( \12931 , \12930 );
buf \U$11049 ( \12932 , \12931 );
and \U$11050 ( \12933 , RI2b5e785496a8_38, \12645 );
and \U$11051 ( \12934 , RI2b5e78538a10_51, \12651 );
and \U$11052 ( \12935 , RI2b5e785383f8_64, \12653 );
and \U$11053 ( \12936 , RI2b5e784a5e80_77, \12655 );
and \U$11054 ( \12937 , RI2b5e784951e8_90, \12657 );
and \U$11055 ( \12938 , RI2b5e78403ce8_103, \12659 );
and \U$11056 ( \12939 , RI2b5e775b1fc8_116, \12661 );
and \U$11057 ( \12940 , RI2b5e775b19b0_129, \12663 );
and \U$11058 ( \12941 , RI2b5e7750b948_142, \12665 );
and \U$11059 ( \12942 , RI2b5e774ff120_155, \12667 );
and \U$11060 ( \12943 , RI2b5e774f6138_168, \12669 );
and \U$11061 ( \12944 , RI2b5e774ea720_181, \12671 );
and \U$11062 ( \12945 , RI2b5e774ddef8_194, \12673 );
and \U$11063 ( \12946 , RI2b5e774d4f10_207, \12675 );
and \U$11064 ( \12947 , RI2b5e785f3e50_220, \12677 );
and \U$11065 ( \12948 , RI2b5e785eb228_233, \12679 );
and \U$11066 ( \12949 , RI2b5e785da3b0_246, \12681 );
or \U$11067 ( \12950 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 );
_DC g342e ( \12951_nG342e , \12950 , \12700 );
buf \U$11068 ( \12952 , \12951_nG342e );
not \U$11069 ( \12953 , \12952 );
and \U$11070 ( \12954 , \12932 , \12953 );
buf \U$11071 ( \12955 , RI2b5e785dab30_26);
buf \U$11074 ( \12956 , \12955 );
and \U$11075 ( \12957 , RI2b5e78549630_39, \12645 );
and \U$11076 ( \12958 , RI2b5e78538998_52, \12651 );
and \U$11077 ( \12959 , RI2b5e78538380_65, \12653 );
and \U$11078 ( \12960 , RI2b5e784a5e08_78, \12655 );
and \U$11079 ( \12961 , RI2b5e78495170_91, \12657 );
and \U$11080 ( \12962 , RI2b5e78403c70_104, \12659 );
and \U$11081 ( \12963 , RI2b5e775b1f50_117, \12661 );
and \U$11082 ( \12964 , RI2b5e775b1938_130, \12663 );
and \U$11083 ( \12965 , RI2b5e7750b8d0_143, \12665 );
and \U$11084 ( \12966 , RI2b5e774ff0a8_156, \12667 );
and \U$11085 ( \12967 , RI2b5e774f60c0_169, \12669 );
and \U$11086 ( \12968 , RI2b5e774ea6a8_182, \12671 );
and \U$11087 ( \12969 , RI2b5e774dde80_195, \12673 );
and \U$11088 ( \12970 , RI2b5e774d4e98_208, \12675 );
and \U$11089 ( \12971 , RI2b5e785f3dd8_221, \12677 );
and \U$11090 ( \12972 , RI2b5e785eb1b0_234, \12679 );
and \U$11091 ( \12973 , RI2b5e785da338_247, \12681 );
or \U$11092 ( \12974 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 );
_DC g3412 ( \12975_nG3412 , \12974 , \12700 );
buf \U$11093 ( \12976 , \12975_nG3412 );
not \U$11094 ( \12977 , \12976 );
or \U$11095 ( \12978 , \12956 , \12977 );
and \U$11096 ( \12979 , \12953 , \12978 );
and \U$11097 ( \12980 , \12932 , \12978 );
or \U$11098 ( \12981 , \12954 , \12979 , \12980 );
and \U$11099 ( \12982 , \12928 , \12981 );
and \U$11100 ( \12983 , \12907 , \12981 );
or \U$11101 ( \12984 , \12929 , \12982 , \12983 );
and \U$11102 ( \12985 , \12903 , \12984 );
and \U$11103 ( \12986 , \12882 , \12984 );
or \U$11104 ( \12987 , \12904 , \12985 , \12986 );
and \U$11105 ( \12988 , \12878 , \12987 );
and \U$11106 ( \12989 , \12857 , \12987 );
or \U$11107 ( \12990 , \12879 , \12988 , \12989 );
and \U$11108 ( \12991 , \12853 , \12990 );
and \U$11109 ( \12992 , \12832 , \12990 );
or \U$11110 ( \12993 , \12854 , \12991 , \12992 );
and \U$11111 ( \12994 , \12828 , \12993 );
and \U$11112 ( \12995 , \12807 , \12993 );
or \U$11113 ( \12996 , \12829 , \12994 , \12995 );
and \U$11114 ( \12997 , \12803 , \12996 );
and \U$11115 ( \12998 , \12782 , \12996 );
or \U$11116 ( \12999 , \12804 , \12997 , \12998 );
and \U$11117 ( \13000 , \12778 , \12999 );
and \U$11118 ( \13001 , \12757 , \12999 );
or \U$11119 ( \13002 , \12779 , \13000 , \13001 );
and \U$11120 ( \13003 , \12753 , \13002 );
and \U$11121 ( \13004 , \12732 , \13002 );
or \U$11122 ( \13005 , \12754 , \13003 , \13004 );
and \U$11123 ( \13006 , \12728 , \13005 );
and \U$11124 ( \13007 , \12707 , \13005 );
or \U$11125 ( \13008 , \12729 , \13006 , \13007 );
xor \U$11126 ( \13009 , \12704 , \13008 );
buf g3b29_GF_PartitionCandidate( \13010_nG3b29 , \13009 );
buf \U$11127 ( \13011 , \13010_nG3b29 );
xor \U$11128 ( \13012 , \12707 , \12728 );
xor \U$11129 ( \13013 , \13012 , \13005 );
buf g3b05_GF_PartitionCandidate( \13014_nG3b05 , \13013 );
buf \U$11130 ( \13015 , \13014_nG3b05 );
xor \U$11131 ( \13016 , \12732 , \12753 );
xor \U$11132 ( \13017 , \13016 , \13002 );
buf g3972_GF_PartitionCandidate( \13018_nG3972 , \13017 );
buf \U$11133 ( \13019 , \13018_nG3972 );
and \U$11134 ( \13020 , \13015 , \13019 );
not \U$11135 ( \13021 , \13020 );
and \U$11136 ( \13022 , \13011 , \13021 );
not \U$11137 ( \13023 , \13022 );
buf \U$11138 ( \13024 , \12595 );
buf \U$11139 ( \13025 , \12616 );
buf \U$11140 ( \13026 , \12620 );
buf \U$11141 ( \13027 , \12624 );
buf \U$11142 ( \13028 , \12628 );
buf \U$11143 ( \13029 , \12632 );
buf \U$11144 ( \13030 , \12636 );
buf \U$11145 ( \13031 , \12640 );
buf \U$11146 ( \13032 , \12644 );
buf \U$11147 ( \13033 , \12611 );
nor \U$11148 ( \13034 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 );
buf \U$11149 ( \13035 , \13034 );
buf \U$11150 ( \13036 , \13035 );
xor \U$11151 ( \13037 , \13024 , \13036 );
buf \U$11152 ( \13038 , \13037 );
buf \U$11153 ( \13039 , \12599 );
and \U$11154 ( \13040 , \13024 , \13036 );
xor \U$11155 ( \13041 , \13039 , \13040 );
buf \U$11156 ( \13042 , \13041 );
buf \U$11157 ( \13043 , \12603 );
and \U$11158 ( \13044 , \13039 , \13040 );
xor \U$11159 ( \13045 , \13043 , \13044 );
buf \U$11160 ( \13046 , \13045 );
buf \U$11161 ( \13047 , \12607 );
and \U$11162 ( \13048 , \13043 , \13044 );
xor \U$11163 ( \13049 , \13047 , \13048 );
buf \U$11164 ( \13050 , \13049 );
buf \U$11165 ( \13051 , \12611 );
and \U$11166 ( \13052 , \13047 , \13048 );
xor \U$11167 ( \13053 , \13051 , \13052 );
buf \U$11168 ( \13054 , \13053 );
not \U$11169 ( \13055 , \13054 );
buf \U$11170 ( \13056 , \12616 );
and \U$11171 ( \13057 , \13051 , \13052 );
xor \U$11172 ( \13058 , \13056 , \13057 );
buf \U$11173 ( \13059 , \13058 );
buf \U$11174 ( \13060 , \12620 );
and \U$11175 ( \13061 , \13056 , \13057 );
xor \U$11176 ( \13062 , \13060 , \13061 );
buf \U$11177 ( \13063 , \13062 );
buf \U$11178 ( \13064 , \12624 );
and \U$11179 ( \13065 , \13060 , \13061 );
xor \U$11180 ( \13066 , \13064 , \13065 );
buf \U$11181 ( \13067 , \13066 );
buf \U$11182 ( \13068 , \12628 );
and \U$11183 ( \13069 , \13064 , \13065 );
xor \U$11184 ( \13070 , \13068 , \13069 );
buf \U$11185 ( \13071 , \13070 );
buf \U$11186 ( \13072 , \12632 );
and \U$11187 ( \13073 , \13068 , \13069 );
xor \U$11188 ( \13074 , \13072 , \13073 );
buf \U$11189 ( \13075 , \13074 );
buf \U$11190 ( \13076 , \12636 );
and \U$11191 ( \13077 , \13072 , \13073 );
xor \U$11192 ( \13078 , \13076 , \13077 );
buf \U$11193 ( \13079 , \13078 );
buf \U$11194 ( \13080 , \12640 );
and \U$11195 ( \13081 , \13076 , \13077 );
xor \U$11196 ( \13082 , \13080 , \13081 );
buf \U$11197 ( \13083 , \13082 );
buf \U$11198 ( \13084 , \12644 );
and \U$11199 ( \13085 , \13080 , \13081 );
xor \U$11200 ( \13086 , \13084 , \13085 );
buf \U$11201 ( \13087 , \13086 );
nor \U$11202 ( \13088 , \13038 , \13042 , \13046 , \13050 , \13055 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11203 ( \13089 , RI2b5e785da248_249, \13088 );
not \U$11204 ( \13090 , \13038 );
not \U$11205 ( \13091 , \13042 );
not \U$11206 ( \13092 , \13046 );
not \U$11207 ( \13093 , \13050 );
nor \U$11208 ( \13094 , \13090 , \13091 , \13092 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11209 ( \13095 , RI2b5e785be750_269, \13094 );
nor \U$11210 ( \13096 , \13038 , \13091 , \13092 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11211 ( \13097 , RI2b5e785bc4a0_289, \13096 );
nor \U$11212 ( \13098 , \13090 , \13042 , \13092 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11213 ( \13099 , RI2b5e785bbb40_309, \13098 );
nor \U$11214 ( \13100 , \13038 , \13042 , \13092 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11215 ( \13101 , RI2b5e785b9c50_329, \13100 );
nor \U$11216 ( \13102 , \13090 , \13091 , \13046 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11217 ( \13103 , RI2b5e785b8120_349, \13102 );
nor \U$11218 ( \13104 , \13038 , \13091 , \13046 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11219 ( \13105 , RI2b5e785b77c0_369, \13104 );
nor \U$11220 ( \13106 , \13090 , \13042 , \13046 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11221 ( \13107 , RI2b5e785b6e60_389, \13106 );
nor \U$11222 ( \13108 , \13038 , \13042 , \13046 , \13093 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11223 ( \13109 , RI2b5e785b56f0_409, \13108 );
nor \U$11224 ( \13110 , \13090 , \13091 , \13092 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11225 ( \13111 , RI2b5e785b4d90_429, \13110 );
nor \U$11226 ( \13112 , \13038 , \13091 , \13092 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11227 ( \13113 , RI2b5e785b39e0_449, \13112 );
nor \U$11228 ( \13114 , \13090 , \13042 , \13092 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11229 ( \13115 , RI2b5e785b3080_469, \13114 );
nor \U$11230 ( \13116 , \13038 , \13042 , \13092 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11231 ( \13117 , RI2b5e785b2720_489, \13116 );
nor \U$11232 ( \13118 , \13090 , \13091 , \13046 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11233 ( \13119 , RI2b5e785b1730_509, \13118 );
nor \U$11234 ( \13120 , \13038 , \13091 , \13046 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11235 ( \13121 , RI2b5e785b0dd0_529, \13120 );
nor \U$11236 ( \13122 , \13090 , \13042 , \13046 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11237 ( \13123 , RI2b5e785b0470_549, \13122 );
nor \U$11238 ( \13124 , \13038 , \13042 , \13046 , \13050 , \13054 , \13059 , \13063 , \13067 , \13071 , \13075 , \13079 , \13083 , \13087 );
and \U$11239 ( \13125 , RI2b5e785af840_569, \13124 );
or \U$11240 ( \13126 , \13089 , \13095 , \13097 , \13099 , \13101 , \13103 , \13105 , \13107 , \13109 , \13111 , \13113 , \13115 , \13117 , \13119 , \13121 , \13123 , \13125 );
buf \U$11241 ( \13127 , \13059 );
buf \U$11242 ( \13128 , \13063 );
buf \U$11243 ( \13129 , \13067 );
buf \U$11244 ( \13130 , \13071 );
buf \U$11245 ( \13131 , \13075 );
buf \U$11246 ( \13132 , \13079 );
buf \U$11247 ( \13133 , \13083 );
buf \U$11248 ( \13134 , \13087 );
buf \U$11249 ( \13135 , \13054 );
buf \U$11250 ( \13136 , \13038 );
buf \U$11251 ( \13137 , \13042 );
buf \U$11252 ( \13138 , \13046 );
buf \U$11253 ( \13139 , \13050 );
or \U$11254 ( \13140 , \13136 , \13137 , \13138 , \13139 );
and \U$11255 ( \13141 , \13135 , \13140 );
or \U$11256 ( \13142 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13141 );
buf \U$11257 ( \13143 , \13142 );
_DC g41fa ( \13144_nG41fa , \13126 , \13143 );
buf \U$11258 ( \13145 , \13144_nG41fa );
buf \U$11259 ( \13146 , RI2b5e785db0d0_14);
and \U$11260 ( \13147 , \12553 , \12572 );
and \U$11261 ( \13148 , \13146 , \13147 );
buf \U$11262 ( \13149 , \13148 );
buf \U$11263 ( \13150 , \13149 );
xor \U$11264 ( \13151 , \13146 , \13147 );
buf \U$11265 ( \13152 , \13151 );
buf \U$11266 ( \13153 , \13152 );
and \U$11267 ( \13154 , RI2b5e785daab8_27, \12645 );
and \U$11268 ( \13155 , RI2b5e785495b8_40, \12651 );
and \U$11269 ( \13156 , RI2b5e78538920_53, \12653 );
and \U$11270 ( \13157 , RI2b5e784a63a8_66, \12655 );
and \U$11271 ( \13158 , RI2b5e78495710_79, \12657 );
and \U$11272 ( \13159 , RI2b5e784950f8_92, \12659 );
and \U$11273 ( \13160 , RI2b5e78403bf8_105, \12661 );
and \U$11274 ( \13161 , RI2b5e775b1ed8_118, \12663 );
and \U$11275 ( \13162 , RI2b5e775b18c0_131, \12665 );
and \U$11276 ( \13163 , RI2b5e7750b858_144, \12667 );
and \U$11277 ( \13164 , RI2b5e774ff030_157, \12669 );
and \U$11278 ( \13165 , RI2b5e774f6048_170, \12671 );
and \U$11279 ( \13166 , RI2b5e774ea630_183, \12673 );
and \U$11280 ( \13167 , RI2b5e774dde08_196, \12675 );
and \U$11281 ( \13168 , RI2b5e774d4e20_209, \12677 );
and \U$11282 ( \13169 , RI2b5e785f3d60_222, \12679 );
and \U$11283 ( \13170 , RI2b5e785eb138_235, \12681 );
or \U$11284 ( \13171 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 );
_DC g3cdb ( \13172_nG3cdb , \13171 , \12700 );
buf \U$11285 ( \13173 , \13172_nG3cdb );
not \U$11286 ( \13174 , \13173 );
and \U$11287 ( \13175 , \13153 , \13174 );
and \U$11288 ( \13176 , \12575 , \12703 );
and \U$11289 ( \13177 , \12703 , \13008 );
and \U$11290 ( \13178 , \12575 , \13008 );
or \U$11291 ( \13179 , \13176 , \13177 , \13178 );
and \U$11292 ( \13180 , \13174 , \13179 );
and \U$11293 ( \13181 , \13153 , \13179 );
or \U$11294 ( \13182 , \13175 , \13180 , \13181 );
xnor \U$11295 ( \13183 , \13150 , \13182 );
buf g3cf0_GF_PartitionCandidate( \13184_nG3cf0 , \13183 );
buf \U$11296 ( \13185 , \13184_nG3cf0 );
xor \U$11297 ( \13186 , \13153 , \13174 );
xor \U$11298 ( \13187 , \13186 , \13179 );
buf g3ce4_GF_PartitionCandidate( \13188_nG3ce4 , \13187 );
buf \U$11299 ( \13189 , \13188_nG3ce4 );
xor \U$11300 ( \13190 , \13185 , \13189 );
xor \U$11301 ( \13191 , \13189 , \13011 );
not \U$11302 ( \13192 , \13191 );
and \U$11303 ( \13193 , \13190 , \13192 );
and \U$11304 ( \13194 , \13145 , \13193 );
and \U$11305 ( \13195 , RI2b5e785da2c0_248, \13088 );
and \U$11306 ( \13196 , RI2b5e785be7c8_268, \13094 );
and \U$11307 ( \13197 , RI2b5e785bc518_288, \13096 );
and \U$11308 ( \13198 , RI2b5e785bbbb8_308, \13098 );
and \U$11309 ( \13199 , RI2b5e785b9cc8_328, \13100 );
and \U$11310 ( \13200 , RI2b5e785b9368_348, \13102 );
and \U$11311 ( \13201 , RI2b5e785b7838_368, \13104 );
and \U$11312 ( \13202 , RI2b5e785b6ed8_388, \13106 );
and \U$11313 ( \13203 , RI2b5e785b5768_408, \13108 );
and \U$11314 ( \13204 , RI2b5e785b4e08_428, \13110 );
and \U$11315 ( \13205 , RI2b5e785b3a58_448, \13112 );
and \U$11316 ( \13206 , RI2b5e785b30f8_468, \13114 );
and \U$11317 ( \13207 , RI2b5e785b2798_488, \13116 );
and \U$11318 ( \13208 , RI2b5e785b17a8_508, \13118 );
and \U$11319 ( \13209 , RI2b5e785b0e48_528, \13120 );
and \U$11320 ( \13210 , RI2b5e785b04e8_548, \13122 );
and \U$11321 ( \13211 , RI2b5e785afb88_568, \13124 );
or \U$11322 ( \13212 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 );
_DC g42ef ( \13213_nG42ef , \13212 , \13143 );
buf \U$11323 ( \13214 , \13213_nG42ef );
and \U$11324 ( \13215 , \13214 , \13191 );
nor \U$11325 ( \13216 , \13194 , \13215 );
and \U$11326 ( \13217 , \13189 , \13011 );
not \U$11327 ( \13218 , \13217 );
and \U$11328 ( \13219 , \13185 , \13218 );
xnor \U$11329 ( \13220 , \13216 , \13219 );
xor \U$11330 ( \13221 , \13023 , \13220 );
and \U$11332 ( \13222 , RI2b5e785da1d0_250, \13088 );
and \U$11333 ( \13223 , RI2b5e785be6d8_270, \13094 );
and \U$11334 ( \13224 , RI2b5e785bc428_290, \13096 );
and \U$11335 ( \13225 , RI2b5e785bbac8_310, \13098 );
and \U$11336 ( \13226 , RI2b5e785b9bd8_330, \13100 );
and \U$11337 ( \13227 , RI2b5e785b80a8_350, \13102 );
and \U$11338 ( \13228 , RI2b5e785b7748_370, \13104 );
and \U$11339 ( \13229 , RI2b5e785b6de8_390, \13106 );
and \U$11340 ( \13230 , RI2b5e785b5678_410, \13108 );
and \U$11341 ( \13231 , RI2b5e785b4d18_430, \13110 );
and \U$11342 ( \13232 , RI2b5e785b3968_450, \13112 );
and \U$11343 ( \13233 , RI2b5e785b3008_470, \13114 );
and \U$11344 ( \13234 , RI2b5e785b26a8_490, \13116 );
and \U$11345 ( \13235 , RI2b5e785b16b8_510, \13118 );
and \U$11346 ( \13236 , RI2b5e785b0d58_530, \13120 );
and \U$11347 ( \13237 , RI2b5e785b03f8_550, \13122 );
and \U$11348 ( \13238 , RI2b5e785af7c8_570, \13124 );
or \U$11349 ( \13239 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 );
_DC g4131 ( \13240_nG4131 , \13239 , \13143 );
buf \U$11350 ( \13241 , \13240_nG4131 );
or \U$11351 ( \13242 , \13150 , \13182 );
not \U$11352 ( \13243 , \13242 );
buf g3eca_GF_PartitionCandidate( \13244_nG3eca , \13243 );
buf \U$11353 ( \13245 , \13244_nG3eca );
xor \U$11354 ( \13246 , \13245 , \13185 );
and \U$11355 ( \13247 , \13241 , \13246 );
nor \U$11356 ( \13248 , 1'b0 , \13247 );
xnor \U$11358 ( \13249 , \13248 , 1'b0 );
xor \U$11359 ( \13250 , \13221 , \13249 );
xor \U$11360 ( \13251 , 1'b0 , \13250 );
xor \U$11362 ( \13252 , \13011 , \13015 );
xor \U$11363 ( \13253 , \13015 , \13019 );
not \U$11364 ( \13254 , \13253 );
and \U$11365 ( \13255 , \13252 , \13254 );
and \U$11366 ( \13256 , \13214 , \13255 );
not \U$11367 ( \13257 , \13256 );
xnor \U$11368 ( \13258 , \13257 , \13022 );
and \U$11369 ( \13259 , \13241 , \13193 );
and \U$11370 ( \13260 , \13145 , \13191 );
nor \U$11371 ( \13261 , \13259 , \13260 );
xnor \U$11372 ( \13262 , \13261 , \13219 );
and \U$11373 ( \13263 , \13258 , \13262 );
or \U$11375 ( \13264 , 1'b0 , \13263 , 1'b0 );
xor \U$11377 ( \13265 , \13264 , 1'b0 );
xor \U$11379 ( \13266 , \13265 , 1'b0 );
and \U$11380 ( \13267 , \13251 , \13266 );
or \U$11381 ( \13268 , 1'b0 , 1'b0 , \13267 );
and \U$11384 ( \13269 , \13214 , \13193 );
not \U$11385 ( \13270 , \13269 );
xnor \U$11386 ( \13271 , \13270 , \13219 );
xor \U$11387 ( \13272 , 1'b0 , \13271 );
and \U$11389 ( \13273 , \13145 , \13246 );
nor \U$11390 ( \13274 , 1'b0 , \13273 );
xnor \U$11391 ( \13275 , \13274 , 1'b0 );
xor \U$11392 ( \13276 , \13272 , \13275 );
xor \U$11393 ( \13277 , 1'b0 , \13276 );
xor \U$11395 ( \13278 , \13277 , 1'b1 );
and \U$11396 ( \13279 , \13023 , \13220 );
and \U$11397 ( \13280 , \13220 , \13249 );
and \U$11398 ( \13281 , \13023 , \13249 );
or \U$11399 ( \13282 , \13279 , \13280 , \13281 );
xor \U$11401 ( \13283 , \13282 , 1'b0 );
xor \U$11403 ( \13284 , \13283 , 1'b0 );
xor \U$11404 ( \13285 , \13278 , \13284 );
and \U$11405 ( \13286 , \13268 , \13285 );
or \U$11407 ( \13287 , 1'b0 , \13286 , 1'b0 );
xor \U$11409 ( \13288 , \13287 , 1'b0 );
and \U$11411 ( \13289 , \13277 , 1'b1 );
and \U$11412 ( \13290 , 1'b1 , \13284 );
and \U$11413 ( \13291 , \13277 , \13284 );
or \U$11414 ( \13292 , \13289 , \13290 , \13291 );
xor \U$11415 ( \13293 , 1'b0 , \13292 );
not \U$11417 ( \13294 , \13219 );
and \U$11419 ( \13295 , \13214 , \13246 );
nor \U$11420 ( \13296 , 1'b0 , \13295 );
xnor \U$11421 ( \13297 , \13296 , 1'b0 );
xor \U$11422 ( \13298 , \13294 , \13297 );
xor \U$11424 ( \13299 , \13298 , 1'b0 );
xor \U$11425 ( \13300 , 1'b0 , \13299 );
xor \U$11427 ( \13301 , \13300 , 1'b0 );
and \U$11429 ( \13302 , \13271 , \13275 );
or \U$11431 ( \13303 , 1'b0 , \13302 , 1'b0 );
xor \U$11433 ( \13304 , \13303 , 1'b0 );
xor \U$11435 ( \13305 , \13304 , 1'b0 );
xor \U$11436 ( \13306 , \13301 , \13305 );
xor \U$11437 ( \13307 , \13293 , \13306 );
xor \U$11438 ( \13308 , \13288 , \13307 );
xor \U$11444 ( \13309 , \12757 , \12778 );
xor \U$11445 ( \13310 , \13309 , \12999 );
buf g394e_GF_PartitionCandidate( \13311_nG394e , \13310 );
buf \U$11446 ( \13312 , \13311_nG394e );
xor \U$11447 ( \13313 , \13019 , \13312 );
xor \U$11448 ( \13314 , \12782 , \12803 );
xor \U$11449 ( \13315 , \13314 , \12996 );
buf g37cf_GF_PartitionCandidate( \13316_nG37cf , \13315 );
buf \U$11450 ( \13317 , \13316_nG37cf );
xor \U$11451 ( \13318 , \13312 , \13317 );
not \U$11452 ( \13319 , \13318 );
and \U$11453 ( \13320 , \13313 , \13319 );
and \U$11454 ( \13321 , \13214 , \13320 );
not \U$11455 ( \13322 , \13321 );
and \U$11456 ( \13323 , \13312 , \13317 );
not \U$11457 ( \13324 , \13323 );
and \U$11458 ( \13325 , \13019 , \13324 );
xnor \U$11459 ( \13326 , \13322 , \13325 );
and \U$11460 ( \13327 , \13241 , \13255 );
and \U$11461 ( \13328 , \13145 , \13253 );
nor \U$11462 ( \13329 , \13327 , \13328 );
xnor \U$11463 ( \13330 , \13329 , \13022 );
and \U$11464 ( \13331 , \13326 , \13330 );
or \U$11466 ( \13332 , 1'b0 , \13331 , 1'b0 );
and \U$11467 ( \13333 , RI2b5e785da0e0_252, \13088 );
and \U$11468 ( \13334 , RI2b5e785be5e8_272, \13094 );
and \U$11469 ( \13335 , RI2b5e785bc338_292, \13096 );
and \U$11470 ( \13336 , RI2b5e785bb9d8_312, \13098 );
and \U$11471 ( \13337 , RI2b5e785b9ae8_332, \13100 );
and \U$11472 ( \13338 , RI2b5e785b7fb8_352, \13102 );
and \U$11473 ( \13339 , RI2b5e785b7658_372, \13104 );
and \U$11474 ( \13340 , RI2b5e785b5ee8_392, \13106 );
and \U$11475 ( \13341 , RI2b5e785b5588_412, \13108 );
and \U$11476 ( \13342 , RI2b5e785b4c28_432, \13110 );
and \U$11477 ( \13343 , RI2b5e785b3878_452, \13112 );
and \U$11478 ( \13344 , RI2b5e785b2f18_472, \13114 );
and \U$11479 ( \13345 , RI2b5e785b25b8_492, \13116 );
and \U$11480 ( \13346 , RI2b5e785b15c8_512, \13118 );
and \U$11481 ( \13347 , RI2b5e785b0c68_532, \13120 );
and \U$11482 ( \13348 , RI2b5e785b0308_552, \13122 );
and \U$11483 ( \13349 , RI2b5e785af6d8_572, \13124 );
or \U$11484 ( \13350 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 );
_DC g3f92 ( \13351_nG3f92 , \13350 , \13143 );
buf \U$11485 ( \13352 , \13351_nG3f92 );
and \U$11486 ( \13353 , \13352 , \13193 );
and \U$11487 ( \13354 , RI2b5e785da158_251, \13088 );
and \U$11488 ( \13355 , RI2b5e785be660_271, \13094 );
and \U$11489 ( \13356 , RI2b5e785bc3b0_291, \13096 );
and \U$11490 ( \13357 , RI2b5e785bba50_311, \13098 );
and \U$11491 ( \13358 , RI2b5e785b9b60_331, \13100 );
and \U$11492 ( \13359 , RI2b5e785b8030_351, \13102 );
and \U$11493 ( \13360 , RI2b5e785b76d0_371, \13104 );
and \U$11494 ( \13361 , RI2b5e785b6d70_391, \13106 );
and \U$11495 ( \13362 , RI2b5e785b5600_411, \13108 );
and \U$11496 ( \13363 , RI2b5e785b4ca0_431, \13110 );
and \U$11497 ( \13364 , RI2b5e785b38f0_451, \13112 );
and \U$11498 ( \13365 , RI2b5e785b2f90_471, \13114 );
and \U$11499 ( \13366 , RI2b5e785b2630_491, \13116 );
and \U$11500 ( \13367 , RI2b5e785b1640_511, \13118 );
and \U$11501 ( \13368 , RI2b5e785b0ce0_531, \13120 );
and \U$11502 ( \13369 , RI2b5e785b0380_551, \13122 );
and \U$11503 ( \13370 , RI2b5e785af750_571, \13124 );
or \U$11504 ( \13371 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 );
_DC g4070 ( \13372_nG4070 , \13371 , \13143 );
buf \U$11505 ( \13373 , \13372_nG4070 );
and \U$11506 ( \13374 , \13373 , \13191 );
nor \U$11507 ( \13375 , \13353 , \13374 );
xnor \U$11508 ( \13376 , \13375 , \13219 );
and \U$11510 ( \13377 , RI2b5e785da068_253, \13088 );
and \U$11511 ( \13378 , RI2b5e785be570_273, \13094 );
and \U$11512 ( \13379 , RI2b5e785bc2c0_293, \13096 );
and \U$11513 ( \13380 , RI2b5e785bb960_313, \13098 );
and \U$11514 ( \13381 , RI2b5e785b9a70_333, \13100 );
and \U$11515 ( \13382 , RI2b5e785b7f40_353, \13102 );
and \U$11516 ( \13383 , RI2b5e785b75e0_373, \13104 );
and \U$11517 ( \13384 , RI2b5e785b5e70_393, \13106 );
and \U$11518 ( \13385 , RI2b5e785b5510_413, \13108 );
and \U$11519 ( \13386 , RI2b5e785b4bb0_433, \13110 );
and \U$11520 ( \13387 , RI2b5e785b3800_453, \13112 );
and \U$11521 ( \13388 , RI2b5e785b2ea0_473, \13114 );
and \U$11522 ( \13389 , RI2b5e785b2540_493, \13116 );
and \U$11523 ( \13390 , RI2b5e785b1550_513, \13118 );
and \U$11524 ( \13391 , RI2b5e785b0bf0_533, \13120 );
and \U$11525 ( \13392 , RI2b5e785b0290_553, \13122 );
and \U$11526 ( \13393 , RI2b5e785af660_573, \13124 );
or \U$11527 ( \13394 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 );
_DC g3ea9 ( \13395_nG3ea9 , \13394 , \13143 );
buf \U$11528 ( \13396 , \13395_nG3ea9 );
and \U$11529 ( \13397 , \13396 , \13246 );
nor \U$11530 ( \13398 , 1'b0 , \13397 );
xnor \U$11531 ( \13399 , \13398 , 1'b0 );
and \U$11532 ( \13400 , \13376 , \13399 );
or \U$11535 ( \13401 , \13400 , 1'b0 , 1'b0 );
and \U$11536 ( \13402 , \13332 , \13401 );
or \U$11539 ( \13403 , \13402 , 1'b0 , 1'b0 );
and \U$11542 ( \13404 , \13352 , \13246 );
nor \U$11543 ( \13405 , 1'b0 , \13404 );
xnor \U$11544 ( \13406 , \13405 , 1'b0 );
xor \U$11546 ( \13407 , \13406 , 1'b0 );
xor \U$11548 ( \13408 , \13407 , 1'b0 );
not \U$11549 ( \13409 , \13325 );
and \U$11550 ( \13410 , \13145 , \13255 );
and \U$11551 ( \13411 , \13214 , \13253 );
nor \U$11552 ( \13412 , \13410 , \13411 );
xnor \U$11553 ( \13413 , \13412 , \13022 );
xor \U$11554 ( \13414 , \13409 , \13413 );
and \U$11555 ( \13415 , \13373 , \13193 );
and \U$11556 ( \13416 , \13241 , \13191 );
nor \U$11557 ( \13417 , \13415 , \13416 );
xnor \U$11558 ( \13418 , \13417 , \13219 );
xor \U$11559 ( \13419 , \13414 , \13418 );
and \U$11560 ( \13420 , \13408 , \13419 );
or \U$11562 ( \13421 , 1'b0 , \13420 , 1'b0 );
and \U$11563 ( \13422 , \13403 , \13421 );
or \U$11564 ( \13423 , 1'b0 , 1'b0 , \13422 );
and \U$11566 ( \13424 , \13373 , \13246 );
nor \U$11567 ( \13425 , 1'b0 , \13424 );
xnor \U$11568 ( \13426 , \13425 , 1'b0 );
xor \U$11570 ( \13427 , \13426 , 1'b0 );
xor \U$11572 ( \13428 , \13427 , 1'b0 );
xor \U$11574 ( \13429 , 1'b0 , \13258 );
xor \U$11575 ( \13430 , \13429 , \13262 );
xor \U$11576 ( \13431 , \13428 , \13430 );
and \U$11578 ( \13432 , \13431 , 1'b1 );
and \U$11579 ( \13433 , \13409 , \13413 );
and \U$11580 ( \13434 , \13413 , \13418 );
and \U$11581 ( \13435 , \13409 , \13418 );
or \U$11582 ( \13436 , \13433 , \13434 , \13435 );
xor \U$11584 ( \13437 , \13436 , 1'b0 );
xor \U$11586 ( \13438 , \13437 , 1'b0 );
and \U$11587 ( \13439 , 1'b1 , \13438 );
and \U$11588 ( \13440 , \13431 , \13438 );
or \U$11589 ( \13441 , \13432 , \13439 , \13440 );
and \U$11590 ( \13442 , \13423 , \13441 );
xor \U$11592 ( \13443 , \13251 , 1'b0 );
xor \U$11593 ( \13444 , \13443 , \13266 );
and \U$11594 ( \13445 , \13441 , \13444 );
and \U$11595 ( \13446 , \13423 , \13444 );
or \U$11596 ( \13447 , \13442 , \13445 , \13446 );
xor \U$11598 ( \13448 , 1'b0 , \13268 );
xor \U$11599 ( \13449 , \13448 , \13285 );
and \U$11600 ( \13450 , \13447 , \13449 );
or \U$11601 ( \13451 , 1'b0 , 1'b0 , \13450 );
nand \U$11602 ( \13452 , \13308 , \13451 );
nor \U$11603 ( \13453 , \13308 , \13451 );
not \U$11604 ( \13454 , \13453 );
nand \U$11605 ( \13455 , \13452 , \13454 );
xor \U$11606 ( \13456 , \12932 , \12953 );
xor \U$11607 ( \13457 , \13456 , \12978 );
buf g3435_GF_PartitionCandidate( \13458_nG3435 , \13457 );
buf \U$11608 ( \13459 , \13458_nG3435 );
xor \U$11609 ( \13460 , \12956 , \12976 );
buf g3415_GF_PartitionCandidate( \13461_nG3415 , \13460 );
buf \U$11610 ( \13462 , \13461_nG3415 );
xor \U$11611 ( \13463 , \13459 , \13462 );
not \U$11612 ( \13464 , \13462 );
and \U$11613 ( \13465 , \13463 , \13464 );
and \U$11614 ( \13466 , \13396 , \13465 );
and \U$11615 ( \13467 , \13352 , \13462 );
nor \U$11616 ( \13468 , \13466 , \13467 );
xnor \U$11617 ( \13469 , \13468 , \13459 );
and \U$11618 ( \13470 , RI2b5e785c2bc0_255, \13088 );
and \U$11619 ( \13471 , RI2b5e785be480_275, \13094 );
and \U$11620 ( \13472 , RI2b5e785bc1d0_295, \13096 );
and \U$11621 ( \13473 , RI2b5e785ba2e0_315, \13098 );
and \U$11622 ( \13474 , RI2b5e785b9980_335, \13100 );
and \U$11623 ( \13475 , RI2b5e785b7e50_355, \13102 );
and \U$11624 ( \13476 , RI2b5e785b74f0_375, \13104 );
and \U$11625 ( \13477 , RI2b5e785b5d80_395, \13106 );
and \U$11626 ( \13478 , RI2b5e785b5420_415, \13108 );
and \U$11627 ( \13479 , RI2b5e785b4ac0_435, \13110 );
and \U$11628 ( \13480 , RI2b5e785b3710_455, \13112 );
and \U$11629 ( \13481 , RI2b5e785b2db0_475, \13114 );
and \U$11630 ( \13482 , RI2b5e785b2450_495, \13116 );
and \U$11631 ( \13483 , RI2b5e785b1460_515, \13118 );
and \U$11632 ( \13484 , RI2b5e785b0b00_535, \13120 );
and \U$11633 ( \13485 , RI2b5e785b01a0_555, \13122 );
and \U$11634 ( \13486 , RI2b5e785af570_575, \13124 );
or \U$11635 ( \13487 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 );
_DC g3d18 ( \13488_nG3d18 , \13487 , \13143 );
buf \U$11636 ( \13489 , \13488_nG3d18 );
xor \U$11637 ( \13490 , \12882 , \12903 );
xor \U$11638 ( \13491 , \13490 , \12984 );
buf g353d_GF_PartitionCandidate( \13492_nG353d , \13491 );
buf \U$11639 ( \13493 , \13492_nG353d );
xor \U$11640 ( \13494 , \12907 , \12928 );
xor \U$11641 ( \13495 , \13494 , \12981 );
buf g3541_GF_PartitionCandidate( \13496_nG3541 , \13495 );
buf \U$11642 ( \13497 , \13496_nG3541 );
xor \U$11643 ( \13498 , \13493 , \13497 );
xor \U$11644 ( \13499 , \13497 , \13459 );
not \U$11645 ( \13500 , \13499 );
and \U$11646 ( \13501 , \13498 , \13500 );
and \U$11647 ( \13502 , \13489 , \13501 );
and \U$11648 ( \13503 , RI2b5e785c2c38_254, \13088 );
and \U$11649 ( \13504 , RI2b5e785be4f8_274, \13094 );
and \U$11650 ( \13505 , RI2b5e785bc248_294, \13096 );
and \U$11651 ( \13506 , RI2b5e785ba358_314, \13098 );
and \U$11652 ( \13507 , RI2b5e785b99f8_334, \13100 );
and \U$11653 ( \13508 , RI2b5e785b7ec8_354, \13102 );
and \U$11654 ( \13509 , RI2b5e785b7568_374, \13104 );
and \U$11655 ( \13510 , RI2b5e785b5df8_394, \13106 );
and \U$11656 ( \13511 , RI2b5e785b5498_414, \13108 );
and \U$11657 ( \13512 , RI2b5e785b4b38_434, \13110 );
and \U$11658 ( \13513 , RI2b5e785b3788_454, \13112 );
and \U$11659 ( \13514 , RI2b5e785b2e28_474, \13114 );
and \U$11660 ( \13515 , RI2b5e785b24c8_494, \13116 );
and \U$11661 ( \13516 , RI2b5e785b14d8_514, \13118 );
and \U$11662 ( \13517 , RI2b5e785b0b78_534, \13120 );
and \U$11663 ( \13518 , RI2b5e785b0218_554, \13122 );
and \U$11664 ( \13519 , RI2b5e785af5e8_574, \13124 );
or \U$11665 ( \13520 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 );
_DC g3dc5 ( \13521_nG3dc5 , \13520 , \13143 );
buf \U$11666 ( \13522 , \13521_nG3dc5 );
and \U$11667 ( \13523 , \13522 , \13499 );
nor \U$11668 ( \13524 , \13502 , \13523 );
and \U$11669 ( \13525 , \13497 , \13459 );
not \U$11670 ( \13526 , \13525 );
and \U$11671 ( \13527 , \13493 , \13526 );
xnor \U$11672 ( \13528 , \13524 , \13527 );
and \U$11673 ( \13529 , \13469 , \13528 );
and \U$11674 ( \13530 , RI2b5e785c0a00_257, \13088 );
and \U$11675 ( \13531 , RI2b5e785be390_277, \13094 );
and \U$11676 ( \13532 , RI2b5e785bc0e0_297, \13096 );
and \U$11677 ( \13533 , RI2b5e785ba1f0_317, \13098 );
and \U$11678 ( \13534 , RI2b5e785b9890_337, \13100 );
and \U$11679 ( \13535 , RI2b5e785b7d60_357, \13102 );
and \U$11680 ( \13536 , RI2b5e785b7400_377, \13104 );
and \U$11681 ( \13537 , RI2b5e785b5c90_397, \13106 );
and \U$11682 ( \13538 , RI2b5e785b5330_417, \13108 );
and \U$11683 ( \13539 , RI2b5e785b49d0_437, \13110 );
and \U$11684 ( \13540 , RI2b5e785b3620_457, \13112 );
and \U$11685 ( \13541 , RI2b5e785b2cc0_477, \13114 );
and \U$11686 ( \13542 , RI2b5e785b2360_497, \13116 );
and \U$11687 ( \13543 , RI2b5e785b1370_517, \13118 );
and \U$11688 ( \13544 , RI2b5e785b0a10_537, \13120 );
and \U$11689 ( \13545 , RI2b5e785b00b0_557, \13122 );
and \U$11690 ( \13546 , RI2b5e785af480_577, \13124 );
or \U$11691 ( \13547 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 );
_DC g3b58 ( \13548_nG3b58 , \13547 , \13143 );
buf \U$11692 ( \13549 , \13548_nG3b58 );
xor \U$11693 ( \13550 , \12832 , \12853 );
xor \U$11694 ( \13551 , \13550 , \12990 );
buf g3660_GF_PartitionCandidate( \13552_nG3660 , \13551 );
buf \U$11695 ( \13553 , \13552_nG3660 );
xor \U$11696 ( \13554 , \12857 , \12878 );
xor \U$11697 ( \13555 , \13554 , \12987 );
buf g363c_GF_PartitionCandidate( \13556_nG363c , \13555 );
buf \U$11698 ( \13557 , \13556_nG363c );
xor \U$11699 ( \13558 , \13553 , \13557 );
xor \U$11700 ( \13559 , \13557 , \13493 );
not \U$11701 ( \13560 , \13559 );
and \U$11702 ( \13561 , \13558 , \13560 );
and \U$11703 ( \13562 , \13549 , \13561 );
and \U$11704 ( \13563 , RI2b5e785c2b48_256, \13088 );
and \U$11705 ( \13564 , RI2b5e785be408_276, \13094 );
and \U$11706 ( \13565 , RI2b5e785bc158_296, \13096 );
and \U$11707 ( \13566 , RI2b5e785ba268_316, \13098 );
and \U$11708 ( \13567 , RI2b5e785b9908_336, \13100 );
and \U$11709 ( \13568 , RI2b5e785b7dd8_356, \13102 );
and \U$11710 ( \13569 , RI2b5e785b7478_376, \13104 );
and \U$11711 ( \13570 , RI2b5e785b5d08_396, \13106 );
and \U$11712 ( \13571 , RI2b5e785b53a8_416, \13108 );
and \U$11713 ( \13572 , RI2b5e785b4a48_436, \13110 );
and \U$11714 ( \13573 , RI2b5e785b3698_456, \13112 );
and \U$11715 ( \13574 , RI2b5e785b2d38_476, \13114 );
and \U$11716 ( \13575 , RI2b5e785b23d8_496, \13116 );
and \U$11717 ( \13576 , RI2b5e785b13e8_516, \13118 );
and \U$11718 ( \13577 , RI2b5e785b0a88_536, \13120 );
and \U$11719 ( \13578 , RI2b5e785b0128_556, \13122 );
and \U$11720 ( \13579 , RI2b5e785af4f8_576, \13124 );
or \U$11721 ( \13580 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 );
_DC g3bf0 ( \13581_nG3bf0 , \13580 , \13143 );
buf \U$11722 ( \13582 , \13581_nG3bf0 );
and \U$11723 ( \13583 , \13582 , \13559 );
nor \U$11724 ( \13584 , \13562 , \13583 );
and \U$11725 ( \13585 , \13557 , \13493 );
not \U$11726 ( \13586 , \13585 );
and \U$11727 ( \13587 , \13553 , \13586 );
xnor \U$11728 ( \13588 , \13584 , \13587 );
and \U$11729 ( \13589 , \13528 , \13588 );
and \U$11730 ( \13590 , \13469 , \13588 );
or \U$11731 ( \13591 , \13529 , \13589 , \13590 );
and \U$11732 ( \13592 , RI2b5e785c0910_259, \13088 );
and \U$11733 ( \13593 , RI2b5e785be2a0_279, \13094 );
and \U$11734 ( \13594 , RI2b5e785bbff0_299, \13096 );
and \U$11735 ( \13595 , RI2b5e785ba100_319, \13098 );
and \U$11736 ( \13596 , RI2b5e785b97a0_339, \13100 );
and \U$11737 ( \13597 , RI2b5e785b7c70_359, \13102 );
and \U$11738 ( \13598 , RI2b5e785b7310_379, \13104 );
and \U$11739 ( \13599 , RI2b5e785b5ba0_399, \13106 );
and \U$11740 ( \13600 , RI2b5e785b5240_419, \13108 );
and \U$11741 ( \13601 , RI2b5e785b48e0_439, \13110 );
and \U$11742 ( \13602 , RI2b5e785b3530_459, \13112 );
and \U$11743 ( \13603 , RI2b5e785b2bd0_479, \13114 );
and \U$11744 ( \13604 , RI2b5e785b2270_499, \13116 );
and \U$11745 ( \13605 , RI2b5e785b1280_519, \13118 );
and \U$11746 ( \13606 , RI2b5e785b0920_539, \13120 );
and \U$11747 ( \13607 , RI2b5e785affc0_559, \13122 );
and \U$11748 ( \13608 , RI2b5e785af390_579, \13124 );
or \U$11749 ( \13609 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 );
_DC g398d ( \13610_nG398d , \13609 , \13143 );
buf \U$11750 ( \13611 , \13610_nG398d );
xor \U$11751 ( \13612 , \12807 , \12828 );
xor \U$11752 ( \13613 , \13612 , \12993 );
buf g37ab_GF_PartitionCandidate( \13614_nG37ab , \13613 );
buf \U$11753 ( \13615 , \13614_nG37ab );
xor \U$11754 ( \13616 , \13317 , \13615 );
xor \U$11755 ( \13617 , \13615 , \13553 );
not \U$11756 ( \13618 , \13617 );
and \U$11757 ( \13619 , \13616 , \13618 );
and \U$11758 ( \13620 , \13611 , \13619 );
and \U$11759 ( \13621 , RI2b5e785c0988_258, \13088 );
and \U$11760 ( \13622 , RI2b5e785be318_278, \13094 );
and \U$11761 ( \13623 , RI2b5e785bc068_298, \13096 );
and \U$11762 ( \13624 , RI2b5e785ba178_318, \13098 );
and \U$11763 ( \13625 , RI2b5e785b9818_338, \13100 );
and \U$11764 ( \13626 , RI2b5e785b7ce8_358, \13102 );
and \U$11765 ( \13627 , RI2b5e785b7388_378, \13104 );
and \U$11766 ( \13628 , RI2b5e785b5c18_398, \13106 );
and \U$11767 ( \13629 , RI2b5e785b52b8_418, \13108 );
and \U$11768 ( \13630 , RI2b5e785b4958_438, \13110 );
and \U$11769 ( \13631 , RI2b5e785b35a8_458, \13112 );
and \U$11770 ( \13632 , RI2b5e785b2c48_478, \13114 );
and \U$11771 ( \13633 , RI2b5e785b22e8_498, \13116 );
and \U$11772 ( \13634 , RI2b5e785b12f8_518, \13118 );
and \U$11773 ( \13635 , RI2b5e785b0998_538, \13120 );
and \U$11774 ( \13636 , RI2b5e785b0038_558, \13122 );
and \U$11775 ( \13637 , RI2b5e785af408_578, \13124 );
or \U$11776 ( \13638 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 );
_DC g3a17 ( \13639_nG3a17 , \13638 , \13143 );
buf \U$11777 ( \13640 , \13639_nG3a17 );
and \U$11778 ( \13641 , \13640 , \13617 );
nor \U$11779 ( \13642 , \13620 , \13641 );
and \U$11780 ( \13643 , \13615 , \13553 );
not \U$11781 ( \13644 , \13643 );
and \U$11782 ( \13645 , \13317 , \13644 );
xnor \U$11783 ( \13646 , \13642 , \13645 );
and \U$11784 ( \13647 , RI2b5e785c0820_261, \13088 );
and \U$11785 ( \13648 , RI2b5e785be1b0_281, \13094 );
and \U$11786 ( \13649 , RI2b5e785bbf00_301, \13096 );
and \U$11787 ( \13650 , RI2b5e785ba010_321, \13098 );
and \U$11788 ( \13651 , RI2b5e785b96b0_341, \13100 );
and \U$11789 ( \13652 , RI2b5e785b7b80_361, \13102 );
and \U$11790 ( \13653 , RI2b5e785b7220_381, \13104 );
and \U$11791 ( \13654 , RI2b5e785b5ab0_401, \13106 );
and \U$11792 ( \13655 , RI2b5e785b5150_421, \13108 );
and \U$11793 ( \13656 , RI2b5e785b47f0_441, \13110 );
and \U$11794 ( \13657 , RI2b5e785b3440_461, \13112 );
and \U$11795 ( \13658 , RI2b5e785b2ae0_481, \13114 );
and \U$11796 ( \13659 , RI2b5e785b2180_501, \13116 );
and \U$11797 ( \13660 , RI2b5e785b1190_521, \13118 );
and \U$11798 ( \13661 , RI2b5e785b0830_541, \13120 );
and \U$11799 ( \13662 , RI2b5e785afed0_561, \13122 );
and \U$11800 ( \13663 , RI2b5e785af2a0_581, \13124 );
or \U$11801 ( \13664 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 );
_DC g37ea ( \13665_nG37ea , \13664 , \13143 );
buf \U$11802 ( \13666 , \13665_nG37ea );
and \U$11803 ( \13667 , \13666 , \13320 );
and \U$11804 ( \13668 , RI2b5e785c0898_260, \13088 );
and \U$11805 ( \13669 , RI2b5e785be228_280, \13094 );
and \U$11806 ( \13670 , RI2b5e785bbf78_300, \13096 );
and \U$11807 ( \13671 , RI2b5e785ba088_320, \13098 );
and \U$11808 ( \13672 , RI2b5e785b9728_340, \13100 );
and \U$11809 ( \13673 , RI2b5e785b7bf8_360, \13102 );
and \U$11810 ( \13674 , RI2b5e785b7298_380, \13104 );
and \U$11811 ( \13675 , RI2b5e785b5b28_400, \13106 );
and \U$11812 ( \13676 , RI2b5e785b51c8_420, \13108 );
and \U$11813 ( \13677 , RI2b5e785b4868_440, \13110 );
and \U$11814 ( \13678 , RI2b5e785b34b8_460, \13112 );
and \U$11815 ( \13679 , RI2b5e785b2b58_480, \13114 );
and \U$11816 ( \13680 , RI2b5e785b21f8_500, \13116 );
and \U$11817 ( \13681 , RI2b5e785b1208_520, \13118 );
and \U$11818 ( \13682 , RI2b5e785b08a8_540, \13120 );
and \U$11819 ( \13683 , RI2b5e785aff48_560, \13122 );
and \U$11820 ( \13684 , RI2b5e785af318_580, \13124 );
or \U$11821 ( \13685 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 );
_DC g385e ( \13686_nG385e , \13685 , \13143 );
buf \U$11822 ( \13687 , \13686_nG385e );
and \U$11823 ( \13688 , \13687 , \13318 );
nor \U$11824 ( \13689 , \13667 , \13688 );
xnor \U$11825 ( \13690 , \13689 , \13325 );
and \U$11826 ( \13691 , \13646 , \13690 );
and \U$11827 ( \13692 , RI2b5e785c0730_263, \13088 );
and \U$11828 ( \13693 , RI2b5e785be0c0_283, \13094 );
and \U$11829 ( \13694 , RI2b5e785bbe10_303, \13096 );
and \U$11830 ( \13695 , RI2b5e785b9f20_323, \13098 );
and \U$11831 ( \13696 , RI2b5e785b95c0_343, \13100 );
and \U$11832 ( \13697 , RI2b5e785b7a90_363, \13102 );
and \U$11833 ( \13698 , RI2b5e785b7130_383, \13104 );
and \U$11834 ( \13699 , RI2b5e785b59c0_403, \13106 );
and \U$11835 ( \13700 , RI2b5e785b5060_423, \13108 );
and \U$11836 ( \13701 , RI2b5e785b3cb0_443, \13110 );
and \U$11837 ( \13702 , RI2b5e785b3350_463, \13112 );
and \U$11838 ( \13703 , RI2b5e785b29f0_483, \13114 );
and \U$11839 ( \13704 , RI2b5e785b1a00_503, \13116 );
and \U$11840 ( \13705 , RI2b5e785b10a0_523, \13118 );
and \U$11841 ( \13706 , RI2b5e785b0740_543, \13120 );
and \U$11842 ( \13707 , RI2b5e785afde0_563, \13122 );
and \U$11843 ( \13708 , RI2b5e785af1b0_583, \13124 );
or \U$11844 ( \13709 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 );
_DC g3679 ( \13710_nG3679 , \13709 , \13143 );
buf \U$11845 ( \13711 , \13710_nG3679 );
and \U$11846 ( \13712 , \13711 , \13255 );
and \U$11847 ( \13713 , RI2b5e785c07a8_262, \13088 );
and \U$11848 ( \13714 , RI2b5e785be138_282, \13094 );
and \U$11849 ( \13715 , RI2b5e785bbe88_302, \13096 );
and \U$11850 ( \13716 , RI2b5e785b9f98_322, \13098 );
and \U$11851 ( \13717 , RI2b5e785b9638_342, \13100 );
and \U$11852 ( \13718 , RI2b5e785b7b08_362, \13102 );
and \U$11853 ( \13719 , RI2b5e785b71a8_382, \13104 );
and \U$11854 ( \13720 , RI2b5e785b5a38_402, \13106 );
and \U$11855 ( \13721 , RI2b5e785b50d8_422, \13108 );
and \U$11856 ( \13722 , RI2b5e785b4778_442, \13110 );
and \U$11857 ( \13723 , RI2b5e785b33c8_462, \13112 );
and \U$11858 ( \13724 , RI2b5e785b2a68_482, \13114 );
and \U$11859 ( \13725 , RI2b5e785b1a78_502, \13116 );
and \U$11860 ( \13726 , RI2b5e785b1118_522, \13118 );
and \U$11861 ( \13727 , RI2b5e785b07b8_542, \13120 );
and \U$11862 ( \13728 , RI2b5e785afe58_562, \13122 );
and \U$11863 ( \13729 , RI2b5e785af228_582, \13124 );
or \U$11864 ( \13730 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 );
_DC g36e0 ( \13731_nG36e0 , \13730 , \13143 );
buf \U$11865 ( \13732 , \13731_nG36e0 );
and \U$11866 ( \13733 , \13732 , \13253 );
nor \U$11867 ( \13734 , \13712 , \13733 );
xnor \U$11868 ( \13735 , \13734 , \13022 );
and \U$11869 ( \13736 , \13690 , \13735 );
and \U$11870 ( \13737 , \13646 , \13735 );
or \U$11871 ( \13738 , \13691 , \13736 , \13737 );
and \U$11872 ( \13739 , \13591 , \13738 );
and \U$11873 ( \13740 , RI2b5e785c0640_265, \13088 );
and \U$11874 ( \13741 , RI2b5e785bdfd0_285, \13094 );
and \U$11875 ( \13742 , RI2b5e785bbd20_305, \13096 );
and \U$11876 ( \13743 , RI2b5e785b9e30_325, \13098 );
and \U$11877 ( \13744 , RI2b5e785b94d0_345, \13100 );
and \U$11878 ( \13745 , RI2b5e785b79a0_365, \13102 );
and \U$11879 ( \13746 , RI2b5e785b7040_385, \13104 );
and \U$11880 ( \13747 , RI2b5e785b58d0_405, \13106 );
and \U$11881 ( \13748 , RI2b5e785b4f70_425, \13108 );
and \U$11882 ( \13749 , RI2b5e785b3bc0_445, \13110 );
and \U$11883 ( \13750 , RI2b5e785b3260_465, \13112 );
and \U$11884 ( \13751 , RI2b5e785b2900_485, \13114 );
and \U$11885 ( \13752 , RI2b5e785b1910_505, \13116 );
and \U$11886 ( \13753 , RI2b5e785b0fb0_525, \13118 );
and \U$11887 ( \13754 , RI2b5e785b0650_545, \13120 );
and \U$11888 ( \13755 , RI2b5e785afcf0_565, \13122 );
and \U$11889 ( \13756 , RI2b5e785af0c0_585, \13124 );
or \U$11890 ( \13757 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 );
_DC g34fb ( \13758_nG34fb , \13757 , \13143 );
buf \U$11891 ( \13759 , \13758_nG34fb );
and \U$11892 ( \13760 , \13759 , \13193 );
and \U$11893 ( \13761 , RI2b5e785c06b8_264, \13088 );
and \U$11894 ( \13762 , RI2b5e785be048_284, \13094 );
and \U$11895 ( \13763 , RI2b5e785bbd98_304, \13096 );
and \U$11896 ( \13764 , RI2b5e785b9ea8_324, \13098 );
and \U$11897 ( \13765 , RI2b5e785b9548_344, \13100 );
and \U$11898 ( \13766 , RI2b5e785b7a18_364, \13102 );
and \U$11899 ( \13767 , RI2b5e785b70b8_384, \13104 );
and \U$11900 ( \13768 , RI2b5e785b5948_404, \13106 );
and \U$11901 ( \13769 , RI2b5e785b4fe8_424, \13108 );
and \U$11902 ( \13770 , RI2b5e785b3c38_444, \13110 );
and \U$11903 ( \13771 , RI2b5e785b32d8_464, \13112 );
and \U$11904 ( \13772 , RI2b5e785b2978_484, \13114 );
and \U$11905 ( \13773 , RI2b5e785b1988_504, \13116 );
and \U$11906 ( \13774 , RI2b5e785b1028_524, \13118 );
and \U$11907 ( \13775 , RI2b5e785b06c8_544, \13120 );
and \U$11908 ( \13776 , RI2b5e785afd68_564, \13122 );
and \U$11909 ( \13777 , RI2b5e785af138_584, \13124 );
or \U$11910 ( \13778 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 );
_DC g358e ( \13779_nG358e , \13778 , \13143 );
buf \U$11911 ( \13780 , \13779_nG358e );
and \U$11912 ( \13781 , \13780 , \13191 );
nor \U$11913 ( \13782 , \13760 , \13781 );
xnor \U$11914 ( \13783 , \13782 , \13219 );
and \U$11916 ( \13784 , RI2b5e785c05c8_266, \13088 );
and \U$11917 ( \13785 , RI2b5e785bdf58_286, \13094 );
and \U$11918 ( \13786 , RI2b5e785bbca8_306, \13096 );
and \U$11919 ( \13787 , RI2b5e785b9db8_326, \13098 );
and \U$11920 ( \13788 , RI2b5e785b9458_346, \13100 );
and \U$11921 ( \13789 , RI2b5e785b7928_366, \13102 );
and \U$11922 ( \13790 , RI2b5e785b6fc8_386, \13104 );
and \U$11923 ( \13791 , RI2b5e785b5858_406, \13106 );
and \U$11924 ( \13792 , RI2b5e785b4ef8_426, \13108 );
and \U$11925 ( \13793 , RI2b5e785b3b48_446, \13110 );
and \U$11926 ( \13794 , RI2b5e785b31e8_466, \13112 );
and \U$11927 ( \13795 , RI2b5e785b2888_486, \13114 );
and \U$11928 ( \13796 , RI2b5e785b1898_506, \13116 );
and \U$11929 ( \13797 , RI2b5e785b0f38_526, \13118 );
and \U$11930 ( \13798 , RI2b5e785b05d8_546, \13120 );
and \U$11931 ( \13799 , RI2b5e785afc78_566, \13122 );
and \U$11932 ( \13800 , RI2b5e785af048_586, \13124 );
or \U$11933 ( \13801 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 );
_DC g3473 ( \13802_nG3473 , \13801 , \13143 );
buf \U$11934 ( \13803 , \13802_nG3473 );
and \U$11935 ( \13804 , \13803 , \13246 );
nor \U$11936 ( \13805 , 1'b0 , \13804 );
xnor \U$11937 ( \13806 , \13805 , 1'b0 );
and \U$11938 ( \13807 , \13783 , \13806 );
and \U$11939 ( \13808 , \13738 , \13807 );
and \U$11940 ( \13809 , \13591 , \13807 );
or \U$11941 ( \13810 , \13739 , \13808 , \13809 );
and \U$11943 ( \13811 , \13732 , \13255 );
and \U$11944 ( \13812 , \13666 , \13253 );
nor \U$11945 ( \13813 , \13811 , \13812 );
xnor \U$11946 ( \13814 , \13813 , \13022 );
and \U$11947 ( \13815 , \13780 , \13193 );
and \U$11948 ( \13816 , \13711 , \13191 );
nor \U$11949 ( \13817 , \13815 , \13816 );
xnor \U$11950 ( \13818 , \13817 , \13219 );
xor \U$11951 ( \13819 , \13814 , \13818 );
and \U$11953 ( \13820 , \13759 , \13246 );
nor \U$11954 ( \13821 , 1'b0 , \13820 );
xnor \U$11955 ( \13822 , \13821 , 1'b0 );
xor \U$11956 ( \13823 , \13819 , \13822 );
and \U$11957 ( \13824 , \13582 , \13561 );
and \U$11958 ( \13825 , \13489 , \13559 );
nor \U$11959 ( \13826 , \13824 , \13825 );
xnor \U$11960 ( \13827 , \13826 , \13587 );
and \U$11961 ( \13828 , \13640 , \13619 );
and \U$11962 ( \13829 , \13549 , \13617 );
nor \U$11963 ( \13830 , \13828 , \13829 );
xnor \U$11964 ( \13831 , \13830 , \13645 );
xor \U$11965 ( \13832 , \13827 , \13831 );
and \U$11966 ( \13833 , \13687 , \13320 );
and \U$11967 ( \13834 , \13611 , \13318 );
nor \U$11968 ( \13835 , \13833 , \13834 );
xnor \U$11969 ( \13836 , \13835 , \13325 );
xor \U$11970 ( \13837 , \13832 , \13836 );
and \U$11971 ( \13838 , \13823 , \13837 );
or \U$11973 ( \13839 , 1'b0 , \13838 , 1'b0 );
xor \U$11974 ( \13840 , \13810 , \13839 );
and \U$11975 ( \13841 , \13711 , \13193 );
and \U$11976 ( \13842 , \13732 , \13191 );
nor \U$11977 ( \13843 , \13841 , \13842 );
xnor \U$11978 ( \13844 , \13843 , \13219 );
and \U$11980 ( \13845 , \13780 , \13246 );
nor \U$11981 ( \13846 , 1'b0 , \13845 );
xnor \U$11982 ( \13847 , \13846 , 1'b0 );
xor \U$11983 ( \13848 , \13844 , \13847 );
xor \U$11985 ( \13849 , \13848 , 1'b0 );
and \U$11986 ( \13850 , \13549 , \13619 );
and \U$11987 ( \13851 , \13582 , \13617 );
nor \U$11988 ( \13852 , \13850 , \13851 );
xnor \U$11989 ( \13853 , \13852 , \13645 );
and \U$11990 ( \13854 , \13611 , \13320 );
and \U$11991 ( \13855 , \13640 , \13318 );
nor \U$11992 ( \13856 , \13854 , \13855 );
xnor \U$11993 ( \13857 , \13856 , \13325 );
xor \U$11994 ( \13858 , \13853 , \13857 );
and \U$11995 ( \13859 , \13666 , \13255 );
and \U$11996 ( \13860 , \13687 , \13253 );
nor \U$11997 ( \13861 , \13859 , \13860 );
xnor \U$11998 ( \13862 , \13861 , \13022 );
xor \U$11999 ( \13863 , \13858 , \13862 );
xor \U$12000 ( \13864 , \13849 , \13863 );
and \U$12001 ( \13865 , \13373 , \13465 );
and \U$12002 ( \13866 , \13241 , \13462 );
nor \U$12003 ( \13867 , \13865 , \13866 );
xnor \U$12004 ( \13868 , \13867 , \13459 );
and \U$12005 ( \13869 , \13396 , \13501 );
and \U$12006 ( \13870 , \13352 , \13499 );
nor \U$12007 ( \13871 , \13869 , \13870 );
xnor \U$12008 ( \13872 , \13871 , \13527 );
xor \U$12009 ( \13873 , \13868 , \13872 );
and \U$12010 ( \13874 , \13489 , \13561 );
and \U$12011 ( \13875 , \13522 , \13559 );
nor \U$12012 ( \13876 , \13874 , \13875 );
xnor \U$12013 ( \13877 , \13876 , \13587 );
xor \U$12014 ( \13878 , \13873 , \13877 );
xor \U$12015 ( \13879 , \13864 , \13878 );
xor \U$12016 ( \13880 , \13840 , \13879 );
and \U$12018 ( \13881 , \13522 , \13465 );
and \U$12019 ( \13882 , \13396 , \13462 );
nor \U$12020 ( \13883 , \13881 , \13882 );
xnor \U$12021 ( \13884 , \13883 , \13459 );
and \U$12022 ( \13885 , \13582 , \13501 );
and \U$12023 ( \13886 , \13489 , \13499 );
nor \U$12024 ( \13887 , \13885 , \13886 );
xnor \U$12025 ( \13888 , \13887 , \13527 );
and \U$12026 ( \13889 , \13884 , \13888 );
or \U$12028 ( \13890 , 1'b0 , \13889 , 1'b0 );
and \U$12029 ( \13891 , \13640 , \13561 );
and \U$12030 ( \13892 , \13549 , \13559 );
nor \U$12031 ( \13893 , \13891 , \13892 );
xnor \U$12032 ( \13894 , \13893 , \13587 );
and \U$12033 ( \13895 , \13687 , \13619 );
and \U$12034 ( \13896 , \13611 , \13617 );
nor \U$12035 ( \13897 , \13895 , \13896 );
xnor \U$12036 ( \13898 , \13897 , \13645 );
and \U$12037 ( \13899 , \13894 , \13898 );
and \U$12038 ( \13900 , \13732 , \13320 );
and \U$12039 ( \13901 , \13666 , \13318 );
nor \U$12040 ( \13902 , \13900 , \13901 );
xnor \U$12041 ( \13903 , \13902 , \13325 );
and \U$12042 ( \13904 , \13898 , \13903 );
and \U$12043 ( \13905 , \13894 , \13903 );
or \U$12044 ( \13906 , \13899 , \13904 , \13905 );
and \U$12045 ( \13907 , \13890 , \13906 );
and \U$12046 ( \13908 , \13780 , \13255 );
and \U$12047 ( \13909 , \13711 , \13253 );
nor \U$12048 ( \13910 , \13908 , \13909 );
xnor \U$12049 ( \13911 , \13910 , \13022 );
and \U$12050 ( \13912 , \13803 , \13193 );
and \U$12051 ( \13913 , \13759 , \13191 );
nor \U$12052 ( \13914 , \13912 , \13913 );
xnor \U$12053 ( \13915 , \13914 , \13219 );
and \U$12054 ( \13916 , \13911 , \13915 );
and \U$12055 ( \13917 , RI2b5e785c0550_267, \13088 );
and \U$12056 ( \13918 , RI2b5e785bc590_287, \13094 );
and \U$12057 ( \13919 , RI2b5e785bbc30_307, \13096 );
and \U$12058 ( \13920 , RI2b5e785b9d40_327, \13098 );
and \U$12059 ( \13921 , RI2b5e785b93e0_347, \13100 );
and \U$12060 ( \13922 , RI2b5e785b78b0_367, \13102 );
and \U$12061 ( \13923 , RI2b5e785b6f50_387, \13104 );
and \U$12062 ( \13924 , RI2b5e785b57e0_407, \13106 );
and \U$12063 ( \13925 , RI2b5e785b4e80_427, \13108 );
and \U$12064 ( \13926 , RI2b5e785b3ad0_447, \13110 );
and \U$12065 ( \13927 , RI2b5e785b3170_467, \13112 );
and \U$12066 ( \13928 , RI2b5e785b2810_487, \13114 );
and \U$12067 ( \13929 , RI2b5e785b1820_507, \13116 );
and \U$12068 ( \13930 , RI2b5e785b0ec0_527, \13118 );
and \U$12069 ( \13931 , RI2b5e785b0560_547, \13120 );
and \U$12070 ( \13932 , RI2b5e785afc00_567, \13122 );
and \U$12071 ( \13933 , RI2b5e785aefd0_587, \13124 );
or \U$12072 ( \13934 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 );
_DC g33d8 ( \13935_nG33d8 , \13934 , \13143 );
buf \U$12073 ( \13936 , \13935_nG33d8 );
nand \U$12074 ( \13937 , \13936 , \13246 );
xnor \U$12075 ( \13938 , \13937 , 1'b0 );
and \U$12076 ( \13939 , \13915 , \13938 );
and \U$12077 ( \13940 , \13911 , \13938 );
or \U$12078 ( \13941 , \13916 , \13939 , \13940 );
and \U$12079 ( \13942 , \13906 , \13941 );
and \U$12080 ( \13943 , \13890 , \13941 );
or \U$12081 ( \13944 , \13907 , \13942 , \13943 );
xor \U$12082 ( \13945 , \13783 , \13806 );
xor \U$12083 ( \13946 , \13646 , \13690 );
xor \U$12084 ( \13947 , \13946 , \13735 );
and \U$12085 ( \13948 , \13945 , \13947 );
xor \U$12086 ( \13949 , \13469 , \13528 );
xor \U$12087 ( \13950 , \13949 , \13588 );
and \U$12088 ( \13951 , \13947 , \13950 );
and \U$12089 ( \13952 , \13945 , \13950 );
or \U$12090 ( \13953 , \13948 , \13951 , \13952 );
and \U$12091 ( \13954 , \13944 , \13953 );
and \U$12093 ( \13955 , \13352 , \13465 );
and \U$12094 ( \13956 , \13373 , \13462 );
nor \U$12095 ( \13957 , \13955 , \13956 );
xnor \U$12096 ( \13958 , \13957 , \13459 );
xor \U$12097 ( \13959 , 1'b0 , \13958 );
and \U$12098 ( \13960 , \13522 , \13501 );
and \U$12099 ( \13961 , \13396 , \13499 );
nor \U$12100 ( \13962 , \13960 , \13961 );
xnor \U$12101 ( \13963 , \13962 , \13527 );
xor \U$12102 ( \13964 , \13959 , \13963 );
and \U$12103 ( \13965 , \13953 , \13964 );
and \U$12104 ( \13966 , \13944 , \13964 );
or \U$12105 ( \13967 , \13954 , \13965 , \13966 );
xor \U$12107 ( \13968 , 1'b0 , \13823 );
xor \U$12108 ( \13969 , \13968 , \13837 );
xor \U$12109 ( \13970 , \13591 , \13738 );
xor \U$12110 ( \13971 , \13970 , \13807 );
and \U$12111 ( \13972 , \13969 , \13971 );
xor \U$12112 ( \13973 , \13967 , \13972 );
and \U$12114 ( \13974 , \13958 , \13963 );
or \U$12116 ( \13975 , 1'b0 , \13974 , 1'b0 );
and \U$12117 ( \13976 , \13827 , \13831 );
and \U$12118 ( \13977 , \13831 , \13836 );
and \U$12119 ( \13978 , \13827 , \13836 );
or \U$12120 ( \13979 , \13976 , \13977 , \13978 );
xor \U$12121 ( \13980 , \13975 , \13979 );
and \U$12122 ( \13981 , \13814 , \13818 );
and \U$12123 ( \13982 , \13818 , \13822 );
and \U$12124 ( \13983 , \13814 , \13822 );
or \U$12125 ( \13984 , \13981 , \13982 , \13983 );
xor \U$12126 ( \13985 , \13980 , \13984 );
xor \U$12127 ( \13986 , \13973 , \13985 );
xor \U$12128 ( \13987 , \13880 , \13986 );
and \U$12129 ( \13988 , \13489 , \13465 );
and \U$12130 ( \13989 , \13522 , \13462 );
nor \U$12131 ( \13990 , \13988 , \13989 );
xnor \U$12132 ( \13991 , \13990 , \13459 );
and \U$12133 ( \13992 , \13549 , \13501 );
and \U$12134 ( \13993 , \13582 , \13499 );
nor \U$12135 ( \13994 , \13992 , \13993 );
xnor \U$12136 ( \13995 , \13994 , \13527 );
and \U$12137 ( \13996 , \13991 , \13995 );
and \U$12138 ( \13997 , \13611 , \13561 );
and \U$12139 ( \13998 , \13640 , \13559 );
nor \U$12140 ( \13999 , \13997 , \13998 );
xnor \U$12141 ( \14000 , \13999 , \13587 );
and \U$12142 ( \14001 , \13995 , \14000 );
and \U$12143 ( \14002 , \13991 , \14000 );
or \U$12144 ( \14003 , \13996 , \14001 , \14002 );
and \U$12145 ( \14004 , \13666 , \13619 );
and \U$12146 ( \14005 , \13687 , \13617 );
nor \U$12147 ( \14006 , \14004 , \14005 );
xnor \U$12148 ( \14007 , \14006 , \13645 );
and \U$12149 ( \14008 , \13711 , \13320 );
and \U$12150 ( \14009 , \13732 , \13318 );
nor \U$12151 ( \14010 , \14008 , \14009 );
xnor \U$12152 ( \14011 , \14010 , \13325 );
and \U$12153 ( \14012 , \14007 , \14011 );
and \U$12154 ( \14013 , \13759 , \13255 );
and \U$12155 ( \14014 , \13780 , \13253 );
nor \U$12156 ( \14015 , \14013 , \14014 );
xnor \U$12157 ( \14016 , \14015 , \13022 );
and \U$12158 ( \14017 , \14011 , \14016 );
and \U$12159 ( \14018 , \14007 , \14016 );
or \U$12160 ( \14019 , \14012 , \14017 , \14018 );
and \U$12161 ( \14020 , \14003 , \14019 );
xor \U$12162 ( \14021 , \13911 , \13915 );
xor \U$12163 ( \14022 , \14021 , \13938 );
and \U$12164 ( \14023 , \14019 , \14022 );
and \U$12165 ( \14024 , \14003 , \14022 );
or \U$12166 ( \14025 , \14020 , \14023 , \14024 );
xor \U$12167 ( \14026 , \13894 , \13898 );
xor \U$12168 ( \14027 , \14026 , \13903 );
xor \U$12169 ( \14028 , 1'b0 , \13884 );
xor \U$12170 ( \14029 , \14028 , \13888 );
and \U$12171 ( \14030 , \14027 , \14029 );
and \U$12172 ( \14031 , \14025 , \14030 );
xor \U$12173 ( \14032 , \13945 , \13947 );
xor \U$12174 ( \14033 , \14032 , \13950 );
and \U$12175 ( \14034 , \14030 , \14033 );
and \U$12176 ( \14035 , \14025 , \14033 );
or \U$12177 ( \14036 , \14031 , \14034 , \14035 );
xor \U$12178 ( \14037 , \13969 , \13971 );
and \U$12179 ( \14038 , \14036 , \14037 );
xor \U$12180 ( \14039 , \13944 , \13953 );
xor \U$12181 ( \14040 , \14039 , \13964 );
and \U$12182 ( \14041 , \14037 , \14040 );
and \U$12183 ( \14042 , \14036 , \14040 );
or \U$12184 ( \14043 , \14038 , \14041 , \14042 );
nor \U$12185 ( \14044 , \13987 , \14043 );
and \U$12186 ( \14045 , \13967 , \13972 );
and \U$12187 ( \14046 , \13972 , \13985 );
and \U$12188 ( \14047 , \13967 , \13985 );
or \U$12189 ( \14048 , \14045 , \14046 , \14047 );
and \U$12190 ( \14049 , \13810 , \13839 );
and \U$12191 ( \14050 , \13839 , \13879 );
and \U$12192 ( \14051 , \13810 , \13879 );
or \U$12193 ( \14052 , \14049 , \14050 , \14051 );
and \U$12195 ( \14053 , \13241 , \13465 );
and \U$12196 ( \14054 , \13145 , \13462 );
nor \U$12197 ( \14055 , \14053 , \14054 );
xnor \U$12198 ( \14056 , \14055 , \13459 );
xor \U$12199 ( \14057 , 1'b0 , \14056 );
and \U$12200 ( \14058 , \13352 , \13501 );
and \U$12201 ( \14059 , \13373 , \13499 );
nor \U$12202 ( \14060 , \14058 , \14059 );
xnor \U$12203 ( \14061 , \14060 , \13527 );
xor \U$12204 ( \14062 , \14057 , \14061 );
and \U$12206 ( \14063 , \13687 , \13255 );
and \U$12207 ( \14064 , \13611 , \13253 );
nor \U$12208 ( \14065 , \14063 , \14064 );
xnor \U$12209 ( \14066 , \14065 , \13022 );
and \U$12210 ( \14067 , \13732 , \13193 );
and \U$12211 ( \14068 , \13666 , \13191 );
nor \U$12212 ( \14069 , \14067 , \14068 );
xnor \U$12213 ( \14070 , \14069 , \13219 );
xor \U$12214 ( \14071 , \14066 , \14070 );
and \U$12216 ( \14072 , \13711 , \13246 );
nor \U$12217 ( \14073 , 1'b0 , \14072 );
xnor \U$12218 ( \14074 , \14073 , 1'b0 );
xor \U$12219 ( \14075 , \14071 , \14074 );
xor \U$12220 ( \14076 , 1'b0 , \14075 );
xor \U$12221 ( \14077 , \14062 , \14076 );
and \U$12222 ( \14078 , \13868 , \13872 );
and \U$12223 ( \14079 , \13872 , \13877 );
and \U$12224 ( \14080 , \13868 , \13877 );
or \U$12225 ( \14081 , \14078 , \14079 , \14080 );
and \U$12226 ( \14082 , \13853 , \13857 );
and \U$12227 ( \14083 , \13857 , \13862 );
and \U$12228 ( \14084 , \13853 , \13862 );
or \U$12229 ( \14085 , \14082 , \14083 , \14084 );
xor \U$12230 ( \14086 , \14081 , \14085 );
and \U$12231 ( \14087 , \13844 , \13847 );
or \U$12234 ( \14088 , \14087 , 1'b0 , 1'b0 );
xor \U$12235 ( \14089 , \14086 , \14088 );
xor \U$12236 ( \14090 , \14077 , \14089 );
xor \U$12237 ( \14091 , \14052 , \14090 );
and \U$12238 ( \14092 , \13975 , \13979 );
and \U$12239 ( \14093 , \13979 , \13984 );
and \U$12240 ( \14094 , \13975 , \13984 );
or \U$12241 ( \14095 , \14092 , \14093 , \14094 );
and \U$12242 ( \14096 , \13849 , \13863 );
and \U$12243 ( \14097 , \13863 , \13878 );
and \U$12244 ( \14098 , \13849 , \13878 );
or \U$12245 ( \14099 , \14096 , \14097 , \14098 );
xor \U$12246 ( \14100 , \14095 , \14099 );
and \U$12247 ( \14101 , \13522 , \13561 );
and \U$12248 ( \14102 , \13396 , \13559 );
nor \U$12249 ( \14103 , \14101 , \14102 );
xnor \U$12250 ( \14104 , \14103 , \13587 );
and \U$12251 ( \14105 , \13582 , \13619 );
and \U$12252 ( \14106 , \13489 , \13617 );
nor \U$12253 ( \14107 , \14105 , \14106 );
xnor \U$12254 ( \14108 , \14107 , \13645 );
xor \U$12255 ( \14109 , \14104 , \14108 );
and \U$12256 ( \14110 , \13640 , \13320 );
and \U$12257 ( \14111 , \13549 , \13318 );
nor \U$12258 ( \14112 , \14110 , \14111 );
xnor \U$12259 ( \14113 , \14112 , \13325 );
xor \U$12260 ( \14114 , \14109 , \14113 );
xor \U$12261 ( \14115 , \14100 , \14114 );
xor \U$12262 ( \14116 , \14091 , \14115 );
xor \U$12263 ( \14117 , \14048 , \14116 );
and \U$12264 ( \14118 , \13880 , \13986 );
nor \U$12265 ( \14119 , \14117 , \14118 );
nor \U$12266 ( \14120 , \14044 , \14119 );
and \U$12267 ( \14121 , \14052 , \14090 );
and \U$12268 ( \14122 , \14090 , \14115 );
and \U$12269 ( \14123 , \14052 , \14115 );
or \U$12270 ( \14124 , \14121 , \14122 , \14123 );
and \U$12272 ( \14125 , \14056 , \14061 );
or \U$12274 ( \14126 , 1'b0 , \14125 , 1'b0 );
and \U$12275 ( \14127 , \14104 , \14108 );
and \U$12276 ( \14128 , \14108 , \14113 );
and \U$12277 ( \14129 , \14104 , \14113 );
or \U$12278 ( \14130 , \14127 , \14128 , \14129 );
xor \U$12279 ( \14131 , \14126 , \14130 );
and \U$12280 ( \14132 , \14066 , \14070 );
and \U$12281 ( \14133 , \14070 , \14074 );
and \U$12282 ( \14134 , \14066 , \14074 );
or \U$12283 ( \14135 , \14132 , \14133 , \14134 );
xor \U$12284 ( \14136 , \14131 , \14135 );
and \U$12285 ( \14137 , \14081 , \14085 );
and \U$12286 ( \14138 , \14085 , \14088 );
and \U$12287 ( \14139 , \14081 , \14088 );
or \U$12288 ( \14140 , \14137 , \14138 , \14139 );
xor \U$12290 ( \14141 , \14140 , 1'b0 );
and \U$12291 ( \14142 , \13145 , \13465 );
and \U$12292 ( \14143 , \13214 , \13462 );
nor \U$12293 ( \14144 , \14142 , \14143 );
xnor \U$12294 ( \14145 , \14144 , \13459 );
and \U$12295 ( \14146 , \13373 , \13501 );
and \U$12296 ( \14147 , \13241 , \13499 );
nor \U$12297 ( \14148 , \14146 , \14147 );
xnor \U$12298 ( \14149 , \14148 , \13527 );
xor \U$12299 ( \14150 , \14145 , \14149 );
and \U$12300 ( \14151 , \13396 , \13561 );
and \U$12301 ( \14152 , \13352 , \13559 );
nor \U$12302 ( \14153 , \14151 , \14152 );
xnor \U$12303 ( \14154 , \14153 , \13587 );
xor \U$12304 ( \14155 , \14150 , \14154 );
xor \U$12305 ( \14156 , \14141 , \14155 );
xor \U$12306 ( \14157 , \14136 , \14156 );
xor \U$12307 ( \14158 , \14124 , \14157 );
and \U$12308 ( \14159 , \14095 , \14099 );
and \U$12309 ( \14160 , \14099 , \14114 );
and \U$12310 ( \14161 , \14095 , \14114 );
or \U$12311 ( \14162 , \14159 , \14160 , \14161 );
and \U$12312 ( \14163 , \14062 , \14076 );
and \U$12313 ( \14164 , \14076 , \14089 );
and \U$12314 ( \14165 , \14062 , \14089 );
or \U$12315 ( \14166 , \14163 , \14164 , \14165 );
xor \U$12316 ( \14167 , \14162 , \14166 );
and \U$12318 ( \14168 , \13666 , \13193 );
and \U$12319 ( \14169 , \13687 , \13191 );
nor \U$12320 ( \14170 , \14168 , \14169 );
xnor \U$12321 ( \14171 , \14170 , \13219 );
and \U$12323 ( \14172 , \13732 , \13246 );
nor \U$12324 ( \14173 , 1'b0 , \14172 );
xnor \U$12325 ( \14174 , \14173 , 1'b0 );
xor \U$12326 ( \14175 , \14171 , \14174 );
xor \U$12328 ( \14176 , \14175 , 1'b0 );
xor \U$12329 ( \14177 , 1'b0 , \14176 );
and \U$12330 ( \14178 , \13489 , \13619 );
and \U$12331 ( \14179 , \13522 , \13617 );
nor \U$12332 ( \14180 , \14178 , \14179 );
xnor \U$12333 ( \14181 , \14180 , \13645 );
and \U$12334 ( \14182 , \13549 , \13320 );
and \U$12335 ( \14183 , \13582 , \13318 );
nor \U$12336 ( \14184 , \14182 , \14183 );
xnor \U$12337 ( \14185 , \14184 , \13325 );
xor \U$12338 ( \14186 , \14181 , \14185 );
and \U$12339 ( \14187 , \13611 , \13255 );
and \U$12340 ( \14188 , \13640 , \13253 );
nor \U$12341 ( \14189 , \14187 , \14188 );
xnor \U$12342 ( \14190 , \14189 , \13022 );
xor \U$12343 ( \14191 , \14186 , \14190 );
xor \U$12344 ( \14192 , \14177 , \14191 );
xor \U$12345 ( \14193 , \14167 , \14192 );
xor \U$12346 ( \14194 , \14158 , \14193 );
and \U$12347 ( \14195 , \14048 , \14116 );
nor \U$12348 ( \14196 , \14194 , \14195 );
and \U$12349 ( \14197 , \14162 , \14166 );
and \U$12350 ( \14198 , \14166 , \14192 );
and \U$12351 ( \14199 , \14162 , \14192 );
or \U$12352 ( \14200 , \14197 , \14198 , \14199 );
and \U$12353 ( \14201 , \14136 , \14156 );
xor \U$12354 ( \14202 , \14200 , \14201 );
and \U$12357 ( \14203 , \14140 , \14155 );
or \U$12358 ( \14204 , 1'b0 , 1'b0 , \14203 );
and \U$12360 ( \14205 , \13640 , \13255 );
and \U$12361 ( \14206 , \13549 , \13253 );
nor \U$12362 ( \14207 , \14205 , \14206 );
xnor \U$12363 ( \14208 , \14207 , \13022 );
and \U$12364 ( \14209 , \13687 , \13193 );
and \U$12365 ( \14210 , \13611 , \13191 );
nor \U$12366 ( \14211 , \14209 , \14210 );
xnor \U$12367 ( \14212 , \14211 , \13219 );
xor \U$12368 ( \14213 , \14208 , \14212 );
and \U$12370 ( \14214 , \13666 , \13246 );
nor \U$12371 ( \14215 , 1'b0 , \14214 );
xnor \U$12372 ( \14216 , \14215 , 1'b0 );
xor \U$12373 ( \14217 , \14213 , \14216 );
xor \U$12374 ( \14218 , 1'b0 , \14217 );
and \U$12375 ( \14219 , \13352 , \13561 );
and \U$12376 ( \14220 , \13373 , \13559 );
nor \U$12377 ( \14221 , \14219 , \14220 );
xnor \U$12378 ( \14222 , \14221 , \13587 );
and \U$12379 ( \14223 , \13522 , \13619 );
and \U$12380 ( \14224 , \13396 , \13617 );
nor \U$12381 ( \14225 , \14223 , \14224 );
xnor \U$12382 ( \14226 , \14225 , \13645 );
xor \U$12383 ( \14227 , \14222 , \14226 );
and \U$12384 ( \14228 , \13582 , \13320 );
and \U$12385 ( \14229 , \13489 , \13318 );
nor \U$12386 ( \14230 , \14228 , \14229 );
xnor \U$12387 ( \14231 , \14230 , \13325 );
xor \U$12388 ( \14232 , \14227 , \14231 );
xor \U$12389 ( \14233 , \14218 , \14232 );
and \U$12390 ( \14234 , \14145 , \14149 );
and \U$12391 ( \14235 , \14149 , \14154 );
and \U$12392 ( \14236 , \14145 , \14154 );
or \U$12393 ( \14237 , \14234 , \14235 , \14236 );
and \U$12394 ( \14238 , \14181 , \14185 );
and \U$12395 ( \14239 , \14185 , \14190 );
and \U$12396 ( \14240 , \14181 , \14190 );
or \U$12397 ( \14241 , \14238 , \14239 , \14240 );
xor \U$12398 ( \14242 , \14237 , \14241 );
and \U$12399 ( \14243 , \14171 , \14174 );
or \U$12402 ( \14244 , \14243 , 1'b0 , 1'b0 );
xor \U$12403 ( \14245 , \14242 , \14244 );
xor \U$12404 ( \14246 , \14233 , \14245 );
xor \U$12405 ( \14247 , \14204 , \14246 );
and \U$12406 ( \14248 , \14126 , \14130 );
and \U$12407 ( \14249 , \14130 , \14135 );
and \U$12408 ( \14250 , \14126 , \14135 );
or \U$12409 ( \14251 , \14248 , \14249 , \14250 );
and \U$12411 ( \14252 , \14176 , \14191 );
or \U$12413 ( \14253 , 1'b0 , \14252 , 1'b0 );
xor \U$12414 ( \14254 , \14251 , \14253 );
and \U$12416 ( \14255 , \13214 , \13465 );
not \U$12417 ( \14256 , \14255 );
xnor \U$12418 ( \14257 , \14256 , \13459 );
xor \U$12419 ( \14258 , 1'b0 , \14257 );
and \U$12420 ( \14259 , \13241 , \13501 );
and \U$12421 ( \14260 , \13145 , \13499 );
nor \U$12422 ( \14261 , \14259 , \14260 );
xnor \U$12423 ( \14262 , \14261 , \13527 );
xor \U$12424 ( \14263 , \14258 , \14262 );
xor \U$12425 ( \14264 , \14254 , \14263 );
xor \U$12426 ( \14265 , \14247 , \14264 );
xor \U$12427 ( \14266 , \14202 , \14265 );
and \U$12428 ( \14267 , \14124 , \14157 );
and \U$12429 ( \14268 , \14157 , \14193 );
and \U$12430 ( \14269 , \14124 , \14193 );
or \U$12431 ( \14270 , \14267 , \14268 , \14269 );
nor \U$12432 ( \14271 , \14266 , \14270 );
nor \U$12433 ( \14272 , \14196 , \14271 );
nand \U$12434 ( \14273 , \14120 , \14272 );
and \U$12435 ( \14274 , \14204 , \14246 );
and \U$12436 ( \14275 , \14246 , \14264 );
and \U$12437 ( \14276 , \14204 , \14264 );
or \U$12438 ( \14277 , \14274 , \14275 , \14276 );
and \U$12439 ( \14278 , \14237 , \14241 );
and \U$12440 ( \14279 , \14241 , \14244 );
and \U$12441 ( \14280 , \14237 , \14244 );
or \U$12442 ( \14281 , \14278 , \14279 , \14280 );
and \U$12444 ( \14282 , \14217 , \14232 );
or \U$12446 ( \14283 , 1'b0 , \14282 , 1'b0 );
xor \U$12447 ( \14284 , \14281 , \14283 );
and \U$12448 ( \14285 , \13396 , \13619 );
and \U$12449 ( \14286 , \13352 , \13617 );
nor \U$12450 ( \14287 , \14285 , \14286 );
xnor \U$12451 ( \14288 , \14287 , \13645 );
and \U$12452 ( \14289 , \13489 , \13320 );
and \U$12453 ( \14290 , \13522 , \13318 );
nor \U$12454 ( \14291 , \14289 , \14290 );
xnor \U$12455 ( \14292 , \14291 , \13325 );
xor \U$12456 ( \14293 , \14288 , \14292 );
and \U$12457 ( \14294 , \13549 , \13255 );
and \U$12458 ( \14295 , \13582 , \13253 );
nor \U$12459 ( \14296 , \14294 , \14295 );
xnor \U$12460 ( \14297 , \14296 , \13022 );
xor \U$12461 ( \14298 , \14293 , \14297 );
xor \U$12462 ( \14299 , \14284 , \14298 );
xor \U$12463 ( \14300 , \14277 , \14299 );
and \U$12464 ( \14301 , \14251 , \14253 );
and \U$12465 ( \14302 , \14253 , \14263 );
and \U$12466 ( \14303 , \14251 , \14263 );
or \U$12467 ( \14304 , \14301 , \14302 , \14303 );
and \U$12468 ( \14305 , \14233 , \14245 );
xor \U$12469 ( \14306 , \14304 , \14305 );
not \U$12470 ( \14307 , \13459 );
and \U$12471 ( \14308 , \13145 , \13501 );
and \U$12472 ( \14309 , \13214 , \13499 );
nor \U$12473 ( \14310 , \14308 , \14309 );
xnor \U$12474 ( \14311 , \14310 , \13527 );
xor \U$12475 ( \14312 , \14307 , \14311 );
and \U$12476 ( \14313 , \13373 , \13561 );
and \U$12477 ( \14314 , \13241 , \13559 );
nor \U$12478 ( \14315 , \14313 , \14314 );
xnor \U$12479 ( \14316 , \14315 , \13587 );
xor \U$12480 ( \14317 , \14312 , \14316 );
and \U$12482 ( \14318 , \13611 , \13193 );
and \U$12483 ( \14319 , \13640 , \13191 );
nor \U$12484 ( \14320 , \14318 , \14319 );
xnor \U$12485 ( \14321 , \14320 , \13219 );
and \U$12487 ( \14322 , \13687 , \13246 );
nor \U$12488 ( \14323 , 1'b0 , \14322 );
xnor \U$12489 ( \14324 , \14323 , 1'b0 );
xor \U$12490 ( \14325 , \14321 , \14324 );
xor \U$12492 ( \14326 , \14325 , 1'b0 );
xor \U$12493 ( \14327 , 1'b1 , \14326 );
xor \U$12494 ( \14328 , \14317 , \14327 );
and \U$12496 ( \14329 , \14257 , \14262 );
or \U$12498 ( \14330 , 1'b0 , \14329 , 1'b0 );
and \U$12499 ( \14331 , \14222 , \14226 );
and \U$12500 ( \14332 , \14226 , \14231 );
and \U$12501 ( \14333 , \14222 , \14231 );
or \U$12502 ( \14334 , \14331 , \14332 , \14333 );
xor \U$12503 ( \14335 , \14330 , \14334 );
and \U$12504 ( \14336 , \14208 , \14212 );
and \U$12505 ( \14337 , \14212 , \14216 );
and \U$12506 ( \14338 , \14208 , \14216 );
or \U$12507 ( \14339 , \14336 , \14337 , \14338 );
xor \U$12508 ( \14340 , \14335 , \14339 );
xor \U$12509 ( \14341 , \14328 , \14340 );
xor \U$12510 ( \14342 , \14306 , \14341 );
xor \U$12511 ( \14343 , \14300 , \14342 );
and \U$12512 ( \14344 , \14200 , \14201 );
and \U$12513 ( \14345 , \14201 , \14265 );
and \U$12514 ( \14346 , \14200 , \14265 );
or \U$12515 ( \14347 , \14344 , \14345 , \14346 );
nor \U$12516 ( \14348 , \14343 , \14347 );
and \U$12517 ( \14349 , \14304 , \14305 );
and \U$12518 ( \14350 , \14305 , \14341 );
and \U$12519 ( \14351 , \14304 , \14341 );
or \U$12520 ( \14352 , \14349 , \14350 , \14351 );
and \U$12521 ( \14353 , \14307 , \14311 );
and \U$12522 ( \14354 , \14311 , \14316 );
and \U$12523 ( \14355 , \14307 , \14316 );
or \U$12524 ( \14356 , \14353 , \14354 , \14355 );
and \U$12525 ( \14357 , \14288 , \14292 );
and \U$12526 ( \14358 , \14292 , \14297 );
and \U$12527 ( \14359 , \14288 , \14297 );
or \U$12528 ( \14360 , \14357 , \14358 , \14359 );
xor \U$12529 ( \14361 , \14356 , \14360 );
and \U$12530 ( \14362 , \14321 , \14324 );
or \U$12533 ( \14363 , \14362 , 1'b0 , 1'b0 );
xor \U$12534 ( \14364 , \14361 , \14363 );
and \U$12535 ( \14365 , \14330 , \14334 );
and \U$12536 ( \14366 , \14334 , \14339 );
and \U$12537 ( \14367 , \14330 , \14339 );
or \U$12538 ( \14368 , \14365 , \14366 , \14367 );
and \U$12541 ( \14369 , 1'b1 , \14326 );
or \U$12543 ( \14370 , 1'b0 , \14369 , 1'b0 );
xor \U$12544 ( \14371 , \14368 , \14370 );
and \U$12545 ( \14372 , \13640 , \13193 );
and \U$12546 ( \14373 , \13549 , \13191 );
nor \U$12547 ( \14374 , \14372 , \14373 );
xnor \U$12548 ( \14375 , \14374 , \13219 );
and \U$12550 ( \14376 , \13611 , \13246 );
nor \U$12551 ( \14377 , 1'b0 , \14376 );
xnor \U$12552 ( \14378 , \14377 , 1'b0 );
xor \U$12553 ( \14379 , \14375 , \14378 );
xor \U$12555 ( \14380 , \14379 , 1'b0 );
and \U$12556 ( \14381 , \13352 , \13619 );
and \U$12557 ( \14382 , \13373 , \13617 );
nor \U$12558 ( \14383 , \14381 , \14382 );
xnor \U$12559 ( \14384 , \14383 , \13645 );
and \U$12560 ( \14385 , \13522 , \13320 );
and \U$12561 ( \14386 , \13396 , \13318 );
nor \U$12562 ( \14387 , \14385 , \14386 );
xnor \U$12563 ( \14388 , \14387 , \13325 );
xor \U$12564 ( \14389 , \14384 , \14388 );
and \U$12565 ( \14390 , \13582 , \13255 );
and \U$12566 ( \14391 , \13489 , \13253 );
nor \U$12567 ( \14392 , \14390 , \14391 );
xnor \U$12568 ( \14393 , \14392 , \13022 );
xor \U$12569 ( \14394 , \14389 , \14393 );
xor \U$12570 ( \14395 , \14380 , \14394 );
and \U$12572 ( \14396 , \13214 , \13501 );
not \U$12573 ( \14397 , \14396 );
xnor \U$12574 ( \14398 , \14397 , \13527 );
xor \U$12575 ( \14399 , 1'b0 , \14398 );
and \U$12576 ( \14400 , \13241 , \13561 );
and \U$12577 ( \14401 , \13145 , \13559 );
nor \U$12578 ( \14402 , \14400 , \14401 );
xnor \U$12579 ( \14403 , \14402 , \13587 );
xor \U$12580 ( \14404 , \14399 , \14403 );
xor \U$12581 ( \14405 , \14395 , \14404 );
xor \U$12582 ( \14406 , \14371 , \14405 );
xor \U$12583 ( \14407 , \14364 , \14406 );
xor \U$12584 ( \14408 , \14352 , \14407 );
and \U$12585 ( \14409 , \14281 , \14283 );
and \U$12586 ( \14410 , \14283 , \14298 );
and \U$12587 ( \14411 , \14281 , \14298 );
or \U$12588 ( \14412 , \14409 , \14410 , \14411 );
and \U$12589 ( \14413 , \14317 , \14327 );
and \U$12590 ( \14414 , \14327 , \14340 );
and \U$12591 ( \14415 , \14317 , \14340 );
or \U$12592 ( \14416 , \14413 , \14414 , \14415 );
xor \U$12593 ( \14417 , \14412 , \14416 );
xor \U$12595 ( \14418 , \14417 , 1'b1 );
xor \U$12596 ( \14419 , \14408 , \14418 );
and \U$12597 ( \14420 , \14277 , \14299 );
and \U$12598 ( \14421 , \14299 , \14342 );
and \U$12599 ( \14422 , \14277 , \14342 );
or \U$12600 ( \14423 , \14420 , \14421 , \14422 );
nor \U$12601 ( \14424 , \14419 , \14423 );
nor \U$12602 ( \14425 , \14348 , \14424 );
and \U$12603 ( \14426 , \14412 , \14416 );
and \U$12604 ( \14427 , \14416 , 1'b1 );
and \U$12605 ( \14428 , \14412 , 1'b1 );
or \U$12606 ( \14429 , \14426 , \14427 , \14428 );
and \U$12607 ( \14430 , \14364 , \14406 );
xor \U$12608 ( \14431 , \14429 , \14430 );
and \U$12609 ( \14432 , \14368 , \14370 );
and \U$12610 ( \14433 , \14370 , \14405 );
and \U$12611 ( \14434 , \14368 , \14405 );
or \U$12612 ( \14435 , \14432 , \14433 , \14434 );
and \U$12614 ( \14436 , \13640 , \13246 );
nor \U$12615 ( \14437 , 1'b0 , \14436 );
xnor \U$12616 ( \14438 , \14437 , 1'b0 );
xor \U$12618 ( \14439 , \14438 , 1'b0 );
xor \U$12620 ( \14440 , \14439 , 1'b0 );
and \U$12621 ( \14441 , \13396 , \13320 );
and \U$12622 ( \14442 , \13352 , \13318 );
nor \U$12623 ( \14443 , \14441 , \14442 );
xnor \U$12624 ( \14444 , \14443 , \13325 );
and \U$12625 ( \14445 , \13489 , \13255 );
and \U$12626 ( \14446 , \13522 , \13253 );
nor \U$12627 ( \14447 , \14445 , \14446 );
xnor \U$12628 ( \14448 , \14447 , \13022 );
xor \U$12629 ( \14449 , \14444 , \14448 );
and \U$12630 ( \14450 , \13549 , \13193 );
and \U$12631 ( \14451 , \13582 , \13191 );
nor \U$12632 ( \14452 , \14450 , \14451 );
xnor \U$12633 ( \14453 , \14452 , \13219 );
xor \U$12634 ( \14454 , \14449 , \14453 );
xor \U$12635 ( \14455 , \14440 , \14454 );
not \U$12636 ( \14456 , \13527 );
and \U$12637 ( \14457 , \13145 , \13561 );
and \U$12638 ( \14458 , \13214 , \13559 );
nor \U$12639 ( \14459 , \14457 , \14458 );
xnor \U$12640 ( \14460 , \14459 , \13587 );
xor \U$12641 ( \14461 , \14456 , \14460 );
and \U$12642 ( \14462 , \13373 , \13619 );
and \U$12643 ( \14463 , \13241 , \13617 );
nor \U$12644 ( \14464 , \14462 , \14463 );
xnor \U$12645 ( \14465 , \14464 , \13645 );
xor \U$12646 ( \14466 , \14461 , \14465 );
xor \U$12647 ( \14467 , \14455 , \14466 );
xor \U$12649 ( \14468 , \14467 , 1'b0 );
and \U$12651 ( \14469 , \14398 , \14403 );
or \U$12653 ( \14470 , 1'b0 , \14469 , 1'b0 );
and \U$12654 ( \14471 , \14384 , \14388 );
and \U$12655 ( \14472 , \14388 , \14393 );
and \U$12656 ( \14473 , \14384 , \14393 );
or \U$12657 ( \14474 , \14471 , \14472 , \14473 );
xor \U$12658 ( \14475 , \14470 , \14474 );
and \U$12659 ( \14476 , \14375 , \14378 );
or \U$12662 ( \14477 , \14476 , 1'b0 , 1'b0 );
xor \U$12663 ( \14478 , \14475 , \14477 );
xor \U$12664 ( \14479 , \14468 , \14478 );
xor \U$12665 ( \14480 , \14435 , \14479 );
and \U$12666 ( \14481 , \14356 , \14360 );
and \U$12667 ( \14482 , \14360 , \14363 );
and \U$12668 ( \14483 , \14356 , \14363 );
or \U$12669 ( \14484 , \14481 , \14482 , \14483 );
xor \U$12671 ( \14485 , \14484 , 1'b0 );
and \U$12672 ( \14486 , \14380 , \14394 );
and \U$12673 ( \14487 , \14394 , \14404 );
and \U$12674 ( \14488 , \14380 , \14404 );
or \U$12675 ( \14489 , \14486 , \14487 , \14488 );
xor \U$12676 ( \14490 , \14485 , \14489 );
xor \U$12677 ( \14491 , \14480 , \14490 );
xor \U$12678 ( \14492 , \14431 , \14491 );
and \U$12679 ( \14493 , \14352 , \14407 );
and \U$12680 ( \14494 , \14407 , \14418 );
and \U$12681 ( \14495 , \14352 , \14418 );
or \U$12682 ( \14496 , \14493 , \14494 , \14495 );
nor \U$12683 ( \14497 , \14492 , \14496 );
and \U$12684 ( \14498 , \14435 , \14479 );
and \U$12685 ( \14499 , \14479 , \14490 );
and \U$12686 ( \14500 , \14435 , \14490 );
or \U$12687 ( \14501 , \14498 , \14499 , \14500 );
and \U$12688 ( \14502 , \14470 , \14474 );
and \U$12689 ( \14503 , \14474 , \14477 );
and \U$12690 ( \14504 , \14470 , \14477 );
or \U$12691 ( \14505 , \14502 , \14503 , \14504 );
xor \U$12693 ( \14506 , \14505 , 1'b0 );
and \U$12694 ( \14507 , \14440 , \14454 );
and \U$12695 ( \14508 , \14454 , \14466 );
and \U$12696 ( \14509 , \14440 , \14466 );
or \U$12697 ( \14510 , \14507 , \14508 , \14509 );
xor \U$12698 ( \14511 , \14506 , \14510 );
xor \U$12699 ( \14512 , \14501 , \14511 );
and \U$12702 ( \14513 , \14484 , \14489 );
or \U$12703 ( \14514 , 1'b0 , 1'b0 , \14513 );
and \U$12706 ( \14515 , \14467 , \14478 );
or \U$12707 ( \14516 , 1'b0 , 1'b0 , \14515 );
xor \U$12708 ( \14517 , \14514 , \14516 );
and \U$12709 ( \14518 , \13352 , \13320 );
and \U$12710 ( \14519 , \13373 , \13318 );
nor \U$12711 ( \14520 , \14518 , \14519 );
xnor \U$12712 ( \14521 , \14520 , \13325 );
and \U$12713 ( \14522 , \13522 , \13255 );
and \U$12714 ( \14523 , \13396 , \13253 );
nor \U$12715 ( \14524 , \14522 , \14523 );
xnor \U$12716 ( \14525 , \14524 , \13022 );
xor \U$12717 ( \14526 , \14521 , \14525 );
and \U$12718 ( \14527 , \13582 , \13193 );
and \U$12719 ( \14528 , \13489 , \13191 );
nor \U$12720 ( \14529 , \14527 , \14528 );
xnor \U$12721 ( \14530 , \14529 , \13219 );
xor \U$12722 ( \14531 , \14526 , \14530 );
and \U$12724 ( \14532 , \13214 , \13561 );
not \U$12725 ( \14533 , \14532 );
xnor \U$12726 ( \14534 , \14533 , \13587 );
xor \U$12727 ( \14535 , 1'b0 , \14534 );
and \U$12728 ( \14536 , \13241 , \13619 );
and \U$12729 ( \14537 , \13145 , \13617 );
nor \U$12730 ( \14538 , \14536 , \14537 );
xnor \U$12731 ( \14539 , \14538 , \13645 );
xor \U$12732 ( \14540 , \14535 , \14539 );
xor \U$12733 ( \14541 , \14531 , \14540 );
and \U$12736 ( \14542 , \13549 , \13246 );
nor \U$12737 ( \14543 , 1'b0 , \14542 );
xnor \U$12738 ( \14544 , \14543 , 1'b0 );
xor \U$12740 ( \14545 , \14544 , 1'b0 );
xor \U$12742 ( \14546 , \14545 , 1'b0 );
xnor \U$12743 ( \14547 , 1'b0 , \14546 );
xor \U$12744 ( \14548 , \14541 , \14547 );
and \U$12745 ( \14549 , \14456 , \14460 );
and \U$12746 ( \14550 , \14460 , \14465 );
and \U$12747 ( \14551 , \14456 , \14465 );
or \U$12748 ( \14552 , \14549 , \14550 , \14551 );
and \U$12749 ( \14553 , \14444 , \14448 );
and \U$12750 ( \14554 , \14448 , \14453 );
and \U$12751 ( \14555 , \14444 , \14453 );
or \U$12752 ( \14556 , \14553 , \14554 , \14555 );
xor \U$12753 ( \14557 , \14552 , \14556 );
xor \U$12755 ( \14558 , \14557 , 1'b0 );
xor \U$12756 ( \14559 , \14548 , \14558 );
xor \U$12757 ( \14560 , \14517 , \14559 );
xor \U$12758 ( \14561 , \14512 , \14560 );
and \U$12759 ( \14562 , \14429 , \14430 );
and \U$12760 ( \14563 , \14430 , \14491 );
and \U$12761 ( \14564 , \14429 , \14491 );
or \U$12762 ( \14565 , \14562 , \14563 , \14564 );
nor \U$12763 ( \14566 , \14561 , \14565 );
nor \U$12764 ( \14567 , \14497 , \14566 );
nand \U$12765 ( \14568 , \14425 , \14567 );
nor \U$12766 ( \14569 , \14273 , \14568 );
and \U$12767 ( \14570 , \14514 , \14516 );
and \U$12768 ( \14571 , \14516 , \14559 );
and \U$12769 ( \14572 , \14514 , \14559 );
or \U$12770 ( \14573 , \14570 , \14571 , \14572 );
and \U$12771 ( \14574 , \14552 , \14556 );
or \U$12774 ( \14575 , \14574 , 1'b0 , 1'b0 );
or \U$12775 ( \14576 , 1'b0 , \14546 );
xor \U$12776 ( \14577 , \14575 , \14576 );
and \U$12777 ( \14578 , \14531 , \14540 );
xor \U$12778 ( \14579 , \14577 , \14578 );
xor \U$12779 ( \14580 , \14573 , \14579 );
and \U$12782 ( \14581 , \14505 , \14510 );
or \U$12783 ( \14582 , 1'b0 , 1'b0 , \14581 );
and \U$12784 ( \14583 , \14541 , \14547 );
and \U$12785 ( \14584 , \14547 , \14558 );
and \U$12786 ( \14585 , \14541 , \14558 );
or \U$12787 ( \14586 , \14583 , \14584 , \14585 );
xor \U$12788 ( \14587 , \14582 , \14586 );
and \U$12790 ( \14588 , \13396 , \13255 );
and \U$12791 ( \14589 , \13352 , \13253 );
nor \U$12792 ( \14590 , \14588 , \14589 );
xnor \U$12793 ( \14591 , \14590 , \13022 );
and \U$12794 ( \14592 , \13489 , \13193 );
and \U$12795 ( \14593 , \13522 , \13191 );
nor \U$12796 ( \14594 , \14592 , \14593 );
xnor \U$12797 ( \14595 , \14594 , \13219 );
xor \U$12798 ( \14596 , \14591 , \14595 );
and \U$12800 ( \14597 , \13582 , \13246 );
nor \U$12801 ( \14598 , 1'b0 , \14597 );
xnor \U$12802 ( \14599 , \14598 , 1'b0 );
xor \U$12803 ( \14600 , \14596 , \14599 );
xor \U$12804 ( \14601 , 1'b0 , \14600 );
not \U$12805 ( \14602 , \13587 );
and \U$12806 ( \14603 , \13145 , \13619 );
and \U$12807 ( \14604 , \13214 , \13617 );
nor \U$12808 ( \14605 , \14603 , \14604 );
xnor \U$12809 ( \14606 , \14605 , \13645 );
xor \U$12810 ( \14607 , \14602 , \14606 );
and \U$12811 ( \14608 , \13373 , \13320 );
and \U$12812 ( \14609 , \13241 , \13318 );
nor \U$12813 ( \14610 , \14608 , \14609 );
xnor \U$12814 ( \14611 , \14610 , \13325 );
xor \U$12815 ( \14612 , \14607 , \14611 );
xor \U$12816 ( \14613 , \14601 , \14612 );
xor \U$12818 ( \14614 , \14613 , 1'b0 );
and \U$12820 ( \14615 , \14534 , \14539 );
or \U$12822 ( \14616 , 1'b0 , \14615 , 1'b0 );
and \U$12823 ( \14617 , \14521 , \14525 );
and \U$12824 ( \14618 , \14525 , \14530 );
and \U$12825 ( \14619 , \14521 , \14530 );
or \U$12826 ( \14620 , \14617 , \14618 , \14619 );
xor \U$12827 ( \14621 , \14616 , \14620 );
xor \U$12829 ( \14622 , \14621 , 1'b0 );
xor \U$12830 ( \14623 , \14614 , \14622 );
xor \U$12831 ( \14624 , \14587 , \14623 );
xor \U$12832 ( \14625 , \14580 , \14624 );
and \U$12833 ( \14626 , \14501 , \14511 );
and \U$12834 ( \14627 , \14511 , \14560 );
and \U$12835 ( \14628 , \14501 , \14560 );
or \U$12836 ( \14629 , \14626 , \14627 , \14628 );
nor \U$12837 ( \14630 , \14625 , \14629 );
and \U$12838 ( \14631 , \14582 , \14586 );
and \U$12839 ( \14632 , \14586 , \14623 );
and \U$12840 ( \14633 , \14582 , \14623 );
or \U$12841 ( \14634 , \14631 , \14632 , \14633 );
and \U$12842 ( \14635 , \14616 , \14620 );
or \U$12845 ( \14636 , \14635 , 1'b0 , 1'b0 );
xor \U$12847 ( \14637 , \14636 , 1'b0 );
and \U$12849 ( \14638 , \14600 , \14612 );
or \U$12851 ( \14639 , 1'b0 , \14638 , 1'b0 );
xor \U$12852 ( \14640 , \14637 , \14639 );
xor \U$12853 ( \14641 , \14634 , \14640 );
and \U$12854 ( \14642 , \14575 , \14576 );
and \U$12855 ( \14643 , \14576 , \14578 );
and \U$12856 ( \14644 , \14575 , \14578 );
or \U$12857 ( \14645 , \14642 , \14643 , \14644 );
and \U$12860 ( \14646 , \14613 , \14622 );
or \U$12861 ( \14647 , 1'b0 , 1'b0 , \14646 );
xor \U$12862 ( \14648 , \14645 , \14647 );
and \U$12863 ( \14649 , \13352 , \13255 );
and \U$12864 ( \14650 , \13373 , \13253 );
nor \U$12865 ( \14651 , \14649 , \14650 );
xnor \U$12866 ( \14652 , \14651 , \13022 );
and \U$12867 ( \14653 , \13522 , \13193 );
and \U$12868 ( \14654 , \13396 , \13191 );
nor \U$12869 ( \14655 , \14653 , \14654 );
xnor \U$12870 ( \14656 , \14655 , \13219 );
xor \U$12871 ( \14657 , \14652 , \14656 );
and \U$12873 ( \14658 , \13489 , \13246 );
nor \U$12874 ( \14659 , 1'b0 , \14658 );
xnor \U$12875 ( \14660 , \14659 , 1'b0 );
xor \U$12876 ( \14661 , \14657 , \14660 );
and \U$12878 ( \14662 , \13214 , \13619 );
not \U$12879 ( \14663 , \14662 );
xnor \U$12880 ( \14664 , \14663 , \13645 );
xor \U$12881 ( \14665 , 1'b0 , \14664 );
and \U$12882 ( \14666 , \13241 , \13320 );
and \U$12883 ( \14667 , \13145 , \13318 );
nor \U$12884 ( \14668 , \14666 , \14667 );
xnor \U$12885 ( \14669 , \14668 , \13325 );
xor \U$12886 ( \14670 , \14665 , \14669 );
xor \U$12887 ( \14671 , \14661 , \14670 );
xor \U$12889 ( \14672 , \14671 , 1'b1 );
and \U$12890 ( \14673 , \14602 , \14606 );
and \U$12891 ( \14674 , \14606 , \14611 );
and \U$12892 ( \14675 , \14602 , \14611 );
or \U$12893 ( \14676 , \14673 , \14674 , \14675 );
and \U$12894 ( \14677 , \14591 , \14595 );
and \U$12895 ( \14678 , \14595 , \14599 );
and \U$12896 ( \14679 , \14591 , \14599 );
or \U$12897 ( \14680 , \14677 , \14678 , \14679 );
xor \U$12898 ( \14681 , \14676 , \14680 );
xor \U$12900 ( \14682 , \14681 , 1'b0 );
xor \U$12901 ( \14683 , \14672 , \14682 );
xor \U$12902 ( \14684 , \14648 , \14683 );
xor \U$12903 ( \14685 , \14641 , \14684 );
and \U$12904 ( \14686 , \14573 , \14579 );
and \U$12905 ( \14687 , \14579 , \14624 );
and \U$12906 ( \14688 , \14573 , \14624 );
or \U$12907 ( \14689 , \14686 , \14687 , \14688 );
nor \U$12908 ( \14690 , \14685 , \14689 );
nor \U$12909 ( \14691 , \14630 , \14690 );
and \U$12910 ( \14692 , \14645 , \14647 );
and \U$12911 ( \14693 , \14647 , \14683 );
and \U$12912 ( \14694 , \14645 , \14683 );
or \U$12913 ( \14695 , \14692 , \14693 , \14694 );
and \U$12914 ( \14696 , \14676 , \14680 );
or \U$12917 ( \14697 , \14696 , 1'b0 , 1'b0 );
xor \U$12919 ( \14698 , \14697 , 1'b0 );
and \U$12920 ( \14699 , \14661 , \14670 );
xor \U$12921 ( \14700 , \14698 , \14699 );
xor \U$12922 ( \14701 , \14695 , \14700 );
and \U$12925 ( \14702 , \14636 , \14639 );
or \U$12926 ( \14703 , 1'b0 , 1'b0 , \14702 );
and \U$12927 ( \14704 , \14671 , 1'b1 );
and \U$12928 ( \14705 , 1'b1 , \14682 );
and \U$12929 ( \14706 , \14671 , \14682 );
or \U$12930 ( \14707 , \14704 , \14705 , \14706 );
xor \U$12931 ( \14708 , \14703 , \14707 );
and \U$12933 ( \14709 , \13396 , \13193 );
and \U$12934 ( \14710 , \13352 , \13191 );
nor \U$12935 ( \14711 , \14709 , \14710 );
xnor \U$12936 ( \14712 , \14711 , \13219 );
and \U$12938 ( \14713 , \13522 , \13246 );
nor \U$12939 ( \14714 , 1'b0 , \14713 );
xnor \U$12940 ( \14715 , \14714 , 1'b0 );
xor \U$12941 ( \14716 , \14712 , \14715 );
xor \U$12943 ( \14717 , \14716 , 1'b0 );
xor \U$12944 ( \14718 , 1'b0 , \14717 );
not \U$12945 ( \14719 , \13645 );
and \U$12946 ( \14720 , \13145 , \13320 );
and \U$12947 ( \14721 , \13214 , \13318 );
nor \U$12948 ( \14722 , \14720 , \14721 );
xnor \U$12949 ( \14723 , \14722 , \13325 );
xor \U$12950 ( \14724 , \14719 , \14723 );
and \U$12951 ( \14725 , \13373 , \13255 );
and \U$12952 ( \14726 , \13241 , \13253 );
nor \U$12953 ( \14727 , \14725 , \14726 );
xnor \U$12954 ( \14728 , \14727 , \13022 );
xor \U$12955 ( \14729 , \14724 , \14728 );
xor \U$12956 ( \14730 , \14718 , \14729 );
xor \U$12958 ( \14731 , \14730 , 1'b0 );
and \U$12960 ( \14732 , \14664 , \14669 );
or \U$12962 ( \14733 , 1'b0 , \14732 , 1'b0 );
and \U$12963 ( \14734 , \14652 , \14656 );
and \U$12964 ( \14735 , \14656 , \14660 );
and \U$12965 ( \14736 , \14652 , \14660 );
or \U$12966 ( \14737 , \14734 , \14735 , \14736 );
xor \U$12967 ( \14738 , \14733 , \14737 );
xor \U$12969 ( \14739 , \14738 , 1'b0 );
xor \U$12970 ( \14740 , \14731 , \14739 );
xor \U$12971 ( \14741 , \14708 , \14740 );
xor \U$12972 ( \14742 , \14701 , \14741 );
and \U$12973 ( \14743 , \14634 , \14640 );
and \U$12974 ( \14744 , \14640 , \14684 );
and \U$12975 ( \14745 , \14634 , \14684 );
or \U$12976 ( \14746 , \14743 , \14744 , \14745 );
nor \U$12977 ( \14747 , \14742 , \14746 );
and \U$12978 ( \14748 , \14703 , \14707 );
and \U$12979 ( \14749 , \14707 , \14740 );
and \U$12980 ( \14750 , \14703 , \14740 );
or \U$12981 ( \14751 , \14748 , \14749 , \14750 );
and \U$12982 ( \14752 , \14733 , \14737 );
or \U$12985 ( \14753 , \14752 , 1'b0 , 1'b0 );
xor \U$12987 ( \14754 , \14753 , 1'b0 );
and \U$12989 ( \14755 , \14717 , \14729 );
or \U$12991 ( \14756 , 1'b0 , \14755 , 1'b0 );
xor \U$12992 ( \14757 , \14754 , \14756 );
xor \U$12993 ( \14758 , \14751 , \14757 );
and \U$12996 ( \14759 , \14697 , \14699 );
or \U$12997 ( \14760 , 1'b0 , 1'b0 , \14759 );
and \U$13000 ( \14761 , \14730 , \14739 );
or \U$13001 ( \14762 , 1'b0 , 1'b0 , \14761 );
xor \U$13002 ( \14763 , \14760 , \14762 );
xor \U$13003 ( \14764 , \13376 , \13399 );
xor \U$13005 ( \14765 , \14764 , 1'b0 );
xor \U$13007 ( \14766 , 1'b0 , \13326 );
xor \U$13008 ( \14767 , \14766 , \13330 );
xor \U$13009 ( \14768 , \14765 , \14767 );
xor \U$13011 ( \14769 , \14768 , 1'b1 );
and \U$13012 ( \14770 , \14719 , \14723 );
and \U$13013 ( \14771 , \14723 , \14728 );
and \U$13014 ( \14772 , \14719 , \14728 );
or \U$13015 ( \14773 , \14770 , \14771 , \14772 );
and \U$13016 ( \14774 , \14712 , \14715 );
or \U$13019 ( \14775 , \14774 , 1'b0 , 1'b0 );
xor \U$13020 ( \14776 , \14773 , \14775 );
xor \U$13022 ( \14777 , \14776 , 1'b0 );
xor \U$13023 ( \14778 , \14769 , \14777 );
xor \U$13024 ( \14779 , \14763 , \14778 );
xor \U$13025 ( \14780 , \14758 , \14779 );
and \U$13026 ( \14781 , \14695 , \14700 );
and \U$13027 ( \14782 , \14700 , \14741 );
and \U$13028 ( \14783 , \14695 , \14741 );
or \U$13029 ( \14784 , \14781 , \14782 , \14783 );
nor \U$13030 ( \14785 , \14780 , \14784 );
nor \U$13031 ( \14786 , \14747 , \14785 );
nand \U$13032 ( \14787 , \14691 , \14786 );
and \U$13033 ( \14788 , \14760 , \14762 );
and \U$13034 ( \14789 , \14762 , \14778 );
and \U$13035 ( \14790 , \14760 , \14778 );
or \U$13036 ( \14791 , \14788 , \14789 , \14790 );
and \U$13037 ( \14792 , \14773 , \14775 );
or \U$13040 ( \14793 , \14792 , 1'b0 , 1'b0 );
xor \U$13042 ( \14794 , \14793 , 1'b0 );
and \U$13043 ( \14795 , \14765 , \14767 );
xor \U$13044 ( \14796 , \14794 , \14795 );
xor \U$13045 ( \14797 , \14791 , \14796 );
and \U$13048 ( \14798 , \14753 , \14756 );
or \U$13049 ( \14799 , 1'b0 , 1'b0 , \14798 );
and \U$13050 ( \14800 , \14768 , 1'b1 );
and \U$13051 ( \14801 , 1'b1 , \14777 );
and \U$13052 ( \14802 , \14768 , \14777 );
or \U$13053 ( \14803 , \14800 , \14801 , \14802 );
xor \U$13054 ( \14804 , \14799 , \14803 );
xor \U$13056 ( \14805 , 1'b0 , \13408 );
xor \U$13057 ( \14806 , \14805 , \13419 );
xor \U$13059 ( \14807 , \14806 , 1'b0 );
xor \U$13060 ( \14808 , \13332 , \13401 );
xor \U$13062 ( \14809 , \14808 , 1'b0 );
xor \U$13063 ( \14810 , \14807 , \14809 );
xor \U$13064 ( \14811 , \14804 , \14810 );
xor \U$13065 ( \14812 , \14797 , \14811 );
and \U$13066 ( \14813 , \14751 , \14757 );
and \U$13067 ( \14814 , \14757 , \14779 );
and \U$13068 ( \14815 , \14751 , \14779 );
or \U$13069 ( \14816 , \14813 , \14814 , \14815 );
nor \U$13070 ( \14817 , \14812 , \14816 );
and \U$13071 ( \14818 , \14799 , \14803 );
and \U$13072 ( \14819 , \14803 , \14810 );
and \U$13073 ( \14820 , \14799 , \14810 );
or \U$13074 ( \14821 , \14818 , \14819 , \14820 );
xor \U$13076 ( \14822 , \13403 , 1'b0 );
xor \U$13077 ( \14823 , \14822 , \13421 );
xor \U$13078 ( \14824 , \14821 , \14823 );
and \U$13081 ( \14825 , \14793 , \14795 );
or \U$13082 ( \14826 , 1'b0 , 1'b0 , \14825 );
and \U$13085 ( \14827 , \14806 , \14809 );
or \U$13086 ( \14828 , 1'b0 , 1'b0 , \14827 );
xor \U$13087 ( \14829 , \14826 , \14828 );
xor \U$13088 ( \14830 , \13431 , 1'b1 );
xor \U$13089 ( \14831 , \14830 , \13438 );
xor \U$13090 ( \14832 , \14829 , \14831 );
xor \U$13091 ( \14833 , \14824 , \14832 );
and \U$13092 ( \14834 , \14791 , \14796 );
and \U$13093 ( \14835 , \14796 , \14811 );
and \U$13094 ( \14836 , \14791 , \14811 );
or \U$13095 ( \14837 , \14834 , \14835 , \14836 );
nor \U$13096 ( \14838 , \14833 , \14837 );
nor \U$13097 ( \14839 , \14817 , \14838 );
and \U$13098 ( \14840 , \14826 , \14828 );
and \U$13099 ( \14841 , \14828 , \14831 );
and \U$13100 ( \14842 , \14826 , \14831 );
or \U$13101 ( \14843 , \14840 , \14841 , \14842 );
and \U$13103 ( \14844 , \13428 , \13430 );
xor \U$13104 ( \14845 , 1'b0 , \14844 );
xor \U$13105 ( \14846 , \14843 , \14845 );
xor \U$13106 ( \14847 , \13423 , \13441 );
xor \U$13107 ( \14848 , \14847 , \13444 );
xor \U$13108 ( \14849 , \14846 , \14848 );
and \U$13109 ( \14850 , \14821 , \14823 );
and \U$13110 ( \14851 , \14823 , \14832 );
and \U$13111 ( \14852 , \14821 , \14832 );
or \U$13112 ( \14853 , \14850 , \14851 , \14852 );
nor \U$13113 ( \14854 , \14849 , \14853 );
xor \U$13115 ( \14855 , \13447 , 1'b0 );
xor \U$13116 ( \14856 , \14855 , \13449 );
and \U$13117 ( \14857 , \14843 , \14845 );
and \U$13118 ( \14858 , \14845 , \14848 );
and \U$13119 ( \14859 , \14843 , \14848 );
or \U$13120 ( \14860 , \14857 , \14858 , \14859 );
nor \U$13121 ( \14861 , \14856 , \14860 );
nor \U$13122 ( \14862 , \14854 , \14861 );
nand \U$13123 ( \14863 , \14839 , \14862 );
nor \U$13124 ( \14864 , \14787 , \14863 );
nand \U$13125 ( \14865 , \14569 , \14864 );
and \U$13126 ( \14866 , \13666 , \13465 );
and \U$13127 ( \14867 , \13687 , \13462 );
nor \U$13128 ( \14868 , \14866 , \14867 );
xnor \U$13129 ( \14869 , \14868 , \13459 );
and \U$13130 ( \14870 , \13711 , \13501 );
and \U$13131 ( \14871 , \13732 , \13499 );
nor \U$13132 ( \14872 , \14870 , \14871 );
xnor \U$13133 ( \14873 , \14872 , \13527 );
and \U$13134 ( \14874 , \14869 , \14873 );
and \U$13135 ( \14875 , \13759 , \13561 );
and \U$13136 ( \14876 , \13780 , \13559 );
nor \U$13137 ( \14877 , \14875 , \14876 );
xnor \U$13138 ( \14878 , \14877 , \13587 );
and \U$13139 ( \14879 , \14873 , \14878 );
and \U$13140 ( \14880 , \14869 , \14878 );
or \U$13141 ( \14881 , \14874 , \14879 , \14880 );
and \U$13142 ( \14882 , \13780 , \13561 );
and \U$13143 ( \14883 , \13711 , \13559 );
nor \U$13144 ( \14884 , \14882 , \14883 );
xnor \U$13145 ( \14885 , \14884 , \13587 );
and \U$13146 ( \14886 , \13803 , \13619 );
and \U$13147 ( \14887 , \13759 , \13617 );
nor \U$13148 ( \14888 , \14886 , \14887 );
xnor \U$13149 ( \14889 , \14888 , \13645 );
xor \U$13150 ( \14890 , \14885 , \14889 );
nand \U$13151 ( \14891 , \13936 , \13318 );
xnor \U$13152 ( \14892 , \14891 , \13325 );
xor \U$13153 ( \14893 , \14890 , \14892 );
and \U$13154 ( \14894 , \14881 , \14893 );
and \U$13155 ( \14895 , \13687 , \13465 );
and \U$13156 ( \14896 , \13611 , \13462 );
nor \U$13157 ( \14897 , \14895 , \14896 );
xnor \U$13158 ( \14898 , \14897 , \13459 );
xor \U$13159 ( \14899 , \13325 , \14898 );
and \U$13160 ( \14900 , \13732 , \13501 );
and \U$13161 ( \14901 , \13666 , \13499 );
nor \U$13162 ( \14902 , \14900 , \14901 );
xnor \U$13163 ( \14903 , \14902 , \13527 );
xor \U$13164 ( \14904 , \14899 , \14903 );
and \U$13165 ( \14905 , \14893 , \14904 );
and \U$13166 ( \14906 , \14881 , \14904 );
or \U$13167 ( \14907 , \14894 , \14905 , \14906 );
and \U$13168 ( \14908 , \13936 , \13320 );
and \U$13169 ( \14909 , \13803 , \13318 );
nor \U$13170 ( \14910 , \14908 , \14909 );
xnor \U$13171 ( \14911 , \14910 , \13325 );
and \U$13172 ( \14912 , \13611 , \13465 );
and \U$13173 ( \14913 , \13640 , \13462 );
nor \U$13174 ( \14914 , \14912 , \14913 );
xnor \U$13175 ( \14915 , \14914 , \13459 );
and \U$13176 ( \14916 , \13666 , \13501 );
and \U$13177 ( \14917 , \13687 , \13499 );
nor \U$13178 ( \14918 , \14916 , \14917 );
xnor \U$13179 ( \14919 , \14918 , \13527 );
xor \U$13180 ( \14920 , \14915 , \14919 );
and \U$13181 ( \14921 , \13711 , \13561 );
and \U$13182 ( \14922 , \13732 , \13559 );
nor \U$13183 ( \14923 , \14921 , \14922 );
xnor \U$13184 ( \14924 , \14923 , \13587 );
xor \U$13185 ( \14925 , \14920 , \14924 );
xor \U$13186 ( \14926 , \14911 , \14925 );
xor \U$13187 ( \14927 , \14907 , \14926 );
and \U$13188 ( \14928 , \13325 , \14898 );
and \U$13189 ( \14929 , \14898 , \14903 );
and \U$13190 ( \14930 , \13325 , \14903 );
or \U$13191 ( \14931 , \14928 , \14929 , \14930 );
and \U$13192 ( \14932 , \14885 , \14889 );
and \U$13193 ( \14933 , \14889 , \14892 );
and \U$13194 ( \14934 , \14885 , \14892 );
or \U$13195 ( \14935 , \14932 , \14933 , \14934 );
xor \U$13196 ( \14936 , \14931 , \14935 );
and \U$13197 ( \14937 , \13759 , \13619 );
and \U$13198 ( \14938 , \13780 , \13617 );
nor \U$13199 ( \14939 , \14937 , \14938 );
xnor \U$13200 ( \14940 , \14939 , \13645 );
xor \U$13201 ( \14941 , \14936 , \14940 );
xor \U$13202 ( \14942 , \14927 , \14941 );
and \U$13203 ( \14943 , \13732 , \13465 );
and \U$13204 ( \14944 , \13666 , \13462 );
nor \U$13205 ( \14945 , \14943 , \14944 );
xnor \U$13206 ( \14946 , \14945 , \13459 );
and \U$13207 ( \14947 , \13645 , \14946 );
and \U$13208 ( \14948 , \13780 , \13501 );
and \U$13209 ( \14949 , \13711 , \13499 );
nor \U$13210 ( \14950 , \14948 , \14949 );
xnor \U$13211 ( \14951 , \14950 , \13527 );
and \U$13212 ( \14952 , \14946 , \14951 );
and \U$13213 ( \14953 , \13645 , \14951 );
or \U$13214 ( \14954 , \14947 , \14952 , \14953 );
and \U$13215 ( \14955 , \13803 , \13561 );
and \U$13216 ( \14956 , \13759 , \13559 );
nor \U$13217 ( \14957 , \14955 , \14956 );
xnor \U$13218 ( \14958 , \14957 , \13587 );
nand \U$13219 ( \14959 , \13936 , \13617 );
xnor \U$13220 ( \14960 , \14959 , \13645 );
and \U$13221 ( \14961 , \14958 , \14960 );
and \U$13222 ( \14962 , \14954 , \14961 );
and \U$13223 ( \14963 , \13936 , \13619 );
and \U$13224 ( \14964 , \13803 , \13617 );
nor \U$13225 ( \14965 , \14963 , \14964 );
xnor \U$13226 ( \14966 , \14965 , \13645 );
and \U$13227 ( \14967 , \14961 , \14966 );
and \U$13228 ( \14968 , \14954 , \14966 );
or \U$13229 ( \14969 , \14962 , \14967 , \14968 );
xor \U$13230 ( \14970 , \14881 , \14893 );
xor \U$13231 ( \14971 , \14970 , \14904 );
and \U$13232 ( \14972 , \14969 , \14971 );
nor \U$13233 ( \14973 , \14942 , \14972 );
and \U$13234 ( \14974 , \14915 , \14919 );
and \U$13235 ( \14975 , \14919 , \14924 );
and \U$13236 ( \14976 , \14915 , \14924 );
or \U$13237 ( \14977 , \14974 , \14975 , \14976 );
nand \U$13238 ( \14978 , \13936 , \13253 );
xnor \U$13239 ( \14979 , \14978 , \13022 );
xor \U$13240 ( \14980 , \14977 , \14979 );
and \U$13241 ( \14981 , \13732 , \13561 );
and \U$13242 ( \14982 , \13666 , \13559 );
nor \U$13243 ( \14983 , \14981 , \14982 );
xnor \U$13244 ( \14984 , \14983 , \13587 );
and \U$13245 ( \14985 , \13780 , \13619 );
and \U$13246 ( \14986 , \13711 , \13617 );
nor \U$13247 ( \14987 , \14985 , \14986 );
xnor \U$13248 ( \14988 , \14987 , \13645 );
xor \U$13249 ( \14989 , \14984 , \14988 );
and \U$13250 ( \14990 , \13803 , \13320 );
and \U$13251 ( \14991 , \13759 , \13318 );
nor \U$13252 ( \14992 , \14990 , \14991 );
xnor \U$13253 ( \14993 , \14992 , \13325 );
xor \U$13254 ( \14994 , \14989 , \14993 );
xor \U$13255 ( \14995 , \14980 , \14994 );
and \U$13256 ( \14996 , \14931 , \14935 );
and \U$13257 ( \14997 , \14935 , \14940 );
and \U$13258 ( \14998 , \14931 , \14940 );
or \U$13259 ( \14999 , \14996 , \14997 , \14998 );
and \U$13260 ( \15000 , \14911 , \14925 );
xor \U$13261 ( \15001 , \14999 , \15000 );
and \U$13262 ( \15002 , \13640 , \13465 );
and \U$13263 ( \15003 , \13549 , \13462 );
nor \U$13264 ( \15004 , \15002 , \15003 );
xnor \U$13265 ( \15005 , \15004 , \13459 );
xor \U$13266 ( \15006 , \13022 , \15005 );
and \U$13267 ( \15007 , \13687 , \13501 );
and \U$13268 ( \15008 , \13611 , \13499 );
nor \U$13269 ( \15009 , \15007 , \15008 );
xnor \U$13270 ( \15010 , \15009 , \13527 );
xor \U$13271 ( \15011 , \15006 , \15010 );
xor \U$13272 ( \15012 , \15001 , \15011 );
xor \U$13273 ( \15013 , \14995 , \15012 );
and \U$13274 ( \15014 , \14907 , \14926 );
and \U$13275 ( \15015 , \14926 , \14941 );
and \U$13276 ( \15016 , \14907 , \14941 );
or \U$13277 ( \15017 , \15014 , \15015 , \15016 );
nor \U$13278 ( \15018 , \15013 , \15017 );
nor \U$13279 ( \15019 , \14973 , \15018 );
and \U$13280 ( \15020 , \14999 , \15000 );
and \U$13281 ( \15021 , \15000 , \15011 );
and \U$13282 ( \15022 , \14999 , \15011 );
or \U$13283 ( \15023 , \15020 , \15021 , \15022 );
and \U$13284 ( \15024 , \14977 , \14979 );
and \U$13285 ( \15025 , \14979 , \14994 );
and \U$13286 ( \15026 , \14977 , \14994 );
or \U$13287 ( \15027 , \15024 , \15025 , \15026 );
and \U$13288 ( \15028 , \13549 , \13465 );
and \U$13289 ( \15029 , \13582 , \13462 );
nor \U$13290 ( \15030 , \15028 , \15029 );
xnor \U$13291 ( \15031 , \15030 , \13459 );
and \U$13292 ( \15032 , \13611 , \13501 );
and \U$13293 ( \15033 , \13640 , \13499 );
nor \U$13294 ( \15034 , \15032 , \15033 );
xnor \U$13295 ( \15035 , \15034 , \13527 );
xor \U$13296 ( \15036 , \15031 , \15035 );
and \U$13297 ( \15037 , \13666 , \13561 );
and \U$13298 ( \15038 , \13687 , \13559 );
nor \U$13299 ( \15039 , \15037 , \15038 );
xnor \U$13300 ( \15040 , \15039 , \13587 );
xor \U$13301 ( \15041 , \15036 , \15040 );
xor \U$13302 ( \15042 , \15027 , \15041 );
and \U$13303 ( \15043 , \13022 , \15005 );
and \U$13304 ( \15044 , \15005 , \15010 );
and \U$13305 ( \15045 , \13022 , \15010 );
or \U$13306 ( \15046 , \15043 , \15044 , \15045 );
and \U$13307 ( \15047 , \14984 , \14988 );
and \U$13308 ( \15048 , \14988 , \14993 );
and \U$13309 ( \15049 , \14984 , \14993 );
or \U$13310 ( \15050 , \15047 , \15048 , \15049 );
xor \U$13311 ( \15051 , \15046 , \15050 );
and \U$13312 ( \15052 , \13711 , \13619 );
and \U$13313 ( \15053 , \13732 , \13617 );
nor \U$13314 ( \15054 , \15052 , \15053 );
xnor \U$13315 ( \15055 , \15054 , \13645 );
and \U$13316 ( \15056 , \13759 , \13320 );
and \U$13317 ( \15057 , \13780 , \13318 );
nor \U$13318 ( \15058 , \15056 , \15057 );
xnor \U$13319 ( \15059 , \15058 , \13325 );
xor \U$13320 ( \15060 , \15055 , \15059 );
and \U$13321 ( \15061 , \13936 , \13255 );
and \U$13322 ( \15062 , \13803 , \13253 );
nor \U$13323 ( \15063 , \15061 , \15062 );
xnor \U$13324 ( \15064 , \15063 , \13022 );
xor \U$13325 ( \15065 , \15060 , \15064 );
xor \U$13326 ( \15066 , \15051 , \15065 );
xor \U$13327 ( \15067 , \15042 , \15066 );
xor \U$13328 ( \15068 , \15023 , \15067 );
and \U$13329 ( \15069 , \14995 , \15012 );
nor \U$13330 ( \15070 , \15068 , \15069 );
and \U$13331 ( \15071 , \15027 , \15041 );
and \U$13332 ( \15072 , \15041 , \15066 );
and \U$13333 ( \15073 , \15027 , \15066 );
or \U$13334 ( \15074 , \15071 , \15072 , \15073 );
and \U$13335 ( \15075 , \15046 , \15050 );
and \U$13336 ( \15076 , \15050 , \15065 );
and \U$13337 ( \15077 , \15046 , \15065 );
or \U$13338 ( \15078 , \15075 , \15076 , \15077 );
nand \U$13339 ( \15079 , \13936 , \13191 );
xnor \U$13340 ( \15080 , \15079 , \13219 );
and \U$13341 ( \15081 , \13687 , \13561 );
and \U$13342 ( \15082 , \13611 , \13559 );
nor \U$13343 ( \15083 , \15081 , \15082 );
xnor \U$13344 ( \15084 , \15083 , \13587 );
and \U$13345 ( \15085 , \13732 , \13619 );
and \U$13346 ( \15086 , \13666 , \13617 );
nor \U$13347 ( \15087 , \15085 , \15086 );
xnor \U$13348 ( \15088 , \15087 , \13645 );
xor \U$13349 ( \15089 , \15084 , \15088 );
and \U$13350 ( \15090 , \13780 , \13320 );
and \U$13351 ( \15091 , \13711 , \13318 );
nor \U$13352 ( \15092 , \15090 , \15091 );
xnor \U$13353 ( \15093 , \15092 , \13325 );
xor \U$13354 ( \15094 , \15089 , \15093 );
xor \U$13355 ( \15095 , \15080 , \15094 );
and \U$13356 ( \15096 , \13582 , \13465 );
and \U$13357 ( \15097 , \13489 , \13462 );
nor \U$13358 ( \15098 , \15096 , \15097 );
xnor \U$13359 ( \15099 , \15098 , \13459 );
xor \U$13360 ( \15100 , \13219 , \15099 );
and \U$13361 ( \15101 , \13640 , \13501 );
and \U$13362 ( \15102 , \13549 , \13499 );
nor \U$13363 ( \15103 , \15101 , \15102 );
xnor \U$13364 ( \15104 , \15103 , \13527 );
xor \U$13365 ( \15105 , \15100 , \15104 );
xor \U$13366 ( \15106 , \15095 , \15105 );
xor \U$13367 ( \15107 , \15078 , \15106 );
and \U$13368 ( \15108 , \15031 , \15035 );
and \U$13369 ( \15109 , \15035 , \15040 );
and \U$13370 ( \15110 , \15031 , \15040 );
or \U$13371 ( \15111 , \15108 , \15109 , \15110 );
and \U$13372 ( \15112 , \15055 , \15059 );
and \U$13373 ( \15113 , \15059 , \15064 );
and \U$13374 ( \15114 , \15055 , \15064 );
or \U$13375 ( \15115 , \15112 , \15113 , \15114 );
xor \U$13376 ( \15116 , \15111 , \15115 );
and \U$13377 ( \15117 , \13803 , \13255 );
and \U$13378 ( \15118 , \13759 , \13253 );
nor \U$13379 ( \15119 , \15117 , \15118 );
xnor \U$13380 ( \15120 , \15119 , \13022 );
xor \U$13381 ( \15121 , \15116 , \15120 );
xor \U$13382 ( \15122 , \15107 , \15121 );
xor \U$13383 ( \15123 , \15074 , \15122 );
and \U$13384 ( \15124 , \15023 , \15067 );
nor \U$13385 ( \15125 , \15123 , \15124 );
nor \U$13386 ( \15126 , \15070 , \15125 );
nand \U$13387 ( \15127 , \15019 , \15126 );
and \U$13388 ( \15128 , \15078 , \15106 );
and \U$13389 ( \15129 , \15106 , \15121 );
and \U$13390 ( \15130 , \15078 , \15121 );
or \U$13391 ( \15131 , \15128 , \15129 , \15130 );
xor \U$13392 ( \15132 , \13991 , \13995 );
xor \U$13393 ( \15133 , \15132 , \14000 );
and \U$13394 ( \15134 , \13219 , \15099 );
and \U$13395 ( \15135 , \15099 , \15104 );
and \U$13396 ( \15136 , \13219 , \15104 );
or \U$13397 ( \15137 , \15134 , \15135 , \15136 );
and \U$13398 ( \15138 , \15084 , \15088 );
and \U$13399 ( \15139 , \15088 , \15093 );
and \U$13400 ( \15140 , \15084 , \15093 );
or \U$13401 ( \15141 , \15138 , \15139 , \15140 );
xor \U$13402 ( \15142 , \15137 , \15141 );
and \U$13403 ( \15143 , \13936 , \13193 );
and \U$13404 ( \15144 , \13803 , \13191 );
nor \U$13405 ( \15145 , \15143 , \15144 );
xnor \U$13406 ( \15146 , \15145 , \13219 );
xor \U$13407 ( \15147 , \15142 , \15146 );
xor \U$13408 ( \15148 , \15133 , \15147 );
xor \U$13409 ( \15149 , \15131 , \15148 );
and \U$13410 ( \15150 , \15111 , \15115 );
and \U$13411 ( \15151 , \15115 , \15120 );
and \U$13412 ( \15152 , \15111 , \15120 );
or \U$13413 ( \15153 , \15150 , \15151 , \15152 );
and \U$13414 ( \15154 , \15080 , \15094 );
and \U$13415 ( \15155 , \15094 , \15105 );
and \U$13416 ( \15156 , \15080 , \15105 );
or \U$13417 ( \15157 , \15154 , \15155 , \15156 );
xor \U$13418 ( \15158 , \15153 , \15157 );
xor \U$13419 ( \15159 , \14007 , \14011 );
xor \U$13420 ( \15160 , \15159 , \14016 );
xor \U$13421 ( \15161 , \15158 , \15160 );
xor \U$13422 ( \15162 , \15149 , \15161 );
and \U$13423 ( \15163 , \15074 , \15122 );
nor \U$13424 ( \15164 , \15162 , \15163 );
and \U$13425 ( \15165 , \15153 , \15157 );
and \U$13426 ( \15166 , \15157 , \15160 );
and \U$13427 ( \15167 , \15153 , \15160 );
or \U$13428 ( \15168 , \15165 , \15166 , \15167 );
and \U$13429 ( \15169 , \15133 , \15147 );
xor \U$13430 ( \15170 , \15168 , \15169 );
and \U$13431 ( \15171 , \15137 , \15141 );
and \U$13432 ( \15172 , \15141 , \15146 );
and \U$13433 ( \15173 , \15137 , \15146 );
or \U$13434 ( \15174 , \15171 , \15172 , \15173 );
xor \U$13435 ( \15175 , \14027 , \14029 );
xor \U$13436 ( \15176 , \15174 , \15175 );
xor \U$13437 ( \15177 , \14003 , \14019 );
xor \U$13438 ( \15178 , \15177 , \14022 );
xor \U$13439 ( \15179 , \15176 , \15178 );
xor \U$13440 ( \15180 , \15170 , \15179 );
and \U$13441 ( \15181 , \15131 , \15148 );
and \U$13442 ( \15182 , \15148 , \15161 );
and \U$13443 ( \15183 , \15131 , \15161 );
or \U$13444 ( \15184 , \15181 , \15182 , \15183 );
nor \U$13445 ( \15185 , \15180 , \15184 );
nor \U$13446 ( \15186 , \15164 , \15185 );
and \U$13447 ( \15187 , \15174 , \15175 );
and \U$13448 ( \15188 , \15175 , \15178 );
and \U$13449 ( \15189 , \15174 , \15178 );
or \U$13450 ( \15190 , \15187 , \15188 , \15189 );
xor \U$13451 ( \15191 , \13890 , \13906 );
xor \U$13452 ( \15192 , \15191 , \13941 );
xor \U$13453 ( \15193 , \15190 , \15192 );
xor \U$13454 ( \15194 , \14025 , \14030 );
xor \U$13455 ( \15195 , \15194 , \14033 );
xor \U$13456 ( \15196 , \15193 , \15195 );
and \U$13457 ( \15197 , \15168 , \15169 );
and \U$13458 ( \15198 , \15169 , \15179 );
and \U$13459 ( \15199 , \15168 , \15179 );
or \U$13460 ( \15200 , \15197 , \15198 , \15199 );
nor \U$13461 ( \15201 , \15196 , \15200 );
xor \U$13462 ( \15202 , \14036 , \14037 );
xor \U$13463 ( \15203 , \15202 , \14040 );
and \U$13464 ( \15204 , \15190 , \15192 );
and \U$13465 ( \15205 , \15192 , \15195 );
and \U$13466 ( \15206 , \15190 , \15195 );
or \U$13467 ( \15207 , \15204 , \15205 , \15206 );
nor \U$13468 ( \15208 , \15203 , \15207 );
nor \U$13469 ( \15209 , \15201 , \15208 );
nand \U$13470 ( \15210 , \15186 , \15209 );
nor \U$13471 ( \15211 , \15127 , \15210 );
and \U$13472 ( \15212 , \13780 , \13465 );
and \U$13473 ( \15213 , \13711 , \13462 );
nor \U$13474 ( \15214 , \15212 , \15213 );
xnor \U$13475 ( \15215 , \15214 , \13459 );
and \U$13476 ( \15216 , \13587 , \15215 );
and \U$13477 ( \15217 , \13803 , \13501 );
and \U$13478 ( \15218 , \13759 , \13499 );
nor \U$13479 ( \15219 , \15217 , \15218 );
xnor \U$13480 ( \15220 , \15219 , \13527 );
and \U$13481 ( \15221 , \15215 , \15220 );
and \U$13482 ( \15222 , \13587 , \15220 );
or \U$13483 ( \15223 , \15216 , \15221 , \15222 );
and \U$13484 ( \15224 , \13711 , \13465 );
and \U$13485 ( \15225 , \13732 , \13462 );
nor \U$13486 ( \15226 , \15224 , \15225 );
xnor \U$13487 ( \15227 , \15226 , \13459 );
and \U$13488 ( \15228 , \13759 , \13501 );
and \U$13489 ( \15229 , \13780 , \13499 );
nor \U$13490 ( \15230 , \15228 , \15229 );
xnor \U$13491 ( \15231 , \15230 , \13527 );
xor \U$13492 ( \15232 , \15227 , \15231 );
and \U$13493 ( \15233 , \13936 , \13561 );
and \U$13494 ( \15234 , \13803 , \13559 );
nor \U$13495 ( \15235 , \15233 , \15234 );
xnor \U$13496 ( \15236 , \15235 , \13587 );
xor \U$13497 ( \15237 , \15232 , \15236 );
xor \U$13498 ( \15238 , \15223 , \15237 );
nand \U$13499 ( \15239 , \13936 , \13559 );
xnor \U$13500 ( \15240 , \15239 , \13587 );
xor \U$13501 ( \15241 , \13587 , \15215 );
xor \U$13502 ( \15242 , \15241 , \15220 );
and \U$13503 ( \15243 , \15240 , \15242 );
nor \U$13504 ( \15244 , \15238 , \15243 );
and \U$13505 ( \15245 , \15227 , \15231 );
and \U$13506 ( \15246 , \15231 , \15236 );
and \U$13507 ( \15247 , \15227 , \15236 );
or \U$13508 ( \15248 , \15245 , \15246 , \15247 );
xor \U$13509 ( \15249 , \14958 , \14960 );
xor \U$13510 ( \15250 , \15248 , \15249 );
xor \U$13511 ( \15251 , \13645 , \14946 );
xor \U$13512 ( \15252 , \15251 , \14951 );
xor \U$13513 ( \15253 , \15250 , \15252 );
and \U$13514 ( \15254 , \15223 , \15237 );
nor \U$13515 ( \15255 , \15253 , \15254 );
nor \U$13516 ( \15256 , \15244 , \15255 );
xor \U$13517 ( \15257 , \14869 , \14873 );
xor \U$13518 ( \15258 , \15257 , \14878 );
xor \U$13519 ( \15259 , \14954 , \14961 );
xor \U$13520 ( \15260 , \15259 , \14966 );
xor \U$13521 ( \15261 , \15258 , \15260 );
and \U$13522 ( \15262 , \15248 , \15249 );
and \U$13523 ( \15263 , \15249 , \15252 );
and \U$13524 ( \15264 , \15248 , \15252 );
or \U$13525 ( \15265 , \15262 , \15263 , \15264 );
nor \U$13526 ( \15266 , \15261 , \15265 );
xor \U$13527 ( \15267 , \14969 , \14971 );
and \U$13528 ( \15268 , \15258 , \15260 );
nor \U$13529 ( \15269 , \15267 , \15268 );
nor \U$13530 ( \15270 , \15266 , \15269 );
nand \U$13531 ( \15271 , \15256 , \15270 );
and \U$13532 ( \15272 , \13759 , \13465 );
and \U$13533 ( \15273 , \13780 , \13462 );
nor \U$13534 ( \15274 , \15272 , \15273 );
xnor \U$13535 ( \15275 , \15274 , \13459 );
and \U$13536 ( \15276 , \13936 , \13501 );
and \U$13537 ( \15277 , \13803 , \13499 );
nor \U$13538 ( \15278 , \15276 , \15277 );
xnor \U$13539 ( \15279 , \15278 , \13527 );
xor \U$13540 ( \15280 , \15275 , \15279 );
and \U$13541 ( \15281 , \13803 , \13465 );
and \U$13542 ( \15282 , \13759 , \13462 );
nor \U$13543 ( \15283 , \15281 , \15282 );
xnor \U$13544 ( \15284 , \15283 , \13459 );
and \U$13545 ( \15285 , \15284 , \13527 );
nor \U$13546 ( \15286 , \15280 , \15285 );
xor \U$13547 ( \15287 , \15240 , \15242 );
and \U$13548 ( \15288 , \15275 , \15279 );
nor \U$13549 ( \15289 , \15287 , \15288 );
nor \U$13550 ( \15290 , \15286 , \15289 );
xor \U$13551 ( \15291 , \15284 , \13527 );
nand \U$13552 ( \15292 , \13936 , \13499 );
xnor \U$13553 ( \15293 , \15292 , \13527 );
nor \U$13554 ( \15294 , \15291 , \15293 );
and \U$13555 ( \15295 , \13936 , \13465 );
and \U$13556 ( \15296 , \13803 , \13462 );
nor \U$13557 ( \15297 , \15295 , \15296 );
xnor \U$13558 ( \15298 , \15297 , \13459 );
nand \U$13559 ( \15299 , \13936 , \13462 );
xnor \U$13560 ( \15300 , \15299 , \13459 );
and \U$13561 ( \15301 , \15300 , \13459 );
nand \U$13562 ( \15302 , \15298 , \15301 );
or \U$13563 ( \15303 , \15294 , \15302 );
nand \U$13564 ( \15304 , \15291 , \15293 );
nand \U$13565 ( \15305 , \15303 , \15304 );
and \U$13566 ( \15306 , \15290 , \15305 );
nand \U$13567 ( \15307 , \15280 , \15285 );
or \U$13568 ( \15308 , \15289 , \15307 );
nand \U$13569 ( \15309 , \15287 , \15288 );
nand \U$13570 ( \15310 , \15308 , \15309 );
nor \U$13571 ( \15311 , \15306 , \15310 );
or \U$13572 ( \15312 , \15271 , \15311 );
nand \U$13573 ( \15313 , \15238 , \15243 );
or \U$13574 ( \15314 , \15255 , \15313 );
nand \U$13575 ( \15315 , \15253 , \15254 );
nand \U$13576 ( \15316 , \15314 , \15315 );
and \U$13577 ( \15317 , \15270 , \15316 );
nand \U$13578 ( \15318 , \15261 , \15265 );
or \U$13579 ( \15319 , \15269 , \15318 );
nand \U$13580 ( \15320 , \15267 , \15268 );
nand \U$13581 ( \15321 , \15319 , \15320 );
nor \U$13582 ( \15322 , \15317 , \15321 );
nand \U$13583 ( \15323 , \15312 , \15322 );
and \U$13584 ( \15324 , \15211 , \15323 );
nand \U$13585 ( \15325 , \14942 , \14972 );
or \U$13586 ( \15326 , \15018 , \15325 );
nand \U$13587 ( \15327 , \15013 , \15017 );
nand \U$13588 ( \15328 , \15326 , \15327 );
and \U$13589 ( \15329 , \15126 , \15328 );
nand \U$13590 ( \15330 , \15068 , \15069 );
or \U$13591 ( \15331 , \15125 , \15330 );
nand \U$13592 ( \15332 , \15123 , \15124 );
nand \U$13593 ( \15333 , \15331 , \15332 );
nor \U$13594 ( \15334 , \15329 , \15333 );
or \U$13595 ( \15335 , \15210 , \15334 );
nand \U$13596 ( \15336 , \15162 , \15163 );
or \U$13597 ( \15337 , \15185 , \15336 );
nand \U$13598 ( \15338 , \15180 , \15184 );
nand \U$13599 ( \15339 , \15337 , \15338 );
and \U$13600 ( \15340 , \15209 , \15339 );
nand \U$13601 ( \15341 , \15196 , \15200 );
or \U$13602 ( \15342 , \15208 , \15341 );
nand \U$13603 ( \15343 , \15203 , \15207 );
nand \U$13604 ( \15344 , \15342 , \15343 );
nor \U$13605 ( \15345 , \15340 , \15344 );
nand \U$13606 ( \15346 , \15335 , \15345 );
nor \U$13607 ( \15347 , \15324 , \15346 );
or \U$13608 ( \15348 , \14865 , \15347 );
nand \U$13609 ( \15349 , \13987 , \14043 );
or \U$13610 ( \15350 , \14119 , \15349 );
nand \U$13611 ( \15351 , \14117 , \14118 );
nand \U$13612 ( \15352 , \15350 , \15351 );
and \U$13613 ( \15353 , \14272 , \15352 );
nand \U$13614 ( \15354 , \14194 , \14195 );
or \U$13615 ( \15355 , \14271 , \15354 );
nand \U$13616 ( \15356 , \14266 , \14270 );
nand \U$13617 ( \15357 , \15355 , \15356 );
nor \U$13618 ( \15358 , \15353 , \15357 );
or \U$13619 ( \15359 , \14568 , \15358 );
nand \U$13620 ( \15360 , \14343 , \14347 );
or \U$13621 ( \15361 , \14424 , \15360 );
nand \U$13622 ( \15362 , \14419 , \14423 );
nand \U$13623 ( \15363 , \15361 , \15362 );
and \U$13624 ( \15364 , \14567 , \15363 );
nand \U$13625 ( \15365 , \14492 , \14496 );
or \U$13626 ( \15366 , \14566 , \15365 );
nand \U$13627 ( \15367 , \14561 , \14565 );
nand \U$13628 ( \15368 , \15366 , \15367 );
nor \U$13629 ( \15369 , \15364 , \15368 );
nand \U$13630 ( \15370 , \15359 , \15369 );
and \U$13631 ( \15371 , \14864 , \15370 );
nand \U$13632 ( \15372 , \14625 , \14629 );
or \U$13633 ( \15373 , \14690 , \15372 );
nand \U$13634 ( \15374 , \14685 , \14689 );
nand \U$13635 ( \15375 , \15373 , \15374 );
and \U$13636 ( \15376 , \14786 , \15375 );
nand \U$13637 ( \15377 , \14742 , \14746 );
or \U$13638 ( \15378 , \14785 , \15377 );
nand \U$13639 ( \15379 , \14780 , \14784 );
nand \U$13640 ( \15380 , \15378 , \15379 );
nor \U$13641 ( \15381 , \15376 , \15380 );
or \U$13642 ( \15382 , \14863 , \15381 );
nand \U$13643 ( \15383 , \14812 , \14816 );
or \U$13644 ( \15384 , \14838 , \15383 );
nand \U$13645 ( \15385 , \14833 , \14837 );
nand \U$13646 ( \15386 , \15384 , \15385 );
and \U$13647 ( \15387 , \14862 , \15386 );
nand \U$13648 ( \15388 , \14849 , \14853 );
or \U$13649 ( \15389 , \14861 , \15388 );
nand \U$13650 ( \15390 , \14856 , \14860 );
nand \U$13651 ( \15391 , \15389 , \15390 );
nor \U$13652 ( \15392 , \15387 , \15391 );
nand \U$13653 ( \15393 , \15382 , \15392 );
nor \U$13654 ( \15394 , \15371 , \15393 );
nand \U$13655 ( \15395 , \15348 , \15394 );
not \U$13656 ( \15396 , \15395 );
xor \U$13657 ( \15397 , \13455 , \15396 );
buf g4ba0_GF_PartitionCandidate( \15398_nG4ba0 , \15397 );
buf \U$13658 ( \15399 , RI2b5e785db0d0_14);
buf \U$13659 ( \15400 , RI2b5e785db058_15);
buf \U$13660 ( \15401 , RI2b5e785dafe0_16);
buf \U$13661 ( \15402 , RI2b5e785daf68_17);
buf \U$13662 ( \15403 , RI2b5e785daef0_18);
buf \U$13663 ( \15404 , RI2b5e785dae78_19);
buf \U$13664 ( \15405 , RI2b5e785dae00_20);
buf \U$13665 ( \15406 , RI2b5e785dad88_21);
buf \U$13666 ( \15407 , RI2b5e785dad10_22);
buf \U$13667 ( \15408 , RI2b5e785dac98_23);
buf \U$13668 ( \15409 , RI2b5e785dac20_24);
buf \U$13669 ( \15410 , RI2b5e785daba8_25);
not \U$13670 ( \15411 , RI2b5e785ae328_614);
buf \U$13671 ( \15412 , \15411 );
and \U$13672 ( \15413 , \15410 , \15412 );
and \U$13673 ( \15414 , \15409 , \15413 );
and \U$13674 ( \15415 , \15408 , \15414 );
and \U$13675 ( \15416 , \15407 , \15415 );
and \U$13676 ( \15417 , \15406 , \15416 );
and \U$13677 ( \15418 , \15405 , \15417 );
and \U$13678 ( \15419 , \15404 , \15418 );
and \U$13679 ( \15420 , \15403 , \15419 );
and \U$13680 ( \15421 , \15402 , \15420 );
and \U$13681 ( \15422 , \15401 , \15421 );
and \U$13682 ( \15423 , \15400 , \15422 );
xor \U$13683 ( \15424 , \15399 , \15423 );
buf \U$13684 ( \15425 , \15424 );
buf \U$13685 ( \15426 , \15425 );
not \U$13686 ( \15427 , \15426 );
nor \U$13687 ( \15428 , \12595 , \12599 , \12603 , \12607 , \12612 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13688 ( \15429 , RI2b5e785daab8_27, \15428 );
nor \U$13689 ( \15430 , \12647 , \12648 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13690 ( \15431 , RI2b5e785495b8_40, \15430 );
nor \U$13691 ( \15432 , \12595 , \12648 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13692 ( \15433 , RI2b5e78538920_53, \15432 );
nor \U$13693 ( \15434 , \12647 , \12599 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13694 ( \15435 , RI2b5e784a63a8_66, \15434 );
nor \U$13695 ( \15436 , \12595 , \12599 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13696 ( \15437 , RI2b5e78495710_79, \15436 );
nor \U$13697 ( \15438 , \12647 , \12648 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13698 ( \15439 , RI2b5e784950f8_92, \15438 );
nor \U$13699 ( \15440 , \12595 , \12648 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13700 ( \15441 , RI2b5e78403bf8_105, \15440 );
nor \U$13701 ( \15442 , \12647 , \12599 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13702 ( \15443 , RI2b5e775b1ed8_118, \15442 );
nor \U$13703 ( \15444 , \12595 , \12599 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13704 ( \15445 , RI2b5e775b18c0_131, \15444 );
nor \U$13705 ( \15446 , \12647 , \12648 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13706 ( \15447 , RI2b5e7750b858_144, \15446 );
nor \U$13707 ( \15448 , \12595 , \12648 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13708 ( \15449 , RI2b5e774ff030_157, \15448 );
nor \U$13709 ( \15450 , \12647 , \12599 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13710 ( \15451 , RI2b5e774f6048_170, \15450 );
nor \U$13711 ( \15452 , \12595 , \12599 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13712 ( \15453 , RI2b5e774ea630_183, \15452 );
nor \U$13713 ( \15454 , \12647 , \12648 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13714 ( \15455 , RI2b5e774dde08_196, \15454 );
nor \U$13715 ( \15456 , \12595 , \12648 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13716 ( \15457 , RI2b5e774d4e20_209, \15456 );
nor \U$13717 ( \15458 , \12647 , \12599 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13718 ( \15459 , RI2b5e785f3d60_222, \15458 );
nor \U$13719 ( \15460 , \12595 , \12599 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$13720 ( \15461 , RI2b5e785eb138_235, \15460 );
or \U$13721 ( \15462 , \15429 , \15431 , \15433 , \15435 , \15437 , \15439 , \15441 , \15443 , \15445 , \15447 , \15449 , \15451 , \15453 , \15455 , \15457 , \15459 , \15461 );
buf \U$13722 ( \15463 , \12616 );
buf \U$13723 ( \15464 , \12620 );
buf \U$13724 ( \15465 , \12624 );
buf \U$13725 ( \15466 , \12628 );
buf \U$13726 ( \15467 , \12632 );
buf \U$13727 ( \15468 , \12636 );
buf \U$13728 ( \15469 , \12640 );
buf \U$13729 ( \15470 , \12644 );
buf \U$13730 ( \15471 , \12611 );
buf \U$13731 ( \15472 , \12595 );
buf \U$13732 ( \15473 , \12599 );
buf \U$13733 ( \15474 , \12603 );
buf \U$13734 ( \15475 , \12607 );
or \U$13735 ( \15476 , \15472 , \15473 , \15474 , \15475 );
and \U$13736 ( \15477 , \15471 , \15476 );
or \U$13737 ( \15478 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15477 );
buf \U$13738 ( \15479 , \15478 );
_DC g1512 ( \15480_nG1512 , \15462 , \15479 );
buf \U$13739 ( \15481 , \15480_nG1512 );
and \U$13740 ( \15482 , \15427 , \15481 );
xor \U$13741 ( \15483 , \15400 , \15422 );
buf \U$13742 ( \15484 , \15483 );
buf \U$13743 ( \15485 , \15484 );
not \U$13744 ( \15486 , \15485 );
and \U$13745 ( \15487 , RI2b5e785daa40_28, \15428 );
and \U$13746 ( \15488 , RI2b5e78549540_41, \15430 );
and \U$13747 ( \15489 , RI2b5e785388a8_54, \15432 );
and \U$13748 ( \15490 , RI2b5e784a6330_67, \15434 );
and \U$13749 ( \15491 , RI2b5e78495698_80, \15436 );
and \U$13750 ( \15492 , RI2b5e78495080_93, \15438 );
and \U$13751 ( \15493 , RI2b5e78403b80_106, \15440 );
and \U$13752 ( \15494 , RI2b5e775b1e60_119, \15442 );
and \U$13753 ( \15495 , RI2b5e7750bdf8_132, \15444 );
and \U$13754 ( \15496 , RI2b5e774ff5d0_145, \15446 );
and \U$13755 ( \15497 , RI2b5e774f65e8_158, \15448 );
and \U$13756 ( \15498 , RI2b5e774eabd0_171, \15450 );
and \U$13757 ( \15499 , RI2b5e774de3a8_184, \15452 );
and \U$13758 ( \15500 , RI2b5e774d53c0_197, \15454 );
and \U$13759 ( \15501 , RI2b5e785f4300_210, \15456 );
and \U$13760 ( \15502 , RI2b5e785f3ce8_223, \15458 );
and \U$13761 ( \15503 , RI2b5e785eb0c0_236, \15460 );
or \U$13762 ( \15504 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 );
_DC g152b ( \15505_nG152b , \15504 , \15479 );
buf \U$13763 ( \15506 , \15505_nG152b );
and \U$13764 ( \15507 , \15486 , \15506 );
xor \U$13765 ( \15508 , \15401 , \15421 );
buf \U$13766 ( \15509 , \15508 );
buf \U$13767 ( \15510 , \15509 );
not \U$13768 ( \15511 , \15510 );
and \U$13769 ( \15512 , RI2b5e785da9c8_29, \15428 );
and \U$13770 ( \15513 , RI2b5e785494c8_42, \15430 );
and \U$13771 ( \15514 , RI2b5e78538830_55, \15432 );
and \U$13772 ( \15515 , RI2b5e784a62b8_68, \15434 );
and \U$13773 ( \15516 , RI2b5e78495620_81, \15436 );
and \U$13774 ( \15517 , RI2b5e78495008_94, \15438 );
and \U$13775 ( \15518 , RI2b5e78403b08_107, \15440 );
and \U$13776 ( \15519 , RI2b5e775b1de8_120, \15442 );
and \U$13777 ( \15520 , RI2b5e7750bd80_133, \15444 );
and \U$13778 ( \15521 , RI2b5e774ff558_146, \15446 );
and \U$13779 ( \15522 , RI2b5e774f6570_159, \15448 );
and \U$13780 ( \15523 , RI2b5e774eab58_172, \15450 );
and \U$13781 ( \15524 , RI2b5e774de330_185, \15452 );
and \U$13782 ( \15525 , RI2b5e774d5348_198, \15454 );
and \U$13783 ( \15526 , RI2b5e785f4288_211, \15456 );
and \U$13784 ( \15527 , RI2b5e785f3658_224, \15458 );
and \U$13785 ( \15528 , RI2b5e785eb048_237, \15460 );
or \U$13786 ( \15529 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 );
_DC g1544 ( \15530_nG1544 , \15529 , \15479 );
buf \U$13787 ( \15531 , \15530_nG1544 );
and \U$13788 ( \15532 , \15511 , \15531 );
xor \U$13789 ( \15533 , \15402 , \15420 );
buf \U$13790 ( \15534 , \15533 );
buf \U$13791 ( \15535 , \15534 );
not \U$13792 ( \15536 , \15535 );
and \U$13793 ( \15537 , RI2b5e785da950_30, \15428 );
and \U$13794 ( \15538 , RI2b5e78549450_43, \15430 );
and \U$13795 ( \15539 , RI2b5e785387b8_56, \15432 );
and \U$13796 ( \15540 , RI2b5e784a6240_69, \15434 );
and \U$13797 ( \15541 , RI2b5e784955a8_82, \15436 );
and \U$13798 ( \15542 , RI2b5e78494f90_95, \15438 );
and \U$13799 ( \15543 , RI2b5e78403a90_108, \15440 );
and \U$13800 ( \15544 , RI2b5e775b1d70_121, \15442 );
and \U$13801 ( \15545 , RI2b5e7750bd08_134, \15444 );
and \U$13802 ( \15546 , RI2b5e774ff4e0_147, \15446 );
and \U$13803 ( \15547 , RI2b5e774f64f8_160, \15448 );
and \U$13804 ( \15548 , RI2b5e774eaae0_173, \15450 );
and \U$13805 ( \15549 , RI2b5e774de2b8_186, \15452 );
and \U$13806 ( \15550 , RI2b5e774d52d0_199, \15454 );
and \U$13807 ( \15551 , RI2b5e785f4210_212, \15456 );
and \U$13808 ( \15552 , RI2b5e785eb5e8_225, \15458 );
and \U$13809 ( \15553 , RI2b5e785e6c50_238, \15460 );
or \U$13810 ( \15554 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 );
_DC g155d ( \15555_nG155d , \15554 , \15479 );
buf \U$13811 ( \15556 , \15555_nG155d );
and \U$13812 ( \15557 , \15536 , \15556 );
xor \U$13813 ( \15558 , \15403 , \15419 );
buf \U$13814 ( \15559 , \15558 );
buf \U$13815 ( \15560 , \15559 );
not \U$13816 ( \15561 , \15560 );
and \U$13817 ( \15562 , RI2b5e785da8d8_31, \15428 );
and \U$13818 ( \15563 , RI2b5e785493d8_44, \15430 );
and \U$13819 ( \15564 , RI2b5e78538740_57, \15432 );
and \U$13820 ( \15565 , RI2b5e784a61c8_70, \15434 );
and \U$13821 ( \15566 , RI2b5e78495530_83, \15436 );
and \U$13822 ( \15567 , RI2b5e78494f18_96, \15438 );
and \U$13823 ( \15568 , RI2b5e78403a18_109, \15440 );
and \U$13824 ( \15569 , RI2b5e775b1cf8_122, \15442 );
and \U$13825 ( \15570 , RI2b5e7750bc90_135, \15444 );
and \U$13826 ( \15571 , RI2b5e774ff468_148, \15446 );
and \U$13827 ( \15572 , RI2b5e774f6480_161, \15448 );
and \U$13828 ( \15573 , RI2b5e774eaa68_174, \15450 );
and \U$13829 ( \15574 , RI2b5e774de240_187, \15452 );
and \U$13830 ( \15575 , RI2b5e774d5258_200, \15454 );
and \U$13831 ( \15576 , RI2b5e785f4198_213, \15456 );
and \U$13832 ( \15577 , RI2b5e785eb570_226, \15458 );
and \U$13833 ( \15578 , RI2b5e785e6bd8_239, \15460 );
or \U$13834 ( \15579 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 );
_DC g1576 ( \15580_nG1576 , \15579 , \15479 );
buf \U$13835 ( \15581 , \15580_nG1576 );
and \U$13836 ( \15582 , \15561 , \15581 );
xor \U$13837 ( \15583 , \15404 , \15418 );
buf \U$13838 ( \15584 , \15583 );
buf \U$13839 ( \15585 , \15584 );
not \U$13840 ( \15586 , \15585 );
and \U$13841 ( \15587 , RI2b5e785da860_32, \15428 );
and \U$13842 ( \15588 , RI2b5e78549360_45, \15430 );
and \U$13843 ( \15589 , RI2b5e785386c8_58, \15432 );
and \U$13844 ( \15590 , RI2b5e784a6150_71, \15434 );
and \U$13845 ( \15591 , RI2b5e784954b8_84, \15436 );
and \U$13846 ( \15592 , RI2b5e78494ea0_97, \15438 );
and \U$13847 ( \15593 , RI2b5e784039a0_110, \15440 );
and \U$13848 ( \15594 , RI2b5e775b1c80_123, \15442 );
and \U$13849 ( \15595 , RI2b5e7750bc18_136, \15444 );
and \U$13850 ( \15596 , RI2b5e774ff3f0_149, \15446 );
and \U$13851 ( \15597 , RI2b5e774f6408_162, \15448 );
and \U$13852 ( \15598 , RI2b5e774ea9f0_175, \15450 );
and \U$13853 ( \15599 , RI2b5e774de1c8_188, \15452 );
and \U$13854 ( \15600 , RI2b5e774d51e0_201, \15454 );
and \U$13855 ( \15601 , RI2b5e785f4120_214, \15456 );
and \U$13856 ( \15602 , RI2b5e785eb4f8_227, \15458 );
and \U$13857 ( \15603 , RI2b5e785e64d0_240, \15460 );
or \U$13858 ( \15604 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 );
_DC g158f ( \15605_nG158f , \15604 , \15479 );
buf \U$13859 ( \15606 , \15605_nG158f );
and \U$13860 ( \15607 , \15586 , \15606 );
xor \U$13861 ( \15608 , \15405 , \15417 );
buf \U$13862 ( \15609 , \15608 );
buf \U$13863 ( \15610 , \15609 );
not \U$13864 ( \15611 , \15610 );
and \U$13865 ( \15612 , RI2b5e78549900_33, \15428 );
and \U$13866 ( \15613 , RI2b5e78538c68_46, \15430 );
and \U$13867 ( \15614 , RI2b5e78538650_59, \15432 );
and \U$13868 ( \15615 , RI2b5e784a60d8_72, \15434 );
and \U$13869 ( \15616 , RI2b5e78495440_85, \15436 );
and \U$13870 ( \15617 , RI2b5e78494e28_98, \15438 );
and \U$13871 ( \15618 , RI2b5e78403928_111, \15440 );
and \U$13872 ( \15619 , RI2b5e775b1c08_124, \15442 );
and \U$13873 ( \15620 , RI2b5e7750bba0_137, \15444 );
and \U$13874 ( \15621 , RI2b5e774ff378_150, \15446 );
and \U$13875 ( \15622 , RI2b5e774f6390_163, \15448 );
and \U$13876 ( \15623 , RI2b5e774ea978_176, \15450 );
and \U$13877 ( \15624 , RI2b5e774de150_189, \15452 );
and \U$13878 ( \15625 , RI2b5e774d5168_202, \15454 );
and \U$13879 ( \15626 , RI2b5e785f40a8_215, \15456 );
and \U$13880 ( \15627 , RI2b5e785eb480_228, \15458 );
and \U$13881 ( \15628 , RI2b5e785da608_241, \15460 );
or \U$13882 ( \15629 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 );
_DC g15a8 ( \15630_nG15a8 , \15629 , \15479 );
buf \U$13883 ( \15631 , \15630_nG15a8 );
and \U$13884 ( \15632 , \15611 , \15631 );
xor \U$13885 ( \15633 , \15406 , \15416 );
buf \U$13886 ( \15634 , \15633 );
buf \U$13887 ( \15635 , \15634 );
not \U$13888 ( \15636 , \15635 );
and \U$13889 ( \15637 , RI2b5e78549888_34, \15428 );
and \U$13890 ( \15638 , RI2b5e78538bf0_47, \15430 );
and \U$13891 ( \15639 , RI2b5e785385d8_60, \15432 );
and \U$13892 ( \15640 , RI2b5e784a6060_73, \15434 );
and \U$13893 ( \15641 , RI2b5e784953c8_86, \15436 );
and \U$13894 ( \15642 , RI2b5e78403ec8_99, \15438 );
and \U$13895 ( \15643 , RI2b5e775b21a8_112, \15440 );
and \U$13896 ( \15644 , RI2b5e775b1b90_125, \15442 );
and \U$13897 ( \15645 , RI2b5e7750bb28_138, \15444 );
and \U$13898 ( \15646 , RI2b5e774ff300_151, \15446 );
and \U$13899 ( \15647 , RI2b5e774f6318_164, \15448 );
and \U$13900 ( \15648 , RI2b5e774ea900_177, \15450 );
and \U$13901 ( \15649 , RI2b5e774de0d8_190, \15452 );
and \U$13902 ( \15650 , RI2b5e774d50f0_203, \15454 );
and \U$13903 ( \15651 , RI2b5e785f4030_216, \15456 );
and \U$13904 ( \15652 , RI2b5e785eb408_229, \15458 );
and \U$13905 ( \15653 , RI2b5e785da590_242, \15460 );
or \U$13906 ( \15654 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 );
_DC g15c1 ( \15655_nG15c1 , \15654 , \15479 );
buf \U$13907 ( \15656 , \15655_nG15c1 );
and \U$13908 ( \15657 , \15636 , \15656 );
xor \U$13909 ( \15658 , \15407 , \15415 );
buf \U$13910 ( \15659 , \15658 );
buf \U$13911 ( \15660 , \15659 );
not \U$13912 ( \15661 , \15660 );
and \U$13913 ( \15662 , RI2b5e78549810_35, \15428 );
and \U$13914 ( \15663 , RI2b5e78538b78_48, \15430 );
and \U$13915 ( \15664 , RI2b5e78538560_61, \15432 );
and \U$13916 ( \15665 , RI2b5e784a5fe8_74, \15434 );
and \U$13917 ( \15666 , RI2b5e78495350_87, \15436 );
and \U$13918 ( \15667 , RI2b5e78403e50_100, \15438 );
and \U$13919 ( \15668 , RI2b5e775b2130_113, \15440 );
and \U$13920 ( \15669 , RI2b5e775b1b18_126, \15442 );
and \U$13921 ( \15670 , RI2b5e7750bab0_139, \15444 );
and \U$13922 ( \15671 , RI2b5e774ff288_152, \15446 );
and \U$13923 ( \15672 , RI2b5e774f62a0_165, \15448 );
and \U$13924 ( \15673 , RI2b5e774ea888_178, \15450 );
and \U$13925 ( \15674 , RI2b5e774de060_191, \15452 );
and \U$13926 ( \15675 , RI2b5e774d5078_204, \15454 );
and \U$13927 ( \15676 , RI2b5e785f3fb8_217, \15456 );
and \U$13928 ( \15677 , RI2b5e785eb390_230, \15458 );
and \U$13929 ( \15678 , RI2b5e785da518_243, \15460 );
or \U$13930 ( \15679 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 );
_DC g15da ( \15680_nG15da , \15679 , \15479 );
buf \U$13931 ( \15681 , \15680_nG15da );
and \U$13932 ( \15682 , \15661 , \15681 );
xor \U$13933 ( \15683 , \15408 , \15414 );
buf \U$13934 ( \15684 , \15683 );
buf \U$13935 ( \15685 , \15684 );
not \U$13936 ( \15686 , \15685 );
and \U$13937 ( \15687 , RI2b5e78549798_36, \15428 );
and \U$13938 ( \15688 , RI2b5e78538b00_49, \15430 );
and \U$13939 ( \15689 , RI2b5e785384e8_62, \15432 );
and \U$13940 ( \15690 , RI2b5e784a5f70_75, \15434 );
and \U$13941 ( \15691 , RI2b5e784952d8_88, \15436 );
and \U$13942 ( \15692 , RI2b5e78403dd8_101, \15438 );
and \U$13943 ( \15693 , RI2b5e775b20b8_114, \15440 );
and \U$13944 ( \15694 , RI2b5e775b1aa0_127, \15442 );
and \U$13945 ( \15695 , RI2b5e7750ba38_140, \15444 );
and \U$13946 ( \15696 , RI2b5e774ff210_153, \15446 );
and \U$13947 ( \15697 , RI2b5e774f6228_166, \15448 );
and \U$13948 ( \15698 , RI2b5e774ea810_179, \15450 );
and \U$13949 ( \15699 , RI2b5e774ddfe8_192, \15452 );
and \U$13950 ( \15700 , RI2b5e774d5000_205, \15454 );
and \U$13951 ( \15701 , RI2b5e785f3f40_218, \15456 );
and \U$13952 ( \15702 , RI2b5e785eb318_231, \15458 );
and \U$13953 ( \15703 , RI2b5e785da4a0_244, \15460 );
or \U$13954 ( \15704 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 );
_DC g15f3 ( \15705_nG15f3 , \15704 , \15479 );
buf \U$13955 ( \15706 , \15705_nG15f3 );
and \U$13956 ( \15707 , \15686 , \15706 );
xor \U$13957 ( \15708 , \15409 , \15413 );
buf \U$13958 ( \15709 , \15708 );
buf \U$13959 ( \15710 , \15709 );
not \U$13960 ( \15711 , \15710 );
and \U$13961 ( \15712 , RI2b5e78549720_37, \15428 );
and \U$13962 ( \15713 , RI2b5e78538a88_50, \15430 );
and \U$13963 ( \15714 , RI2b5e78538470_63, \15432 );
and \U$13964 ( \15715 , RI2b5e784a5ef8_76, \15434 );
and \U$13965 ( \15716 , RI2b5e78495260_89, \15436 );
and \U$13966 ( \15717 , RI2b5e78403d60_102, \15438 );
and \U$13967 ( \15718 , RI2b5e775b2040_115, \15440 );
and \U$13968 ( \15719 , RI2b5e775b1a28_128, \15442 );
and \U$13969 ( \15720 , RI2b5e7750b9c0_141, \15444 );
and \U$13970 ( \15721 , RI2b5e774ff198_154, \15446 );
and \U$13971 ( \15722 , RI2b5e774f61b0_167, \15448 );
and \U$13972 ( \15723 , RI2b5e774ea798_180, \15450 );
and \U$13973 ( \15724 , RI2b5e774ddf70_193, \15452 );
and \U$13974 ( \15725 , RI2b5e774d4f88_206, \15454 );
and \U$13975 ( \15726 , RI2b5e785f3ec8_219, \15456 );
and \U$13976 ( \15727 , RI2b5e785eb2a0_232, \15458 );
and \U$13977 ( \15728 , RI2b5e785da428_245, \15460 );
or \U$13978 ( \15729 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 );
_DC g160c ( \15730_nG160c , \15729 , \15479 );
buf \U$13979 ( \15731 , \15730_nG160c );
and \U$13980 ( \15732 , \15711 , \15731 );
xor \U$13981 ( \15733 , \15410 , \15412 );
buf \U$13982 ( \15734 , \15733 );
buf \U$13983 ( \15735 , \15734 );
not \U$13984 ( \15736 , \15735 );
and \U$13985 ( \15737 , RI2b5e785496a8_38, \15428 );
and \U$13986 ( \15738 , RI2b5e78538a10_51, \15430 );
and \U$13987 ( \15739 , RI2b5e785383f8_64, \15432 );
and \U$13988 ( \15740 , RI2b5e784a5e80_77, \15434 );
and \U$13989 ( \15741 , RI2b5e784951e8_90, \15436 );
and \U$13990 ( \15742 , RI2b5e78403ce8_103, \15438 );
and \U$13991 ( \15743 , RI2b5e775b1fc8_116, \15440 );
and \U$13992 ( \15744 , RI2b5e775b19b0_129, \15442 );
and \U$13993 ( \15745 , RI2b5e7750b948_142, \15444 );
and \U$13994 ( \15746 , RI2b5e774ff120_155, \15446 );
and \U$13995 ( \15747 , RI2b5e774f6138_168, \15448 );
and \U$13996 ( \15748 , RI2b5e774ea720_181, \15450 );
and \U$13997 ( \15749 , RI2b5e774ddef8_194, \15452 );
and \U$13998 ( \15750 , RI2b5e774d4f10_207, \15454 );
and \U$13999 ( \15751 , RI2b5e785f3e50_220, \15456 );
and \U$14000 ( \15752 , RI2b5e785eb228_233, \15458 );
and \U$14001 ( \15753 , RI2b5e785da3b0_246, \15460 );
or \U$14002 ( \15754 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 );
_DC g1625 ( \15755_nG1625 , \15754 , \15479 );
buf \U$14003 ( \15756 , \15755_nG1625 );
and \U$14004 ( \15757 , \15736 , \15756 );
buf \U$14005 ( \15758 , RI2b5e785dab30_26);
buf \U$14008 ( \15759 , \15758 );
not \U$14009 ( \15760 , \15759 );
and \U$14010 ( \15761 , RI2b5e78549630_39, \15428 );
and \U$14011 ( \15762 , RI2b5e78538998_52, \15430 );
and \U$14012 ( \15763 , RI2b5e78538380_65, \15432 );
and \U$14013 ( \15764 , RI2b5e784a5e08_78, \15434 );
and \U$14014 ( \15765 , RI2b5e78495170_91, \15436 );
and \U$14015 ( \15766 , RI2b5e78403c70_104, \15438 );
and \U$14016 ( \15767 , RI2b5e775b1f50_117, \15440 );
and \U$14017 ( \15768 , RI2b5e775b1938_130, \15442 );
and \U$14018 ( \15769 , RI2b5e7750b8d0_143, \15444 );
and \U$14019 ( \15770 , RI2b5e774ff0a8_156, \15446 );
and \U$14020 ( \15771 , RI2b5e774f60c0_169, \15448 );
and \U$14021 ( \15772 , RI2b5e774ea6a8_182, \15450 );
and \U$14022 ( \15773 , RI2b5e774dde80_195, \15452 );
and \U$14023 ( \15774 , RI2b5e774d4e98_208, \15454 );
and \U$14024 ( \15775 , RI2b5e785f3dd8_221, \15456 );
and \U$14025 ( \15776 , RI2b5e785eb1b0_234, \15458 );
and \U$14026 ( \15777 , RI2b5e785da338_247, \15460 );
or \U$14027 ( \15778 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 );
_DC g163f ( \15779_nG163f , \15778 , \15479 );
buf \U$14028 ( \15780 , \15779_nG163f );
and \U$14029 ( \15781 , \15760 , \15780 );
xnor \U$14030 ( \15782 , \15735 , \15756 );
and \U$14031 ( \15783 , \15781 , \15782 );
or \U$14032 ( \15784 , \15757 , \15783 );
xnor \U$14033 ( \15785 , \15710 , \15731 );
and \U$14034 ( \15786 , \15784 , \15785 );
or \U$14035 ( \15787 , \15732 , \15786 );
xnor \U$14036 ( \15788 , \15685 , \15706 );
and \U$14037 ( \15789 , \15787 , \15788 );
or \U$14038 ( \15790 , \15707 , \15789 );
xnor \U$14039 ( \15791 , \15660 , \15681 );
and \U$14040 ( \15792 , \15790 , \15791 );
or \U$14041 ( \15793 , \15682 , \15792 );
xnor \U$14042 ( \15794 , \15635 , \15656 );
and \U$14043 ( \15795 , \15793 , \15794 );
or \U$14044 ( \15796 , \15657 , \15795 );
xnor \U$14045 ( \15797 , \15610 , \15631 );
and \U$14046 ( \15798 , \15796 , \15797 );
or \U$14047 ( \15799 , \15632 , \15798 );
xnor \U$14048 ( \15800 , \15585 , \15606 );
and \U$14049 ( \15801 , \15799 , \15800 );
or \U$14050 ( \15802 , \15607 , \15801 );
xnor \U$14051 ( \15803 , \15560 , \15581 );
and \U$14052 ( \15804 , \15802 , \15803 );
or \U$14053 ( \15805 , \15582 , \15804 );
xnor \U$14054 ( \15806 , \15535 , \15556 );
and \U$14055 ( \15807 , \15805 , \15806 );
or \U$14056 ( \15808 , \15557 , \15807 );
xnor \U$14057 ( \15809 , \15510 , \15531 );
and \U$14058 ( \15810 , \15808 , \15809 );
or \U$14059 ( \15811 , \15532 , \15810 );
xnor \U$14060 ( \15812 , \15485 , \15506 );
and \U$14061 ( \15813 , \15811 , \15812 );
or \U$14062 ( \15814 , \15507 , \15813 );
xnor \U$14063 ( \15815 , \15426 , \15481 );
and \U$14064 ( \15816 , \15814 , \15815 );
or \U$14065 ( \15817 , \15482 , \15816 );
not \U$14066 ( \15818 , \15817 );
buf \U$14067 ( \15819 , \15818 );
buf \U$14068 ( \15820 , RI2b5e785ae580_609);
buf \U$14069 ( \15821 , RI2b5e785ae5f8_608);
buf \U$14070 ( \15822 , RI2b5e785ae670_607);
buf \U$14071 ( \15823 , RI2b5e785ae6e8_606);
buf \U$14072 ( \15824 , RI2b5e785ae760_605);
buf \U$14073 ( \15825 , RI2b5e785ae7d8_604);
buf \U$14074 ( \15826 , RI2b5e785ae850_603);
buf \U$14075 ( \15827 , RI2b5e785ae8c8_602);
buf \U$14076 ( \15828 , RI2b5e785ae940_601);
buf \U$14077 ( \15829 , RI2b5e785ae3a0_613);
buf \U$14078 ( \15830 , RI2b5e785ae418_612);
buf \U$14079 ( \15831 , RI2b5e785ae490_611);
buf \U$14080 ( \15832 , RI2b5e785ae508_610);
and \U$14081 ( \15833 , \15829 , \15830 , \15831 , \15832 );
nor \U$14082 ( \15834 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15833 );
buf \U$14083 ( \15835 , \15834 );
and \U$14084 ( \15836 , \15819 , \15835 );
nor \U$14085 ( \15837 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9798 , RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14086 ( \15838 , RI2b5e785daab8_27, \15837 );
nor \U$14087 ( \15839 , \9801 , \9802 , \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14088 ( \15840 , RI2b5e785495b8_40, \15839 );
nor \U$14089 ( \15841 , RI2b5e785ae3a0_613, \9802 , \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14090 ( \15842 , RI2b5e78538920_53, \15841 );
nor \U$14091 ( \15843 , \9801 , RI2b5e785ae418_612, \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14092 ( \15844 , RI2b5e784a63a8_66, \15843 );
nor \U$14093 ( \15845 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9803 , \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14094 ( \15846 , RI2b5e78495710_79, \15845 );
nor \U$14095 ( \15847 , \9801 , \9802 , RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14096 ( \15848 , RI2b5e784950f8_92, \15847 );
nor \U$14097 ( \15849 , RI2b5e785ae3a0_613, \9802 , RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14098 ( \15850 , RI2b5e78403bf8_105, \15849 );
nor \U$14099 ( \15851 , \9801 , RI2b5e785ae418_612, RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14100 ( \15852 , RI2b5e775b1ed8_118, \15851 );
nor \U$14101 ( \15853 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, \9804 , RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14102 ( \15854 , RI2b5e775b18c0_131, \15853 );
nor \U$14103 ( \15855 , \9801 , \9802 , \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14104 ( \15856 , RI2b5e7750b858_144, \15855 );
nor \U$14105 ( \15857 , RI2b5e785ae3a0_613, \9802 , \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14106 ( \15858 , RI2b5e774ff030_157, \15857 );
nor \U$14107 ( \15859 , \9801 , RI2b5e785ae418_612, \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14108 ( \15860 , RI2b5e774f6048_170, \15859 );
nor \U$14109 ( \15861 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9803 , RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14110 ( \15862 , RI2b5e774ea630_183, \15861 );
nor \U$14111 ( \15863 , \9801 , \9802 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14112 ( \15864 , RI2b5e774dde08_196, \15863 );
nor \U$14113 ( \15865 , RI2b5e785ae3a0_613, \9802 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14114 ( \15866 , RI2b5e774d4e20_209, \15865 );
nor \U$14115 ( \15867 , \9801 , RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14116 ( \15868 , RI2b5e785f3d60_222, \15867 );
nor \U$14117 ( \15869 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609, RI2b5e785ae5f8_608, RI2b5e785ae670_607, RI2b5e785ae6e8_606, RI2b5e785ae760_605, RI2b5e785ae7d8_604, RI2b5e785ae850_603, RI2b5e785ae8c8_602, RI2b5e785ae940_601);
and \U$14118 ( \15870 , RI2b5e785eb138_235, \15869 );
or \U$14119 ( \15871 , \15838 , \15840 , \15842 , \15844 , \15846 , \15848 , \15850 , \15852 , \15854 , \15856 , \15858 , \15860 , \15862 , \15864 , \15866 , \15868 , \15870 );
buf \U$14120 ( \15872 , RI2b5e785ae5f8_608);
buf \U$14121 ( \15873 , RI2b5e785ae670_607);
buf \U$14122 ( \15874 , RI2b5e785ae6e8_606);
buf \U$14123 ( \15875 , RI2b5e785ae760_605);
buf \U$14124 ( \15876 , RI2b5e785ae7d8_604);
buf \U$14125 ( \15877 , RI2b5e785ae850_603);
buf \U$14126 ( \15878 , RI2b5e785ae8c8_602);
buf \U$14127 ( \15879 , RI2b5e785ae940_601);
buf \U$14128 ( \15880 , RI2b5e785ae580_609);
buf \U$14129 ( \15881 , RI2b5e785ae3a0_613);
buf \U$14130 ( \15882 , RI2b5e785ae418_612);
buf \U$14131 ( \15883 , RI2b5e785ae490_611);
buf \U$14132 ( \15884 , RI2b5e785ae508_610);
or \U$14133 ( \15885 , \15881 , \15882 , \15883 , \15884 );
and \U$14134 ( \15886 , \15880 , \15885 );
or \U$14135 ( \15887 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15886 );
buf \U$14136 ( \15888 , \15887 );
_DC g16b2 ( \15889_nG16b2 , \15871 , \15888 );
buf \U$14137 ( \15890 , \15889_nG16b2 );
not \U$14138 ( \15891 , \15890 );
nor \U$14139 ( \15892 , \12595 , \12599 , \12603 , \12607 , \12612 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14140 ( \15893 , RI2b5e785daab8_27, \15892 );
nor \U$14141 ( \15894 , \12647 , \12648 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14142 ( \15895 , RI2b5e785495b8_40, \15894 );
nor \U$14143 ( \15896 , \12595 , \12648 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14144 ( \15897 , RI2b5e78538920_53, \15896 );
nor \U$14145 ( \15898 , \12647 , \12599 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14146 ( \15899 , RI2b5e784a63a8_66, \15898 );
nor \U$14147 ( \15900 , \12595 , \12599 , \12649 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14148 ( \15901 , RI2b5e78495710_79, \15900 );
nor \U$14149 ( \15902 , \12647 , \12648 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14150 ( \15903 , RI2b5e784950f8_92, \15902 );
nor \U$14151 ( \15904 , \12595 , \12648 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14152 ( \15905 , RI2b5e78403bf8_105, \15904 );
nor \U$14153 ( \15906 , \12647 , \12599 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14154 ( \15907 , RI2b5e775b1ed8_118, \15906 );
nor \U$14155 ( \15908 , \12595 , \12599 , \12603 , \12650 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14156 ( \15909 , RI2b5e775b18c0_131, \15908 );
nor \U$14157 ( \15910 , \12647 , \12648 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14158 ( \15911 , RI2b5e7750b858_144, \15910 );
nor \U$14159 ( \15912 , \12595 , \12648 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14160 ( \15913 , RI2b5e774ff030_157, \15912 );
nor \U$14161 ( \15914 , \12647 , \12599 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14162 ( \15915 , RI2b5e774f6048_170, \15914 );
nor \U$14163 ( \15916 , \12595 , \12599 , \12649 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14164 ( \15917 , RI2b5e774ea630_183, \15916 );
nor \U$14165 ( \15918 , \12647 , \12648 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14166 ( \15919 , RI2b5e774dde08_196, \15918 );
nor \U$14167 ( \15920 , \12595 , \12648 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14168 ( \15921 , RI2b5e774d4e20_209, \15920 );
nor \U$14169 ( \15922 , \12647 , \12599 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14170 ( \15923 , RI2b5e785f3d60_222, \15922 );
nor \U$14171 ( \15924 , \12595 , \12599 , \12603 , \12607 , \12611 , \12616 , \12620 , \12624 , \12628 , \12632 , \12636 , \12640 , \12644 );
and \U$14172 ( \15925 , RI2b5e785eb138_235, \15924 );
or \U$14173 ( \15926 , \15893 , \15895 , \15897 , \15899 , \15901 , \15903 , \15905 , \15907 , \15909 , \15911 , \15913 , \15915 , \15917 , \15919 , \15921 , \15923 , \15925 );
buf \U$14174 ( \15927 , \12616 );
buf \U$14175 ( \15928 , \12620 );
buf \U$14176 ( \15929 , \12624 );
buf \U$14177 ( \15930 , \12628 );
buf \U$14178 ( \15931 , \12632 );
buf \U$14179 ( \15932 , \12636 );
buf \U$14180 ( \15933 , \12640 );
buf \U$14181 ( \15934 , \12644 );
buf \U$14182 ( \15935 , \12611 );
buf \U$14183 ( \15936 , \12595 );
buf \U$14184 ( \15937 , \12599 );
buf \U$14185 ( \15938 , \12603 );
buf \U$14186 ( \15939 , \12607 );
or \U$14187 ( \15940 , \15936 , \15937 , \15938 , \15939 );
and \U$14188 ( \15941 , \15935 , \15940 );
or \U$14189 ( \15942 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15941 );
buf \U$14190 ( \15943 , \15942 );
_DC g16e9 ( \15944_nG16e9 , \15926 , \15943 );
buf \U$14191 ( \15945 , \15944_nG16e9 );
and \U$14192 ( \15946 , \15891 , \15945 );
and \U$14193 ( \15947 , RI2b5e785daa40_28, \15837 );
and \U$14194 ( \15948 , RI2b5e78549540_41, \15839 );
and \U$14195 ( \15949 , RI2b5e785388a8_54, \15841 );
and \U$14196 ( \15950 , RI2b5e784a6330_67, \15843 );
and \U$14197 ( \15951 , RI2b5e78495698_80, \15845 );
and \U$14198 ( \15952 , RI2b5e78495080_93, \15847 );
and \U$14199 ( \15953 , RI2b5e78403b80_106, \15849 );
and \U$14200 ( \15954 , RI2b5e775b1e60_119, \15851 );
and \U$14201 ( \15955 , RI2b5e7750bdf8_132, \15853 );
and \U$14202 ( \15956 , RI2b5e774ff5d0_145, \15855 );
and \U$14203 ( \15957 , RI2b5e774f65e8_158, \15857 );
and \U$14204 ( \15958 , RI2b5e774eabd0_171, \15859 );
and \U$14205 ( \15959 , RI2b5e774de3a8_184, \15861 );
and \U$14206 ( \15960 , RI2b5e774d53c0_197, \15863 );
and \U$14207 ( \15961 , RI2b5e785f4300_210, \15865 );
and \U$14208 ( \15962 , RI2b5e785f3ce8_223, \15867 );
and \U$14209 ( \15963 , RI2b5e785eb0c0_236, \15869 );
or \U$14210 ( \15964 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 );
_DC g16fe ( \15965_nG16fe , \15964 , \15888 );
buf \U$14211 ( \15966 , \15965_nG16fe );
not \U$14212 ( \15967 , \15966 );
and \U$14213 ( \15968 , RI2b5e785daa40_28, \15892 );
and \U$14214 ( \15969 , RI2b5e78549540_41, \15894 );
and \U$14215 ( \15970 , RI2b5e785388a8_54, \15896 );
and \U$14216 ( \15971 , RI2b5e784a6330_67, \15898 );
and \U$14217 ( \15972 , RI2b5e78495698_80, \15900 );
and \U$14218 ( \15973 , RI2b5e78495080_93, \15902 );
and \U$14219 ( \15974 , RI2b5e78403b80_106, \15904 );
and \U$14220 ( \15975 , RI2b5e775b1e60_119, \15906 );
and \U$14221 ( \15976 , RI2b5e7750bdf8_132, \15908 );
and \U$14222 ( \15977 , RI2b5e774ff5d0_145, \15910 );
and \U$14223 ( \15978 , RI2b5e774f65e8_158, \15912 );
and \U$14224 ( \15979 , RI2b5e774eabd0_171, \15914 );
and \U$14225 ( \15980 , RI2b5e774de3a8_184, \15916 );
and \U$14226 ( \15981 , RI2b5e774d53c0_197, \15918 );
and \U$14227 ( \15982 , RI2b5e785f4300_210, \15920 );
and \U$14228 ( \15983 , RI2b5e785f3ce8_223, \15922 );
and \U$14229 ( \15984 , RI2b5e785eb0c0_236, \15924 );
or \U$14230 ( \15985 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 );
_DC g1713 ( \15986_nG1713 , \15985 , \15943 );
buf \U$14231 ( \15987 , \15986_nG1713 );
and \U$14232 ( \15988 , \15967 , \15987 );
and \U$14233 ( \15989 , RI2b5e785da9c8_29, \15837 );
and \U$14234 ( \15990 , RI2b5e785494c8_42, \15839 );
and \U$14235 ( \15991 , RI2b5e78538830_55, \15841 );
and \U$14236 ( \15992 , RI2b5e784a62b8_68, \15843 );
and \U$14237 ( \15993 , RI2b5e78495620_81, \15845 );
and \U$14238 ( \15994 , RI2b5e78495008_94, \15847 );
and \U$14239 ( \15995 , RI2b5e78403b08_107, \15849 );
and \U$14240 ( \15996 , RI2b5e775b1de8_120, \15851 );
and \U$14241 ( \15997 , RI2b5e7750bd80_133, \15853 );
and \U$14242 ( \15998 , RI2b5e774ff558_146, \15855 );
and \U$14243 ( \15999 , RI2b5e774f6570_159, \15857 );
and \U$14244 ( \16000 , RI2b5e774eab58_172, \15859 );
and \U$14245 ( \16001 , RI2b5e774de330_185, \15861 );
and \U$14246 ( \16002 , RI2b5e774d5348_198, \15863 );
and \U$14247 ( \16003 , RI2b5e785f4288_211, \15865 );
and \U$14248 ( \16004 , RI2b5e785f3658_224, \15867 );
and \U$14249 ( \16005 , RI2b5e785eb048_237, \15869 );
or \U$14250 ( \16006 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 );
_DC g1728 ( \16007_nG1728 , \16006 , \15888 );
buf \U$14251 ( \16008 , \16007_nG1728 );
not \U$14252 ( \16009 , \16008 );
and \U$14253 ( \16010 , RI2b5e785da9c8_29, \15892 );
and \U$14254 ( \16011 , RI2b5e785494c8_42, \15894 );
and \U$14255 ( \16012 , RI2b5e78538830_55, \15896 );
and \U$14256 ( \16013 , RI2b5e784a62b8_68, \15898 );
and \U$14257 ( \16014 , RI2b5e78495620_81, \15900 );
and \U$14258 ( \16015 , RI2b5e78495008_94, \15902 );
and \U$14259 ( \16016 , RI2b5e78403b08_107, \15904 );
and \U$14260 ( \16017 , RI2b5e775b1de8_120, \15906 );
and \U$14261 ( \16018 , RI2b5e7750bd80_133, \15908 );
and \U$14262 ( \16019 , RI2b5e774ff558_146, \15910 );
and \U$14263 ( \16020 , RI2b5e774f6570_159, \15912 );
and \U$14264 ( \16021 , RI2b5e774eab58_172, \15914 );
and \U$14265 ( \16022 , RI2b5e774de330_185, \15916 );
and \U$14266 ( \16023 , RI2b5e774d5348_198, \15918 );
and \U$14267 ( \16024 , RI2b5e785f4288_211, \15920 );
and \U$14268 ( \16025 , RI2b5e785f3658_224, \15922 );
and \U$14269 ( \16026 , RI2b5e785eb048_237, \15924 );
or \U$14270 ( \16027 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 );
_DC g173d ( \16028_nG173d , \16027 , \15943 );
buf \U$14271 ( \16029 , \16028_nG173d );
and \U$14272 ( \16030 , \16009 , \16029 );
and \U$14273 ( \16031 , RI2b5e785da950_30, \15837 );
and \U$14274 ( \16032 , RI2b5e78549450_43, \15839 );
and \U$14275 ( \16033 , RI2b5e785387b8_56, \15841 );
and \U$14276 ( \16034 , RI2b5e784a6240_69, \15843 );
and \U$14277 ( \16035 , RI2b5e784955a8_82, \15845 );
and \U$14278 ( \16036 , RI2b5e78494f90_95, \15847 );
and \U$14279 ( \16037 , RI2b5e78403a90_108, \15849 );
and \U$14280 ( \16038 , RI2b5e775b1d70_121, \15851 );
and \U$14281 ( \16039 , RI2b5e7750bd08_134, \15853 );
and \U$14282 ( \16040 , RI2b5e774ff4e0_147, \15855 );
and \U$14283 ( \16041 , RI2b5e774f64f8_160, \15857 );
and \U$14284 ( \16042 , RI2b5e774eaae0_173, \15859 );
and \U$14285 ( \16043 , RI2b5e774de2b8_186, \15861 );
and \U$14286 ( \16044 , RI2b5e774d52d0_199, \15863 );
and \U$14287 ( \16045 , RI2b5e785f4210_212, \15865 );
and \U$14288 ( \16046 , RI2b5e785eb5e8_225, \15867 );
and \U$14289 ( \16047 , RI2b5e785e6c50_238, \15869 );
or \U$14290 ( \16048 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 );
_DC g1752 ( \16049_nG1752 , \16048 , \15888 );
buf \U$14291 ( \16050 , \16049_nG1752 );
not \U$14292 ( \16051 , \16050 );
and \U$14293 ( \16052 , RI2b5e785da950_30, \15892 );
and \U$14294 ( \16053 , RI2b5e78549450_43, \15894 );
and \U$14295 ( \16054 , RI2b5e785387b8_56, \15896 );
and \U$14296 ( \16055 , RI2b5e784a6240_69, \15898 );
and \U$14297 ( \16056 , RI2b5e784955a8_82, \15900 );
and \U$14298 ( \16057 , RI2b5e78494f90_95, \15902 );
and \U$14299 ( \16058 , RI2b5e78403a90_108, \15904 );
and \U$14300 ( \16059 , RI2b5e775b1d70_121, \15906 );
and \U$14301 ( \16060 , RI2b5e7750bd08_134, \15908 );
and \U$14302 ( \16061 , RI2b5e774ff4e0_147, \15910 );
and \U$14303 ( \16062 , RI2b5e774f64f8_160, \15912 );
and \U$14304 ( \16063 , RI2b5e774eaae0_173, \15914 );
and \U$14305 ( \16064 , RI2b5e774de2b8_186, \15916 );
and \U$14306 ( \16065 , RI2b5e774d52d0_199, \15918 );
and \U$14307 ( \16066 , RI2b5e785f4210_212, \15920 );
and \U$14308 ( \16067 , RI2b5e785eb5e8_225, \15922 );
and \U$14309 ( \16068 , RI2b5e785e6c50_238, \15924 );
or \U$14310 ( \16069 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 );
_DC g1767 ( \16070_nG1767 , \16069 , \15943 );
buf \U$14311 ( \16071 , \16070_nG1767 );
and \U$14312 ( \16072 , \16051 , \16071 );
and \U$14313 ( \16073 , RI2b5e785da8d8_31, \15837 );
and \U$14314 ( \16074 , RI2b5e785493d8_44, \15839 );
and \U$14315 ( \16075 , RI2b5e78538740_57, \15841 );
and \U$14316 ( \16076 , RI2b5e784a61c8_70, \15843 );
and \U$14317 ( \16077 , RI2b5e78495530_83, \15845 );
and \U$14318 ( \16078 , RI2b5e78494f18_96, \15847 );
and \U$14319 ( \16079 , RI2b5e78403a18_109, \15849 );
and \U$14320 ( \16080 , RI2b5e775b1cf8_122, \15851 );
and \U$14321 ( \16081 , RI2b5e7750bc90_135, \15853 );
and \U$14322 ( \16082 , RI2b5e774ff468_148, \15855 );
and \U$14323 ( \16083 , RI2b5e774f6480_161, \15857 );
and \U$14324 ( \16084 , RI2b5e774eaa68_174, \15859 );
and \U$14325 ( \16085 , RI2b5e774de240_187, \15861 );
and \U$14326 ( \16086 , RI2b5e774d5258_200, \15863 );
and \U$14327 ( \16087 , RI2b5e785f4198_213, \15865 );
and \U$14328 ( \16088 , RI2b5e785eb570_226, \15867 );
and \U$14329 ( \16089 , RI2b5e785e6bd8_239, \15869 );
or \U$14330 ( \16090 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 );
_DC g177c ( \16091_nG177c , \16090 , \15888 );
buf \U$14331 ( \16092 , \16091_nG177c );
not \U$14332 ( \16093 , \16092 );
and \U$14333 ( \16094 , RI2b5e785da8d8_31, \15892 );
and \U$14334 ( \16095 , RI2b5e785493d8_44, \15894 );
and \U$14335 ( \16096 , RI2b5e78538740_57, \15896 );
and \U$14336 ( \16097 , RI2b5e784a61c8_70, \15898 );
and \U$14337 ( \16098 , RI2b5e78495530_83, \15900 );
and \U$14338 ( \16099 , RI2b5e78494f18_96, \15902 );
and \U$14339 ( \16100 , RI2b5e78403a18_109, \15904 );
and \U$14340 ( \16101 , RI2b5e775b1cf8_122, \15906 );
and \U$14341 ( \16102 , RI2b5e7750bc90_135, \15908 );
and \U$14342 ( \16103 , RI2b5e774ff468_148, \15910 );
and \U$14343 ( \16104 , RI2b5e774f6480_161, \15912 );
and \U$14344 ( \16105 , RI2b5e774eaa68_174, \15914 );
and \U$14345 ( \16106 , RI2b5e774de240_187, \15916 );
and \U$14346 ( \16107 , RI2b5e774d5258_200, \15918 );
and \U$14347 ( \16108 , RI2b5e785f4198_213, \15920 );
and \U$14348 ( \16109 , RI2b5e785eb570_226, \15922 );
and \U$14349 ( \16110 , RI2b5e785e6bd8_239, \15924 );
or \U$14350 ( \16111 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 );
_DC g1791 ( \16112_nG1791 , \16111 , \15943 );
buf \U$14351 ( \16113 , \16112_nG1791 );
and \U$14352 ( \16114 , \16093 , \16113 );
and \U$14353 ( \16115 , RI2b5e785da860_32, \15837 );
and \U$14354 ( \16116 , RI2b5e78549360_45, \15839 );
and \U$14355 ( \16117 , RI2b5e785386c8_58, \15841 );
and \U$14356 ( \16118 , RI2b5e784a6150_71, \15843 );
and \U$14357 ( \16119 , RI2b5e784954b8_84, \15845 );
and \U$14358 ( \16120 , RI2b5e78494ea0_97, \15847 );
and \U$14359 ( \16121 , RI2b5e784039a0_110, \15849 );
and \U$14360 ( \16122 , RI2b5e775b1c80_123, \15851 );
and \U$14361 ( \16123 , RI2b5e7750bc18_136, \15853 );
and \U$14362 ( \16124 , RI2b5e774ff3f0_149, \15855 );
and \U$14363 ( \16125 , RI2b5e774f6408_162, \15857 );
and \U$14364 ( \16126 , RI2b5e774ea9f0_175, \15859 );
and \U$14365 ( \16127 , RI2b5e774de1c8_188, \15861 );
and \U$14366 ( \16128 , RI2b5e774d51e0_201, \15863 );
and \U$14367 ( \16129 , RI2b5e785f4120_214, \15865 );
and \U$14368 ( \16130 , RI2b5e785eb4f8_227, \15867 );
and \U$14369 ( \16131 , RI2b5e785e64d0_240, \15869 );
or \U$14370 ( \16132 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 );
_DC g17a6 ( \16133_nG17a6 , \16132 , \15888 );
buf \U$14371 ( \16134 , \16133_nG17a6 );
not \U$14372 ( \16135 , \16134 );
and \U$14373 ( \16136 , RI2b5e785da860_32, \15892 );
and \U$14374 ( \16137 , RI2b5e78549360_45, \15894 );
and \U$14375 ( \16138 , RI2b5e785386c8_58, \15896 );
and \U$14376 ( \16139 , RI2b5e784a6150_71, \15898 );
and \U$14377 ( \16140 , RI2b5e784954b8_84, \15900 );
and \U$14378 ( \16141 , RI2b5e78494ea0_97, \15902 );
and \U$14379 ( \16142 , RI2b5e784039a0_110, \15904 );
and \U$14380 ( \16143 , RI2b5e775b1c80_123, \15906 );
and \U$14381 ( \16144 , RI2b5e7750bc18_136, \15908 );
and \U$14382 ( \16145 , RI2b5e774ff3f0_149, \15910 );
and \U$14383 ( \16146 , RI2b5e774f6408_162, \15912 );
and \U$14384 ( \16147 , RI2b5e774ea9f0_175, \15914 );
and \U$14385 ( \16148 , RI2b5e774de1c8_188, \15916 );
and \U$14386 ( \16149 , RI2b5e774d51e0_201, \15918 );
and \U$14387 ( \16150 , RI2b5e785f4120_214, \15920 );
and \U$14388 ( \16151 , RI2b5e785eb4f8_227, \15922 );
and \U$14389 ( \16152 , RI2b5e785e64d0_240, \15924 );
or \U$14390 ( \16153 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 );
_DC g17bb ( \16154_nG17bb , \16153 , \15943 );
buf \U$14391 ( \16155 , \16154_nG17bb );
and \U$14392 ( \16156 , \16135 , \16155 );
and \U$14393 ( \16157 , RI2b5e78549900_33, \15837 );
and \U$14394 ( \16158 , RI2b5e78538c68_46, \15839 );
and \U$14395 ( \16159 , RI2b5e78538650_59, \15841 );
and \U$14396 ( \16160 , RI2b5e784a60d8_72, \15843 );
and \U$14397 ( \16161 , RI2b5e78495440_85, \15845 );
and \U$14398 ( \16162 , RI2b5e78494e28_98, \15847 );
and \U$14399 ( \16163 , RI2b5e78403928_111, \15849 );
and \U$14400 ( \16164 , RI2b5e775b1c08_124, \15851 );
and \U$14401 ( \16165 , RI2b5e7750bba0_137, \15853 );
and \U$14402 ( \16166 , RI2b5e774ff378_150, \15855 );
and \U$14403 ( \16167 , RI2b5e774f6390_163, \15857 );
and \U$14404 ( \16168 , RI2b5e774ea978_176, \15859 );
and \U$14405 ( \16169 , RI2b5e774de150_189, \15861 );
and \U$14406 ( \16170 , RI2b5e774d5168_202, \15863 );
and \U$14407 ( \16171 , RI2b5e785f40a8_215, \15865 );
and \U$14408 ( \16172 , RI2b5e785eb480_228, \15867 );
and \U$14409 ( \16173 , RI2b5e785da608_241, \15869 );
or \U$14410 ( \16174 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 );
_DC g17d0 ( \16175_nG17d0 , \16174 , \15888 );
buf \U$14411 ( \16176 , \16175_nG17d0 );
not \U$14412 ( \16177 , \16176 );
and \U$14413 ( \16178 , RI2b5e78549900_33, \15892 );
and \U$14414 ( \16179 , RI2b5e78538c68_46, \15894 );
and \U$14415 ( \16180 , RI2b5e78538650_59, \15896 );
and \U$14416 ( \16181 , RI2b5e784a60d8_72, \15898 );
and \U$14417 ( \16182 , RI2b5e78495440_85, \15900 );
and \U$14418 ( \16183 , RI2b5e78494e28_98, \15902 );
and \U$14419 ( \16184 , RI2b5e78403928_111, \15904 );
and \U$14420 ( \16185 , RI2b5e775b1c08_124, \15906 );
and \U$14421 ( \16186 , RI2b5e7750bba0_137, \15908 );
and \U$14422 ( \16187 , RI2b5e774ff378_150, \15910 );
and \U$14423 ( \16188 , RI2b5e774f6390_163, \15912 );
and \U$14424 ( \16189 , RI2b5e774ea978_176, \15914 );
and \U$14425 ( \16190 , RI2b5e774de150_189, \15916 );
and \U$14426 ( \16191 , RI2b5e774d5168_202, \15918 );
and \U$14427 ( \16192 , RI2b5e785f40a8_215, \15920 );
and \U$14428 ( \16193 , RI2b5e785eb480_228, \15922 );
and \U$14429 ( \16194 , RI2b5e785da608_241, \15924 );
or \U$14430 ( \16195 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 );
_DC g17e5 ( \16196_nG17e5 , \16195 , \15943 );
buf \U$14431 ( \16197 , \16196_nG17e5 );
and \U$14432 ( \16198 , \16177 , \16197 );
and \U$14433 ( \16199 , RI2b5e78549888_34, \15837 );
and \U$14434 ( \16200 , RI2b5e78538bf0_47, \15839 );
and \U$14435 ( \16201 , RI2b5e785385d8_60, \15841 );
and \U$14436 ( \16202 , RI2b5e784a6060_73, \15843 );
and \U$14437 ( \16203 , RI2b5e784953c8_86, \15845 );
and \U$14438 ( \16204 , RI2b5e78403ec8_99, \15847 );
and \U$14439 ( \16205 , RI2b5e775b21a8_112, \15849 );
and \U$14440 ( \16206 , RI2b5e775b1b90_125, \15851 );
and \U$14441 ( \16207 , RI2b5e7750bb28_138, \15853 );
and \U$14442 ( \16208 , RI2b5e774ff300_151, \15855 );
and \U$14443 ( \16209 , RI2b5e774f6318_164, \15857 );
and \U$14444 ( \16210 , RI2b5e774ea900_177, \15859 );
and \U$14445 ( \16211 , RI2b5e774de0d8_190, \15861 );
and \U$14446 ( \16212 , RI2b5e774d50f0_203, \15863 );
and \U$14447 ( \16213 , RI2b5e785f4030_216, \15865 );
and \U$14448 ( \16214 , RI2b5e785eb408_229, \15867 );
and \U$14449 ( \16215 , RI2b5e785da590_242, \15869 );
or \U$14450 ( \16216 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 );
_DC g17fa ( \16217_nG17fa , \16216 , \15888 );
buf \U$14451 ( \16218 , \16217_nG17fa );
not \U$14452 ( \16219 , \16218 );
and \U$14453 ( \16220 , RI2b5e78549888_34, \15892 );
and \U$14454 ( \16221 , RI2b5e78538bf0_47, \15894 );
and \U$14455 ( \16222 , RI2b5e785385d8_60, \15896 );
and \U$14456 ( \16223 , RI2b5e784a6060_73, \15898 );
and \U$14457 ( \16224 , RI2b5e784953c8_86, \15900 );
and \U$14458 ( \16225 , RI2b5e78403ec8_99, \15902 );
and \U$14459 ( \16226 , RI2b5e775b21a8_112, \15904 );
and \U$14460 ( \16227 , RI2b5e775b1b90_125, \15906 );
and \U$14461 ( \16228 , RI2b5e7750bb28_138, \15908 );
and \U$14462 ( \16229 , RI2b5e774ff300_151, \15910 );
and \U$14463 ( \16230 , RI2b5e774f6318_164, \15912 );
and \U$14464 ( \16231 , RI2b5e774ea900_177, \15914 );
and \U$14465 ( \16232 , RI2b5e774de0d8_190, \15916 );
and \U$14466 ( \16233 , RI2b5e774d50f0_203, \15918 );
and \U$14467 ( \16234 , RI2b5e785f4030_216, \15920 );
and \U$14468 ( \16235 , RI2b5e785eb408_229, \15922 );
and \U$14469 ( \16236 , RI2b5e785da590_242, \15924 );
or \U$14470 ( \16237 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 );
_DC g180f ( \16238_nG180f , \16237 , \15943 );
buf \U$14471 ( \16239 , \16238_nG180f );
and \U$14472 ( \16240 , \16219 , \16239 );
and \U$14473 ( \16241 , RI2b5e78549810_35, \15837 );
and \U$14474 ( \16242 , RI2b5e78538b78_48, \15839 );
and \U$14475 ( \16243 , RI2b5e78538560_61, \15841 );
and \U$14476 ( \16244 , RI2b5e784a5fe8_74, \15843 );
and \U$14477 ( \16245 , RI2b5e78495350_87, \15845 );
and \U$14478 ( \16246 , RI2b5e78403e50_100, \15847 );
and \U$14479 ( \16247 , RI2b5e775b2130_113, \15849 );
and \U$14480 ( \16248 , RI2b5e775b1b18_126, \15851 );
and \U$14481 ( \16249 , RI2b5e7750bab0_139, \15853 );
and \U$14482 ( \16250 , RI2b5e774ff288_152, \15855 );
and \U$14483 ( \16251 , RI2b5e774f62a0_165, \15857 );
and \U$14484 ( \16252 , RI2b5e774ea888_178, \15859 );
and \U$14485 ( \16253 , RI2b5e774de060_191, \15861 );
and \U$14486 ( \16254 , RI2b5e774d5078_204, \15863 );
and \U$14487 ( \16255 , RI2b5e785f3fb8_217, \15865 );
and \U$14488 ( \16256 , RI2b5e785eb390_230, \15867 );
and \U$14489 ( \16257 , RI2b5e785da518_243, \15869 );
or \U$14490 ( \16258 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 );
_DC g1824 ( \16259_nG1824 , \16258 , \15888 );
buf \U$14491 ( \16260 , \16259_nG1824 );
not \U$14492 ( \16261 , \16260 );
and \U$14493 ( \16262 , RI2b5e78549810_35, \15892 );
and \U$14494 ( \16263 , RI2b5e78538b78_48, \15894 );
and \U$14495 ( \16264 , RI2b5e78538560_61, \15896 );
and \U$14496 ( \16265 , RI2b5e784a5fe8_74, \15898 );
and \U$14497 ( \16266 , RI2b5e78495350_87, \15900 );
and \U$14498 ( \16267 , RI2b5e78403e50_100, \15902 );
and \U$14499 ( \16268 , RI2b5e775b2130_113, \15904 );
and \U$14500 ( \16269 , RI2b5e775b1b18_126, \15906 );
and \U$14501 ( \16270 , RI2b5e7750bab0_139, \15908 );
and \U$14502 ( \16271 , RI2b5e774ff288_152, \15910 );
and \U$14503 ( \16272 , RI2b5e774f62a0_165, \15912 );
and \U$14504 ( \16273 , RI2b5e774ea888_178, \15914 );
and \U$14505 ( \16274 , RI2b5e774de060_191, \15916 );
and \U$14506 ( \16275 , RI2b5e774d5078_204, \15918 );
and \U$14507 ( \16276 , RI2b5e785f3fb8_217, \15920 );
and \U$14508 ( \16277 , RI2b5e785eb390_230, \15922 );
and \U$14509 ( \16278 , RI2b5e785da518_243, \15924 );
or \U$14510 ( \16279 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 );
_DC g1839 ( \16280_nG1839 , \16279 , \15943 );
buf \U$14511 ( \16281 , \16280_nG1839 );
and \U$14512 ( \16282 , \16261 , \16281 );
and \U$14513 ( \16283 , RI2b5e78549798_36, \15837 );
and \U$14514 ( \16284 , RI2b5e78538b00_49, \15839 );
and \U$14515 ( \16285 , RI2b5e785384e8_62, \15841 );
and \U$14516 ( \16286 , RI2b5e784a5f70_75, \15843 );
and \U$14517 ( \16287 , RI2b5e784952d8_88, \15845 );
and \U$14518 ( \16288 , RI2b5e78403dd8_101, \15847 );
and \U$14519 ( \16289 , RI2b5e775b20b8_114, \15849 );
and \U$14520 ( \16290 , RI2b5e775b1aa0_127, \15851 );
and \U$14521 ( \16291 , RI2b5e7750ba38_140, \15853 );
and \U$14522 ( \16292 , RI2b5e774ff210_153, \15855 );
and \U$14523 ( \16293 , RI2b5e774f6228_166, \15857 );
and \U$14524 ( \16294 , RI2b5e774ea810_179, \15859 );
and \U$14525 ( \16295 , RI2b5e774ddfe8_192, \15861 );
and \U$14526 ( \16296 , RI2b5e774d5000_205, \15863 );
and \U$14527 ( \16297 , RI2b5e785f3f40_218, \15865 );
and \U$14528 ( \16298 , RI2b5e785eb318_231, \15867 );
and \U$14529 ( \16299 , RI2b5e785da4a0_244, \15869 );
or \U$14530 ( \16300 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 );
_DC g184e ( \16301_nG184e , \16300 , \15888 );
buf \U$14531 ( \16302 , \16301_nG184e );
not \U$14532 ( \16303 , \16302 );
and \U$14533 ( \16304 , RI2b5e78549798_36, \15892 );
and \U$14534 ( \16305 , RI2b5e78538b00_49, \15894 );
and \U$14535 ( \16306 , RI2b5e785384e8_62, \15896 );
and \U$14536 ( \16307 , RI2b5e784a5f70_75, \15898 );
and \U$14537 ( \16308 , RI2b5e784952d8_88, \15900 );
and \U$14538 ( \16309 , RI2b5e78403dd8_101, \15902 );
and \U$14539 ( \16310 , RI2b5e775b20b8_114, \15904 );
and \U$14540 ( \16311 , RI2b5e775b1aa0_127, \15906 );
and \U$14541 ( \16312 , RI2b5e7750ba38_140, \15908 );
and \U$14542 ( \16313 , RI2b5e774ff210_153, \15910 );
and \U$14543 ( \16314 , RI2b5e774f6228_166, \15912 );
and \U$14544 ( \16315 , RI2b5e774ea810_179, \15914 );
and \U$14545 ( \16316 , RI2b5e774ddfe8_192, \15916 );
and \U$14546 ( \16317 , RI2b5e774d5000_205, \15918 );
and \U$14547 ( \16318 , RI2b5e785f3f40_218, \15920 );
and \U$14548 ( \16319 , RI2b5e785eb318_231, \15922 );
and \U$14549 ( \16320 , RI2b5e785da4a0_244, \15924 );
or \U$14550 ( \16321 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 );
_DC g1863 ( \16322_nG1863 , \16321 , \15943 );
buf \U$14551 ( \16323 , \16322_nG1863 );
and \U$14552 ( \16324 , \16303 , \16323 );
and \U$14553 ( \16325 , RI2b5e78549720_37, \15837 );
and \U$14554 ( \16326 , RI2b5e78538a88_50, \15839 );
and \U$14555 ( \16327 , RI2b5e78538470_63, \15841 );
and \U$14556 ( \16328 , RI2b5e784a5ef8_76, \15843 );
and \U$14557 ( \16329 , RI2b5e78495260_89, \15845 );
and \U$14558 ( \16330 , RI2b5e78403d60_102, \15847 );
and \U$14559 ( \16331 , RI2b5e775b2040_115, \15849 );
and \U$14560 ( \16332 , RI2b5e775b1a28_128, \15851 );
and \U$14561 ( \16333 , RI2b5e7750b9c0_141, \15853 );
and \U$14562 ( \16334 , RI2b5e774ff198_154, \15855 );
and \U$14563 ( \16335 , RI2b5e774f61b0_167, \15857 );
and \U$14564 ( \16336 , RI2b5e774ea798_180, \15859 );
and \U$14565 ( \16337 , RI2b5e774ddf70_193, \15861 );
and \U$14566 ( \16338 , RI2b5e774d4f88_206, \15863 );
and \U$14567 ( \16339 , RI2b5e785f3ec8_219, \15865 );
and \U$14568 ( \16340 , RI2b5e785eb2a0_232, \15867 );
and \U$14569 ( \16341 , RI2b5e785da428_245, \15869 );
or \U$14570 ( \16342 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 );
_DC g1878 ( \16343_nG1878 , \16342 , \15888 );
buf \U$14571 ( \16344 , \16343_nG1878 );
not \U$14572 ( \16345 , \16344 );
and \U$14573 ( \16346 , RI2b5e78549720_37, \15892 );
and \U$14574 ( \16347 , RI2b5e78538a88_50, \15894 );
and \U$14575 ( \16348 , RI2b5e78538470_63, \15896 );
and \U$14576 ( \16349 , RI2b5e784a5ef8_76, \15898 );
and \U$14577 ( \16350 , RI2b5e78495260_89, \15900 );
and \U$14578 ( \16351 , RI2b5e78403d60_102, \15902 );
and \U$14579 ( \16352 , RI2b5e775b2040_115, \15904 );
and \U$14580 ( \16353 , RI2b5e775b1a28_128, \15906 );
and \U$14581 ( \16354 , RI2b5e7750b9c0_141, \15908 );
and \U$14582 ( \16355 , RI2b5e774ff198_154, \15910 );
and \U$14583 ( \16356 , RI2b5e774f61b0_167, \15912 );
and \U$14584 ( \16357 , RI2b5e774ea798_180, \15914 );
and \U$14585 ( \16358 , RI2b5e774ddf70_193, \15916 );
and \U$14586 ( \16359 , RI2b5e774d4f88_206, \15918 );
and \U$14587 ( \16360 , RI2b5e785f3ec8_219, \15920 );
and \U$14588 ( \16361 , RI2b5e785eb2a0_232, \15922 );
and \U$14589 ( \16362 , RI2b5e785da428_245, \15924 );
or \U$14590 ( \16363 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 );
_DC g188d ( \16364_nG188d , \16363 , \15943 );
buf \U$14591 ( \16365 , \16364_nG188d );
and \U$14592 ( \16366 , \16345 , \16365 );
and \U$14593 ( \16367 , RI2b5e785496a8_38, \15837 );
and \U$14594 ( \16368 , RI2b5e78538a10_51, \15839 );
and \U$14595 ( \16369 , RI2b5e785383f8_64, \15841 );
and \U$14596 ( \16370 , RI2b5e784a5e80_77, \15843 );
and \U$14597 ( \16371 , RI2b5e784951e8_90, \15845 );
and \U$14598 ( \16372 , RI2b5e78403ce8_103, \15847 );
and \U$14599 ( \16373 , RI2b5e775b1fc8_116, \15849 );
and \U$14600 ( \16374 , RI2b5e775b19b0_129, \15851 );
and \U$14601 ( \16375 , RI2b5e7750b948_142, \15853 );
and \U$14602 ( \16376 , RI2b5e774ff120_155, \15855 );
and \U$14603 ( \16377 , RI2b5e774f6138_168, \15857 );
and \U$14604 ( \16378 , RI2b5e774ea720_181, \15859 );
and \U$14605 ( \16379 , RI2b5e774ddef8_194, \15861 );
and \U$14606 ( \16380 , RI2b5e774d4f10_207, \15863 );
and \U$14607 ( \16381 , RI2b5e785f3e50_220, \15865 );
and \U$14608 ( \16382 , RI2b5e785eb228_233, \15867 );
and \U$14609 ( \16383 , RI2b5e785da3b0_246, \15869 );
or \U$14610 ( \16384 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 );
_DC g18a2 ( \16385_nG18a2 , \16384 , \15888 );
buf \U$14611 ( \16386 , \16385_nG18a2 );
not \U$14612 ( \16387 , \16386 );
and \U$14613 ( \16388 , RI2b5e785496a8_38, \15892 );
and \U$14614 ( \16389 , RI2b5e78538a10_51, \15894 );
and \U$14615 ( \16390 , RI2b5e785383f8_64, \15896 );
and \U$14616 ( \16391 , RI2b5e784a5e80_77, \15898 );
and \U$14617 ( \16392 , RI2b5e784951e8_90, \15900 );
and \U$14618 ( \16393 , RI2b5e78403ce8_103, \15902 );
and \U$14619 ( \16394 , RI2b5e775b1fc8_116, \15904 );
and \U$14620 ( \16395 , RI2b5e775b19b0_129, \15906 );
and \U$14621 ( \16396 , RI2b5e7750b948_142, \15908 );
and \U$14622 ( \16397 , RI2b5e774ff120_155, \15910 );
and \U$14623 ( \16398 , RI2b5e774f6138_168, \15912 );
and \U$14624 ( \16399 , RI2b5e774ea720_181, \15914 );
and \U$14625 ( \16400 , RI2b5e774ddef8_194, \15916 );
and \U$14626 ( \16401 , RI2b5e774d4f10_207, \15918 );
and \U$14627 ( \16402 , RI2b5e785f3e50_220, \15920 );
and \U$14628 ( \16403 , RI2b5e785eb228_233, \15922 );
and \U$14629 ( \16404 , RI2b5e785da3b0_246, \15924 );
or \U$14630 ( \16405 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 );
_DC g18b7 ( \16406_nG18b7 , \16405 , \15943 );
buf \U$14631 ( \16407 , \16406_nG18b7 );
and \U$14632 ( \16408 , \16387 , \16407 );
and \U$14633 ( \16409 , RI2b5e78549630_39, \15837 );
and \U$14634 ( \16410 , RI2b5e78538998_52, \15839 );
and \U$14635 ( \16411 , RI2b5e78538380_65, \15841 );
and \U$14636 ( \16412 , RI2b5e784a5e08_78, \15843 );
and \U$14637 ( \16413 , RI2b5e78495170_91, \15845 );
and \U$14638 ( \16414 , RI2b5e78403c70_104, \15847 );
and \U$14639 ( \16415 , RI2b5e775b1f50_117, \15849 );
and \U$14640 ( \16416 , RI2b5e775b1938_130, \15851 );
and \U$14641 ( \16417 , RI2b5e7750b8d0_143, \15853 );
and \U$14642 ( \16418 , RI2b5e774ff0a8_156, \15855 );
and \U$14643 ( \16419 , RI2b5e774f60c0_169, \15857 );
and \U$14644 ( \16420 , RI2b5e774ea6a8_182, \15859 );
and \U$14645 ( \16421 , RI2b5e774dde80_195, \15861 );
and \U$14646 ( \16422 , RI2b5e774d4e98_208, \15863 );
and \U$14647 ( \16423 , RI2b5e785f3dd8_221, \15865 );
and \U$14648 ( \16424 , RI2b5e785eb1b0_234, \15867 );
and \U$14649 ( \16425 , RI2b5e785da338_247, \15869 );
or \U$14650 ( \16426 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 );
_DC g18cc ( \16427_nG18cc , \16426 , \15888 );
buf \U$14651 ( \16428 , \16427_nG18cc );
not \U$14652 ( \16429 , \16428 );
and \U$14653 ( \16430 , RI2b5e78549630_39, \15892 );
and \U$14654 ( \16431 , RI2b5e78538998_52, \15894 );
and \U$14655 ( \16432 , RI2b5e78538380_65, \15896 );
and \U$14656 ( \16433 , RI2b5e784a5e08_78, \15898 );
and \U$14657 ( \16434 , RI2b5e78495170_91, \15900 );
and \U$14658 ( \16435 , RI2b5e78403c70_104, \15902 );
and \U$14659 ( \16436 , RI2b5e775b1f50_117, \15904 );
and \U$14660 ( \16437 , RI2b5e775b1938_130, \15906 );
and \U$14661 ( \16438 , RI2b5e7750b8d0_143, \15908 );
and \U$14662 ( \16439 , RI2b5e774ff0a8_156, \15910 );
and \U$14663 ( \16440 , RI2b5e774f60c0_169, \15912 );
and \U$14664 ( \16441 , RI2b5e774ea6a8_182, \15914 );
and \U$14665 ( \16442 , RI2b5e774dde80_195, \15916 );
and \U$14666 ( \16443 , RI2b5e774d4e98_208, \15918 );
and \U$14667 ( \16444 , RI2b5e785f3dd8_221, \15920 );
and \U$14668 ( \16445 , RI2b5e785eb1b0_234, \15922 );
and \U$14669 ( \16446 , RI2b5e785da338_247, \15924 );
or \U$14670 ( \16447 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 );
_DC g18e1 ( \16448_nG18e1 , \16447 , \15943 );
buf \U$14671 ( \16449 , \16448_nG18e1 );
and \U$14672 ( \16450 , \16429 , \16449 );
xnor \U$14673 ( \16451 , \16407 , \16386 );
and \U$14674 ( \16452 , \16450 , \16451 );
or \U$14675 ( \16453 , \16408 , \16452 );
xnor \U$14676 ( \16454 , \16365 , \16344 );
and \U$14677 ( \16455 , \16453 , \16454 );
or \U$14678 ( \16456 , \16366 , \16455 );
xnor \U$14679 ( \16457 , \16323 , \16302 );
and \U$14680 ( \16458 , \16456 , \16457 );
or \U$14681 ( \16459 , \16324 , \16458 );
xnor \U$14682 ( \16460 , \16281 , \16260 );
and \U$14683 ( \16461 , \16459 , \16460 );
or \U$14684 ( \16462 , \16282 , \16461 );
xnor \U$14685 ( \16463 , \16239 , \16218 );
and \U$14686 ( \16464 , \16462 , \16463 );
or \U$14687 ( \16465 , \16240 , \16464 );
xnor \U$14688 ( \16466 , \16197 , \16176 );
and \U$14689 ( \16467 , \16465 , \16466 );
or \U$14690 ( \16468 , \16198 , \16467 );
xnor \U$14691 ( \16469 , \16155 , \16134 );
and \U$14692 ( \16470 , \16468 , \16469 );
or \U$14693 ( \16471 , \16156 , \16470 );
xnor \U$14694 ( \16472 , \16113 , \16092 );
and \U$14695 ( \16473 , \16471 , \16472 );
or \U$14696 ( \16474 , \16114 , \16473 );
xnor \U$14697 ( \16475 , \16071 , \16050 );
and \U$14698 ( \16476 , \16474 , \16475 );
or \U$14699 ( \16477 , \16072 , \16476 );
xnor \U$14700 ( \16478 , \16029 , \16008 );
and \U$14701 ( \16479 , \16477 , \16478 );
or \U$14702 ( \16480 , \16030 , \16479 );
xnor \U$14703 ( \16481 , \15987 , \15966 );
and \U$14704 ( \16482 , \16480 , \16481 );
or \U$14705 ( \16483 , \15988 , \16482 );
xnor \U$14706 ( \16484 , \15945 , \15890 );
and \U$14707 ( \16485 , \16483 , \16484 );
or \U$14708 ( \16486 , \15946 , \16485 );
buf \U$14709 ( \16487 , \16486 );
and \U$14710 ( \16488 , \15836 , \16487 );
_HMUX g4ba1_GF_PartitionCandidate ( \16489_nG4ba1 , \12552_nG4b72 , \15398_nG4ba0 , \16488 );
buf \U$14711 ( \16490 , \16489_nG4ba1 );
not \U$14712 ( \16491 , \12015 );
nand \U$14713 ( \16492 , \12544 , \16491 );
nor \U$14714 ( \16493 , \12362 , \11198 );
nor \U$14715 ( \16494 , \11273 , \11350 );
nand \U$14716 ( \16495 , \16493 , \16494 );
nor \U$14717 ( \16496 , \11425 , \11502 );
nor \U$14718 ( \16497 , \11578 , \11651 );
nand \U$14719 ( \16498 , \16496 , \16497 );
nor \U$14720 ( \16499 , \16495 , \16498 );
nor \U$14721 ( \16500 , \11720 , \11784 );
nor \U$14722 ( \16501 , \11844 , \11901 );
nand \U$14723 ( \16502 , \16500 , \16501 );
nor \U$14724 ( \16503 , \11939 , \11971 );
nor \U$14725 ( \16504 , \11992 , \12008 );
nand \U$14726 ( \16505 , \16503 , \16504 );
nor \U$14727 ( \16506 , \16502 , \16505 );
nand \U$14728 ( \16507 , \16499 , \16506 );
nor \U$14729 ( \16508 , \12423 , \12127 );
nor \U$14730 ( \16509 , \12172 , \12224 );
nand \U$14731 ( \16510 , \16508 , \16509 );
nor \U$14732 ( \16511 , \12279 , \12318 );
nor \U$14733 ( \16512 , \12339 , \12355 );
nand \U$14734 ( \16513 , \16511 , \16512 );
nor \U$14735 ( \16514 , \16510 , \16513 );
nor \U$14736 ( \16515 , \12443 , \12398 );
nor \U$14737 ( \16516 , \12409 , \12420 );
nand \U$14738 ( \16517 , \16515 , \16516 );
nor \U$14739 ( \16518 , \12448 , \12440 );
not \U$14740 ( \16519 , \12456 );
and \U$14741 ( \16520 , \16518 , \16519 );
or \U$14742 ( \16521 , \12440 , \12458 );
nand \U$14743 ( \16522 , \16521 , \12461 );
nor \U$14744 ( \16523 , \16520 , \16522 );
or \U$14745 ( \16524 , \16517 , \16523 );
or \U$14746 ( \16525 , \12398 , \12463 );
nand \U$14747 ( \16526 , \16525 , \12467 );
and \U$14748 ( \16527 , \16516 , \16526 );
or \U$14749 ( \16528 , \12420 , \12469 );
nand \U$14750 ( \16529 , \16528 , \12472 );
nor \U$14751 ( \16530 , \16527 , \16529 );
nand \U$14752 ( \16531 , \16524 , \16530 );
and \U$14753 ( \16532 , \16514 , \16531 );
or \U$14754 ( \16533 , \12127 , \12474 );
nand \U$14755 ( \16534 , \16533 , \12479 );
and \U$14756 ( \16535 , \16509 , \16534 );
or \U$14757 ( \16536 , \12224 , \12481 );
nand \U$14758 ( \16537 , \16536 , \12484 );
nor \U$14759 ( \16538 , \16535 , \16537 );
or \U$14760 ( \16539 , \16513 , \16538 );
or \U$14761 ( \16540 , \12318 , \12486 );
nand \U$14762 ( \16541 , \16540 , \12490 );
and \U$14763 ( \16542 , \16512 , \16541 );
or \U$14764 ( \16543 , \12355 , \12492 );
nand \U$14765 ( \16544 , \16543 , \12495 );
nor \U$14766 ( \16545 , \16542 , \16544 );
nand \U$14767 ( \16546 , \16539 , \16545 );
nor \U$14768 ( \16547 , \16532 , \16546 );
or \U$14769 ( \16548 , \16507 , \16547 );
or \U$14770 ( \16549 , \11198 , \12497 );
nand \U$14771 ( \16550 , \16549 , \12503 );
and \U$14772 ( \16551 , \16494 , \16550 );
or \U$14773 ( \16552 , \11350 , \12505 );
nand \U$14774 ( \16553 , \16552 , \12508 );
nor \U$14775 ( \16554 , \16551 , \16553 );
or \U$14776 ( \16555 , \16498 , \16554 );
or \U$14777 ( \16556 , \11502 , \12510 );
nand \U$14778 ( \16557 , \16556 , \12514 );
and \U$14779 ( \16558 , \16497 , \16557 );
or \U$14780 ( \16559 , \11651 , \12516 );
nand \U$14781 ( \16560 , \16559 , \12519 );
nor \U$14782 ( \16561 , \16558 , \16560 );
nand \U$14783 ( \16562 , \16555 , \16561 );
and \U$14784 ( \16563 , \16506 , \16562 );
or \U$14785 ( \16564 , \11784 , \12521 );
nand \U$14786 ( \16565 , \16564 , \12526 );
and \U$14787 ( \16566 , \16501 , \16565 );
or \U$14788 ( \16567 , \11901 , \12528 );
nand \U$14789 ( \16568 , \16567 , \12531 );
nor \U$14790 ( \16569 , \16566 , \16568 );
or \U$14791 ( \16570 , \16505 , \16569 );
or \U$14792 ( \16571 , \11971 , \12533 );
nand \U$14793 ( \16572 , \16571 , \12537 );
and \U$14794 ( \16573 , \16504 , \16572 );
or \U$14795 ( \16574 , \12008 , \12539 );
nand \U$14796 ( \16575 , \16574 , \12542 );
nor \U$14797 ( \16576 , \16573 , \16575 );
nand \U$14798 ( \16577 , \16570 , \16576 );
nor \U$14799 ( \16578 , \16563 , \16577 );
nand \U$14800 ( \16579 , \16548 , \16578 );
not \U$14801 ( \16580 , \16579 );
xor \U$14802 ( \16581 , \16492 , \16580 );
buf g4b0f_GF_PartitionCandidate( \16582_nG4b0f , \16581 );
not \U$14803 ( \16583 , \14861 );
nand \U$14804 ( \16584 , \15390 , \16583 );
nor \U$14805 ( \16585 , \15208 , \14044 );
nor \U$14806 ( \16586 , \14119 , \14196 );
nand \U$14807 ( \16587 , \16585 , \16586 );
nor \U$14808 ( \16588 , \14271 , \14348 );
nor \U$14809 ( \16589 , \14424 , \14497 );
nand \U$14810 ( \16590 , \16588 , \16589 );
nor \U$14811 ( \16591 , \16587 , \16590 );
nor \U$14812 ( \16592 , \14566 , \14630 );
nor \U$14813 ( \16593 , \14690 , \14747 );
nand \U$14814 ( \16594 , \16592 , \16593 );
nor \U$14815 ( \16595 , \14785 , \14817 );
nor \U$14816 ( \16596 , \14838 , \14854 );
nand \U$14817 ( \16597 , \16595 , \16596 );
nor \U$14818 ( \16598 , \16594 , \16597 );
nand \U$14819 ( \16599 , \16591 , \16598 );
nor \U$14820 ( \16600 , \15269 , \14973 );
nor \U$14821 ( \16601 , \15018 , \15070 );
nand \U$14822 ( \16602 , \16600 , \16601 );
nor \U$14823 ( \16603 , \15125 , \15164 );
nor \U$14824 ( \16604 , \15185 , \15201 );
nand \U$14825 ( \16605 , \16603 , \16604 );
nor \U$14826 ( \16606 , \16602 , \16605 );
nor \U$14827 ( \16607 , \15289 , \15244 );
nor \U$14828 ( \16608 , \15255 , \15266 );
nand \U$14829 ( \16609 , \16607 , \16608 );
nor \U$14830 ( \16610 , \15294 , \15286 );
not \U$14831 ( \16611 , \15302 );
and \U$14832 ( \16612 , \16610 , \16611 );
or \U$14833 ( \16613 , \15286 , \15304 );
nand \U$14834 ( \16614 , \16613 , \15307 );
nor \U$14835 ( \16615 , \16612 , \16614 );
or \U$14836 ( \16616 , \16609 , \16615 );
or \U$14837 ( \16617 , \15244 , \15309 );
nand \U$14838 ( \16618 , \16617 , \15313 );
and \U$14839 ( \16619 , \16608 , \16618 );
or \U$14840 ( \16620 , \15266 , \15315 );
nand \U$14841 ( \16621 , \16620 , \15318 );
nor \U$14842 ( \16622 , \16619 , \16621 );
nand \U$14843 ( \16623 , \16616 , \16622 );
and \U$14844 ( \16624 , \16606 , \16623 );
or \U$14845 ( \16625 , \14973 , \15320 );
nand \U$14846 ( \16626 , \16625 , \15325 );
and \U$14847 ( \16627 , \16601 , \16626 );
or \U$14848 ( \16628 , \15070 , \15327 );
nand \U$14849 ( \16629 , \16628 , \15330 );
nor \U$14850 ( \16630 , \16627 , \16629 );
or \U$14851 ( \16631 , \16605 , \16630 );
or \U$14852 ( \16632 , \15164 , \15332 );
nand \U$14853 ( \16633 , \16632 , \15336 );
and \U$14854 ( \16634 , \16604 , \16633 );
or \U$14855 ( \16635 , \15201 , \15338 );
nand \U$14856 ( \16636 , \16635 , \15341 );
nor \U$14857 ( \16637 , \16634 , \16636 );
nand \U$14858 ( \16638 , \16631 , \16637 );
nor \U$14859 ( \16639 , \16624 , \16638 );
or \U$14860 ( \16640 , \16599 , \16639 );
or \U$14861 ( \16641 , \14044 , \15343 );
nand \U$14862 ( \16642 , \16641 , \15349 );
and \U$14863 ( \16643 , \16586 , \16642 );
or \U$14864 ( \16644 , \14196 , \15351 );
nand \U$14865 ( \16645 , \16644 , \15354 );
nor \U$14866 ( \16646 , \16643 , \16645 );
or \U$14867 ( \16647 , \16590 , \16646 );
or \U$14868 ( \16648 , \14348 , \15356 );
nand \U$14869 ( \16649 , \16648 , \15360 );
and \U$14870 ( \16650 , \16589 , \16649 );
or \U$14871 ( \16651 , \14497 , \15362 );
nand \U$14872 ( \16652 , \16651 , \15365 );
nor \U$14873 ( \16653 , \16650 , \16652 );
nand \U$14874 ( \16654 , \16647 , \16653 );
and \U$14875 ( \16655 , \16598 , \16654 );
or \U$14876 ( \16656 , \14630 , \15367 );
nand \U$14877 ( \16657 , \16656 , \15372 );
and \U$14878 ( \16658 , \16593 , \16657 );
or \U$14879 ( \16659 , \14747 , \15374 );
nand \U$14880 ( \16660 , \16659 , \15377 );
nor \U$14881 ( \16661 , \16658 , \16660 );
or \U$14882 ( \16662 , \16597 , \16661 );
or \U$14883 ( \16663 , \14817 , \15379 );
nand \U$14884 ( \16664 , \16663 , \15383 );
and \U$14885 ( \16665 , \16596 , \16664 );
or \U$14886 ( \16666 , \14854 , \15385 );
nand \U$14887 ( \16667 , \16666 , \15388 );
nor \U$14888 ( \16668 , \16665 , \16667 );
nand \U$14889 ( \16669 , \16662 , \16668 );
nor \U$14890 ( \16670 , \16655 , \16669 );
nand \U$14891 ( \16671 , \16640 , \16670 );
not \U$14892 ( \16672 , \16671 );
xor \U$14893 ( \16673 , \16584 , \16672 );
buf g4b43_GF_PartitionCandidate( \16674_nG4b43 , \16673 );
_HMUX g4b44_GF_PartitionCandidate ( \16675_nG4b44 , \16582_nG4b0f , \16674_nG4b43 , \16488 );
buf \U$14894 ( \16676 , \16675_nG4b44 );
not \U$14895 ( \16677 , \12008 );
nand \U$14896 ( \16678 , \12542 , \16677 );
nand \U$14897 ( \16679 , \12363 , \11274 );
nand \U$14898 ( \16680 , \11426 , \11579 );
nor \U$14899 ( \16681 , \16679 , \16680 );
nand \U$14900 ( \16682 , \11721 , \11845 );
nand \U$14901 ( \16683 , \11940 , \11993 );
nor \U$14902 ( \16684 , \16682 , \16683 );
nand \U$14903 ( \16685 , \16681 , \16684 );
nand \U$14904 ( \16686 , \12424 , \12173 );
nand \U$14905 ( \16687 , \12280 , \12340 );
nor \U$14906 ( \16688 , \16686 , \16687 );
nand \U$14907 ( \16689 , \12444 , \12410 );
not \U$14908 ( \16690 , \12459 );
or \U$14909 ( \16691 , \16689 , \16690 );
and \U$14910 ( \16692 , \12410 , \12464 );
nor \U$14911 ( \16693 , \16692 , \12470 );
nand \U$14912 ( \16694 , \16691 , \16693 );
and \U$14913 ( \16695 , \16688 , \16694 );
and \U$14914 ( \16696 , \12173 , \12475 );
nor \U$14915 ( \16697 , \16696 , \12482 );
or \U$14916 ( \16698 , \16687 , \16697 );
and \U$14917 ( \16699 , \12340 , \12487 );
nor \U$14918 ( \16700 , \16699 , \12493 );
nand \U$14919 ( \16701 , \16698 , \16700 );
nor \U$14920 ( \16702 , \16695 , \16701 );
or \U$14921 ( \16703 , \16685 , \16702 );
and \U$14922 ( \16704 , \11274 , \12498 );
nor \U$14923 ( \16705 , \16704 , \12506 );
or \U$14924 ( \16706 , \16680 , \16705 );
and \U$14925 ( \16707 , \11579 , \12511 );
nor \U$14926 ( \16708 , \16707 , \12517 );
nand \U$14927 ( \16709 , \16706 , \16708 );
and \U$14928 ( \16710 , \16684 , \16709 );
and \U$14929 ( \16711 , \11845 , \12522 );
nor \U$14930 ( \16712 , \16711 , \12529 );
or \U$14931 ( \16713 , \16683 , \16712 );
and \U$14932 ( \16714 , \11993 , \12534 );
nor \U$14933 ( \16715 , \16714 , \12540 );
nand \U$14934 ( \16716 , \16713 , \16715 );
nor \U$14935 ( \16717 , \16710 , \16716 );
nand \U$14936 ( \16718 , \16703 , \16717 );
not \U$14937 ( \16719 , \16718 );
xor \U$14938 ( \16720 , \16678 , \16719 );
buf g4aa0_GF_PartitionCandidate( \16721_nG4aa0 , \16720 );
not \U$14939 ( \16722 , \14854 );
nand \U$14940 ( \16723 , \15388 , \16722 );
nand \U$14941 ( \16724 , \15209 , \14120 );
nand \U$14942 ( \16725 , \14272 , \14425 );
nor \U$14943 ( \16726 , \16724 , \16725 );
nand \U$14944 ( \16727 , \14567 , \14691 );
nand \U$14945 ( \16728 , \14786 , \14839 );
nor \U$14946 ( \16729 , \16727 , \16728 );
nand \U$14947 ( \16730 , \16726 , \16729 );
nand \U$14948 ( \16731 , \15270 , \15019 );
nand \U$14949 ( \16732 , \15126 , \15186 );
nor \U$14950 ( \16733 , \16731 , \16732 );
nand \U$14951 ( \16734 , \15290 , \15256 );
not \U$14952 ( \16735 , \15305 );
or \U$14953 ( \16736 , \16734 , \16735 );
and \U$14954 ( \16737 , \15256 , \15310 );
nor \U$14955 ( \16738 , \16737 , \15316 );
nand \U$14956 ( \16739 , \16736 , \16738 );
and \U$14957 ( \16740 , \16733 , \16739 );
and \U$14958 ( \16741 , \15019 , \15321 );
nor \U$14959 ( \16742 , \16741 , \15328 );
or \U$14960 ( \16743 , \16732 , \16742 );
and \U$14961 ( \16744 , \15186 , \15333 );
nor \U$14962 ( \16745 , \16744 , \15339 );
nand \U$14963 ( \16746 , \16743 , \16745 );
nor \U$14964 ( \16747 , \16740 , \16746 );
or \U$14965 ( \16748 , \16730 , \16747 );
and \U$14966 ( \16749 , \14120 , \15344 );
nor \U$14967 ( \16750 , \16749 , \15352 );
or \U$14968 ( \16751 , \16725 , \16750 );
and \U$14969 ( \16752 , \14425 , \15357 );
nor \U$14970 ( \16753 , \16752 , \15363 );
nand \U$14971 ( \16754 , \16751 , \16753 );
and \U$14972 ( \16755 , \16729 , \16754 );
and \U$14973 ( \16756 , \14691 , \15368 );
nor \U$14974 ( \16757 , \16756 , \15375 );
or \U$14975 ( \16758 , \16728 , \16757 );
and \U$14976 ( \16759 , \14839 , \15380 );
nor \U$14977 ( \16760 , \16759 , \15386 );
nand \U$14978 ( \16761 , \16758 , \16760 );
nor \U$14979 ( \16762 , \16755 , \16761 );
nand \U$14980 ( \16763 , \16748 , \16762 );
not \U$14981 ( \16764 , \16763 );
xor \U$14982 ( \16765 , \16723 , \16764 );
buf g4ada_GF_PartitionCandidate( \16766_nG4ada , \16765 );
_HMUX g4adb_GF_PartitionCandidate ( \16767_nG4adb , \16721_nG4aa0 , \16766_nG4ada , \16488 );
buf \U$14983 ( \16768 , \16767_nG4adb );
not \U$14984 ( \16769 , \11992 );
nand \U$14985 ( \16770 , \12539 , \16769 );
nand \U$14986 ( \16771 , \16512 , \16493 );
nand \U$14987 ( \16772 , \16494 , \16496 );
nor \U$14988 ( \16773 , \16771 , \16772 );
nand \U$14989 ( \16774 , \16497 , \16500 );
nand \U$14990 ( \16775 , \16501 , \16503 );
nor \U$14991 ( \16776 , \16774 , \16775 );
nand \U$14992 ( \16777 , \16773 , \16776 );
nand \U$14993 ( \16778 , \16516 , \16508 );
nand \U$14994 ( \16779 , \16509 , \16511 );
nor \U$14995 ( \16780 , \16778 , \16779 );
nand \U$14996 ( \16781 , \16518 , \16515 );
or \U$14997 ( \16782 , \16781 , \12456 );
and \U$14998 ( \16783 , \16515 , \16522 );
nor \U$14999 ( \16784 , \16783 , \16526 );
nand \U$15000 ( \16785 , \16782 , \16784 );
and \U$15001 ( \16786 , \16780 , \16785 );
and \U$15002 ( \16787 , \16508 , \16529 );
nor \U$15003 ( \16788 , \16787 , \16534 );
or \U$15004 ( \16789 , \16779 , \16788 );
and \U$15005 ( \16790 , \16511 , \16537 );
nor \U$15006 ( \16791 , \16790 , \16541 );
nand \U$15007 ( \16792 , \16789 , \16791 );
nor \U$15008 ( \16793 , \16786 , \16792 );
or \U$15009 ( \16794 , \16777 , \16793 );
and \U$15010 ( \16795 , \16493 , \16544 );
nor \U$15011 ( \16796 , \16795 , \16550 );
or \U$15012 ( \16797 , \16772 , \16796 );
and \U$15013 ( \16798 , \16496 , \16553 );
nor \U$15014 ( \16799 , \16798 , \16557 );
nand \U$15015 ( \16800 , \16797 , \16799 );
and \U$15016 ( \16801 , \16776 , \16800 );
and \U$15017 ( \16802 , \16500 , \16560 );
nor \U$15018 ( \16803 , \16802 , \16565 );
or \U$15019 ( \16804 , \16775 , \16803 );
and \U$15020 ( \16805 , \16503 , \16568 );
nor \U$15021 ( \16806 , \16805 , \16572 );
nand \U$15022 ( \16807 , \16804 , \16806 );
nor \U$15023 ( \16808 , \16801 , \16807 );
nand \U$15024 ( \16809 , \16794 , \16808 );
not \U$15025 ( \16810 , \16809 );
xor \U$15026 ( \16811 , \16770 , \16810 );
buf g4a23_GF_PartitionCandidate( \16812_nG4a23 , \16811 );
not \U$15027 ( \16813 , \14838 );
nand \U$15028 ( \16814 , \15385 , \16813 );
nand \U$15029 ( \16815 , \16604 , \16585 );
nand \U$15030 ( \16816 , \16586 , \16588 );
nor \U$15031 ( \16817 , \16815 , \16816 );
nand \U$15032 ( \16818 , \16589 , \16592 );
nand \U$15033 ( \16819 , \16593 , \16595 );
nor \U$15034 ( \16820 , \16818 , \16819 );
nand \U$15035 ( \16821 , \16817 , \16820 );
nand \U$15036 ( \16822 , \16608 , \16600 );
nand \U$15037 ( \16823 , \16601 , \16603 );
nor \U$15038 ( \16824 , \16822 , \16823 );
nand \U$15039 ( \16825 , \16610 , \16607 );
or \U$15040 ( \16826 , \16825 , \15302 );
and \U$15041 ( \16827 , \16607 , \16614 );
nor \U$15042 ( \16828 , \16827 , \16618 );
nand \U$15043 ( \16829 , \16826 , \16828 );
and \U$15044 ( \16830 , \16824 , \16829 );
and \U$15045 ( \16831 , \16600 , \16621 );
nor \U$15046 ( \16832 , \16831 , \16626 );
or \U$15047 ( \16833 , \16823 , \16832 );
and \U$15048 ( \16834 , \16603 , \16629 );
nor \U$15049 ( \16835 , \16834 , \16633 );
nand \U$15050 ( \16836 , \16833 , \16835 );
nor \U$15051 ( \16837 , \16830 , \16836 );
or \U$15052 ( \16838 , \16821 , \16837 );
and \U$15053 ( \16839 , \16585 , \16636 );
nor \U$15054 ( \16840 , \16839 , \16642 );
or \U$15055 ( \16841 , \16816 , \16840 );
and \U$15056 ( \16842 , \16588 , \16645 );
nor \U$15057 ( \16843 , \16842 , \16649 );
nand \U$15058 ( \16844 , \16841 , \16843 );
and \U$15059 ( \16845 , \16820 , \16844 );
and \U$15060 ( \16846 , \16592 , \16652 );
nor \U$15061 ( \16847 , \16846 , \16657 );
or \U$15062 ( \16848 , \16819 , \16847 );
and \U$15063 ( \16849 , \16595 , \16660 );
nor \U$15064 ( \16850 , \16849 , \16664 );
nand \U$15065 ( \16851 , \16848 , \16850 );
nor \U$15066 ( \16852 , \16845 , \16851 );
nand \U$15067 ( \16853 , \16838 , \16852 );
not \U$15068 ( \16854 , \16853 );
xor \U$15069 ( \16855 , \16814 , \16854 );
buf g4a65_GF_PartitionCandidate( \16856_nG4a65 , \16855 );
_HMUX g4a66_GF_PartitionCandidate ( \16857_nG4a66 , \16812_nG4a23 , \16856_nG4a65 , \16488 );
buf \U$15070 ( \16858 , \16857_nG4a66 );
not \U$15071 ( \16859 , \11971 );
nand \U$15072 ( \16860 , \12537 , \16859 );
nor \U$15073 ( \16861 , \12364 , \11427 );
nor \U$15074 ( \16862 , \11722 , \11941 );
nand \U$15075 ( \16863 , \16861 , \16862 );
nor \U$15076 ( \16864 , \12425 , \12281 );
not \U$15077 ( \16865 , \12465 );
and \U$15078 ( \16866 , \16864 , \16865 );
or \U$15079 ( \16867 , \12281 , \12476 );
nand \U$15080 ( \16868 , \16867 , \12488 );
nor \U$15081 ( \16869 , \16866 , \16868 );
or \U$15082 ( \16870 , \16863 , \16869 );
or \U$15083 ( \16871 , \11427 , \12499 );
nand \U$15084 ( \16872 , \16871 , \12512 );
and \U$15085 ( \16873 , \16862 , \16872 );
or \U$15086 ( \16874 , \11941 , \12523 );
nand \U$15087 ( \16875 , \16874 , \12535 );
nor \U$15088 ( \16876 , \16873 , \16875 );
nand \U$15089 ( \16877 , \16870 , \16876 );
not \U$15090 ( \16878 , \16877 );
xor \U$15091 ( \16879 , \16860 , \16878 );
buf g499a_GF_PartitionCandidate( \16880_nG499a , \16879 );
not \U$15092 ( \16881 , \14817 );
nand \U$15093 ( \16882 , \15383 , \16881 );
nor \U$15094 ( \16883 , \15210 , \14273 );
nor \U$15095 ( \16884 , \14568 , \14787 );
nand \U$15096 ( \16885 , \16883 , \16884 );
nor \U$15097 ( \16886 , \15271 , \15127 );
not \U$15098 ( \16887 , \15311 );
and \U$15099 ( \16888 , \16886 , \16887 );
or \U$15100 ( \16889 , \15127 , \15322 );
nand \U$15101 ( \16890 , \16889 , \15334 );
nor \U$15102 ( \16891 , \16888 , \16890 );
or \U$15103 ( \16892 , \16885 , \16891 );
or \U$15104 ( \16893 , \14273 , \15345 );
nand \U$15105 ( \16894 , \16893 , \15358 );
and \U$15106 ( \16895 , \16884 , \16894 );
or \U$15107 ( \16896 , \14787 , \15369 );
nand \U$15108 ( \16897 , \16896 , \15381 );
nor \U$15109 ( \16898 , \16895 , \16897 );
nand \U$15110 ( \16899 , \16892 , \16898 );
not \U$15111 ( \16900 , \16899 );
xor \U$15112 ( \16901 , \16882 , \16900 );
buf g49e0_GF_PartitionCandidate( \16902_nG49e0 , \16901 );
_HMUX g49e1_GF_PartitionCandidate ( \16903_nG49e1 , \16880_nG499a , \16902_nG49e0 , \16488 );
buf \U$15113 ( \16904 , \16903_nG49e1 );
not \U$15114 ( \16905 , \11939 );
nand \U$15115 ( \16906 , \12533 , \16905 );
nor \U$15116 ( \16907 , \16513 , \16495 );
nor \U$15117 ( \16908 , \16498 , \16502 );
nand \U$15118 ( \16909 , \16907 , \16908 );
nor \U$15119 ( \16910 , \16517 , \16510 );
not \U$15120 ( \16911 , \16523 );
and \U$15121 ( \16912 , \16910 , \16911 );
or \U$15122 ( \16913 , \16510 , \16530 );
nand \U$15123 ( \16914 , \16913 , \16538 );
nor \U$15124 ( \16915 , \16912 , \16914 );
or \U$15125 ( \16916 , \16909 , \16915 );
or \U$15126 ( \16917 , \16495 , \16545 );
nand \U$15127 ( \16918 , \16917 , \16554 );
and \U$15128 ( \16919 , \16908 , \16918 );
or \U$15129 ( \16920 , \16502 , \16561 );
nand \U$15130 ( \16921 , \16920 , \16569 );
nor \U$15131 ( \16922 , \16919 , \16921 );
nand \U$15132 ( \16923 , \16916 , \16922 );
not \U$15133 ( \16924 , \16923 );
xor \U$15134 ( \16925 , \16906 , \16924 );
buf g490b_GF_PartitionCandidate( \16926_nG490b , \16925 );
not \U$15135 ( \16927 , \14785 );
nand \U$15136 ( \16928 , \15379 , \16927 );
nor \U$15137 ( \16929 , \16605 , \16587 );
nor \U$15138 ( \16930 , \16590 , \16594 );
nand \U$15139 ( \16931 , \16929 , \16930 );
nor \U$15140 ( \16932 , \16609 , \16602 );
not \U$15141 ( \16933 , \16615 );
and \U$15142 ( \16934 , \16932 , \16933 );
or \U$15143 ( \16935 , \16602 , \16622 );
nand \U$15144 ( \16936 , \16935 , \16630 );
nor \U$15145 ( \16937 , \16934 , \16936 );
or \U$15146 ( \16938 , \16931 , \16937 );
or \U$15147 ( \16939 , \16587 , \16637 );
nand \U$15148 ( \16940 , \16939 , \16646 );
and \U$15149 ( \16941 , \16930 , \16940 );
or \U$15150 ( \16942 , \16594 , \16653 );
nand \U$15151 ( \16943 , \16942 , \16661 );
nor \U$15152 ( \16944 , \16941 , \16943 );
nand \U$15153 ( \16945 , \16938 , \16944 );
not \U$15154 ( \16946 , \16945 );
xor \U$15155 ( \16947 , \16928 , \16946 );
buf g4953_GF_PartitionCandidate( \16948_nG4953 , \16947 );
_HMUX g4954_GF_PartitionCandidate ( \16949_nG4954 , \16926_nG490b , \16948_nG4953 , \16488 );
buf \U$15156 ( \16950 , \16949_nG4954 );
not \U$15157 ( \16951 , \11901 );
nand \U$15158 ( \16952 , \12531 , \16951 );
nor \U$15159 ( \16953 , \16687 , \16679 );
nor \U$15160 ( \16954 , \16680 , \16682 );
nand \U$15161 ( \16955 , \16953 , \16954 );
nor \U$15162 ( \16956 , \16689 , \16686 );
and \U$15163 ( \16957 , \16956 , \12459 );
or \U$15164 ( \16958 , \16686 , \16693 );
nand \U$15165 ( \16959 , \16958 , \16697 );
nor \U$15166 ( \16960 , \16957 , \16959 );
or \U$15167 ( \16961 , \16955 , \16960 );
or \U$15168 ( \16962 , \16679 , \16700 );
nand \U$15169 ( \16963 , \16962 , \16705 );
and \U$15170 ( \16964 , \16954 , \16963 );
or \U$15171 ( \16965 , \16682 , \16708 );
nand \U$15172 ( \16966 , \16965 , \16712 );
nor \U$15173 ( \16967 , \16964 , \16966 );
nand \U$15174 ( \16968 , \16961 , \16967 );
not \U$15175 ( \16969 , \16968 );
xor \U$15176 ( \16970 , \16952 , \16969 );
buf g4876_GF_PartitionCandidate( \16971_nG4876 , \16970 );
not \U$15177 ( \16972 , \14747 );
nand \U$15178 ( \16973 , \15377 , \16972 );
nor \U$15179 ( \16974 , \16732 , \16724 );
nor \U$15180 ( \16975 , \16725 , \16727 );
nand \U$15181 ( \16976 , \16974 , \16975 );
nor \U$15182 ( \16977 , \16734 , \16731 );
and \U$15183 ( \16978 , \16977 , \15305 );
or \U$15184 ( \16979 , \16731 , \16738 );
nand \U$15185 ( \16980 , \16979 , \16742 );
nor \U$15186 ( \16981 , \16978 , \16980 );
or \U$15187 ( \16982 , \16976 , \16981 );
or \U$15188 ( \16983 , \16724 , \16745 );
nand \U$15189 ( \16984 , \16983 , \16750 );
and \U$15190 ( \16985 , \16975 , \16984 );
or \U$15191 ( \16986 , \16727 , \16753 );
nand \U$15192 ( \16987 , \16986 , \16757 );
nor \U$15193 ( \16988 , \16985 , \16987 );
nand \U$15194 ( \16989 , \16982 , \16988 );
not \U$15195 ( \16990 , \16989 );
xor \U$15196 ( \16991 , \16973 , \16990 );
buf g48c2_GF_PartitionCandidate( \16992_nG48c2 , \16991 );
_HMUX g48c3_GF_PartitionCandidate ( \16993_nG48c3 , \16971_nG4876 , \16992_nG48c2 , \16488 );
buf \U$15197 ( \16994 , \16993_nG48c3 );
not \U$15198 ( \16995 , \11844 );
nand \U$15199 ( \16996 , \12528 , \16995 );
nor \U$15200 ( \16997 , \16779 , \16771 );
nor \U$15201 ( \16998 , \16772 , \16774 );
nand \U$15202 ( \16999 , \16997 , \16998 );
nor \U$15203 ( \17000 , \16781 , \16778 );
and \U$15204 ( \17001 , \17000 , \16519 );
or \U$15205 ( \17002 , \16778 , \16784 );
nand \U$15206 ( \17003 , \17002 , \16788 );
nor \U$15207 ( \17004 , \17001 , \17003 );
or \U$15208 ( \17005 , \16999 , \17004 );
or \U$15209 ( \17006 , \16771 , \16791 );
nand \U$15210 ( \17007 , \17006 , \16796 );
and \U$15211 ( \17008 , \16998 , \17007 );
or \U$15212 ( \17009 , \16774 , \16799 );
nand \U$15213 ( \17010 , \17009 , \16803 );
nor \U$15214 ( \17011 , \17008 , \17010 );
nand \U$15215 ( \17012 , \17005 , \17011 );
not \U$15216 ( \17013 , \17012 );
xor \U$15217 ( \17014 , \16996 , \17013 );
buf g47d9_GF_PartitionCandidate( \17015_nG47d9 , \17014 );
not \U$15218 ( \17016 , \14690 );
nand \U$15219 ( \17017 , \15374 , \17016 );
nor \U$15220 ( \17018 , \16823 , \16815 );
nor \U$15221 ( \17019 , \16816 , \16818 );
nand \U$15222 ( \17020 , \17018 , \17019 );
nor \U$15223 ( \17021 , \16825 , \16822 );
and \U$15224 ( \17022 , \17021 , \16611 );
or \U$15225 ( \17023 , \16822 , \16828 );
nand \U$15226 ( \17024 , \17023 , \16832 );
nor \U$15227 ( \17025 , \17022 , \17024 );
or \U$15228 ( \17026 , \17020 , \17025 );
or \U$15229 ( \17027 , \16815 , \16835 );
nand \U$15230 ( \17028 , \17027 , \16840 );
and \U$15231 ( \17029 , \17019 , \17028 );
or \U$15232 ( \17030 , \16818 , \16843 );
nand \U$15233 ( \17031 , \17030 , \16847 );
nor \U$15234 ( \17032 , \17029 , \17031 );
nand \U$15235 ( \17033 , \17026 , \17032 );
not \U$15236 ( \17034 , \17033 );
xor \U$15237 ( \17035 , \17017 , \17034 );
buf g4829_GF_PartitionCandidate( \17036_nG4829 , \17035 );
_HMUX g482a_GF_PartitionCandidate ( \17037_nG482a , \17015_nG47d9 , \17036_nG4829 , \16488 );
buf \U$15238 ( \17038 , \17037_nG482a );
not \U$15239 ( \17039 , \11784 );
nand \U$15240 ( \17040 , \12526 , \17039 );
nand \U$15241 ( \17041 , \12365 , \11723 );
not \U$15242 ( \17042 , \12477 );
or \U$15243 ( \17043 , \17041 , \17042 );
and \U$15244 ( \17044 , \11723 , \12500 );
nor \U$15245 ( \17045 , \17044 , \12524 );
nand \U$15246 ( \17046 , \17043 , \17045 );
not \U$15247 ( \17047 , \17046 );
xor \U$15248 ( \17048 , \17040 , \17047 );
buf g4737_GF_PartitionCandidate( \17049_nG4737 , \17048 );
not \U$15249 ( \17050 , \14630 );
nand \U$15250 ( \17051 , \15372 , \17050 );
nand \U$15251 ( \17052 , \15211 , \14569 );
not \U$15252 ( \17053 , \15323 );
or \U$15253 ( \17054 , \17052 , \17053 );
and \U$15254 ( \17055 , \14569 , \15346 );
nor \U$15255 ( \17056 , \17055 , \15370 );
nand \U$15256 ( \17057 , \17054 , \17056 );
not \U$15257 ( \17058 , \17057 );
xor \U$15258 ( \17059 , \17051 , \17058 );
buf g4788_GF_PartitionCandidate( \17060_nG4788 , \17059 );
_HMUX g4789_GF_PartitionCandidate ( \17061_nG4789 , \17049_nG4737 , \17060_nG4788 , \16488 );
buf \U$15259 ( \17062 , \17061_nG4789 );
not \U$15260 ( \17063 , \11720 );
nand \U$15261 ( \17064 , \12521 , \17063 );
nand \U$15262 ( \17065 , \16514 , \16499 );
not \U$15263 ( \17066 , \16531 );
or \U$15264 ( \17067 , \17065 , \17066 );
and \U$15265 ( \17068 , \16499 , \16546 );
nor \U$15266 ( \17069 , \17068 , \16562 );
nand \U$15267 ( \17070 , \17067 , \17069 );
not \U$15268 ( \17071 , \17070 );
xor \U$15269 ( \17072 , \17064 , \17071 );
buf g468c_GF_PartitionCandidate( \17073_nG468c , \17072 );
not \U$15270 ( \17074 , \14566 );
nand \U$15271 ( \17075 , \15367 , \17074 );
nand \U$15272 ( \17076 , \16606 , \16591 );
not \U$15273 ( \17077 , \16623 );
or \U$15274 ( \17078 , \17076 , \17077 );
and \U$15275 ( \17079 , \16591 , \16638 );
nor \U$15276 ( \17080 , \17079 , \16654 );
nand \U$15277 ( \17081 , \17078 , \17080 );
not \U$15278 ( \17082 , \17081 );
xor \U$15279 ( \17083 , \17075 , \17082 );
buf g46e5_GF_PartitionCandidate( \17084_nG46e5 , \17083 );
_HMUX g46e6_GF_PartitionCandidate ( \17085_nG46e6 , \17073_nG468c , \17084_nG46e5 , \16488 );
buf \U$15280 ( \17086 , \17085_nG46e6 );
not \U$15281 ( \17087 , \11651 );
nand \U$15282 ( \17088 , \12519 , \17087 );
nand \U$15283 ( \17089 , \16688 , \16681 );
not \U$15284 ( \17090 , \16694 );
or \U$15285 ( \17091 , \17089 , \17090 );
and \U$15286 ( \17092 , \16681 , \16701 );
nor \U$15287 ( \17093 , \17092 , \16709 );
nand \U$15288 ( \17094 , \17091 , \17093 );
not \U$15289 ( \17095 , \17094 );
xor \U$15290 ( \17096 , \17088 , \17095 );
buf g45d6_GF_PartitionCandidate( \17097_nG45d6 , \17096 );
not \U$15291 ( \17098 , \14497 );
nand \U$15292 ( \17099 , \15365 , \17098 );
nand \U$15293 ( \17100 , \16733 , \16726 );
not \U$15294 ( \17101 , \16739 );
or \U$15295 ( \17102 , \17100 , \17101 );
and \U$15296 ( \17103 , \16726 , \16746 );
nor \U$15297 ( \17104 , \17103 , \16754 );
nand \U$15298 ( \17105 , \17102 , \17104 );
not \U$15299 ( \17106 , \17105 );
xor \U$15300 ( \17107 , \17099 , \17106 );
buf g4632_GF_PartitionCandidate( \17108_nG4632 , \17107 );
_HMUX g4633_GF_PartitionCandidate ( \17109_nG4633 , \17097_nG45d6 , \17108_nG4632 , \16488 );
buf \U$15301 ( \17110 , \17109_nG4633 );
not \U$15302 ( \17111 , \11578 );
nand \U$15303 ( \17112 , \12516 , \17111 );
nand \U$15304 ( \17113 , \16780 , \16773 );
not \U$15305 ( \17114 , \16785 );
or \U$15306 ( \17115 , \17113 , \17114 );
and \U$15307 ( \17116 , \16773 , \16792 );
nor \U$15308 ( \17117 , \17116 , \16800 );
nand \U$15309 ( \17118 , \17115 , \17117 );
not \U$15310 ( \17119 , \17118 );
xor \U$15311 ( \17120 , \17112 , \17119 );
buf g4519_GF_PartitionCandidate( \17121_nG4519 , \17120 );
not \U$15312 ( \17122 , \14424 );
nand \U$15313 ( \17123 , \15362 , \17122 );
nand \U$15314 ( \17124 , \16824 , \16817 );
not \U$15315 ( \17125 , \16829 );
or \U$15316 ( \17126 , \17124 , \17125 );
and \U$15317 ( \17127 , \16817 , \16836 );
nor \U$15318 ( \17128 , \17127 , \16844 );
nand \U$15319 ( \17129 , \17126 , \17128 );
not \U$15320 ( \17130 , \17129 );
xor \U$15321 ( \17131 , \17123 , \17130 );
buf g4579_GF_PartitionCandidate( \17132_nG4579 , \17131 );
_HMUX g457a_GF_PartitionCandidate ( \17133_nG457a , \17121_nG4519 , \17132_nG4579 , \16488 );
buf \U$15322 ( \17134 , \17133_nG457a );
not \U$15323 ( \17135 , \11502 );
nand \U$15324 ( \17136 , \12514 , \17135 );
nand \U$15325 ( \17137 , \16864 , \16861 );
or \U$15326 ( \17138 , \17137 , \12465 );
and \U$15327 ( \17139 , \16861 , \16868 );
nor \U$15328 ( \17140 , \17139 , \16872 );
nand \U$15329 ( \17141 , \17138 , \17140 );
not \U$15330 ( \17142 , \17141 );
xor \U$15331 ( \17143 , \17136 , \17142 );
buf g4459_GF_PartitionCandidate( \17144_nG4459 , \17143 );
not \U$15332 ( \17145 , \14348 );
nand \U$15333 ( \17146 , \15360 , \17145 );
nand \U$15334 ( \17147 , \16886 , \16883 );
or \U$15335 ( \17148 , \17147 , \15311 );
and \U$15336 ( \17149 , \16883 , \16890 );
nor \U$15337 ( \17150 , \17149 , \16894 );
nand \U$15338 ( \17151 , \17148 , \17150 );
not \U$15339 ( \17152 , \17151 );
xor \U$15340 ( \17153 , \17146 , \17152 );
buf g44b8_GF_PartitionCandidate( \17154_nG44b8 , \17153 );
_HMUX g44b9_GF_PartitionCandidate ( \17155_nG44b9 , \17144_nG4459 , \17154_nG44b8 , \16488 );
buf \U$15341 ( \17156 , \17155_nG44b9 );
not \U$15342 ( \17157 , \11425 );
nand \U$15343 ( \17158 , \12510 , \17157 );
nand \U$15344 ( \17159 , \16910 , \16907 );
or \U$15345 ( \17160 , \17159 , \16523 );
and \U$15346 ( \17161 , \16907 , \16914 );
nor \U$15347 ( \17162 , \17161 , \16918 );
nand \U$15348 ( \17163 , \17160 , \17162 );
not \U$15349 ( \17164 , \17163 );
xor \U$15350 ( \17165 , \17158 , \17164 );
buf g439a_GF_PartitionCandidate( \17166_nG439a , \17165 );
not \U$15351 ( \17167 , \14271 );
nand \U$15352 ( \17168 , \15356 , \17167 );
nand \U$15353 ( \17169 , \16932 , \16929 );
or \U$15354 ( \17170 , \17169 , \16615 );
and \U$15355 ( \17171 , \16929 , \16936 );
nor \U$15356 ( \17172 , \17171 , \16940 );
nand \U$15357 ( \17173 , \17170 , \17172 );
not \U$15358 ( \17174 , \17173 );
xor \U$15359 ( \17175 , \17168 , \17174 );
buf g43f9_GF_PartitionCandidate( \17176_nG43f9 , \17175 );
_HMUX g43fa_GF_PartitionCandidate ( \17177_nG43fa , \17166_nG439a , \17176_nG43f9 , \16488 );
buf \U$15360 ( \17178 , \17177_nG43fa );
not \U$15361 ( \17179 , \11350 );
nand \U$15362 ( \17180 , \12508 , \17179 );
nand \U$15363 ( \17181 , \16956 , \16953 );
or \U$15364 ( \17182 , \17181 , \16690 );
and \U$15365 ( \17183 , \16953 , \16959 );
nor \U$15366 ( \17184 , \17183 , \16963 );
nand \U$15367 ( \17185 , \17182 , \17184 );
not \U$15368 ( \17186 , \17185 );
xor \U$15369 ( \17187 , \17180 , \17186 );
buf g42c6_GF_PartitionCandidate( \17188_nG42c6 , \17187 );
not \U$15370 ( \17189 , \14196 );
nand \U$15371 ( \17190 , \15354 , \17189 );
nand \U$15372 ( \17191 , \16977 , \16974 );
or \U$15373 ( \17192 , \17191 , \16735 );
and \U$15374 ( \17193 , \16974 , \16980 );
nor \U$15375 ( \17194 , \17193 , \16984 );
nand \U$15376 ( \17195 , \17192 , \17194 );
not \U$15377 ( \17196 , \17195 );
xor \U$15378 ( \17197 , \17190 , \17196 );
buf g433a_GF_PartitionCandidate( \17198_nG433a , \17197 );
_HMUX g433b_GF_PartitionCandidate ( \17199_nG433b , \17188_nG42c6 , \17198_nG433a , \16488 );
buf \U$15379 ( \17200 , \17199_nG433b );
not \U$15380 ( \17201 , \11273 );
nand \U$15381 ( \17202 , \12505 , \17201 );
nand \U$15382 ( \17203 , \17000 , \16997 );
or \U$15383 ( \17204 , \17203 , \12456 );
and \U$15384 ( \17205 , \16997 , \17003 );
nor \U$15385 ( \17206 , \17205 , \17007 );
nand \U$15386 ( \17207 , \17204 , \17206 );
not \U$15387 ( \17208 , \17207 );
xor \U$15388 ( \17209 , \17202 , \17208 );
buf g41de_GF_PartitionCandidate( \17210_nG41de , \17209 );
not \U$15389 ( \17211 , \14119 );
nand \U$15390 ( \17212 , \15351 , \17211 );
nand \U$15391 ( \17213 , \17021 , \17018 );
or \U$15392 ( \17214 , \17213 , \15302 );
and \U$15393 ( \17215 , \17018 , \17024 );
nor \U$15394 ( \17216 , \17215 , \17028 );
nand \U$15395 ( \17217 , \17214 , \17216 );
not \U$15396 ( \17218 , \17217 );
xor \U$15397 ( \17219 , \17212 , \17218 );
buf g4251_GF_PartitionCandidate( \17220_nG4251 , \17219 );
_HMUX g4252_GF_PartitionCandidate ( \17221_nG4252 , \17210_nG41de , \17220_nG4251 , \16488 );
buf \U$15398 ( \17222 , \17221_nG4252 );
not \U$15399 ( \17223 , \11198 );
nand \U$15400 ( \17224 , \12503 , \17223 );
xor \U$15401 ( \17225 , \17224 , \12501 );
buf g40fe_GF_PartitionCandidate( \17226_nG40fe , \17225 );
not \U$15402 ( \17227 , \14044 );
nand \U$15403 ( \17228 , \15349 , \17227 );
xor \U$15404 ( \17229 , \17228 , \15347 );
buf g416a_GF_PartitionCandidate( \17230_nG416a , \17229 );
_HMUX g416b_GF_PartitionCandidate ( \17231_nG416b , \17226_nG40fe , \17230_nG416a , \16488 );
buf \U$15405 ( \17232 , \17231_nG416b );
not \U$15406 ( \17233 , \12362 );
nand \U$15407 ( \17234 , \12497 , \17233 );
xor \U$15408 ( \17235 , \17234 , \16547 );
buf g4025_GF_PartitionCandidate( \17236_nG4025 , \17235 );
not \U$15409 ( \17237 , \15208 );
nand \U$15410 ( \17238 , \15343 , \17237 );
xor \U$15411 ( \17239 , \17238 , \16639 );
buf g4091_GF_PartitionCandidate( \17240_nG4091 , \17239 );
_HMUX g4092_GF_PartitionCandidate ( \17241_nG4092 , \17236_nG4025 , \17240_nG4091 , \16488 );
buf \U$15412 ( \17242 , \17241_nG4092 );
not \U$15413 ( \17243 , \12355 );
nand \U$15414 ( \17244 , \12495 , \17243 );
xor \U$15415 ( \17245 , \17244 , \16702 );
buf g3f50_GF_PartitionCandidate( \17246_nG3f50 , \17245 );
not \U$15416 ( \17247 , \15201 );
nand \U$15417 ( \17248 , \15341 , \17247 );
xor \U$15418 ( \17249 , \17248 , \16747 );
buf g3fb8_GF_PartitionCandidate( \17250_nG3fb8 , \17249 );
_HMUX g3fb9_GF_PartitionCandidate ( \17251_nG3fb9 , \17246_nG3f50 , \17250_nG3fb8 , \16488 );
buf \U$15419 ( \17252 , \17251_nG3fb9 );
not \U$15420 ( \17253 , \12339 );
nand \U$15421 ( \17254 , \12492 , \17253 );
xor \U$15422 ( \17255 , \17254 , \16793 );
buf g3e7d_GF_PartitionCandidate( \17256_nG3e7d , \17255 );
not \U$15423 ( \17257 , \15185 );
nand \U$15424 ( \17258 , \15338 , \17257 );
xor \U$15425 ( \17259 , \17258 , \16837 );
buf g3ee7_GF_PartitionCandidate( \17260_nG3ee7 , \17259 );
_HMUX g3ee8_GF_PartitionCandidate ( \17261_nG3ee8 , \17256_nG3e7d , \17260_nG3ee7 , \16488 );
buf \U$15426 ( \17262 , \17261_nG3ee8 );
not \U$15427 ( \17263 , \12318 );
nand \U$15428 ( \17264 , \12490 , \17263 );
xor \U$15429 ( \17265 , \17264 , \16869 );
buf g3dad_GF_PartitionCandidate( \17266_nG3dad , \17265 );
not \U$15430 ( \17267 , \15164 );
nand \U$15431 ( \17268 , \15336 , \17267 );
xor \U$15432 ( \17269 , \17268 , \16891 );
buf g3e12_GF_PartitionCandidate( \17270_nG3e12 , \17269 );
_HMUX g3e13_GF_PartitionCandidate ( \17271_nG3e13 , \17266_nG3dad , \17270_nG3e12 , \16488 );
buf \U$15433 ( \17272 , \17271_nG3e13 );
not \U$15434 ( \17273 , \12279 );
nand \U$15435 ( \17274 , \12486 , \17273 );
xor \U$15436 ( \17275 , \17274 , \16915 );
buf g3cbb_GF_PartitionCandidate( \17276_nG3cbb , \17275 );
not \U$15437 ( \17277 , \15125 );
nand \U$15438 ( \17278 , \15332 , \17277 );
xor \U$15439 ( \17279 , \17278 , \16937 );
buf g3d47_GF_PartitionCandidate( \17280_nG3d47 , \17279 );
_HMUX g3d48_GF_PartitionCandidate ( \17281_nG3d48 , \17276_nG3cbb , \17280_nG3d47 , \16488 );
buf \U$15440 ( \17282 , \17281_nG3d48 );
not \U$15441 ( \17283 , \12224 );
nand \U$15442 ( \17284 , \12484 , \17283 );
xor \U$15443 ( \17285 , \17284 , \16960 );
buf g3bd4_GF_PartitionCandidate( \17286_nG3bd4 , \17285 );
not \U$15444 ( \17287 , \15070 );
nand \U$15445 ( \17288 , \15330 , \17287 );
xor \U$15446 ( \17289 , \17288 , \16981 );
buf g3c2e_GF_PartitionCandidate( \17290_nG3c2e , \17289 );
_HMUX g3c2f_GF_PartitionCandidate ( \17291_nG3c2f , \17286_nG3bd4 , \17290_nG3c2e , \16488 );
buf \U$15447 ( \17292 , \17291_nG3c2f );
not \U$15448 ( \17293 , \12172 );
nand \U$15449 ( \17294 , \12481 , \17293 );
xor \U$15450 ( \17295 , \17294 , \17004 );
buf g3ae0_GF_PartitionCandidate( \17296_nG3ae0 , \17295 );
not \U$15451 ( \17297 , \15018 );
nand \U$15452 ( \17298 , \15327 , \17297 );
xor \U$15453 ( \17299 , \17298 , \17025 );
buf g3b79_GF_PartitionCandidate( \17300_nG3b79 , \17299 );
_HMUX g3b7a_GF_PartitionCandidate ( \17301_nG3b7a , \17296_nG3ae0 , \17300_nG3b79 , \16488 );
buf \U$15454 ( \17302 , \17301_nG3b7a );
not \U$15455 ( \17303 , \12127 );
nand \U$15456 ( \17304 , \12479 , \17303 );
xor \U$15457 ( \17305 , \17304 , \17042 );
buf g39f8_GF_PartitionCandidate( \17306_nG39f8 , \17305 );
not \U$15458 ( \17307 , \14973 );
nand \U$15459 ( \17308 , \15325 , \17307 );
xor \U$15460 ( \17309 , \17308 , \17053 );
buf g3a46_GF_PartitionCandidate( \17310_nG3a46 , \17309 );
_HMUX g3a47_GF_PartitionCandidate ( \17311_nG3a47 , \17306_nG39f8 , \17310_nG3a46 , \16488 );
buf \U$15461 ( \17312 , \17311_nG3a47 );
not \U$15462 ( \17313 , \12423 );
nand \U$15463 ( \17314 , \12474 , \17313 );
xor \U$15464 ( \17315 , \17314 , \17066 );
buf g391c_GF_PartitionCandidate( \17316_nG391c , \17315 );
not \U$15465 ( \17317 , \15269 );
nand \U$15466 ( \17318 , \15320 , \17317 );
xor \U$15467 ( \17319 , \17318 , \17077 );
buf g39a9_GF_PartitionCandidate( \17320_nG39a9 , \17319 );
_HMUX g39aa_GF_PartitionCandidate ( \17321_nG39aa , \17316_nG391c , \17320_nG39a9 , \16488 );
buf \U$15468 ( \17322 , \17321_nG39aa );
not \U$15469 ( \17323 , \12420 );
nand \U$15470 ( \17324 , \12472 , \17323 );
xor \U$15471 ( \17325 , \17324 , \17090 );
buf g384a_GF_PartitionCandidate( \17326_nG384a , \17325 );
not \U$15472 ( \17327 , \15266 );
nand \U$15473 ( \17328 , \15318 , \17327 );
xor \U$15474 ( \17329 , \17328 , \17101 );
buf g388e_GF_PartitionCandidate( \17330_nG388e , \17329 );
_HMUX g388f_GF_PartitionCandidate ( \17331_nG388f , \17326_nG384a , \17330_nG388e , \16488 );
buf \U$15475 ( \17332 , \17331_nG388f );
not \U$15476 ( \17333 , \12409 );
nand \U$15477 ( \17334 , \12469 , \17333 );
xor \U$15478 ( \17335 , \17334 , \17114 );
buf g3782_GF_PartitionCandidate( \17336_nG3782 , \17335 );
not \U$15479 ( \17337 , \15255 );
nand \U$15480 ( \17338 , \15315 , \17337 );
xor \U$15481 ( \17339 , \17338 , \17125 );
buf g3805_GF_PartitionCandidate( \17340_nG3805 , \17339 );
_HMUX g3806_GF_PartitionCandidate ( \17341_nG3806 , \17336_nG3782 , \17340_nG3805 , \16488 );
buf \U$15482 ( \17342 , \17341_nG3806 );
not \U$15483 ( \17343 , \12398 );
nand \U$15484 ( \17344 , \12467 , \17343 );
xor \U$15485 ( \17345 , \17344 , \12465 );
buf g36c8_GF_PartitionCandidate( \17346_nG36c8 , \17345 );
not \U$15486 ( \17347 , \15244 );
nand \U$15487 ( \17348 , \15313 , \17347 );
xor \U$15488 ( \17349 , \17348 , \15311 );
buf g36fe_GF_PartitionCandidate( \17350_nG36fe , \17349 );
_HMUX g36ff_GF_PartitionCandidate ( \17351_nG36ff , \17346_nG36c8 , \17350_nG36fe , \16488 );
buf \U$15489 ( \17352 , \17351_nG36ff );
not \U$15490 ( \17353 , \12443 );
nand \U$15491 ( \17354 , \12463 , \17353 );
xor \U$15492 ( \17355 , \17354 , \16523 );
buf g361b_GF_PartitionCandidate( \17356_nG361b , \17355 );
not \U$15493 ( \17357 , \15289 );
nand \U$15494 ( \17358 , \15309 , \17357 );
xor \U$15495 ( \17359 , \17358 , \16615 );
buf g3691_GF_PartitionCandidate( \17360_nG3691 , \17359 );
_HMUX g3692_GF_PartitionCandidate ( \17361_nG3692 , \17356_nG361b , \17360_nG3691 , \16488 );
buf \U$15496 ( \17362 , \17361_nG3692 );
not \U$15497 ( \17363 , \12440 );
nand \U$15498 ( \17364 , \12461 , \17363 );
xor \U$15499 ( \17365 , \17364 , \16690 );
buf g357a_GF_PartitionCandidate( \17366_nG357a , \17365 );
not \U$15500 ( \17367 , \15286 );
nand \U$15501 ( \17368 , \15307 , \17367 );
xor \U$15502 ( \17369 , \17368 , \16735 );
buf g35a4_GF_PartitionCandidate( \17370_nG35a4 , \17369 );
_HMUX g35a5_GF_PartitionCandidate ( \17371_nG35a5 , \17366_nG357a , \17370_nG35a4 , \16488 );
buf \U$15503 ( \17372 , \17371_nG35a5 );
not \U$15504 ( \17373 , \12448 );
nand \U$15505 ( \17374 , \12458 , \17373 );
xor \U$15506 ( \17375 , \17374 , \12456 );
buf g34e7_GF_PartitionCandidate( \17376_nG34e7 , \17375 );
not \U$15507 ( \17377 , \15294 );
nand \U$15508 ( \17378 , \15304 , \17377 );
xor \U$15509 ( \17379 , \17378 , \15302 );
buf g354f_GF_PartitionCandidate( \17380_nG354f , \17379 );
_HMUX g3550_GF_PartitionCandidate ( \17381_nG3550 , \17376_nG34e7 , \17380_nG354f , \16488 );
buf \U$15510 ( \17382 , \17381_nG3550 );
nor \U$15511 ( \17383 , \12452 , \12455 );
not \U$15512 ( \17384 , \17383 );
nand \U$15513 ( \17385 , \12456 , \17384 );
not \U$15514 ( \17386 , \17385 );
buf g345c_GF_PartitionCandidate( \17387_nG345c , \17386 );
nor \U$15515 ( \17388 , \15298 , \15301 );
not \U$15516 ( \17389 , \17388 );
nand \U$15517 ( \17390 , \15302 , \17389 );
not \U$15518 ( \17391 , \17390 );
buf g347e_GF_PartitionCandidate( \17392_nG347e , \17391 );
_HMUX g347f_GF_PartitionCandidate ( \17393_nG347f , \17387_nG345c , \17392_nG347e , \16488 );
buf \U$15519 ( \17394 , \17393_nG347f );
xor \U$15520 ( \17395 , \12454 , \10613 );
buf g339e_GF_PartitionCandidate( \17396_nG339e , \17395 );
xor \U$15521 ( \17397 , \15300 , \13459 );
buf g3439_GF_PartitionCandidate( \17398_nG3439 , \17397 );
_HMUX g343a_GF_PartitionCandidate ( \17399_nG343a , \17396_nG339e , \17398_nG3439 , \16488 );
buf \U$15522 ( \17400 , \17399_nG343a );
endmodule

