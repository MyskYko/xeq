//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RIc2257b0_65,RIc2275b0_1,RIc227538_2,RIc2274c0_3,RIc225738_66,RIc227448_4,RIc2273d0_5,RIc2256c0_67,RIc225648_68,
        RIc227358_6,RIc2272e0_7,RIc2255d0_69,RIc225558_70,RIc227268_8,RIc2271f0_9,RIc2254e0_71,RIc225468_72,RIc227178_10,RIc227100_11,
        RIc2253f0_73,RIc225378_74,RIc227088_12,RIc227010_13,RIc225300_75,RIc225288_76,RIc226f98_14,RIc226f20_15,RIc225210_77,RIc225198_78,
        RIc226ea8_16,RIc226e30_17,RIc225120_79,RIc2250a8_80,RIc226db8_18,RIc226d40_19,RIc225030_81,RIc226cc8_20,RIc226c50_21,RIc224fb8_82,
        RIc224f40_83,RIc224ec8_84,RIc226bd8_22,RIc226b60_23,RIc224e50_85,RIc224dd8_86,RIc226ae8_24,RIc226a70_25,RIc224d60_87,RIc224ce8_88,
        RIc2269f8_26,RIc226980_27,RIc224c70_89,RIc224bf8_90,RIc226908_28,RIc226890_29,RIc224b80_91,RIc224b08_92,RIc226818_30,RIc2267a0_31,
        RIc224a90_93,RIc224a18_94,RIc226728_32,RIc2266b0_33,RIc2249a0_95,RIc224928_96,RIc226638_34,RIc2265c0_35,RIc2248b0_97,RIc224838_98,
        RIc226548_36,RIc2264d0_37,RIc2247c0_99,RIc226458_38,RIc2263e0_39,RIc224748_100,RIc2246d0_101,RIc224658_102,RIc226368_40,RIc2262f0_41,
        RIc2245e0_103,RIc224568_104,RIc226278_42,RIc226200_43,RIc2244f0_105,RIc224478_106,RIc226188_44,RIc226110_45,RIc224400_107,RIc224388_108,
        RIc226098_46,RIc226020_47,RIc224310_109,RIc224298_110,RIc225fa8_48,RIc225f30_49,RIc224220_111,RIc2241a8_112,RIc225eb8_50,RIc225e40_51,
        RIc224130_113,RIc2240b8_114,RIc225dc8_52,RIc225d50_53,RIc224040_115,RIc223fc8_116,RIc225cd8_54,RIc225c60_55,RIc223f50_117,RIc225be8_56,
        RIc225b70_57,RIc223ed8_118,RIc223e60_119,RIc223de8_120,RIc225af8_58,RIc225a80_59,RIc223d70_121,RIc223cf8_122,RIc225a08_60,RIc225990_61,
        RIc223c80_123,RIc223c08_124,RIc225918_62,RIc2258a0_63,RIc223b90_125,RIc223b18_126,RIc2294a0_127,RIc225828_64,RIc229518_128,RIc229590_129,
        RIc229608_130,RIc229680_131,RIc2296f8_132,RIc229770_133,RIc2297e8_134,RIc229860_135,RIc2298d8_136,RIc229950_137,RIc2299c8_138,RIc229a40_139,
        RIc229ab8_140,RIc229b30_141,RIc229ba8_142,RIc229c20_143,RIc229c98_144,RIc229d10_145,RIc229d88_146,RIc229e00_147,RIc229e78_148,RIc229ef0_149,
        RIc229f68_150,RIc229fe0_151,RIc22a058_152,RIc22a0d0_153,RIc22a148_154,RIc22a1c0_155,RIc22a238_156,RIc22a2b0_157,RIc22a328_158,RIc22a3a0_159,
        RIc22a418_160,RIc22a490_161,RIc22a508_162,RIc22a580_163,RIc22a5f8_164,RIc22a670_165,RIc22a6e8_166,RIc22a760_167,RIc22a7d8_168,RIc22a850_169,
        RIc22a8c8_170,RIc22a940_171,RIc22a9b8_172,RIc22aa30_173,RIc22aaa8_174,RIc22ab20_175,RIc22ab98_176,RIc22ac10_177,RIc22ac88_178,RIc22ad00_179,
        RIc22ad78_180,RIc22adf0_181,RIc22ae68_182,RIc22aee0_183,RIc22af58_184,RIc22afd0_185,RIc22b048_186,RIc22b0c0_187,RIc22b138_188,RIc22b1b0_189,
        RIc22b228_190,RIc22b2a0_191,RIc22b318_192,RIc22b390_193,RIc22b408_194,RIc22b480_195,RIc22b4f8_196,RIc22b570_197,RIc22b5e8_198,RIc22b660_199,
        RIc22b6d8_200,RIc22b750_201,RIc22b7c8_202,RIc22b840_203,RIc22b8b8_204,RIc22b930_205,RIc22b9a8_206,RIc22ba20_207,RIc22ba98_208,RIc22bb10_209,
        RIc22bb88_210,RIc22bc00_211,RIc22bc78_212,RIc22bcf0_213,RIc22bd68_214,RIc22bde0_215,RIc22be58_216,RIc22bed0_217,RIc22bf48_218,RIc22bfc0_219,
        RIc22c038_220,RIc22c0b0_221,RIc22c128_222,RIc22c1a0_223,RIc22c218_224,RIc22c290_225,RIc22c308_226,RIc22c380_227,RIc22c3f8_228,RIc22c470_229,
        RIc22c4e8_230,RIc22c560_231,RIc22c5d8_232,RIc22c650_233,RIc22c6c8_234,RIc22c740_235,RIc22c7b8_236,RIc22c830_237,RIc22c8a8_238,RIc22c920_239,
        RIc22c998_240,RIc22ca10_241,RIc22ca88_242,RIc22cb00_243,RIc22cb78_244,RIc22cbf0_245,RIc22cc68_246,RIc22cce0_247,RIc22cd58_248,RIc22cdd0_249,
        RIc22ce48_250,RIc22cec0_251,RIc22cf38_252,RIc22cfb0_253,RIc22d028_254,RIc22d0a0_255,RIc22d118_256,R_101_9cd3d68,R_102_9cd3e10,R_103_9cd3eb8,
        R_104_9cd3f60,R_105_9cd4008,R_106_9cd40b0,R_107_9cd4158,R_108_9cd4200,R_109_9cd42a8,R_10a_9cd4350,R_10b_9cd43f8,R_10c_9cd44a0,R_10d_9cd4548,
        R_10e_9cd45f0,R_10f_9cd4698,R_110_9cd4740,R_111_9cd47e8,R_112_9cd4890,R_113_9cd4938,R_114_9cd49e0,R_115_9cd4a88,R_116_9cd4b30,R_117_9cd4bd8,
        R_118_9cd4c80,R_119_9cd4d28,R_11a_9cd4dd0,R_11b_9cd4e78,R_11c_9cd4f20,R_11d_9cd4fc8,R_11e_9cd5070,R_11f_9cd5118,R_120_9cd51c0,R_121_9cd5268,
        R_122_9cd5310,R_123_9cd53b8,R_124_9cd5460,R_125_9cd5508,R_126_9cd55b0,R_127_9cd5658,R_128_9cd5700,R_129_9cd57a8,R_12a_9cd5850,R_12b_9cd58f8,
        R_12c_9cd59a0,R_12d_9cd5a48,R_12e_9cd5af0,R_12f_9cd5b98,R_130_9cd5c40,R_131_9cd5ce8,R_132_9cd5d90,R_133_9cd5e38,R_134_9cd5ee0,R_135_9cd5f88,
        R_136_9cd6030,R_137_9cd60d8,R_138_9cd6180,R_139_9cd6228,R_13a_9cd62d0,R_13b_9cd6378,R_13c_9cd6420,R_13d_9cd64c8,R_13e_9cd6570,R_13f_9cd6618,
        R_140_9cd66c0,R_141_9cd6768,R_142_9cd6810,R_143_9cd68b8,R_144_9cd6960,R_145_9cd6a08,R_146_9cd6ab0,R_147_9cd6b58,R_148_9cd6c00,R_149_9cd6ca8,
        R_14a_9cd6d50,R_14b_9cd6df8,R_14c_9cd6ea0,R_14d_9cd6f48,R_14e_9cd6ff0,R_14f_9cd7098,R_150_9cd7140,R_151_9cd71e8,R_152_9cd7290,R_153_9cd7338,
        R_154_9cd73e0,R_155_9cd7488,R_156_9cd7530,R_157_9cd75d8,R_158_9cd7680,R_159_9cd7728,R_15a_9cd77d0,R_15b_9cd7878,R_15c_9cd7920,R_15d_9cd79c8,
        R_15e_9cd7a70,R_15f_9cd7b18,R_160_9cd7bc0,R_161_9cd7c68,R_162_9cd7d10,R_163_9cd7db8,R_164_9cd7e60,R_165_9cd7f08,R_166_9cd7fb0,R_167_9cd8058,
        R_168_9cd8100,R_169_9cd81a8,R_16a_9cd8250,R_16b_9cd82f8,R_16c_9cd83a0,R_16d_9cd8448,R_16e_9cd84f0,R_16f_9cd8598,R_170_9cd8640,R_171_9cd86e8,
        R_172_9cd8790,R_173_9cd8838,R_174_9cd88e0,R_175_9cd8988,R_176_9cd8a30,R_177_9cd8ad8);
input RIc2257b0_65,RIc2275b0_1,RIc227538_2,RIc2274c0_3,RIc225738_66,RIc227448_4,RIc2273d0_5,RIc2256c0_67,RIc225648_68,
        RIc227358_6,RIc2272e0_7,RIc2255d0_69,RIc225558_70,RIc227268_8,RIc2271f0_9,RIc2254e0_71,RIc225468_72,RIc227178_10,RIc227100_11,
        RIc2253f0_73,RIc225378_74,RIc227088_12,RIc227010_13,RIc225300_75,RIc225288_76,RIc226f98_14,RIc226f20_15,RIc225210_77,RIc225198_78,
        RIc226ea8_16,RIc226e30_17,RIc225120_79,RIc2250a8_80,RIc226db8_18,RIc226d40_19,RIc225030_81,RIc226cc8_20,RIc226c50_21,RIc224fb8_82,
        RIc224f40_83,RIc224ec8_84,RIc226bd8_22,RIc226b60_23,RIc224e50_85,RIc224dd8_86,RIc226ae8_24,RIc226a70_25,RIc224d60_87,RIc224ce8_88,
        RIc2269f8_26,RIc226980_27,RIc224c70_89,RIc224bf8_90,RIc226908_28,RIc226890_29,RIc224b80_91,RIc224b08_92,RIc226818_30,RIc2267a0_31,
        RIc224a90_93,RIc224a18_94,RIc226728_32,RIc2266b0_33,RIc2249a0_95,RIc224928_96,RIc226638_34,RIc2265c0_35,RIc2248b0_97,RIc224838_98,
        RIc226548_36,RIc2264d0_37,RIc2247c0_99,RIc226458_38,RIc2263e0_39,RIc224748_100,RIc2246d0_101,RIc224658_102,RIc226368_40,RIc2262f0_41,
        RIc2245e0_103,RIc224568_104,RIc226278_42,RIc226200_43,RIc2244f0_105,RIc224478_106,RIc226188_44,RIc226110_45,RIc224400_107,RIc224388_108,
        RIc226098_46,RIc226020_47,RIc224310_109,RIc224298_110,RIc225fa8_48,RIc225f30_49,RIc224220_111,RIc2241a8_112,RIc225eb8_50,RIc225e40_51,
        RIc224130_113,RIc2240b8_114,RIc225dc8_52,RIc225d50_53,RIc224040_115,RIc223fc8_116,RIc225cd8_54,RIc225c60_55,RIc223f50_117,RIc225be8_56,
        RIc225b70_57,RIc223ed8_118,RIc223e60_119,RIc223de8_120,RIc225af8_58,RIc225a80_59,RIc223d70_121,RIc223cf8_122,RIc225a08_60,RIc225990_61,
        RIc223c80_123,RIc223c08_124,RIc225918_62,RIc2258a0_63,RIc223b90_125,RIc223b18_126,RIc2294a0_127,RIc225828_64,RIc229518_128,RIc229590_129,
        RIc229608_130,RIc229680_131,RIc2296f8_132,RIc229770_133,RIc2297e8_134,RIc229860_135,RIc2298d8_136,RIc229950_137,RIc2299c8_138,RIc229a40_139,
        RIc229ab8_140,RIc229b30_141,RIc229ba8_142,RIc229c20_143,RIc229c98_144,RIc229d10_145,RIc229d88_146,RIc229e00_147,RIc229e78_148,RIc229ef0_149,
        RIc229f68_150,RIc229fe0_151,RIc22a058_152,RIc22a0d0_153,RIc22a148_154,RIc22a1c0_155,RIc22a238_156,RIc22a2b0_157,RIc22a328_158,RIc22a3a0_159,
        RIc22a418_160,RIc22a490_161,RIc22a508_162,RIc22a580_163,RIc22a5f8_164,RIc22a670_165,RIc22a6e8_166,RIc22a760_167,RIc22a7d8_168,RIc22a850_169,
        RIc22a8c8_170,RIc22a940_171,RIc22a9b8_172,RIc22aa30_173,RIc22aaa8_174,RIc22ab20_175,RIc22ab98_176,RIc22ac10_177,RIc22ac88_178,RIc22ad00_179,
        RIc22ad78_180,RIc22adf0_181,RIc22ae68_182,RIc22aee0_183,RIc22af58_184,RIc22afd0_185,RIc22b048_186,RIc22b0c0_187,RIc22b138_188,RIc22b1b0_189,
        RIc22b228_190,RIc22b2a0_191,RIc22b318_192,RIc22b390_193,RIc22b408_194,RIc22b480_195,RIc22b4f8_196,RIc22b570_197,RIc22b5e8_198,RIc22b660_199,
        RIc22b6d8_200,RIc22b750_201,RIc22b7c8_202,RIc22b840_203,RIc22b8b8_204,RIc22b930_205,RIc22b9a8_206,RIc22ba20_207,RIc22ba98_208,RIc22bb10_209,
        RIc22bb88_210,RIc22bc00_211,RIc22bc78_212,RIc22bcf0_213,RIc22bd68_214,RIc22bde0_215,RIc22be58_216,RIc22bed0_217,RIc22bf48_218,RIc22bfc0_219,
        RIc22c038_220,RIc22c0b0_221,RIc22c128_222,RIc22c1a0_223,RIc22c218_224,RIc22c290_225,RIc22c308_226,RIc22c380_227,RIc22c3f8_228,RIc22c470_229,
        RIc22c4e8_230,RIc22c560_231,RIc22c5d8_232,RIc22c650_233,RIc22c6c8_234,RIc22c740_235,RIc22c7b8_236,RIc22c830_237,RIc22c8a8_238,RIc22c920_239,
        RIc22c998_240,RIc22ca10_241,RIc22ca88_242,RIc22cb00_243,RIc22cb78_244,RIc22cbf0_245,RIc22cc68_246,RIc22cce0_247,RIc22cd58_248,RIc22cdd0_249,
        RIc22ce48_250,RIc22cec0_251,RIc22cf38_252,RIc22cfb0_253,RIc22d028_254,RIc22d0a0_255,RIc22d118_256;
output R_101_9cd3d68,R_102_9cd3e10,R_103_9cd3eb8,R_104_9cd3f60,R_105_9cd4008,R_106_9cd40b0,R_107_9cd4158,R_108_9cd4200,R_109_9cd42a8,
        R_10a_9cd4350,R_10b_9cd43f8,R_10c_9cd44a0,R_10d_9cd4548,R_10e_9cd45f0,R_10f_9cd4698,R_110_9cd4740,R_111_9cd47e8,R_112_9cd4890,R_113_9cd4938,
        R_114_9cd49e0,R_115_9cd4a88,R_116_9cd4b30,R_117_9cd4bd8,R_118_9cd4c80,R_119_9cd4d28,R_11a_9cd4dd0,R_11b_9cd4e78,R_11c_9cd4f20,R_11d_9cd4fc8,
        R_11e_9cd5070,R_11f_9cd5118,R_120_9cd51c0,R_121_9cd5268,R_122_9cd5310,R_123_9cd53b8,R_124_9cd5460,R_125_9cd5508,R_126_9cd55b0,R_127_9cd5658,
        R_128_9cd5700,R_129_9cd57a8,R_12a_9cd5850,R_12b_9cd58f8,R_12c_9cd59a0,R_12d_9cd5a48,R_12e_9cd5af0,R_12f_9cd5b98,R_130_9cd5c40,R_131_9cd5ce8,
        R_132_9cd5d90,R_133_9cd5e38,R_134_9cd5ee0,R_135_9cd5f88,R_136_9cd6030,R_137_9cd60d8,R_138_9cd6180,R_139_9cd6228,R_13a_9cd62d0,R_13b_9cd6378,
        R_13c_9cd6420,R_13d_9cd64c8,R_13e_9cd6570,R_13f_9cd6618,R_140_9cd66c0,R_141_9cd6768,R_142_9cd6810,R_143_9cd68b8,R_144_9cd6960,R_145_9cd6a08,
        R_146_9cd6ab0,R_147_9cd6b58,R_148_9cd6c00,R_149_9cd6ca8,R_14a_9cd6d50,R_14b_9cd6df8,R_14c_9cd6ea0,R_14d_9cd6f48,R_14e_9cd6ff0,R_14f_9cd7098,
        R_150_9cd7140,R_151_9cd71e8,R_152_9cd7290,R_153_9cd7338,R_154_9cd73e0,R_155_9cd7488,R_156_9cd7530,R_157_9cd75d8,R_158_9cd7680,R_159_9cd7728,
        R_15a_9cd77d0,R_15b_9cd7878,R_15c_9cd7920,R_15d_9cd79c8,R_15e_9cd7a70,R_15f_9cd7b18,R_160_9cd7bc0,R_161_9cd7c68,R_162_9cd7d10,R_163_9cd7db8,
        R_164_9cd7e60,R_165_9cd7f08,R_166_9cd7fb0,R_167_9cd8058,R_168_9cd8100,R_169_9cd81a8,R_16a_9cd8250,R_16b_9cd82f8,R_16c_9cd83a0,R_16d_9cd8448,
        R_16e_9cd84f0,R_16f_9cd8598,R_170_9cd8640,R_171_9cd86e8,R_172_9cd8790,R_173_9cd8838,R_174_9cd88e0,R_175_9cd8988,R_176_9cd8a30,R_177_9cd8ad8;

wire \376_ZERO , \377_ONE , \378 , \379 , \380 , \381 , \382 , \383 , \384 ,
         \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 ,
         \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 ,
         \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 ,
         \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 ,
         \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 ,
         \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 ,
         \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 ,
         \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 ,
         \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 ,
         \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 ,
         \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 ,
         \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 ,
         \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 ,
         \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 ,
         \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 ,
         \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 ,
         \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 ,
         \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 ,
         \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 ,
         \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 ,
         \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 ,
         \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 ,
         \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 ,
         \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 ,
         \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 ,
         \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 ,
         \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 ,
         \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 ,
         \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 ,
         \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 ,
         \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 ,
         \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 ,
         \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 ,
         \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 ,
         \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 ,
         \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 ,
         \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 ,
         \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 ,
         \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 ,
         \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 ,
         \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 ,
         \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 ,
         \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 ,
         \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 ,
         \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 ,
         \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 ,
         \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 ,
         \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 ,
         \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 ,
         \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 ,
         \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 ,
         \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 ,
         \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 ,
         \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 ,
         \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 ,
         \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 ,
         \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 ,
         \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 ,
         \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 ,
         \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 ,
         \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 ,
         \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 ,
         \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 ,
         \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 ,
         \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 ,
         \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 ,
         \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 ,
         \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 ,
         \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 ,
         \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 ,
         \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 ,
         \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 ,
         \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 ,
         \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 ,
         \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 ,
         \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 ,
         \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 ,
         \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 ,
         \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 ,
         \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 ,
         \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 ,
         \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 ,
         \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 ,
         \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 ,
         \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 ,
         \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 ,
         \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 ,
         \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 ,
         \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 ,
         \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 ,
         \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 ,
         \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 ,
         \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 ,
         \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 ,
         \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 ,
         \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 ,
         \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 ,
         \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 ,
         \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 ,
         \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 ,
         \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 ,
         \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 ,
         \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 ,
         \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 ,
         \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 ,
         \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 ,
         \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 ,
         \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 ,
         \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 ,
         \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 ,
         \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 ,
         \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 ,
         \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 ,
         \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 ,
         \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 ,
         \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 ,
         \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 ,
         \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 ,
         \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 ,
         \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 ,
         \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 ,
         \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 ,
         \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 ,
         \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 ,
         \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 ,
         \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 ,
         \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 ,
         \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 ,
         \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 ,
         \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 ,
         \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 ,
         \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 ,
         \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 ,
         \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 ,
         \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 ,
         \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 ,
         \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 ,
         \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 ,
         \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 ,
         \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 ,
         \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 ,
         \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 ,
         \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 ,
         \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 ,
         \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 ,
         \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 ,
         \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 ,
         \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 ,
         \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 ,
         \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 ,
         \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 ,
         \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 ,
         \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 ,
         \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 ,
         \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 ,
         \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 ,
         \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 ,
         \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 ,
         \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 ,
         \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 ,
         \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 ,
         \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 ,
         \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 ,
         \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 ,
         \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 ,
         \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 ,
         \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 ,
         \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 ,
         \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 ,
         \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 ,
         \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 ,
         \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 ,
         \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 ,
         \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 ,
         \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 ,
         \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 ,
         \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 ,
         \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 ,
         \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 ,
         \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 ,
         \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 ,
         \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 ,
         \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 ,
         \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 ,
         \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 ,
         \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 ,
         \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 ,
         \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 ,
         \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 ,
         \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 ,
         \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 ,
         \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 ,
         \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 ,
         \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 ,
         \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 ,
         \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 ,
         \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 ,
         \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 ,
         \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 ,
         \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 ,
         \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 ,
         \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 ,
         \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 ,
         \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 ,
         \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 ,
         \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 ,
         \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 ,
         \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 ,
         \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 ,
         \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 ,
         \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 ,
         \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 ,
         \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 ,
         \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 ,
         \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 ,
         \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 ,
         \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 ,
         \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 ,
         \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 ,
         \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 ,
         \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 ,
         \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 ,
         \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 ,
         \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 ,
         \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 ,
         \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 ,
         \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 ,
         \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 ,
         \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 ,
         \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 ,
         \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 ,
         \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 ,
         \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 ,
         \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 ,
         \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 ,
         \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 ,
         \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 ,
         \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 ,
         \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 ,
         \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 ,
         \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 ,
         \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 ,
         \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 ,
         \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 ,
         \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 ,
         \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 ,
         \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 ,
         \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 ,
         \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 ,
         \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 ,
         \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 ,
         \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 ,
         \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 ,
         \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 ,
         \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 ,
         \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 ,
         \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 ,
         \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 ,
         \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 ,
         \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 ,
         \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 ,
         \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 ,
         \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 ,
         \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 ,
         \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 ,
         \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 ,
         \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 ,
         \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 ,
         \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 ,
         \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 ,
         \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 ,
         \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 ,
         \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 ,
         \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 ,
         \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 ,
         \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 ,
         \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 ,
         \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 ,
         \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 ,
         \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 ,
         \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 ,
         \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 ,
         \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 ,
         \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 ,
         \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 ,
         \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 ,
         \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 ,
         \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 ,
         \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 ,
         \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 ,
         \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 ,
         \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 ,
         \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 ,
         \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 ,
         \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 ,
         \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 ,
         \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 ,
         \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 ,
         \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 ,
         \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 ,
         \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 ,
         \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 ,
         \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 ,
         \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 ,
         \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 ,
         \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 ,
         \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 ,
         \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 ,
         \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 ,
         \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 ,
         \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 ,
         \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 ,
         \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 ,
         \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 ,
         \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 ,
         \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 ,
         \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 ,
         \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 ,
         \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 ,
         \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 ,
         \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 ,
         \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 ,
         \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 ,
         \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 ,
         \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 ,
         \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 ,
         \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 ,
         \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 ,
         \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 ,
         \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 ,
         \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 ,
         \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 ,
         \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 ,
         \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 ,
         \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 ,
         \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 ,
         \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 ,
         \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 ,
         \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 ,
         \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 ,
         \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 ,
         \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 ,
         \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 ,
         \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 ,
         \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 ,
         \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 ,
         \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 ,
         \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 ,
         \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 ,
         \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 ,
         \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 ,
         \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 ,
         \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 ,
         \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 ,
         \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 ,
         \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 ,
         \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 ,
         \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 ,
         \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 ,
         \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 ,
         \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 ,
         \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 ,
         \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 ,
         \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 ,
         \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 ,
         \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 ,
         \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 ,
         \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 ,
         \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 ,
         \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 ,
         \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 ,
         \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 ,
         \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 ,
         \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 ,
         \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 ,
         \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 ,
         \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 ,
         \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 ,
         \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 ,
         \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 ,
         \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 ,
         \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 ,
         \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 ,
         \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 ,
         \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 ,
         \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 ,
         \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 ,
         \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 ,
         \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 ,
         \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 ,
         \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 ,
         \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 ,
         \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 ,
         \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 ,
         \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 ,
         \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 ,
         \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 ,
         \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 ,
         \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 ,
         \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 ,
         \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 ,
         \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 ,
         \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 ,
         \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 ,
         \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 ,
         \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 ,
         \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 ,
         \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 ,
         \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 ,
         \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 ,
         \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 ,
         \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 ,
         \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 ,
         \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 ,
         \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 ,
         \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 ,
         \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 ,
         \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 ,
         \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 ,
         \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 ,
         \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 ,
         \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 ,
         \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 ,
         \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 ,
         \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 ,
         \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 ,
         \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 ,
         \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 ,
         \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 ,
         \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 ,
         \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 ,
         \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 ,
         \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 ,
         \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 ,
         \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 ,
         \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 ,
         \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 ,
         \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 ,
         \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 ,
         \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 ,
         \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 ,
         \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 ,
         \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 ,
         \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 ,
         \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 ,
         \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 ,
         \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 ,
         \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 ,
         \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 ,
         \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 ,
         \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 ,
         \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 ,
         \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 ,
         \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 ,
         \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 ,
         \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 ,
         \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 ,
         \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 ,
         \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 ,
         \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 ,
         \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 ,
         \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 ,
         \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 ,
         \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 ,
         \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 ,
         \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 ,
         \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 ,
         \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 ,
         \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 ,
         \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 ,
         \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 ,
         \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 ,
         \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 ,
         \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 ,
         \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 ,
         \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 ,
         \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 ,
         \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 ,
         \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 ,
         \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 ,
         \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 ,
         \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 ,
         \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 ,
         \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 ,
         \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 ,
         \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 ,
         \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 ,
         \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 ,
         \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 ,
         \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 ,
         \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 ,
         \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 ,
         \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 ,
         \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 ,
         \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 ,
         \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 ,
         \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 ,
         \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 ,
         \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 ,
         \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 ,
         \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 ,
         \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 ,
         \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 ,
         \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 ,
         \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 ,
         \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 ,
         \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 ,
         \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 ,
         \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 ,
         \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 ,
         \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 ,
         \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 ,
         \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 ,
         \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 ,
         \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 ,
         \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 ,
         \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 ,
         \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 ,
         \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 ,
         \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 ,
         \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 ,
         \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 ,
         \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 ,
         \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 ,
         \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 ,
         \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 ,
         \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 ,
         \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 ,
         \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 ,
         \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 ,
         \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 ,
         \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 ,
         \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 ,
         \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 ,
         \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 ,
         \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 ,
         \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 ,
         \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 ,
         \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 ,
         \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 ,
         \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 ,
         \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 ,
         \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 ,
         \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 ,
         \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 ,
         \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 ,
         \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 ,
         \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 ,
         \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 ,
         \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 ,
         \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 ,
         \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 ,
         \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 ,
         \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 ,
         \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 ,
         \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 ,
         \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 ,
         \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 ,
         \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 ,
         \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 ,
         \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 ,
         \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 ,
         \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 ,
         \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 ,
         \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 ,
         \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 ,
         \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 ,
         \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 ,
         \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 ,
         \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 ,
         \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 ,
         \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 ,
         \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 ,
         \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 ,
         \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 ,
         \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 ,
         \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 ,
         \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 ,
         \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 ,
         \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 ,
         \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 ,
         \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 ,
         \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 ,
         \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 ,
         \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 ,
         \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 ,
         \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 ,
         \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 ,
         \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 ,
         \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 ,
         \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 ,
         \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 ,
         \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 ,
         \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 ,
         \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 ,
         \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 ,
         \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 ,
         \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 ,
         \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 ,
         \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 ,
         \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 ,
         \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 ,
         \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 ,
         \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 ,
         \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 ,
         \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 ,
         \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 ,
         \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 ,
         \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 ,
         \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 ,
         \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 ,
         \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 ,
         \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 ,
         \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 ,
         \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 ,
         \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 ,
         \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 ,
         \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 ,
         \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 ,
         \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 ,
         \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 ,
         \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 ,
         \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 ,
         \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 ,
         \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 ,
         \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 ,
         \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 ,
         \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 ,
         \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 ,
         \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 ,
         \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 ,
         \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 ,
         \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 ,
         \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 ,
         \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 ,
         \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 ,
         \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 ,
         \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 ,
         \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 ,
         \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 ,
         \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 ,
         \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 ,
         \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 ,
         \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 ,
         \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 ,
         \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 ,
         \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 ,
         \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 ,
         \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 ,
         \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 ,
         \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 ,
         \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 ,
         \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 ,
         \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 ,
         \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 ,
         \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 ,
         \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 ,
         \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 ,
         \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 ,
         \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 ,
         \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 ,
         \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 ,
         \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 ,
         \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 ,
         \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 ,
         \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 ,
         \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 ,
         \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 ,
         \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 ,
         \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 ,
         \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 ,
         \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 ,
         \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 ,
         \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 ,
         \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 ,
         \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 ,
         \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 ,
         \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 ,
         \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 ,
         \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 ,
         \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 ,
         \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 ,
         \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 ,
         \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 ,
         \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 ,
         \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 ,
         \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 ,
         \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 ,
         \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 ,
         \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 ,
         \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 ,
         \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 ,
         \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 ,
         \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 ,
         \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 ,
         \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 ,
         \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 ,
         \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 ,
         \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 ,
         \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 ,
         \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 ,
         \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 ,
         \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 ,
         \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 ,
         \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 ,
         \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 ,
         \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 ,
         \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 ,
         \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 ,
         \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 ,
         \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 ,
         \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 ,
         \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 ,
         \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 ,
         \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 ,
         \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 ,
         \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 ,
         \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 ,
         \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 ,
         \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 ,
         \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 ,
         \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 ,
         \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 ,
         \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 ,
         \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 ,
         \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 ,
         \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 ,
         \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 ,
         \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 ,
         \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 ,
         \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 ,
         \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 ,
         \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 ,
         \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 ,
         \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 ,
         \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 ,
         \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 ,
         \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 ,
         \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 ,
         \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 ,
         \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 ,
         \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 ,
         \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 ,
         \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 ,
         \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 ,
         \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 ,
         \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 ,
         \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 ,
         \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 ,
         \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 ,
         \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 ,
         \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 ,
         \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 ,
         \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 ,
         \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 ,
         \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 ,
         \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 ,
         \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 ,
         \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 ,
         \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 ,
         \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 ,
         \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 ,
         \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 ,
         \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 ,
         \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 ,
         \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 ,
         \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 ,
         \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 ,
         \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 ,
         \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 ,
         \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 ,
         \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 ,
         \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 ,
         \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 ,
         \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 ,
         \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 ,
         \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 ,
         \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 ,
         \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 ,
         \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 ,
         \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 ,
         \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 ,
         \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 ,
         \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 ,
         \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 ,
         \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 ,
         \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 ,
         \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 ,
         \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 ,
         \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 ,
         \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 ,
         \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 ,
         \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 ,
         \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 ,
         \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 ,
         \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 ,
         \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 ,
         \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 ,
         \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 ,
         \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 ,
         \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 ,
         \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 ,
         \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 ,
         \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 ,
         \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 ,
         \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 ,
         \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 ,
         \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 ,
         \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 ,
         \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 ,
         \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 ,
         \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 ,
         \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 ,
         \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 ,
         \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 ,
         \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 ,
         \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 ,
         \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 ,
         \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 ,
         \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 ,
         \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 ,
         \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 ,
         \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 ,
         \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 ,
         \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 ,
         \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 ,
         \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 ,
         \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 ,
         \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 ,
         \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 ,
         \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 ,
         \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 ,
         \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 ,
         \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 ,
         \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 ,
         \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 ,
         \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 ,
         \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 ,
         \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 ,
         \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 ,
         \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 ,
         \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 ,
         \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 ,
         \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 ,
         \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 ,
         \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 ,
         \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 ,
         \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 ,
         \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 ,
         \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 ,
         \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 ,
         \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 ,
         \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 ,
         \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 ,
         \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 ,
         \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 ,
         \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 ,
         \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 ,
         \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 ,
         \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 ,
         \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 ,
         \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 ,
         \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 ,
         \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 ,
         \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 ,
         \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 ,
         \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 ,
         \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 ,
         \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 ,
         \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 ,
         \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 ,
         \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 ,
         \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 ,
         \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 ,
         \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 ,
         \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 ,
         \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 ,
         \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 ,
         \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 ,
         \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 ,
         \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 ,
         \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 ,
         \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 ,
         \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 ,
         \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 ,
         \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 ,
         \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 ,
         \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 ,
         \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 ,
         \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 ,
         \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 ,
         \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 ,
         \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 ,
         \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 ,
         \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 ,
         \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 ,
         \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 ,
         \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 ,
         \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 ,
         \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 ,
         \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 ,
         \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 ,
         \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 ,
         \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 ,
         \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 ,
         \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 ,
         \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 ,
         \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 ,
         \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 ,
         \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 ,
         \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 ,
         \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 ,
         \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 ,
         \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 ,
         \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 ,
         \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 ,
         \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 ,
         \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 ,
         \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 ,
         \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 ,
         \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 ,
         \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 ,
         \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 ,
         \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 ,
         \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 ,
         \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 ,
         \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 ,
         \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 ,
         \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 ,
         \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 ,
         \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 ,
         \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 ,
         \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 ,
         \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 ,
         \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 ,
         \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 ,
         \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 ,
         \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 ,
         \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 ,
         \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 ,
         \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 ,
         \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 ,
         \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 ,
         \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 ,
         \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 ,
         \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 ,
         \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 ,
         \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 ,
         \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 ,
         \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 ,
         \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 ,
         \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 ,
         \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 ,
         \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 ,
         \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 ,
         \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 ,
         \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 ,
         \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 ,
         \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 ,
         \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 ,
         \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 ,
         \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 ,
         \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 ,
         \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 ,
         \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 ,
         \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 ,
         \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 ,
         \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 ,
         \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 ,
         \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 ,
         \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 ,
         \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 ,
         \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 ,
         \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 ,
         \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 ,
         \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 ,
         \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 ,
         \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 ,
         \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 ,
         \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 ,
         \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 ,
         \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 ,
         \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 ,
         \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 ,
         \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 ,
         \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 ,
         \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 ,
         \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 ,
         \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 ,
         \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 ,
         \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 ,
         \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 ,
         \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 ,
         \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 ,
         \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 ,
         \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 ,
         \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 ,
         \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 ,
         \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 ,
         \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 ,
         \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 ,
         \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 ,
         \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 ,
         \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 ,
         \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 ,
         \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 ,
         \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 ,
         \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 ,
         \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 ,
         \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 ,
         \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 ,
         \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 ,
         \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 ,
         \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 ,
         \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 ,
         \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 ,
         \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 ,
         \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 ,
         \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 ,
         \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 ,
         \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 ,
         \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 ,
         \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 ,
         \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 ,
         \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 ,
         \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 ,
         \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 ,
         \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 ,
         \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 ,
         \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 ,
         \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 ,
         \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 ,
         \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 ,
         \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 ,
         \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 ,
         \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 ,
         \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 ,
         \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 ,
         \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 ,
         \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 ,
         \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 ,
         \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 ,
         \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 ,
         \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 ,
         \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 ,
         \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 ,
         \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 ,
         \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 ,
         \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 ,
         \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 ,
         \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 ,
         \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 ,
         \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 ,
         \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 ,
         \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 ,
         \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 ,
         \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 ,
         \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 ,
         \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 ,
         \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 ,
         \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 ,
         \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 ,
         \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 ,
         \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 ,
         \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 ,
         \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 ,
         \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 ,
         \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 ,
         \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 ,
         \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 ,
         \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 ,
         \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 ,
         \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 ,
         \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 ,
         \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 ,
         \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 ,
         \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 ,
         \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 ,
         \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 ,
         \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 ,
         \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 ,
         \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 ,
         \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 ,
         \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 ,
         \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 ,
         \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 ,
         \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 ,
         \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 ,
         \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 ,
         \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 ,
         \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 ,
         \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 ,
         \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 ,
         \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 ,
         \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 ,
         \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 ,
         \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 ,
         \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 ,
         \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 ,
         \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 ,
         \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 ,
         \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 ,
         \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 ,
         \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 ,
         \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 ,
         \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 ,
         \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 ,
         \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 ,
         \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 ,
         \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 ,
         \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 ,
         \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 ,
         \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 ,
         \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 ,
         \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 ,
         \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 ,
         \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 ,
         \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 ,
         \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 ,
         \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 ,
         \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 ,
         \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 ,
         \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 ,
         \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 ,
         \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 ,
         \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 ,
         \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 ,
         \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 ,
         \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 ,
         \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 ,
         \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 ,
         \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 ,
         \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 ,
         \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 ,
         \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 ,
         \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 ,
         \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 ,
         \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 ,
         \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 ,
         \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 ,
         \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 ,
         \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 ,
         \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 ,
         \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 ,
         \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 ,
         \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 ,
         \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 ,
         \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 ,
         \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 ,
         \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 ,
         \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 ,
         \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 ,
         \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 ,
         \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 ,
         \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 ,
         \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 ,
         \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 ,
         \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 ,
         \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 ,
         \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 ,
         \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 ,
         \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 ,
         \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 ,
         \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 ,
         \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 ,
         \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 ,
         \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 ,
         \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 ,
         \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 ,
         \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 ,
         \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 ,
         \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 ,
         \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 ,
         \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 ,
         \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 ,
         \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 ,
         \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 ,
         \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 ,
         \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 ,
         \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 ,
         \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 ,
         \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 ,
         \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 ,
         \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 ,
         \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 ,
         \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 ,
         \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 ,
         \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 ,
         \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 ,
         \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 ,
         \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 ,
         \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 ,
         \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 ,
         \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 ,
         \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 ,
         \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 ,
         \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 ,
         \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 ,
         \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 ,
         \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 ,
         \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 ,
         \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 ,
         \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 ,
         \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 ,
         \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 ,
         \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 ,
         \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 ,
         \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 ,
         \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 ,
         \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 ,
         \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 ,
         \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 ,
         \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 ,
         \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 ,
         \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 ,
         \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 ,
         \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 ,
         \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 ,
         \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 ,
         \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 ,
         \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 ,
         \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 ,
         \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 ,
         \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 ,
         \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 ,
         \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 ,
         \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 ,
         \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 ,
         \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 ,
         \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 ,
         \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 ,
         \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 ,
         \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 ,
         \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 ,
         \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 ,
         \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 ,
         \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 ,
         \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 ,
         \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 ,
         \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 ,
         \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 ,
         \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 ,
         \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 ,
         \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 ,
         \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 ,
         \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 ,
         \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 ,
         \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 ,
         \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 ,
         \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 ,
         \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 ,
         \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 ,
         \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 ,
         \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 ,
         \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 ,
         \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 ,
         \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 ,
         \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 ,
         \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 ,
         \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 ,
         \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 ,
         \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 ,
         \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 ,
         \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 ,
         \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 ,
         \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 ,
         \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 ,
         \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 ,
         \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 ,
         \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 ,
         \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 ,
         \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 ,
         \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 ,
         \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 ,
         \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 ,
         \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 ,
         \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 ,
         \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 ,
         \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 ,
         \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 ,
         \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 ,
         \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 ,
         \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 ,
         \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 ,
         \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 ,
         \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 ,
         \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 ,
         \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 ,
         \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 ,
         \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 ,
         \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 ,
         \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 ,
         \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 ,
         \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 ,
         \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 ,
         \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 ,
         \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 ,
         \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 ,
         \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 ,
         \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 ,
         \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 ,
         \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 ,
         \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 ,
         \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 ,
         \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 ,
         \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 ,
         \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 ,
         \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 ,
         \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 ,
         \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 ,
         \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 ,
         \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 ,
         \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 ,
         \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 ,
         \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 ,
         \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 ,
         \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 ,
         \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 ,
         \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 ,
         \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 ,
         \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 ,
         \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 ,
         \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 ,
         \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 ,
         \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 ,
         \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 ,
         \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 ,
         \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 ,
         \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 ,
         \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 ,
         \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 ,
         \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 ,
         \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 ,
         \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 ,
         \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 ,
         \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 ,
         \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 ,
         \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 ,
         \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 ,
         \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 ,
         \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 ,
         \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 ,
         \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 ,
         \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 ,
         \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 ,
         \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 ,
         \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 ,
         \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 ,
         \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 ,
         \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 ,
         \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 ,
         \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 ,
         \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 ,
         \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 ,
         \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 ,
         \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 ,
         \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 ,
         \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 ,
         \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 ,
         \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 ,
         \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 ,
         \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 ,
         \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 ,
         \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 ,
         \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 ,
         \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 ,
         \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 ,
         \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 ,
         \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 ,
         \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 ,
         \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 ,
         \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 ,
         \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 ,
         \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 ,
         \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 ,
         \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 ,
         \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 ,
         \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 ,
         \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 ,
         \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 ,
         \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 ,
         \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 ,
         \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 ,
         \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 ,
         \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 ,
         \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 ,
         \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 ,
         \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 ,
         \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 ,
         \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 ,
         \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 ,
         \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 ,
         \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 ,
         \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 ,
         \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 ,
         \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 ,
         \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 ,
         \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 ,
         \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 ,
         \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 ,
         \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 ,
         \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 ,
         \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 ,
         \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 ,
         \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 ,
         \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 ,
         \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 ,
         \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 ,
         \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 ,
         \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 ,
         \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 ,
         \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 ,
         \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 ,
         \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 ,
         \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 ,
         \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 ,
         \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 ,
         \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 ,
         \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 ,
         \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 ,
         \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 ,
         \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 ,
         \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 ,
         \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 ,
         \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 ,
         \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 ,
         \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 ,
         \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 ,
         \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 ,
         \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 ,
         \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 ,
         \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 ,
         \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 ,
         \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 ,
         \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 ,
         \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 ,
         \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 ,
         \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 ,
         \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 ,
         \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 ,
         \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 ,
         \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 ,
         \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 ,
         \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 ,
         \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 ,
         \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 ,
         \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 ,
         \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 ,
         \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 ,
         \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 ,
         \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 ,
         \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 ,
         \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 ,
         \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 ,
         \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 ,
         \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 ,
         \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 ,
         \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 ,
         \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 ,
         \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 ,
         \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 ,
         \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 ,
         \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 ,
         \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 ,
         \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 ,
         \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 ,
         \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 ,
         \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 ,
         \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 ,
         \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 ,
         \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 ,
         \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 ,
         \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 ,
         \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 ,
         \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 ,
         \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 ,
         \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 ,
         \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 ,
         \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 ,
         \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 ,
         \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 ,
         \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 ,
         \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 ,
         \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 ,
         \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 ,
         \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 ,
         \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 ,
         \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 ,
         \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 ,
         \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 ,
         \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 ,
         \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 ,
         \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 ,
         \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 ,
         \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 ,
         \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 ,
         \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 ,
         \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 ,
         \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 ,
         \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 ,
         \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 ,
         \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 ,
         \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 ,
         \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 ,
         \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 ,
         \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 ,
         \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 ,
         \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 ,
         \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 ,
         \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 ,
         \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 ,
         \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 ,
         \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 ,
         \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 ,
         \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 ,
         \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 ,
         \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 ,
         \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 ,
         \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 ,
         \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 ,
         \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 ,
         \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 ,
         \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 ,
         \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 ,
         \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 ,
         \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 ,
         \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 ,
         \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 ,
         \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 ,
         \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 ,
         \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 ,
         \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 ,
         \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 ,
         \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 ,
         \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 ,
         \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 ,
         \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 ,
         \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 ,
         \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 ,
         \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 ,
         \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 ,
         \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 ,
         \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 ,
         \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 ,
         \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 ,
         \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 ,
         \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 ,
         \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 ,
         \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 ,
         \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 ,
         \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 ,
         \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 ,
         \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 ,
         \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 ,
         \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 ,
         \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 ,
         \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 ,
         \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 ,
         \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 ,
         \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 ,
         \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 ,
         \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 ,
         \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 ,
         \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 ,
         \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 ,
         \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 ,
         \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 ,
         \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 ,
         \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 ,
         \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 ,
         \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 ,
         \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 ,
         \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 ,
         \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 ,
         \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 ,
         \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 ,
         \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 ,
         \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 ,
         \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 ,
         \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 ,
         \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 ,
         \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 ,
         \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 ,
         \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 ,
         \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 ,
         \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 ,
         \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 ,
         \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 ,
         \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 ,
         \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 ,
         \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 ,
         \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 ,
         \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 ,
         \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 ,
         \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 ,
         \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 ,
         \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 ,
         \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 ,
         \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 ,
         \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 ,
         \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 ,
         \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 ,
         \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 ,
         \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 ,
         \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 ,
         \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 ,
         \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 ,
         \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 ,
         \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 ,
         \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 ,
         \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 ,
         \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 ,
         \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 ,
         \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 ,
         \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 ,
         \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 ,
         \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 ,
         \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 ,
         \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 ,
         \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 ,
         \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 ,
         \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 ,
         \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 ,
         \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 ,
         \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 ,
         \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 ,
         \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 ,
         \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 ,
         \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 ,
         \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 ,
         \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 ,
         \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 ,
         \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 ,
         \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 ,
         \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 ,
         \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 ,
         \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 ,
         \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 ,
         \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 ,
         \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 ,
         \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 ,
         \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 ,
         \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 ,
         \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 ,
         \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 ,
         \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 ,
         \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 ,
         \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 ,
         \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 ,
         \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 ,
         \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 ,
         \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 ,
         \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 ,
         \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 ,
         \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 ,
         \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 ,
         \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 ,
         \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 ,
         \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 ,
         \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 ,
         \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 ,
         \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 ,
         \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 ,
         \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 ,
         \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 ,
         \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 ,
         \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 ,
         \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 ,
         \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 ,
         \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 ,
         \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 ,
         \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 ,
         \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 ,
         \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 ,
         \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 ,
         \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 ,
         \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 ,
         \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 ,
         \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 ,
         \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 ,
         \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 ,
         \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 ,
         \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 ,
         \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 ,
         \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 ,
         \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 ,
         \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 ,
         \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 ,
         \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 ,
         \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 ,
         \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 ,
         \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 ,
         \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 ,
         \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 ,
         \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 ,
         \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 ,
         \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 ,
         \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 ,
         \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 ,
         \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 ,
         \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 ,
         \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 ,
         \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 ,
         \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 ,
         \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 ,
         \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 ,
         \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 ,
         \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 ,
         \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 ,
         \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 ,
         \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 ,
         \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 ,
         \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 ,
         \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 ,
         \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 ,
         \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 ,
         \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 ,
         \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 ,
         \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 ,
         \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 ,
         \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 ,
         \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 ,
         \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 ,
         \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 ,
         \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 ,
         \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 ,
         \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 ,
         \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 ,
         \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 ,
         \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 ,
         \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 ,
         \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 ,
         \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 ,
         \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 ,
         \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 ,
         \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 ,
         \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 ,
         \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 ,
         \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 ,
         \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 ,
         \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 ,
         \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 ,
         \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 ,
         \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 ,
         \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 ,
         \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 ,
         \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 ,
         \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 ,
         \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 ,
         \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 ,
         \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 ,
         \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 ,
         \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 ,
         \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 ,
         \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 ,
         \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 ,
         \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 ,
         \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 ,
         \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 ,
         \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 ,
         \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 ,
         \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 ,
         \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 ,
         \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 ,
         \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 ,
         \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 ,
         \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 ,
         \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 ,
         \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 ,
         \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 ,
         \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 ,
         \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 ,
         \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 ,
         \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 ,
         \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 ,
         \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 ,
         \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 ,
         \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 ,
         \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 ,
         \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 ,
         \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 ,
         \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 ,
         \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 ,
         \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 ,
         \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 ,
         \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 ,
         \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 ,
         \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 ,
         \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 ,
         \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 ,
         \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 ,
         \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 ,
         \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 ,
         \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 ,
         \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 ,
         \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 ,
         \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 ,
         \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 ,
         \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 ,
         \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 ,
         \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 ,
         \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 ,
         \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 ,
         \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 ,
         \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 ,
         \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 ,
         \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 ,
         \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 ,
         \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 ,
         \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 ,
         \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 ,
         \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 ,
         \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 ,
         \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651_nGaed4 , \21652 , \21653 , \21654 ,
         \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 ,
         \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 ,
         \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 ,
         \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 ,
         \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 ,
         \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 ,
         \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 ,
         \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 ,
         \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 ,
         \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 ,
         \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 ,
         \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 ,
         \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 ,
         \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 ,
         \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 ,
         \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 ,
         \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 ,
         \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 ,
         \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 ,
         \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 ,
         \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 ,
         \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 ,
         \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 ,
         \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 ,
         \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 ,
         \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 ,
         \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 ,
         \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 ,
         \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 ,
         \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 ,
         \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 ,
         \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 ,
         \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 ,
         \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 ,
         \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 ,
         \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 ,
         \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 ,
         \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 ,
         \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 ,
         \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 ,
         \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 ,
         \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 ,
         \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 ,
         \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 , \22093 , \22094 ,
         \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 , \22103 , \22104 ,
         \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 ,
         \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 ,
         \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 , \22133 , \22134 ,
         \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 ,
         \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 ,
         \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 ,
         \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 ,
         \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 ,
         \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194 ,
         \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 ,
         \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 ,
         \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 ,
         \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 ,
         \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 ,
         \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 ,
         \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 ,
         \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 ,
         \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 ,
         \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 ,
         \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 ,
         \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 ,
         \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 ,
         \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 ,
         \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 ,
         \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 ,
         \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 ,
         \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 ,
         \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 ,
         \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 ,
         \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 ,
         \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 ,
         \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 ,
         \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 ,
         \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 ,
         \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 ,
         \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 ,
         \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 ,
         \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 ,
         \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 ,
         \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 ,
         \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 ,
         \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 ,
         \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 ,
         \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 ,
         \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553 , \22554 ,
         \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 ,
         \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 ,
         \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 ,
         \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 ,
         \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 ,
         \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 ,
         \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 ,
         \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 , \22633 , \22634 ,
         \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 ,
         \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 ,
         \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 ,
         \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 ,
         \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 ,
         \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 ,
         \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 ,
         \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 ,
         \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 ,
         \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 ,
         \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 ,
         \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 ,
         \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 ,
         \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 ,
         \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 , \22783 , \22784 ,
         \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 ,
         \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 ,
         \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 ,
         \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 ,
         \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 ,
         \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 ,
         \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 ,
         \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 ,
         \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 ,
         \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 ,
         \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 ,
         \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 ,
         \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914 ,
         \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 ,
         \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 ,
         \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 ,
         \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 ,
         \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 ,
         \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 ,
         \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 ,
         \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 ,
         \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 ,
         \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 ,
         \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 ,
         \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 ,
         \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 ,
         \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 ,
         \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 ,
         \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 ,
         \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 ,
         \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 ,
         \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 ,
         \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 ,
         \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 ,
         \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 ,
         \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 ,
         \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 ,
         \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 ,
         \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 ,
         \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 , \23183 , \23184 ,
         \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 , \23193 , \23194 ,
         \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 ,
         \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 ,
         \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 ,
         \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 ,
         \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 ,
         \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 ,
         \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 ,
         \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 ,
         \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 ,
         \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 ,
         \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 ,
         \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 ,
         \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 ,
         \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 ,
         \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 ,
         \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 ,
         \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 ,
         \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 ,
         \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 ,
         \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 ,
         \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 ,
         \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 ,
         \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 ,
         \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 ,
         \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 ,
         \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 ,
         \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 ,
         \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 ,
         \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483 , \23484 ,
         \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 ,
         \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 ,
         \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 ,
         \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 ,
         \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 ,
         \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 ,
         \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 ,
         \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 ,
         \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 ,
         \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 ,
         \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 ,
         \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 ,
         \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 ,
         \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 ,
         \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 ,
         \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 ,
         \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 ,
         \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 ,
         \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 ,
         \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 ,
         \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 ,
         \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 ,
         \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 ,
         \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 ,
         \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 ,
         \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 ,
         \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 ,
         \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 ,
         \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 ,
         \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 ,
         \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 ,
         \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 ,
         \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 ,
         \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 ,
         \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 ,
         \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 ,
         \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 ,
         \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 ,
         \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 ,
         \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 ,
         \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 ,
         \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 ,
         \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 ,
         \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 ,
         \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 ,
         \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 ,
         \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 ,
         \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 ,
         \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 ,
         \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 ,
         \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 ,
         \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 , \24003 , \24004 ,
         \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 ,
         \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 ,
         \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 ,
         \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 ,
         \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 ,
         \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 ,
         \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 ,
         \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 ,
         \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 ,
         \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 ,
         \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 ,
         \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 ,
         \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133 , \24134 ,
         \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 ,
         \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 ,
         \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 ,
         \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 ,
         \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 ,
         \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 ,
         \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 ,
         \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 ,
         \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 ,
         \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 ,
         \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 ,
         \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 ,
         \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 ,
         \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 ,
         \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 ,
         \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 ,
         \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 ,
         \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 ,
         \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 ,
         \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 ,
         \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 ,
         \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 ,
         \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 ,
         \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 , \24373 , \24374 ,
         \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 ,
         \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 ,
         \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 ,
         \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 ,
         \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 ,
         \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 ,
         \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 ,
         \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 ,
         \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 ,
         \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 ,
         \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 ,
         \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 ,
         \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 ,
         \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 ,
         \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 ,
         \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 ,
         \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 ,
         \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 ,
         \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 ,
         \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 ,
         \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 ,
         \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 ,
         \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 ,
         \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 ,
         \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 ,
         \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 ,
         \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 , \24643 , \24644 ,
         \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 ,
         \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 ,
         \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 ,
         \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 ,
         \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 ,
         \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 ,
         \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 ,
         \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 ,
         \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 ,
         \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 ,
         \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 ,
         \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 ,
         \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 , \24773 , \24774 ,
         \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783 , \24784 ,
         \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 ,
         \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 ,
         \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 ,
         \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 ,
         \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 ,
         \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 ,
         \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 ,
         \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 ,
         \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 ,
         \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 ,
         \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 ,
         \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 ,
         \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 ,
         \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 ,
         \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 ,
         \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 ,
         \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 ,
         \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 ,
         \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 ,
         \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 ,
         \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 ,
         \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 ,
         \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 ,
         \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 ,
         \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 ,
         \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 ,
         \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 ,
         \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 ,
         \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 ,
         \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 ,
         \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 ,
         \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 ,
         \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 ,
         \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 ,
         \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 , \25133 , \25134 ,
         \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 ,
         \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 ,
         \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 ,
         \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 ,
         \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 ,
         \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 ,
         \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 ,
         \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 ,
         \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 ,
         \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 ,
         \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 ,
         \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 ,
         \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 , \25263 , \25264 ,
         \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 , \25273 , \25274 ,
         \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 ,
         \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 ,
         \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 ,
         \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 ,
         \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 ,
         \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 ,
         \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 ,
         \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 ,
         \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 ,
         \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 ,
         \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 ,
         \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 ,
         \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 ,
         \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 ,
         \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 ,
         \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 ,
         \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 ,
         \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 ,
         \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 ,
         \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 ,
         \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 ,
         \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 ,
         \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 ,
         \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 ,
         \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 ,
         \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 ,
         \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 ,
         \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 ,
         \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 ,
         \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 ,
         \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 ,
         \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 ,
         \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 ,
         \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 ,
         \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 ,
         \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 ,
         \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 ,
         \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 ,
         \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 ,
         \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 ,
         \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 ,
         \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 ,
         \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 ,
         \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 ,
         \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 ,
         \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 ,
         \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 ,
         \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 ,
         \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 ,
         \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 , \25773 , \25774 ,
         \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 ,
         \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 ,
         \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 ,
         \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 , \25813 , \25814 ,
         \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 ,
         \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 ,
         \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 ,
         \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 ,
         \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 , \25863 , \25864 ,
         \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 ,
         \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 ,
         \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 ,
         \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 ,
         \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 ,
         \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 ,
         \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 ,
         \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 ,
         \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 ,
         \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 ,
         \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 ,
         \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 ,
         \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 ,
         \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 ,
         \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 , \26013 , \26014 ,
         \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 ,
         \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 ,
         \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 ,
         \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 ,
         \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 ,
         \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 ,
         \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 ,
         \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 ,
         \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 ,
         \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 ,
         \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 ,
         \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 ,
         \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144 ,
         \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 ,
         \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 ,
         \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 ,
         \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 ,
         \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 ,
         \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 ,
         \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 ,
         \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 ,
         \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 ,
         \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 ,
         \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 ,
         \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 ,
         \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 ,
         \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 ,
         \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 ,
         \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 ,
         \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 ,
         \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 ,
         \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 ,
         \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 ,
         \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 ,
         \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 ,
         \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 ,
         \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 ,
         \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 ,
         \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 ,
         \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 , \26413 , \26414 ,
         \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 , \26423 , \26424 ,
         \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434 ,
         \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 ,
         \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 ,
         \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 ,
         \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 ,
         \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 ,
         \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 ,
         \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504 ,
         \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 ,
         \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 ,
         \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533 , \26534 ,
         \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 ,
         \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 ,
         \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 ,
         \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 ,
         \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 ,
         \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 ,
         \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 ,
         \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 ,
         \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 ,
         \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 ,
         \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 ,
         \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 ,
         \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 ,
         \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 , \26673 , \26674 ,
         \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 ,
         \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 ,
         \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 ,
         \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 ,
         \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 ,
         \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 ,
         \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 ,
         \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 ,
         \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 ,
         \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 ,
         \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 ,
         \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 ,
         \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804 ,
         \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 ,
         \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 ,
         \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 ,
         \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 ,
         \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 ,
         \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 ,
         \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 ,
         \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 ,
         \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 ,
         \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 ,
         \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 ,
         \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 ,
         \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 ,
         \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 ,
         \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 ,
         \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 ,
         \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 ,
         \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 ,
         \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 ,
         \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 ,
         \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 ,
         \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 ,
         \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 ,
         \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 ,
         \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 ,
         \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 ,
         \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 ,
         \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 ,
         \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 ,
         \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 ,
         \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 ,
         \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 ,
         \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 ,
         \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 ,
         \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 ,
         \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 ,
         \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 ,
         \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 ,
         \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 ,
         \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 ,
         \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 ,
         \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 ,
         \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 ,
         \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 ,
         \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 ,
         \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 ,
         \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 ,
         \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 ,
         \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 , \27293 , \27294 ,
         \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 ,
         \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 , \27313 , \27314 ,
         \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 ,
         \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 ,
         \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 ,
         \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 ,
         \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 ,
         \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 ,
         \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 ,
         \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 ,
         \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 ,
         \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 ,
         \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 ,
         \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 ,
         \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 ,
         \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 ,
         \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 ,
         \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 ,
         \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 ,
         \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 ,
         \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 ,
         \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 ,
         \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 ,
         \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 ,
         \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 ,
         \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 ,
         \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 ,
         \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 ,
         \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 ,
         \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 ,
         \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 ,
         \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 ,
         \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 ,
         \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 ,
         \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 ,
         \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 ,
         \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 ,
         \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 ,
         \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 ,
         \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 ,
         \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 ,
         \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 ,
         \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 ,
         \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 ,
         \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 ,
         \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 ,
         \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 ,
         \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 ,
         \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 ,
         \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 ,
         \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 ,
         \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 ,
         \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 ,
         \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 , \27833 , \27834 ,
         \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 ,
         \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 ,
         \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 ,
         \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 ,
         \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 ,
         \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 ,
         \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 ,
         \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 ,
         \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 ,
         \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 ,
         \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 ,
         \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 ,
         \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 ,
         \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 ,
         \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 ,
         \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 ,
         \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 ,
         \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 ,
         \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 ,
         \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 ,
         \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 ,
         \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 ,
         \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 ,
         \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 ,
         \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 ,
         \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 ,
         \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 ,
         \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 , \28113 , \28114 ,
         \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 ,
         \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 ,
         \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 ,
         \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 ,
         \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 ,
         \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 ,
         \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 ,
         \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 ,
         \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 ,
         \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 ,
         \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 ,
         \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 ,
         \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 ,
         \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 ,
         \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 ,
         \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 ,
         \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 ,
         \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 ,
         \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 ,
         \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 ,
         \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 ,
         \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 ,
         \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 ,
         \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 ,
         \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 ,
         \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 ,
         \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 ,
         \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 , \28393 , \28394 ,
         \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 ,
         \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 ,
         \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 ,
         \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 ,
         \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 ,
         \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 ,
         \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 ,
         \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 ,
         \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 ,
         \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 ,
         \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 ,
         \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 ,
         \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523 , \28524 ,
         \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 , \28533 , \28534 ,
         \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 ,
         \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 ,
         \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 ,
         \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 ,
         \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 ,
         \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 ,
         \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 , \28603 , \28604 ,
         \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 ,
         \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 ,
         \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 ,
         \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 ,
         \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 ,
         \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 ,
         \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 ,
         \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 ,
         \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 ,
         \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 ,
         \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 ,
         \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 ,
         \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 ,
         \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 ,
         \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 ,
         \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 ,
         \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 ,
         \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 ,
         \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 ,
         \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 ,
         \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 ,
         \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 ,
         \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 ,
         \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 ,
         \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 ,
         \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 ,
         \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 ,
         \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 ,
         \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 ,
         \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 ,
         \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 ,
         \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 ,
         \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933 , \28934 ,
         \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 ,
         \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 ,
         \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 ,
         \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 ,
         \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 ,
         \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 ,
         \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 ,
         \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 ,
         \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 ,
         \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 ,
         \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 ,
         \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 ,
         \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 ,
         \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 ,
         \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 , \29083 , \29084 ,
         \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 ,
         \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 ,
         \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 ,
         \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 ,
         \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 ,
         \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 ,
         \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 ,
         \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 ,
         \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 ,
         \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 , \29183 , \29184 ,
         \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 ,
         \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 ,
         \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 ,
         \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 ,
         \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 ,
         \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 ,
         \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 ,
         \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 ,
         \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 ,
         \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 ,
         \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 ,
         \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 ,
         \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 ,
         \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 ,
         \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 ,
         \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 ,
         \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 ,
         \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 ,
         \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 ,
         \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 ,
         \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 ,
         \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 ,
         \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 ,
         \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 ,
         \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433 , \29434 ,
         \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 ,
         \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 ,
         \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 ,
         \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 ,
         \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 ,
         \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 ,
         \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 ,
         \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 ,
         \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 ,
         \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 ,
         \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 ,
         \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 ,
         \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 ,
         \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 ,
         \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 ,
         \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 ,
         \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 ,
         \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 ,
         \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 ,
         \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 ,
         \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 ,
         \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 ,
         \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 ,
         \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 ,
         \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 ,
         \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 ,
         \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 , \29703 , \29704 ,
         \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 ,
         \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 ,
         \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 ,
         \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 ,
         \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 ,
         \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 ,
         \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 ,
         \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 ,
         \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 ,
         \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 ,
         \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 ,
         \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 ,
         \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833 , \29834 ,
         \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844 ,
         \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 ,
         \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 ,
         \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 ,
         \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 ,
         \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 ,
         \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 ,
         \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 ,
         \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 ,
         \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 ,
         \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 ,
         \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 ,
         \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 ,
         \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 ,
         \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 ,
         \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 ,
         \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 ,
         \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 ,
         \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 ,
         \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 ,
         \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 ,
         \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 ,
         \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 ,
         \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 ,
         \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 ,
         \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 ,
         \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 ,
         \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 , \30113 , \30114 ,
         \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 ,
         \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 ,
         \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 ,
         \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 ,
         \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 ,
         \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 ,
         \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 ,
         \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 ,
         \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 ,
         \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 ,
         \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 ,
         \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 ,
         \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243 , \30244 ,
         \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 ,
         \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 ,
         \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 ,
         \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 ,
         \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 ,
         \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 ,
         \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 ,
         \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 ,
         \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 ,
         \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 ,
         \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 ,
         \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 ,
         \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 ,
         \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 ,
         \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 ,
         \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 ,
         \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 ,
         \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 ,
         \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 ,
         \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 ,
         \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 ,
         \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 ,
         \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 ,
         \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 ,
         \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 ,
         \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 ,
         \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 ,
         \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 ,
         \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 ,
         \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 ,
         \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 ,
         \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 ,
         \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 ,
         \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 ,
         \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 ,
         \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 ,
         \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 ,
         \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 ,
         \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 ,
         \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 ,
         \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 ,
         \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 ,
         \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 ,
         \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 ,
         \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 ,
         \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 ,
         \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 ,
         \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 ,
         \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 ,
         \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 ,
         \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 ,
         \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 ,
         \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 ,
         \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 ,
         \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 ,
         \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 , \30803 , \30804 ,
         \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 , \30813 , \30814 ,
         \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 ,
         \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 ,
         \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 ,
         \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 ,
         \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 ,
         \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874 ,
         \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 ,
         \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 , \30893 , \30894 ,
         \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 ,
         \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 ,
         \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 ,
         \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 ,
         \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 , \30943 , \30944 ,
         \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 ,
         \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 ,
         \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 ,
         \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 ,
         \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 ,
         \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 ,
         \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 ,
         \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 ,
         \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 ,
         \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 ,
         \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 ,
         \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 ,
         \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 ,
         \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 , \31083 , \31084 ,
         \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 ,
         \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 ,
         \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 ,
         \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 ,
         \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 ,
         \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 ,
         \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 ,
         \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 ,
         \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 ,
         \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 ,
         \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 ,
         \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 ,
         \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 ,
         \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 ,
         \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 ,
         \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 ,
         \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 ,
         \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 ,
         \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 ,
         \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 ,
         \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 ,
         \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 ,
         \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 ,
         \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 ,
         \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 ,
         \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 ,
         \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 , \31353 , \31354 ,
         \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 ,
         \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 ,
         \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 ,
         \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 ,
         \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 ,
         \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 ,
         \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 ,
         \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 ,
         \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 ,
         \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 ,
         \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 ,
         \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 ,
         \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483 , \31484 ,
         \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 ,
         \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 ,
         \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 ,
         \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 ,
         \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 ,
         \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 ,
         \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 ,
         \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 ,
         \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 ,
         \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 ,
         \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 ,
         \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 ,
         \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 ,
         \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 ,
         \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 , \31633 , \31634 ,
         \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 ,
         \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 ,
         \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 ,
         \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 ,
         \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 ,
         \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 ,
         \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 ,
         \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 ,
         \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 ,
         \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 ,
         \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 ,
         \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 ,
         \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 ,
         \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 ,
         \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 ,
         \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 ,
         \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 ,
         \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 ,
         \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 ,
         \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 ,
         \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 ,
         \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 ,
         \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 ,
         \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 ,
         \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 ,
         \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 ,
         \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 ,
         \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 ,
         \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 , \31923 , \31924 ,
         \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 ,
         \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 ,
         \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 ,
         \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 ,
         \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 ,
         \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 ,
         \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 ,
         \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 ,
         \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 ,
         \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 ,
         \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 ,
         \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 ,
         \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 , \32053 , \32054 ,
         \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063 , \32064 ,
         \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 ,
         \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 ,
         \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 ,
         \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 ,
         \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 ,
         \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 ,
         \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 ,
         \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 ,
         \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 ,
         \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 ,
         \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 ,
         \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 , \32183 , \32184 ,
         \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 ,
         \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 ,
         \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 ,
         \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 ,
         \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 ,
         \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 ,
         \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 ,
         \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 ,
         \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 ,
         \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 ,
         \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 ,
         \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 , \32303 , \32304 ,
         \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 ,
         \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 ,
         \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 ,
         \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 ,
         \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 ,
         \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 ,
         \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 ,
         \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 ,
         \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 ,
         \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 ,
         \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 ,
         \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 ,
         \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 ,
         \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 ,
         \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 ,
         \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 ,
         \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 ,
         \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 ,
         \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 ,
         \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 ,
         \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 ,
         \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 ,
         \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 ,
         \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 ,
         \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 ,
         \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 ,
         \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 ,
         \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 ,
         \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 ,
         \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 ,
         \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 ,
         \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 ,
         \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 ,
         \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 ,
         \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 ,
         \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 , \32663 , \32664 ,
         \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 ,
         \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 ,
         \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 ,
         \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 ,
         \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 ,
         \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 ,
         \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 ,
         \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 ,
         \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 ,
         \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 ,
         \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 ,
         \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 ,
         \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 , \32793 , \32794 ,
         \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 , \32803 , \32804 ,
         \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 ,
         \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 ,
         \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 ,
         \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 ,
         \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 ,
         \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 ,
         \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 ,
         \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 ,
         \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 ,
         \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 ,
         \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 ,
         \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 ,
         \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 ,
         \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 ,
         \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 ,
         \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 ,
         \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 ,
         \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 ,
         \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 ,
         \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 ,
         \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 ,
         \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 ,
         \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 ,
         \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 ,
         \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 ,
         \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 ,
         \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 ,
         \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 ,
         \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 ,
         \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 , \33103 , \33104 ,
         \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 ,
         \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 , \33123 , \33124 ,
         \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 ,
         \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 , \33143 , \33144 ,
         \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 ,
         \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 ,
         \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 ,
         \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 , \33183 , \33184 ,
         \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 ,
         \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 ,
         \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 ,
         \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 ,
         \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 ,
         \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 ,
         \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 ,
         \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 ,
         \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 ,
         \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 ,
         \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 ,
         \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 ,
         \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 ,
         \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 ,
         \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 ,
         \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 ,
         \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 ,
         \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 ,
         \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 ,
         \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 ,
         \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 ,
         \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 ,
         \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 ,
         \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 ,
         \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 ,
         \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 ,
         \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 ,
         \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 ,
         \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 ,
         \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 ,
         \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 ,
         \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 ,
         \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 ,
         \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 ,
         \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 ,
         \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 ,
         \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 ,
         \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 ,
         \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 ,
         \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 ,
         \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 ,
         \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 ,
         \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613 , \33614 ,
         \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 ,
         \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 ,
         \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 ,
         \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 ,
         \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 ,
         \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 ,
         \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 ,
         \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 ,
         \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 ,
         \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 ,
         \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 ,
         \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 ,
         \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 ,
         \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 ,
         \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 ,
         \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 ,
         \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 ,
         \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 ,
         \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 ,
         \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 ,
         \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 ,
         \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 ,
         \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 ,
         \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 ,
         \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 ,
         \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 ,
         \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 ,
         \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 ,
         \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 ,
         \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 ,
         \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 ,
         \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 ,
         \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 ,
         \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 ,
         \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 ,
         \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 ,
         \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 ,
         \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 ,
         \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 ,
         \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 ,
         \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 ,
         \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 ,
         \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 , \34043 , \34044 ,
         \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 ,
         \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 , \34063 , \34064 ,
         \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 ,
         \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 ,
         \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 ,
         \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 ,
         \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 ,
         \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 ,
         \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 ,
         \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 ,
         \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 ,
         \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 ,
         \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 ,
         \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 ,
         \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 ,
         \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 ,
         \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 ,
         \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 ,
         \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 ,
         \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 ,
         \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 ,
         \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 ,
         \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 ,
         \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 ,
         \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294 ,
         \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 ,
         \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 ,
         \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 ,
         \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 ,
         \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 ,
         \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 ,
         \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 ,
         \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 ,
         \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 ,
         \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 ,
         \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 ,
         \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 ,
         \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 ,
         \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 ,
         \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 ,
         \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 ,
         \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 ,
         \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 ,
         \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 ,
         \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 ,
         \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 ,
         \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 ,
         \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 ,
         \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 ,
         \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 ,
         \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 ,
         \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 ,
         \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 , \34573 , \34574 ,
         \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 ,
         \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 ,
         \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 ,
         \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 ,
         \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 ,
         \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 ,
         \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643 , \34644 ,
         \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 ,
         \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 ,
         \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 ,
         \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 ,
         \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 ,
         \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 ,
         \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 ,
         \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 ,
         \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 ,
         \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 ,
         \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 ,
         \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 ,
         \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 ,
         \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 ,
         \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 ,
         \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 ,
         \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 ,
         \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 ,
         \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 ,
         \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 ,
         \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 ,
         \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 ,
         \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 ,
         \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 ,
         \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 ,
         \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 ,
         \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 ,
         \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 ,
         \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 ,
         \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 ,
         \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 ,
         \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 ,
         \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 ,
         \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 ,
         \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 ,
         \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 ,
         \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 ,
         \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 ,
         \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 ,
         \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 ,
         \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 ,
         \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 ,
         \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 ,
         \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 ,
         \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094 ,
         \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 ,
         \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 ,
         \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 ,
         \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 ,
         \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 ,
         \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 ,
         \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 ,
         \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 ,
         \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 ,
         \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 ,
         \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 ,
         \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 ,
         \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 ,
         \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 ,
         \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 ,
         \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 ,
         \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 ,
         \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 ,
         \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 ,
         \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 ,
         \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 ,
         \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 ,
         \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 ,
         \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 ,
         \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 ,
         \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 ,
         \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 ,
         \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 ,
         \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 ,
         \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394 ,
         \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 ,
         \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 , \35413 , \35414 ,
         \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 ,
         \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 ,
         \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 ,
         \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 ,
         \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 ,
         \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 ,
         \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 ,
         \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 ,
         \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 ,
         \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 ,
         \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 ,
         \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 ,
         \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 ,
         \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 ,
         \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 ,
         \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 , \35573 , \35574 ,
         \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 ,
         \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 ,
         \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 , \35603 , \35604 ,
         \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 ,
         \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 ,
         \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 ,
         \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 ,
         \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 ,
         \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 ,
         \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 ,
         \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684 ,
         \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 ,
         \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 ,
         \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 ,
         \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 ,
         \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 ,
         \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 ,
         \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 ,
         \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 ,
         \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 ,
         \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 ,
         \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 ,
         \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 , \35803 , \35804 ,
         \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 ,
         \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 ,
         \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 ,
         \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 ,
         \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 ,
         \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 ,
         \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 ,
         \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 ,
         \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 ,
         \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 ,
         \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 ,
         \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 ,
         \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 ,
         \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 ,
         \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 ,
         \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 ,
         \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 ,
         \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 ,
         \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 ,
         \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 ,
         \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 ,
         \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 ,
         \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 ,
         \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 ,
         \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 ,
         \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 ,
         \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 ,
         \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 ,
         \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 ,
         \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 ,
         \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 ,
         \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 ,
         \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 ,
         \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 ,
         \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 ,
         \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 ,
         \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 , \36173 , \36174 ,
         \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 ,
         \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 ,
         \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 ,
         \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 ,
         \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 ,
         \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 ,
         \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 ,
         \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 ,
         \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 ,
         \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 ,
         \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 ,
         \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 ,
         \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 ,
         \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 ,
         \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 ,
         \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 ,
         \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 ,
         \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 ,
         \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 ,
         \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 ,
         \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 ,
         \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 ,
         \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 ,
         \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 ,
         \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 ,
         \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 ,
         \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 ,
         \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 ,
         \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 ,
         \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 ,
         \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 ,
         \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 ,
         \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 ,
         \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 ,
         \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 ,
         \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 ,
         \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 ,
         \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 ,
         \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 ,
         \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 ,
         \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 ,
         \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 , \36593 , \36594 ,
         \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 ,
         \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 ,
         \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 ,
         \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 ,
         \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 ,
         \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 ,
         \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 ,
         \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 ,
         \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 ,
         \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 ,
         \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 ,
         \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 ,
         \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 ,
         \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 ,
         \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 ,
         \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 ,
         \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 ,
         \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 ,
         \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 ,
         \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 ,
         \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 ,
         \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 ,
         \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 ,
         \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 ,
         \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 ,
         \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 ,
         \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 ,
         \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 ,
         \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 ,
         \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 ,
         \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 , \36903 , \36904 ,
         \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 ,
         \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 ,
         \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 ,
         \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943 , \36944 ,
         \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 ,
         \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 ,
         \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 ,
         \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 ,
         \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 ,
         \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 ,
         \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 , \37013 , \37014 ,
         \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 ,
         \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 ,
         \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 ,
         \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 ,
         \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 ,
         \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 ,
         \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 ,
         \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 ,
         \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 ,
         \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 ,
         \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 ,
         \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 ,
         \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 ,
         \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 ,
         \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 ,
         \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 ,
         \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 ,
         \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 ,
         \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 ,
         \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 ,
         \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 ,
         \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 ,
         \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 ,
         \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 , \37253 , \37254 ,
         \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 ,
         \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 ,
         \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 ,
         \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 ,
         \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 ,
         \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 ,
         \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 ,
         \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 ,
         \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 ,
         \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 ,
         \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 ,
         \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 ,
         \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 ,
         \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 ,
         \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 ,
         \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 ,
         \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 ,
         \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 ,
         \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 ,
         \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 ,
         \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 ,
         \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 ,
         \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 ,
         \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 ,
         \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 ,
         \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 ,
         \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 ,
         \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 ,
         \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 ,
         \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 ,
         \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 ,
         \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 ,
         \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 ,
         \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 , \37593 , \37594 ,
         \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 ,
         \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 ,
         \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 ,
         \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634 ,
         \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 ,
         \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 ,
         \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 ,
         \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 ,
         \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 ,
         \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 ,
         \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 ,
         \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 ,
         \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 ,
         \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 ,
         \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 ,
         \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 ,
         \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 ,
         \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 ,
         \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 ,
         \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 ,
         \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 ,
         \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 ,
         \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 ,
         \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 ,
         \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 ,
         \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 ,
         \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 ,
         \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 ,
         \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 ,
         \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 ,
         \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 ,
         \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 ,
         \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 ,
         \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 ,
         \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 ,
         \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 ,
         \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 ,
         \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974 ,
         \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 ,
         \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 ,
         \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 ,
         \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 ,
         \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 ,
         \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 ,
         \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 ,
         \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 ,
         \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 ,
         \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 ,
         \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 ,
         \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 ,
         \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 ,
         \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 ,
         \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 ,
         \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 ,
         \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 ,
         \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 ,
         \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 ,
         \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 ,
         \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 ,
         \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 ,
         \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 ,
         \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 ,
         \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 ,
         \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 ,
         \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 ,
         \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 ,
         \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 ,
         \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 ,
         \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 ,
         \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 ,
         \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 ,
         \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 ,
         \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 ,
         \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 ,
         \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 ,
         \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 ,
         \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 ,
         \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 ,
         \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 ,
         \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 ,
         \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 ,
         \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 ,
         \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 ,
         \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 ,
         \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 ,
         \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 ,
         \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 ,
         \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 ,
         \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 ,
         \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 ,
         \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 ,
         \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 ,
         \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 ,
         \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 ,
         \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 ,
         \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 ,
         \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 ,
         \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 ,
         \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 ,
         \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 ,
         \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 ,
         \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 ,
         \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 ,
         \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 ,
         \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 ,
         \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 ,
         \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663 , \38664 ,
         \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 ,
         \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 ,
         \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 ,
         \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 ,
         \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 ,
         \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 ,
         \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 ,
         \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 ,
         \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 ,
         \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 ,
         \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 ,
         \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 ,
         \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 ,
         \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 ,
         \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 ,
         \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 ,
         \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 ,
         \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 ,
         \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 ,
         \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 ,
         \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 ,
         \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 ,
         \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 ,
         \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 ,
         \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 ,
         \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 ,
         \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 ,
         \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 ,
         \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 ,
         \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 ,
         \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 ,
         \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 ,
         \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 ,
         \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 ,
         \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 ,
         \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 ,
         \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 ,
         \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 ,
         \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 ,
         \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 ,
         \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 ,
         \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 ,
         \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 ,
         \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 ,
         \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 ,
         \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 ,
         \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 ,
         \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 ,
         \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 ,
         \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 , \39163 , \39164 ,
         \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 ,
         \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183 , \39184 ,
         \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 ,
         \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 ,
         \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 ,
         \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 ,
         \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 ,
         \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 ,
         \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 ,
         \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 ,
         \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 ,
         \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 ,
         \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 ,
         \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 ,
         \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 ,
         \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 ,
         \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334 ,
         \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 ,
         \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 ,
         \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 ,
         \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 ,
         \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 ,
         \39385 , \39386 , \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 ,
         \39395 , \39396 , \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 ,
         \39405 , \39406 , \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 ,
         \39415 , \39416 , \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 ,
         \39425 , \39426 , \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 ,
         \39435 , \39436 , \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 ,
         \39445 , \39446 , \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 ,
         \39455 , \39456 , \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 ,
         \39465 , \39466 , \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 ,
         \39475 , \39476 , \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 ,
         \39485 , \39486 , \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 ,
         \39495 , \39496 , \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 ,
         \39505 , \39506 , \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 ,
         \39515 , \39516 , \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 ,
         \39525 , \39526 , \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 ,
         \39535 , \39536 , \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 ,
         \39545 , \39546 , \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 ,
         \39555 , \39556 , \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 ,
         \39565 , \39566 , \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 ,
         \39575 , \39576 , \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 ,
         \39585 , \39586 , \39587 , \39588 , \39589 , \39590 , \39591 , \39592 , \39593 , \39594 ,
         \39595 , \39596 , \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 ,
         \39605 , \39606 , \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 ,
         \39615 , \39616 , \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 ,
         \39625 , \39626 , \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 ,
         \39635 , \39636 , \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 ,
         \39645 , \39646 , \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 ,
         \39655 , \39656 , \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 ,
         \39665 , \39666 , \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 ,
         \39675 , \39676 , \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 ,
         \39685 , \39686 , \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 ,
         \39695 , \39696 , \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 ,
         \39705 , \39706 , \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 ,
         \39715 , \39716 , \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 ,
         \39725 , \39726 , \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 ,
         \39735 , \39736 , \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 ,
         \39745 , \39746 , \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 ,
         \39755 , \39756 , \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 ,
         \39765 , \39766 , \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 ,
         \39775 , \39776 , \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 ,
         \39785 , \39786 , \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 ,
         \39795 , \39796 , \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 ,
         \39805 , \39806 , \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 ,
         \39815 , \39816 , \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 ,
         \39825 , \39826 , \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 ,
         \39835 , \39836 , \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 ,
         \39845 , \39846 , \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 ,
         \39855 , \39856 , \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 ,
         \39865 , \39866 , \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 ,
         \39875 , \39876 , \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 ,
         \39885 , \39886 , \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 ,
         \39895 , \39896 , \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 ,
         \39905 , \39906 , \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 ,
         \39915 , \39916 , \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 ,
         \39925 , \39926 , \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 ,
         \39935 , \39936 , \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 ,
         \39945 , \39946 , \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 ,
         \39955 , \39956 , \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963 , \39964 ,
         \39965 , \39966 , \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 ,
         \39975 , \39976 , \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 ,
         \39985 , \39986 , \39987 , \39988 , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 ,
         \39995 , \39996 , \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 ,
         \40005 , \40006 , \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 ,
         \40015 , \40016 , \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 ,
         \40025 , \40026 , \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 ,
         \40035 , \40036 , \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 ,
         \40045 , \40046 , \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 ,
         \40055 , \40056 , \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 ,
         \40065 , \40066 , \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 ,
         \40075 , \40076 , \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 ,
         \40085 , \40086 , \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 ,
         \40095 , \40096 , \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 ,
         \40105 , \40106 , \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 ,
         \40115 , \40116 , \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 ,
         \40125 , \40126 , \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 ,
         \40135 , \40136 , \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 ,
         \40145 , \40146 , \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 ,
         \40155 , \40156 , \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 ,
         \40165 , \40166 , \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 ,
         \40175 , \40176 , \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 ,
         \40185 , \40186 , \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 ,
         \40195 , \40196 , \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204 ,
         \40205 , \40206 , \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 ,
         \40215 , \40216 , \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 ,
         \40225 , \40226 , \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 ,
         \40235 , \40236 , \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 ,
         \40245 , \40246 , \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 ,
         \40255 , \40256 , \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 ,
         \40265 , \40266 , \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 ,
         \40275 , \40276 , \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 ,
         \40285 , \40286 , \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 ,
         \40295 , \40296 , \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 ,
         \40305 , \40306 , \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 ,
         \40315 , \40316 , \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 ,
         \40325 , \40326 , \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 ,
         \40335 , \40336 , \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 ,
         \40345 , \40346 , \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 ,
         \40355 , \40356 , \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 ,
         \40365 , \40366 , \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 ,
         \40375 , \40376 , \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 ,
         \40385 , \40386 , \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 ,
         \40395 , \40396 , \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404 ,
         \40405 , \40406 , \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 ,
         \40415 , \40416 , \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 ,
         \40425 , \40426 , \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 ,
         \40435 , \40436 , \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 ,
         \40445 , \40446 , \40447 , \40448 , \40449 , \40450 , \40451 , \40452 , \40453 , \40454 ,
         \40455 , \40456 , \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 ,
         \40465 , \40466 , \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 ,
         \40475 , \40476 , \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 ,
         \40485 , \40486 , \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 ,
         \40495 , \40496 , \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 ,
         \40505 , \40506 , \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 ,
         \40515 , \40516 , \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 ,
         \40525 , \40526 , \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 ,
         \40535 , \40536 , \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 ,
         \40545 , \40546 , \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 ,
         \40555 , \40556 , \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 ,
         \40565 , \40566 , \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 ,
         \40575 , \40576 , \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 ,
         \40585 , \40586 , \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 ,
         \40595 , \40596 , \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 ,
         \40605 , \40606 , \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 ,
         \40615 , \40616 , \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 ,
         \40625 , \40626 , \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 ,
         \40635 , \40636 , \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 ,
         \40645 , \40646 , \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 ,
         \40655 , \40656 , \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 ,
         \40665 , \40666 , \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 ,
         \40675 , \40676 , \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 ,
         \40685 , \40686 , \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 ,
         \40695 , \40696 , \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 ,
         \40705 , \40706 , \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 ,
         \40715 , \40716 , \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 ,
         \40725 , \40726 , \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 ,
         \40735 , \40736 , \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 ,
         \40745 , \40746 , \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 ,
         \40755 , \40756 , \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 ,
         \40765 , \40766 , \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 ,
         \40775 , \40776 , \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 ,
         \40785 , \40786 , \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 ,
         \40795 , \40796 , \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 ,
         \40805 , \40806 , \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 ,
         \40815 , \40816 , \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 ,
         \40825 , \40826 , \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 ,
         \40835 , \40836 , \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843 , \40844 ,
         \40845 , \40846 , \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 ,
         \40855 , \40856 , \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 ,
         \40865 , \40866 , \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 ,
         \40875 , \40876 , \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 ,
         \40885 , \40886 , \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 ,
         \40895 , \40896 , \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 ,
         \40905 , \40906 , \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 ,
         \40915 , \40916 , \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 ,
         \40925 , \40926 , \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 ,
         \40935 , \40936 , \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 ,
         \40945 , \40946 , \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 ,
         \40955 , \40956 , \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 ,
         \40965 , \40966 , \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 ,
         \40975 , \40976 , \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 ,
         \40985 , \40986 , \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 ,
         \40995 , \40996 , \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 ,
         \41005 , \41006 , \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 ,
         \41015 , \41016 , \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 ,
         \41025 , \41026 , \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 ,
         \41035 , \41036 , \41037 , \41038 , \41039 , \41040 , \41041 , \41042 , \41043 , \41044 ,
         \41045 , \41046 , \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 ,
         \41055 , \41056 , \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 ,
         \41065 , \41066 , \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 ,
         \41075 , \41076 , \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 ,
         \41085 , \41086 , \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 ,
         \41095 , \41096 , \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 ,
         \41105 , \41106 , \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 ,
         \41115 , \41116 , \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 ,
         \41125 , \41126 , \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 ,
         \41135 , \41136 , \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 ,
         \41145 , \41146 , \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 ,
         \41155 , \41156 , \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 ,
         \41165 , \41166 , \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 ,
         \41175 , \41176 , \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 ,
         \41185 , \41186 , \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 ,
         \41195 , \41196 , \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 ,
         \41205 , \41206 , \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 ,
         \41215 , \41216 , \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 ,
         \41225 , \41226 , \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 ,
         \41235 , \41236 , \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 ,
         \41245 , \41246 , \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 ,
         \41255 , \41256 , \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 ,
         \41265 , \41266 , \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 ,
         \41275 , \41276 , \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 ,
         \41285 , \41286 , \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 ,
         \41295 , \41296 , \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 ,
         \41305 , \41306 , \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 ,
         \41315 , \41316 , \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 ,
         \41325 , \41326 , \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 ,
         \41335 , \41336 , \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 ,
         \41345 , \41346 , \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 ,
         \41355 , \41356 , \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 ,
         \41365 , \41366 , \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 ,
         \41375 , \41376 , \41377 , \41378 , \41379 , \41380 , \41381 , \41382 , \41383 , \41384 ,
         \41385 , \41386 , \41387 , \41388 , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 ,
         \41395 , \41396 , \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 ,
         \41405 , \41406 , \41407 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 ,
         \41415 , \41416 , \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 ,
         \41425 , \41426 , \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 ,
         \41435 , \41436 , \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 ,
         \41445 , \41446 , \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 ,
         \41455 , \41456 , \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 ,
         \41465 , \41466 , \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 ,
         \41475 , \41476 , \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 ,
         \41485 , \41486 , \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493 , \41494 ,
         \41495 , \41496 , \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 ,
         \41505 , \41506 , \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 ,
         \41515 , \41516 , \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 ,
         \41525 , \41526 , \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 ,
         \41535 , \41536 , \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 ,
         \41545 , \41546 , \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 ,
         \41555 , \41556 , \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 ,
         \41565 , \41566 , \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 ,
         \41575 , \41576 , \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 ,
         \41585 , \41586 , \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 ,
         \41595 , \41596 , \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 ,
         \41605 , \41606 , \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 ,
         \41615 , \41616 , \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 ,
         \41625 , \41626 , \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 ,
         \41635 , \41636 , \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 ,
         \41645 , \41646 , \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 ,
         \41655 , \41656 , \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 ,
         \41665 , \41666 , \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 ,
         \41675 , \41676 , \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 ,
         \41685 , \41686 , \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 ,
         \41695 , \41696 , \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 ,
         \41705 , \41706 , \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 ,
         \41715 , \41716 , \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 ,
         \41725 , \41726 , \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 ,
         \41735 , \41736 , \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 ,
         \41745 , \41746 , \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 ,
         \41755 , \41756 , \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 ,
         \41765 , \41766 , \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 ,
         \41775 , \41776 , \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 ,
         \41785 , \41786 , \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 ,
         \41795 , \41796 , \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 ,
         \41805 , \41806 , \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 ,
         \41815 , \41816 , \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 ,
         \41825 , \41826 , \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 ,
         \41835 , \41836 , \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 ,
         \41845 , \41846 , \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 ,
         \41855 , \41856 , \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 ,
         \41865 , \41866 , \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 ,
         \41875 , \41876 , \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 ,
         \41885 , \41886 , \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 ,
         \41895 , \41896 , \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 ,
         \41905 , \41906 , \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 ,
         \41915 , \41916 , \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 ,
         \41925 , \41926 , \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 ,
         \41935 , \41936 , \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 ,
         \41945 , \41946 , \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 ,
         \41955 , \41956 , \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963 , \41964 ,
         \41965 , \41966 , \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 ,
         \41975 , \41976 , \41977 , \41978 , \41979 , \41980 , \41981 , \41982 , \41983 , \41984 ,
         \41985 , \41986 , \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 ,
         \41995 , \41996 , \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 ,
         \42005 , \42006 , \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 ,
         \42015 , \42016 , \42017 , \42018 , \42019 , \42020 , \42021 , \42022 , \42023 , \42024 ,
         \42025 , \42026 , \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 ,
         \42035 , \42036 , \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 ,
         \42045 , \42046 , \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 ,
         \42055 , \42056 , \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 ,
         \42065 , \42066 , \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 ,
         \42075 , \42076 , \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084 ,
         \42085 , \42086 , \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 ,
         \42095 , \42096 , \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 ,
         \42105 , \42106 , \42107 , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 ,
         \42115 , \42116 , \42117 , \42118 , \42119 , \42120 , \42121 , \42122 , \42123 , \42124 ,
         \42125 , \42126 , \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 ,
         \42135 , \42136 , \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 ,
         \42145 , \42146 , \42147 , \42148 , \42149 , \42150 , \42151 , \42152 , \42153 , \42154 ,
         \42155 , \42156 , \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163 , \42164 ,
         \42165 , \42166 , \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 ,
         \42175 , \42176 , \42177 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 ,
         \42185 , \42186 , \42187 , \42188 , \42189 , \42190 , \42191 , \42192 , \42193 , \42194 ,
         \42195 , \42196 , \42197 , \42198 , \42199 , \42200 , \42201 , \42202 , \42203 , \42204 ,
         \42205 , \42206 , \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 ,
         \42215 , \42216 , \42217 , \42218 , \42219 , \42220 , \42221 , \42222 , \42223 , \42224 ,
         \42225 , \42226 , \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233 , \42234 ,
         \42235 , \42236 , \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 ,
         \42245 , \42246 , \42247 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 ,
         \42255 , \42256 , \42257 , \42258 , \42259 , \42260 , \42261 , \42262 , \42263 , \42264 ,
         \42265 , \42266 , \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 ,
         \42275 , \42276 , \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 ,
         \42285 , \42286 , \42287 , \42288 , \42289 , \42290 , \42291 , \42292 , \42293 , \42294 ,
         \42295 , \42296 , \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303 , \42304 ,
         \42305 , \42306 , \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 ,
         \42315 , \42316 , \42317 , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 ,
         \42325 , \42326 , \42327 , \42328 , \42329 , \42330 , \42331 , \42332 , \42333 , \42334 ,
         \42335 , \42336 , \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 ,
         \42345 , \42346 , \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 ,
         \42355 , \42356 , \42357 , \42358 , \42359 , \42360 , \42361 , \42362 , \42363 , \42364 ,
         \42365 , \42366 , \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 ,
         \42375 , \42376 , \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 ,
         \42385 , \42386 , \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 ,
         \42395 , \42396 , \42397 , \42398 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 ,
         \42405 , \42406 , \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 ,
         \42415 , \42416 , \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 ,
         \42425 , \42426 , \42427 , \42428 , \42429 , \42430 , \42431 , \42432 , \42433 , \42434 ,
         \42435 , \42436 , \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443 , \42444 ,
         \42445 , \42446 , \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 ,
         \42455 , \42456 , \42457 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 ,
         \42465 , \42466 , \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 ,
         \42475 , \42476 , \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 ,
         \42485 , \42486 , \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 ,
         \42495 , \42496 , \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504 ,
         \42505 , \42506 , \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513 , \42514 ,
         \42515 , \42516 , \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 ,
         \42525 , \42526 , \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533 , \42534 ,
         \42535 , \42536 , \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 ,
         \42545 , \42546 , \42547 , \42548 , \42549 , \42550 , \42551 , \42552 , \42553 , \42554 ,
         \42555 , \42556 , \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 ,
         \42565 , \42566 , \42567 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 ,
         \42575 , \42576 , \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584 ,
         \42585 , \42586 , \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 ,
         \42595 , \42596 , \42597 , \42598 , \42599 , \42600 , \42601 , \42602 , \42603 , \42604 ,
         \42605 , \42606 , \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 ,
         \42615 , \42616 , \42617 , \42618 , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 ,
         \42625 , \42626 , \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 ,
         \42635 , \42636 , \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 ,
         \42645 , \42646 , \42647 , \42648 , \42649 , \42650 , \42651 , \42652 , \42653 , \42654 ,
         \42655 , \42656 , \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 ,
         \42665 , \42666 , \42667 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 ,
         \42675 , \42676 , \42677 , \42678 , \42679 , \42680 , \42681 , \42682 , \42683 , \42684 ,
         \42685 , \42686 , \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 ,
         \42695 , \42696 , \42697 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 ,
         \42705 , \42706 , \42707 , \42708 , \42709 , \42710 , \42711 , \42712 , \42713 , \42714 ,
         \42715 , \42716 , \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 ,
         \42725 , \42726 , \42727 , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 ,
         \42735 , \42736 , \42737 , \42738 , \42739 , \42740 , \42741 , \42742 , \42743 , \42744 ,
         \42745 , \42746 , \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 ,
         \42755 , \42756 , \42757 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 ,
         \42765 , \42766 , \42767 , \42768 , \42769 , \42770 , \42771 , \42772 , \42773 , \42774 ,
         \42775 , \42776 , \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 ,
         \42785 , \42786 , \42787 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 ,
         \42795 , \42796 , \42797 , \42798 , \42799 , \42800 , \42801 , \42802 , \42803 , \42804 ,
         \42805 , \42806 , \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 ,
         \42815 , \42816 , \42817 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 ,
         \42825 , \42826 , \42827 , \42828 , \42829 , \42830 , \42831 , \42832 , \42833 , \42834 ,
         \42835 , \42836 , \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 ,
         \42845 , \42846 , \42847 , \42848 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 ,
         \42855 , \42856 , \42857 , \42858 , \42859 , \42860 , \42861 , \42862 , \42863 , \42864 ,
         \42865 , \42866 , \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 ,
         \42875 , \42876 , \42877 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 ,
         \42885 , \42886 , \42887 , \42888 , \42889 , \42890 , \42891 , \42892 , \42893 , \42894 ,
         \42895 , \42896 , \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 ,
         \42905 , \42906 , \42907 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 ,
         \42915 , \42916 , \42917 , \42918 , \42919 , \42920 , \42921 , \42922 , \42923 , \42924 ,
         \42925 , \42926_nGaee1 , \42927 , \42928 , \42929 , \42930_nGaeaa , \42931 , \42932 , \42933_nGaebf , \42934 ,
         \42935 , \42936 , \42937_nGae73 , \42938 , \42939 , \42940_nGae8d , \42941 , \42942 , \42943 , \42944_nGae30 ,
         \42945 , \42946 , \42947_nGae51 , \42948 , \42949 , \42950 , \42951_nGade1 , \42952 , \42953 , \42954_nGae07 ,
         \42955 , \42956 , \42957 , \42958_nGad8a , \42959 , \42960 , \42961_nGadb3 , \42962 , \42963 , \42964 ,
         \42965_nGad2b , \42966 , \42967 , \42968_nGad59 , \42969 , \42970 , \42971 , \42972_nGacc0 , \42973 , \42974 ,
         \42975_nGacf5 , \42976 , \42977 , \42978 , \42979_nGac4c , \42980 , \42981 , \42982_nGac83 , \42983 , \42984 ,
         \42985 , \42986_nGabce , \42987 , \42988 , \42989_nGac0d , \42990 , \42991 , \42992 , \42993_nGab43 , \42994 ,
         \42995 , \42996_nGab87 , \42997 , \42998 , \42999 , \43000_nGaab0 , \43001 , \43002 , \43003_nGaaf7 , \43004 ,
         \43005 , \43006 , \43007_nGaa15 , \43008 , \43009 , \43010_nGaa61 , \43011 , \43012 , \43013 , \43014_nGa96e ,
         \43015 , \43016 , \43017_nGa9c1 , \43018 , \43019 , \43020 , \43021_nGa8be , \43022 , \43023 , \43024_nGa913 ,
         \43025 , \43026 , \43027 , \43028_nGa804 , \43029 , \43030 , \43031_nGa861 , \43032 , \43033 , \43034 ,
         \43035_nGa740 , \43036 , \43037 , \43038_nGa79f , \43039 , \43040 , \43041 , \43042_nGa672 , \43043 , \43044 ,
         \43045_nGa6d9 , \43046 , \43047 , \43048 , \43049_nGa59a , \43050 , \43051 , \43052_nGa603 , \43053 , \43054 ,
         \43055 , \43056_nGa4bb , \43057 , \43058 , \43059_nGa529 , \43060 , \43061 , \43062 , \43063_nGa3d1 , \43064 ,
         \43065 , \43066_nGa445 , \43067 , \43068 , \43069 , \43070_nGa2da , \43071 , \43072 , \43073_nGa355 , \43074 ,
         \43075 , \43076 , \43077_nGa1d7 , \43078 , \43079 , \43080_nGa257 , \43081 , \43082 , \43083 , \43084_nGa0c9 ,
         \43085 , \43086 , \43087_nGa14f , \43088 , \43089 , \43090 , \43091_nG9fb4 , \43092 , \43093 , \43094_nGa03b ,
         \43095 , \43096 , \43097 , \43098_nG9e96 , \43099 , \43100 , \43101_nG9f25 , \43102 , \43103 , \43104 ,
         \43105_nG9d6b , \43106 , \43107 , \43108_nG9dff , \43109 , \43110 , \43111 , \43112_nG9c34 , \43113 , \43114 ,
         \43115_nG9ccf , \43116 , \43117 , \43118 , \43119_nG9af1 , \43120 , \43121 , \43122_nG9b91 , \43123 , \43124 ,
         \43125 , \43126_nG99a6 , \43127 , \43128 , \43129_nG9a49 , \43130 , \43131 , \43132 , \43133_nG9856 , \43134 ,
         \43135 , \43136_nG98fb , \43137 , \43138 , \43139 , \43140_nG96ff , \43141 , \43142 , \43143_nG97a9 , \43144 ,
         \43145 , \43146 , \43147_nG95a0 , \43148 , \43149 , \43150_nG964d , \43151 , \43152 , \43153 , \43154_nG9436 ,
         \43155 , \43156 , \43157_nG94eb , \43158 , \43159 , \43160 , \43161_nG92bf , \43162 , \43163 , \43164_nG9379 ,
         \43165 , \43166 , \43167 , \43168_nG913c , \43169 , \43170 , \43171_nG91fd , \43172 , \43173 , \43174 ,
         \43175_nG8fb0 , \43176 , \43177 , \43178_nG9073 , \43179 , \43180 , \43181 , \43182_nG8e1a , \43183 , \43184 ,
         \43185_nG8ee5 , \43186 , \43187 , \43188 , \43189_nG8c7a , \43190 , \43191 , \43192_nG8d47 , \43193 , \43194 ,
         \43195 , \43196_nG8ad0 , \43197 , \43198 , \43199_nG8ba5 , \43200 , \43201 , \43202 , \43203_nG8919 , \43204 ,
         \43205 , \43206_nG89f3 , \43207 , \43208 , \43209 , \43210_nG8757 , \43211 , \43212 , \43213_nG8837 , \43214 ,
         \43215 , \43216 , \43217_nG858b , \43218 , \43219 , \43220_nG866f , \43221 , \43222 , \43223 , \43224_nG83b4 ,
         \43225 , \43226 , \43227_nG849f , \43228 , \43229 , \43230 , \43231_nG81d4 , \43232 , \43233 , \43234_nG82c1 ,
         \43235 , \43236 , \43237 , \43238_nG7fea , \43239 , \43240 , \43241_nG80df , \43242 , \43243 , \43244 ,
         \43245_nG7df3 , \43246 , \43247 , \43248_nG7eed , \43249 , \43250 , \43251 , \43252_nG7bf4 , \43253 , \43254 ,
         \43255_nG7cf1 , \43256 , \43257 , \43258 , \43259_nG79f0 , \43260 , \43261 , \43262_nG7aef , \43263 , \43264 ,
         \43265 , \43266_nG77e5 , \43267 , \43268 , \43269_nG78e9 , \43270 , \43271 , \43272 , \43273_nG75cf , \43274 ,
         \43275 , \43276_nG76d9 , \43277 , \43278 , \43279 , \43280_nG73af , \43281 , \43282 , \43283_nG74bd , \43284 ,
         \43285 , \43286 , \43287_nG7188 , \43288 , \43289 , \43290_nG7299 , \43291 , \43292 , \43293 , \43294_nG6f56 ,
         \43295 , \43296 , \43297_nG706f , \43298 , \43299 , \43300 , \43301_nG6d1a , \43302 , \43303 , \43304_nG6e35 ,
         \43305 , \43306 , \43307 , \43308_nG6ad4 , \43309 , \43310 , \43311_nG6bf7 , \43312 , \43313 , \43314 ,
         \43315_nG6881 , \43316 , \43317 , \43318_nG69a9 , \43319 , \43320 , \43321 , \43322_nG6622 , \43323 , \43324 ,
         \43325_nG6751 , \43326 , \43327 , \43328 , \43329_nG63b7 , \43330 , \43331 , \43332_nG64eb , \43333 , \43334 ,
         \43335 , \43336_nG6144 , \43337 , \43338 , \43339_nG627b , \43340 , \43341 , \43342 , \43343_nG5ec9 , \43344 ,
         \43345 , \43346_nG6005 , \43347 , \43348 , \43349 , \43350_nG5c48 , \43351 , \43352 , \43353_nG5d85 , \43354 ,
         \43355 , \43356 , \43357_nG59c5 , \43358 , \43359 , \43360_nG5b03 , \43361 , \43362 , \43363 , \43364_nG5740 ,
         \43365 , \43366 , \43367_nG587f , \43368 , \43369 , \43370 , \43371_nG54b8 , \43372 , \43373 , \43374_nG55f9 ,
         \43375 , \43376 , \43377 , \43378_nG5231 , \43379 , \43380 , \43381_nG536f , \43382 , \43383 , \43384 ,
         \43385_nG4fb4 , \43386 , \43387 , \43388_nG50eb , \43389 , \43390 , \43391 , \43392_nG4d41 , \43393 , \43394 ,
         \43395_nG4e75 , \43396 , \43397 , \43398 , \43399_nG4ad8 , \43400 , \43401 , \43402_nG4c05 , \43403 , \43404 ,
         \43405 , \43406_nG4879 , \43407 , \43408 , \43409_nG49a3 , \43410 , \43411 , \43412 , \43413_nG4624 , \43414 ,
         \43415 , \43416_nG4747 , \43417 , \43418 , \43419 , \43420_nG43d9 , \43421 , \43422 , \43423_nG44f9 , \43424 ,
         \43425 , \43426 , \43427_nG4198 , \43428 , \43429 , \43430_nG42b1 , \43431 , \43432 , \43433 , \43434_nG3f61 ,
         \43435 , \43436 , \43437_nG4077 , \43438 , \43439 , \43440 , \43441_nG3d34 , \43442 , \43443 , \43444_nG3e43 ,
         \43445 , \43446 , \43447 , \43448_nG3b11 , \43449 , \43450 , \43451_nG3c1d , \43452 , \43453 , \43454 ,
         \43455_nG38f8 , \43456 , \43457 , \43458_nG39fd , \43459 , \43460 , \43461 , \43462_nG36e9 , \43463 , \43464 ,
         \43465_nG37eb , \43466 , \43467 , \43468 , \43469_nG34e4 , \43470 , \43471 , \43472_nG35df , \43473 , \43474 ,
         \43475 , \43476_nG32e9 , \43477 , \43478 , \43479_nG33e1 , \43480 , \43481 , \43482 , \43483_nG30f8 , \43484 ,
         \43485 , \43486_nG31e9 , \43487 , \43488 , \43489 , \43490_nG2f11 , \43491 , \43492 , \43493_nG2fff , \43494 ,
         \43495 , \43496 , \43497_nG2d34 , \43498 , \43499 , \43500_nG2e1b , \43501 , \43502 , \43503 , \43504_nG2b5e ,
         \43505 , \43506 , \43507_nG2c45 , \43508 , \43509 , \43510 , \43511_nG2993 , \43512 , \43513 , \43514_nG2a6f ,
         \43515 , \43516 , \43517 , \43518_nG27d5 , \43519 , \43520 , \43521_nG28af , \43522 , \43523 , \43524 ,
         \43525_nG2620 , \43526 , \43527 , \43528_nG26f3 , \43529 , \43530 , \43531 , \43532_nG2475 , \43533 , \43534 ,
         \43535_nG2545 , \43536 , \43537 , \43538 , \43539_nG22d4 , \43540 , \43541 , \43542_nG239d , \43543 , \43544 ,
         \43545 , \43546_nG213d , \43547 , \43548 , \43549_nG2203 , \43550 , \43551 , \43552 , \43553_nG1fb0 , \43554 ,
         \43555 , \43556_nG206f , \43557 , \43558 , \43559 , \43560_nG1e2d , \43561 , \43562 , \43563_nG1ee9 , \43564 ,
         \43565 , \43566 , \43567_nG1cb4 , \43568 , \43569 , \43570_nG1d69 , \43571 , \43572 , \43573 , \43574_nG1b45 ,
         \43575 , \43576 , \43577_nG1bf7 , \43578 , \43579 , \43580 , \43581_nG19e0 , \43582 , \43583 , \43584_nG1a8b ,
         \43585 , \43586 , \43587 , \43588_nG1885 , \43589 , \43590 , \43591_nG192d , \43592 , \43593 , \43594 ,
         \43595_nG1734 , \43596 , \43597 , \43598_nG17d5 , \43599 , \43600 , \43601 , \43602_nG15ed , \43603 , \43604 ,
         \43605_nG168b , \43606 , \43607 , \43608 , \43609_nG14b0 , \43610 , \43611 , \43612_nG1547 , \43613 , \43614 ,
         \43615 , \43616_nG137d , \43617 , \43618 , \43619_nG1411 , \43620 , \43621 , \43622 , \43623_nG1254 , \43624 ,
         \43625 , \43626_nG12e1 , \43627 , \43628 , \43629 , \43630_nG1135 , \43631 , \43632 , \43633_nG11bf , \43634 ,
         \43635 , \43636 , \43637_nG1020 , \43638 , \43639 , \43640_nG10a3 , \43641 , \43642 , \43643 , \43644_nGf15 ,
         \43645 , \43646 , \43647_nGf95 , \43648 , \43649 , \43650 , \43651_nGe14 , \43652 , \43653 , \43654_nGe8d ,
         \43655 , \43656 , \43657 , \43658_nGd1d , \43659 , \43660 , \43661_nGd93 , \43662 , \43663 , \43664 ,
         \43665_nGc30 , \43666 , \43667 , \43668_nGc9f , \43669 , \43670 , \43671 , \43672_nGb4d , \43673 , \43674 ,
         \43675_nGbb9 , \43676 , \43677 , \43678 , \43679_nGa74 , \43680 , \43681 , \43682_nGad9 , \43683 , \43684 ,
         \43685 , \43686_nG9a5 , \43687 , \43688 , \43689_nGa07 , \43690 , \43691 , \43692 , \43693_nG8e0 , \43694 ,
         \43695 , \43696_nG93b , \43697 , \43698 , \43699 , \43700_nG825 , \43701 , \43702 , \43703_nG87d , \43704 ,
         \43705 , \43706 , \43707_nG774 , \43708 , \43709 , \43710_nG7c5 , \43711 , \43712 , \43713 , \43714_nG6cd ,
         \43715 , \43716 , \43717_nG71b , \43718 , \43719 , \43720 , \43721_nG630 , \43722 , \43723 , \43724_nG677 ,
         \43725 , \43726 , \43727 , \43728_nG59d , \43729 , \43730 , \43731_nG5e1 , \43732 , \43733 , \43734 ,
         \43735_nG514 , \43736 , \43737 , \43738_nG551 , \43739 , \43740 , \43741 , \43742_nG495 , \43743 , \43744 ,
         \43745_nG4cf , \43746 , \43747 , \43748 , \43749_nG420 , \43750 , \43751 , \43752_nG453 , \43753 , \43754 ,
         \43755 , \43756_nG3b5 , \43757 , \43758 , \43759_nG3e5 , \43760 , \43761 , \43762 , \43763_nG354 , \43764 ,
         \43765 , \43766_nG37d , \43767 , \43768 , \43769 , \43770_nG2fd , \43771 , \43772 , \43773_nG323 , \43774 ,
         \43775 , \43776 , \43777_nG2b0 , \43778 , \43779 , \43780_nG2cf , \43781 , \43782 , \43783 , \43784_nG26d ,
         \43785 , \43786 , \43787_nG289 , \43788 , \43789 , \43790 , \43791_nG234 , \43792 , \43793 , \43794_nG249 ,
         \43795 , \43796 , \43797 , \43798_nG204 , \43799 , \43800 , \43801_nG217 , \43802 , \43803 , \43804 ,
         \43805_nG1e0 , \43806 , \43807 , \43808_nG1ec , \43809 , \43810 , \43811 , \43812_nG189 , \43813 , \43814 ,
         \43815_nG191 , \43816 , \43817 , \43818 , \43819 , \43820 , \43821 , \43822 , \43823 , \43824 ,
         \43825 , \43826 , \43827 , \43828 , \43829 , \43830 , \43831 , \43832 , \43833 , \43834 ,
         \43835 , \43836 , \43837 , \43838 , \43839 , \43840 , \43841 , \43842 , \43843 , \43844 ,
         \43845 , \43846 , \43847 , \43848 , \43849 , \43850 , \43851 , \43852 , \43853 , \43854 ,
         \43855 , \43856 , \43857 , \43858 , \43859 , \43860 , \43861 , \43862 , \43863 , \43864 ,
         \43865 , \43866 , \43867 , \43868 , \43869 , \43870 , \43871 , \43872 , \43873 , \43874 ,
         \43875 , \43876 , \43877 , \43878 , \43879 , \43880 , \43881 , \43882 , \43883 , \43884 ,
         \43885 , \43886 , \43887 , \43888 , \43889 , \43890 , \43891 , \43892 , \43893 , \43894 ,
         \43895 , \43896 , \43897 , \43898 , \43899 , \43900 , \43901 , \43902 , \43903 , \43904 ,
         \43905 , \43906 , \43907 , \43908 , \43909 , \43910 , \43911 , \43912 , \43913 , \43914 ,
         \43915 , \43916 , \43917 , \43918 , \43919 , \43920 , \43921 , \43922 , \43923 , \43924 ,
         \43925 , \43926 , \43927 , \43928 , \43929 , \43930 , \43931 , \43932 , \43933 , \43934 ,
         \43935 , \43936 , \43937 , \43938 , \43939 , \43940 , \43941 , \43942 , \43943 , \43944 ,
         \43945 , \43946 , \43947 , \43948 , \43949 , \43950 , \43951 , \43952 , \43953 , \43954 ,
         \43955 , \43956 , \43957 , \43958 , \43959 , \43960 , \43961 , \43962 , \43963 , \43964 ,
         \43965 , \43966 , \43967 , \43968 , \43969 , \43970 , \43971 , \43972 , \43973 , \43974 ,
         \43975 , \43976 , \43977 , \43978 , \43979 , \43980 , \43981 , \43982 , \43983 , \43984 ,
         \43985 , \43986 , \43987 , \43988 , \43989 , \43990 , \43991 , \43992 , \43993 , \43994 ,
         \43995 , \43996 , \43997 , \43998 , \43999 , \44000 , \44001 , \44002 , \44003 , \44004 ,
         \44005 , \44006 , \44007 , \44008 , \44009 , \44010 , \44011 , \44012 , \44013 , \44014 ,
         \44015 , \44016 , \44017 , \44018 , \44019 , \44020 , \44021 , \44022 , \44023 , \44024 ,
         \44025 , \44026 , \44027 , \44028 , \44029 , \44030 , \44031 , \44032 , \44033 , \44034 ,
         \44035 , \44036 , \44037 , \44038 , \44039 , \44040 , \44041 , \44042 , \44043 , \44044 ,
         \44045 , \44046 , \44047 , \44048 , \44049 , \44050 , \44051 , \44052 , \44053 , \44054 ,
         \44055 , \44056 , \44057 , \44058 , \44059 , \44060 , \44061 , \44062 , \44063 , \44064 ,
         \44065 , \44066 , \44067 , \44068 , \44069 , \44070 , \44071 , \44072 , \44073 , \44074 ,
         \44075 , \44076 , \44077 , \44078 , \44079 , \44080 , \44081 , \44082 , \44083 , \44084 ,
         \44085 , \44086 , \44087 , \44088 , \44089 , \44090 , \44091 , \44092 , \44093 , \44094 ,
         \44095 , \44096 , \44097 , \44098 , \44099 , \44100 , \44101 , \44102 , \44103 , \44104 ,
         \44105 , \44106 , \44107 , \44108 , \44109 , \44110 , \44111 , \44112 , \44113 , \44114 ,
         \44115 , \44116 , \44117 , \44118 , \44119 , \44120 , \44121 , \44122 , \44123 , \44124 ,
         \44125 , \44126 , \44127 , \44128 , \44129 , \44130 , \44131 , \44132 , \44133 , \44134 ,
         \44135 , \44136 , \44137 , \44138 , \44139 , \44140 , \44141 , \44142 , \44143 , \44144 ,
         \44145 , \44146 , \44147 , \44148 , \44149 , \44150 , \44151 , \44152 , \44153 , \44154 ,
         \44155 , \44156 , \44157 , \44158 , \44159 , \44160 , \44161 , \44162 , \44163 , \44164 ,
         \44165 , \44166 , \44167 , \44168 , \44169 , \44170 , \44171 , \44172 , \44173 , \44174 ,
         \44175 , \44176 , \44177 , \44178 , \44179 , \44180 , \44181 , \44182 , \44183 , \44184 ,
         \44185 , \44186 , \44187 , \44188 , \44189 , \44190 , \44191 , \44192 , \44193 , \44194 ,
         \44195 , \44196 , \44197_nGaee9 , \44198 , \44199 , \44200 , \44201 , \44202 , \44203 , \44204 ,
         \44205 , \44206 , \44207 , \44208 , \44209 , \44210 , \44211 , \44212 , \44213 , \44214 ,
         \44215 , \44216 , \44217 , \44218 , \44219 , \44220 , \44221 , \44222 , \44223 , \44224 ,
         \44225 , \44226 , \44227 , \44228 , \44229 , \44230 , \44231 , \44232 , \44233 , \44234 ,
         \44235 , \44236 , \44237 , \44238 , \44239 , \44240 , \44241 , \44242 , \44243 , \44244 ,
         \44245 , \44246 , \44247 , \44248 , \44249 , \44250 , \44251 , \44252 , \44253 , \44254 ,
         \44255 , \44256 , \44257 , \44258 , \44259 , \44260 , \44261 , \44262_nGaeea , \44263 , \44264 ,
         \44265 , \44266_nGaec7 , \44267_nGaec8 , \44268 , \44269 , \44270 , \44271_nGae95 , \44272_nGae96 , \44273 , \44274 ,
         \44275 , \44276_nGae59 , \44277_nGae5a , \44278 , \44279 , \44280 , \44281_nGae0f , \44282_nGae10 , \44283 , \44284 ,
         \44285 , \44286_nGadbb , \44287_nGadbc , \44288 , \44289 , \44290 , \44291_nGad61 , \44292_nGad62 , \44293 , \44294 ,
         \44295 , \44296_nGacfd , \44297_nGacfe , \44298 , \44299 , \44300 , \44301_nGac8b , \44302_nGac8c , \44303 , \44304 ,
         \44305 , \44306_nGac15 , \44307_nGac16 , \44308 , \44309 , \44310 , \44311_nGab8f , \44312_nGab90 , \44313 , \44314 ,
         \44315 , \44316_nGaaff , \44317_nGab00 , \44318 , \44319 , \44320 , \44321_nGaa69 , \44322_nGaa6a , \44323 , \44324 ,
         \44325 , \44326_nGa9c9 , \44327_nGa9ca , \44328 , \44329 , \44330 , \44331_nGa91b , \44332_nGa91c , \44333 , \44334 ,
         \44335 , \44336_nGa869 , \44337_nGa86a , \44338 , \44339 , \44340 , \44341_nGa7a7 , \44342_nGa7a8 , \44343 , \44344 ,
         \44345 , \44346_nGa6e1 , \44347_nGa6e2 , \44348 , \44349 , \44350 , \44351_nGa60b , \44352_nGa60c , \44353 , \44354 ,
         \44355 , \44356_nGa531 , \44357_nGa532 , \44358 , \44359 , \44360 , \44361_nGa44d , \44362_nGa44e , \44363 , \44364 ,
         \44365 , \44366_nGa35d , \44367_nGa35e , \44368 , \44369 , \44370 , \44371_nGa25f , \44372_nGa260 , \44373 , \44374 ,
         \44375 , \44376_nGa157 , \44377_nGa158 , \44378 , \44379 , \44380 , \44381_nGa043 , \44382_nGa044 , \44383 , \44384 ,
         \44385 , \44386_nG9f2d , \44387_nG9f2e , \44388 , \44389 , \44390 , \44391_nG9e07 , \44392_nG9e08 , \44393 , \44394 ,
         \44395 , \44396_nG9cd7 , \44397_nG9cd8 , \44398 , \44399 , \44400 , \44401_nG9b99 , \44402_nG9b9a , \44403 , \44404 ,
         \44405 , \44406_nG9a51 , \44407_nG9a52 , \44408 , \44409 , \44410 , \44411_nG9903 , \44412_nG9904 , \44413 , \44414 ,
         \44415 , \44416_nG97b1 , \44417_nG97b2 , \44418 , \44419 , \44420 , \44421_nG9655 , \44422_nG9656 , \44423 , \44424 ,
         \44425 , \44426_nG94f3 , \44427_nG94f4 , \44428 , \44429 , \44430 , \44431_nG9381 , \44432_nG9382 , \44433 , \44434 ,
         \44435 , \44436_nG9205 , \44437_nG9206 , \44438 , \44439 , \44440 , \44441_nG907b , \44442_nG907c , \44443 , \44444 ,
         \44445 , \44446_nG8eed , \44447_nG8eee , \44448 , \44449 , \44450 , \44451_nG8d4f , \44452_nG8d50 , \44453 , \44454 ,
         \44455 , \44456_nG8bad , \44457_nG8bae , \44458 , \44459 , \44460 , \44461_nG89fb , \44462_nG89fc , \44463 , \44464 ,
         \44465 , \44466_nG883f , \44467_nG8840 , \44468 , \44469 , \44470 , \44471_nG8677 , \44472_nG8678 , \44473 , \44474 ,
         \44475 , \44476_nG84a7 , \44477_nG84a8 , \44478 , \44479 , \44480 , \44481_nG82c9 , \44482_nG82ca , \44483 , \44484 ,
         \44485 , \44486_nG80e7 , \44487_nG80e8 , \44488 , \44489 , \44490 , \44491_nG7ef5 , \44492_nG7ef6 , \44493 , \44494 ,
         \44495 , \44496_nG7cf9 , \44497_nG7cfa , \44498 , \44499 , \44500 , \44501_nG7af7 , \44502_nG7af8 , \44503 , \44504 ,
         \44505 , \44506_nG78f1 , \44507_nG78f2 , \44508 , \44509 , \44510 , \44511_nG76e1 , \44512_nG76e2 , \44513 , \44514 ,
         \44515 , \44516_nG74c5 , \44517_nG74c6 , \44518 , \44519 , \44520 , \44521_nG72a1 , \44522_nG72a2 , \44523 , \44524 ,
         \44525 , \44526_nG7077 , \44527_nG7078 , \44528 , \44529 , \44530 , \44531_nG6e3d , \44532_nG6e3e , \44533 , \44534 ,
         \44535 , \44536_nG6bff , \44537_nG6c00 , \44538 , \44539 , \44540 , \44541_nG69b1 , \44542_nG69b2 , \44543 , \44544 ,
         \44545 , \44546_nG6759 , \44547_nG675a , \44548 , \44549 , \44550 , \44551_nG64f3 , \44552_nG64f4 , \44553 , \44554 ,
         \44555 , \44556_nG6283 , \44557_nG6284 , \44558 , \44559 , \44560 , \44561_nG600d , \44562_nG600e , \44563 , \44564 ,
         \44565 , \44566_nG5d8d , \44567_nG5d8e , \44568 , \44569 , \44570 , \44571_nG5b0b , \44572_nG5b0c , \44573 , \44574 ,
         \44575 , \44576_nG5887 , \44577_nG5888 , \44578 , \44579 , \44580 , \44581_nG5601 , \44582_nG5602 , \44583 , \44584 ,
         \44585 , \44586_nG5377 , \44587_nG5378 , \44588 , \44589 , \44590 , \44591_nG50f3 , \44592_nG50f4 , \44593 , \44594 ,
         \44595 , \44596_nG4e7d , \44597_nG4e7e , \44598 , \44599 , \44600 , \44601_nG4c0d , \44602_nG4c0e , \44603 , \44604 ,
         \44605 , \44606_nG49ab , \44607_nG49ac , \44608 , \44609 , \44610 , \44611_nG474f , \44612_nG4750 , \44613 , \44614 ,
         \44615 , \44616_nG4501 , \44617_nG4502 , \44618 , \44619 , \44620 , \44621_nG42b9 , \44622_nG42ba , \44623 , \44624 ,
         \44625 , \44626_nG407f , \44627_nG4080 , \44628 , \44629 , \44630 , \44631_nG3e4b , \44632_nG3e4c , \44633 , \44634 ,
         \44635 , \44636_nG3c25 , \44637_nG3c26 , \44638 , \44639 , \44640 , \44641_nG3a05 , \44642_nG3a06 , \44643 , \44644 ,
         \44645 , \44646_nG37f3 , \44647_nG37f4 , \44648 , \44649 , \44650 , \44651_nG35e7 , \44652_nG35e8 , \44653 , \44654 ,
         \44655 , \44656_nG33e9 , \44657_nG33ea , \44658 , \44659 , \44660 , \44661_nG31f1 , \44662_nG31f2 , \44663 , \44664 ,
         \44665 , \44666_nG3007 , \44667_nG3008 , \44668 , \44669 , \44670 , \44671_nG2e23 , \44672_nG2e24 , \44673 , \44674 ,
         \44675 , \44676_nG2c4d , \44677_nG2c4e , \44678 , \44679 , \44680 , \44681_nG2a77 , \44682_nG2a78 , \44683 , \44684 ,
         \44685 , \44686_nG28b7 , \44687_nG28b8 , \44688 , \44689 , \44690 , \44691_nG26fb , \44692_nG26fc , \44693 , \44694 ,
         \44695 , \44696_nG254d , \44697_nG254e , \44698 , \44699 , \44700 , \44701_nG23a5 , \44702_nG23a6 , \44703 , \44704 ,
         \44705 , \44706_nG220b , \44707_nG220c , \44708 , \44709 , \44710 , \44711_nG2077 , \44712_nG2078 , \44713 , \44714 ,
         \44715 , \44716_nG1ef1 , \44717_nG1ef2 , \44718 , \44719 , \44720 , \44721_nG1d71 , \44722_nG1d72 , \44723 , \44724 ,
         \44725 , \44726_nG1bff , \44727_nG1c00 , \44728 , \44729 , \44730 , \44731_nG1a93 , \44732_nG1a94 , \44733 , \44734 ,
         \44735 , \44736_nG1935 , \44737_nG1936 , \44738 , \44739 , \44740 , \44741_nG17dd , \44742_nG17de , \44743 , \44744 ,
         \44745 , \44746_nG1693 , \44747_nG1694 , \44748 , \44749 , \44750 , \44751_nG154f , \44752_nG1550 , \44753 , \44754 ,
         \44755 , \44756_nG1419 , \44757_nG141a , \44758 , \44759 , \44760 , \44761_nG12e9 , \44762_nG12ea , \44763 , \44764 ,
         \44765 , \44766_nG11c7 , \44767_nG11c8 , \44768 , \44769 , \44770 , \44771_nG10ab , \44772_nG10ac , \44773 , \44774 ,
         \44775 , \44776_nGf9d , \44777_nGf9e , \44778 , \44779 , \44780 , \44781_nGe95 , \44782_nGe96 , \44783 , \44784 ,
         \44785 , \44786_nGd9b , \44787_nGd9c , \44788 , \44789 , \44790 , \44791_nGca7 , \44792_nGca8 , \44793 , \44794 ,
         \44795 , \44796_nGbc1 , \44797_nGbc2 , \44798 , \44799 , \44800 , \44801_nGae1 , \44802_nGae2 , \44803 , \44804 ,
         \44805 , \44806_nGa0f , \44807_nGa10 , \44808 , \44809 , \44810 , \44811_nG943 , \44812_nG944 , \44813 , \44814 ,
         \44815 , \44816_nG885 , \44817_nG886 , \44818 , \44819 , \44820 , \44821_nG7cd , \44822_nG7ce , \44823 , \44824 ,
         \44825 , \44826_nG723 , \44827_nG724 , \44828 , \44829 , \44830 , \44831_nG67f , \44832_nG680 , \44833 , \44834 ,
         \44835 , \44836_nG5e9 , \44837_nG5ea , \44838 , \44839 , \44840 , \44841_nG559 , \44842_nG55a , \44843 , \44844 ,
         \44845 , \44846_nG4d7 , \44847_nG4d8 , \44848 , \44849 , \44850 , \44851_nG45b , \44852_nG45c , \44853 ;
buf \U$labaj4529 ( R_101_9cd3d68, \44263 );
buf \U$labaj4530 ( R_102_9cd3e10, \44268 );
buf \U$labaj4531 ( R_103_9cd3eb8, \44273 );
buf \U$labaj4532 ( R_104_9cd3f60, \44278 );
buf \U$labaj4533 ( R_105_9cd4008, \44283 );
buf \U$labaj4534 ( R_106_9cd40b0, \44288 );
buf \U$labaj4535 ( R_107_9cd4158, \44293 );
buf \U$labaj4536 ( R_108_9cd4200, \44298 );
buf \U$labaj4537 ( R_109_9cd42a8, \44303 );
buf \U$labaj4538 ( R_10a_9cd4350, \44308 );
buf \U$labaj4539 ( R_10b_9cd43f8, \44313 );
buf \U$labaj4540 ( R_10c_9cd44a0, \44318 );
buf \U$labaj4541 ( R_10d_9cd4548, \44323 );
buf \U$labaj4542 ( R_10e_9cd45f0, \44328 );
buf \U$labaj4543 ( R_10f_9cd4698, \44333 );
buf \U$labaj4544 ( R_110_9cd4740, \44338 );
buf \U$labaj4545 ( R_111_9cd47e8, \44343 );
buf \U$labaj4546 ( R_112_9cd4890, \44348 );
buf \U$labaj4547 ( R_113_9cd4938, \44353 );
buf \U$labaj4548 ( R_114_9cd49e0, \44358 );
buf \U$labaj4549 ( R_115_9cd4a88, \44363 );
buf \U$labaj4550 ( R_116_9cd4b30, \44368 );
buf \U$labaj4551 ( R_117_9cd4bd8, \44373 );
buf \U$labaj4552 ( R_118_9cd4c80, \44378 );
buf \U$labaj4553 ( R_119_9cd4d28, \44383 );
buf \U$labaj4554 ( R_11a_9cd4dd0, \44388 );
buf \U$labaj4555 ( R_11b_9cd4e78, \44393 );
buf \U$labaj4556 ( R_11c_9cd4f20, \44398 );
buf \U$labaj4557 ( R_11d_9cd4fc8, \44403 );
buf \U$labaj4558 ( R_11e_9cd5070, \44408 );
buf \U$labaj4559 ( R_11f_9cd5118, \44413 );
buf \U$labaj4560 ( R_120_9cd51c0, \44418 );
buf \U$labaj4561 ( R_121_9cd5268, \44423 );
buf \U$labaj4562 ( R_122_9cd5310, \44428 );
buf \U$labaj4563 ( R_123_9cd53b8, \44433 );
buf \U$labaj4564 ( R_124_9cd5460, \44438 );
buf \U$labaj4565 ( R_125_9cd5508, \44443 );
buf \U$labaj4566 ( R_126_9cd55b0, \44448 );
buf \U$labaj4567 ( R_127_9cd5658, \44453 );
buf \U$labaj4568 ( R_128_9cd5700, \44458 );
buf \U$labaj4569 ( R_129_9cd57a8, \44463 );
buf \U$labaj4570 ( R_12a_9cd5850, \44468 );
buf \U$labaj4571 ( R_12b_9cd58f8, \44473 );
buf \U$labaj4572 ( R_12c_9cd59a0, \44478 );
buf \U$labaj4573 ( R_12d_9cd5a48, \44483 );
buf \U$labaj4574 ( R_12e_9cd5af0, \44488 );
buf \U$labaj4575 ( R_12f_9cd5b98, \44493 );
buf \U$labaj4576 ( R_130_9cd5c40, \44498 );
buf \U$labaj4577 ( R_131_9cd5ce8, \44503 );
buf \U$labaj4578 ( R_132_9cd5d90, \44508 );
buf \U$labaj4579 ( R_133_9cd5e38, \44513 );
buf \U$labaj4580 ( R_134_9cd5ee0, \44518 );
buf \U$labaj4581 ( R_135_9cd5f88, \44523 );
buf \U$labaj4582 ( R_136_9cd6030, \44528 );
buf \U$labaj4583 ( R_137_9cd60d8, \44533 );
buf \U$labaj4584 ( R_138_9cd6180, \44538 );
buf \U$labaj4585 ( R_139_9cd6228, \44543 );
buf \U$labaj4586 ( R_13a_9cd62d0, \44548 );
buf \U$labaj4587 ( R_13b_9cd6378, \44553 );
buf \U$labaj4588 ( R_13c_9cd6420, \44558 );
buf \U$labaj4589 ( R_13d_9cd64c8, \44563 );
buf \U$labaj4590 ( R_13e_9cd6570, \44568 );
buf \U$labaj4591 ( R_13f_9cd6618, \44573 );
buf \U$labaj4592 ( R_140_9cd66c0, \44578 );
buf \U$labaj4593 ( R_141_9cd6768, \44583 );
buf \U$labaj4594 ( R_142_9cd6810, \44588 );
buf \U$labaj4595 ( R_143_9cd68b8, \44593 );
buf \U$labaj4596 ( R_144_9cd6960, \44598 );
buf \U$labaj4597 ( R_145_9cd6a08, \44603 );
buf \U$labaj4598 ( R_146_9cd6ab0, \44608 );
buf \U$labaj4599 ( R_147_9cd6b58, \44613 );
buf \U$labaj4600 ( R_148_9cd6c00, \44618 );
buf \U$labaj4601 ( R_149_9cd6ca8, \44623 );
buf \U$labaj4602 ( R_14a_9cd6d50, \44628 );
buf \U$labaj4603 ( R_14b_9cd6df8, \44633 );
buf \U$labaj4604 ( R_14c_9cd6ea0, \44638 );
buf \U$labaj4605 ( R_14d_9cd6f48, \44643 );
buf \U$labaj4606 ( R_14e_9cd6ff0, \44648 );
buf \U$labaj4607 ( R_14f_9cd7098, \44653 );
buf \U$labaj4608 ( R_150_9cd7140, \44658 );
buf \U$labaj4609 ( R_151_9cd71e8, \44663 );
buf \U$labaj4610 ( R_152_9cd7290, \44668 );
buf \U$labaj4611 ( R_153_9cd7338, \44673 );
buf \U$labaj4612 ( R_154_9cd73e0, \44678 );
buf \U$labaj4613 ( R_155_9cd7488, \44683 );
buf \U$labaj4614 ( R_156_9cd7530, \44688 );
buf \U$labaj4615 ( R_157_9cd75d8, \44693 );
buf \U$labaj4616 ( R_158_9cd7680, \44698 );
buf \U$labaj4617 ( R_159_9cd7728, \44703 );
buf \U$labaj4618 ( R_15a_9cd77d0, \44708 );
buf \U$labaj4619 ( R_15b_9cd7878, \44713 );
buf \U$labaj4620 ( R_15c_9cd7920, \44718 );
buf \U$labaj4621 ( R_15d_9cd79c8, \44723 );
buf \U$labaj4622 ( R_15e_9cd7a70, \44728 );
buf \U$labaj4623 ( R_15f_9cd7b18, \44733 );
buf \U$labaj4624 ( R_160_9cd7bc0, \44738 );
buf \U$labaj4625 ( R_161_9cd7c68, \44743 );
buf \U$labaj4626 ( R_162_9cd7d10, \44748 );
buf \U$labaj4627 ( R_163_9cd7db8, \44753 );
buf \U$labaj4628 ( R_164_9cd7e60, \44758 );
buf \U$labaj4629 ( R_165_9cd7f08, \44763 );
buf \U$labaj4630 ( R_166_9cd7fb0, \44768 );
buf \U$labaj4631 ( R_167_9cd8058, \44773 );
buf \U$labaj4632 ( R_168_9cd8100, \44778 );
buf \U$labaj4633 ( R_169_9cd81a8, \44783 );
buf \U$labaj4634 ( R_16a_9cd8250, \44788 );
buf \U$labaj4635 ( R_16b_9cd82f8, \44793 );
buf \U$labaj4636 ( R_16c_9cd83a0, \44798 );
buf \U$labaj4637 ( R_16d_9cd8448, \44803 );
buf \U$labaj4638 ( R_16e_9cd84f0, \44808 );
buf \U$labaj4639 ( R_16f_9cd8598, \44813 );
buf \U$labaj4640 ( R_170_9cd8640, \44818 );
buf \U$labaj4641 ( R_171_9cd86e8, \44823 );
buf \U$labaj4642 ( R_172_9cd8790, \44828 );
buf \U$labaj4643 ( R_173_9cd8838, \44833 );
buf \U$labaj4644 ( R_174_9cd88e0, \44838 );
buf \U$labaj4645 ( R_175_9cd8988, \44843 );
buf \U$labaj4646 ( R_176_9cd8a30, \44848 );
buf \U$labaj4647 ( R_177_9cd8ad8, \44853 );
buf \U$1 ( \378 , RIc2257b0_65);
buf \U$2 ( \379 , RIc2275b0_1);
buf \U$3 ( \380 , RIc227538_2);
xor \U$4 ( \381 , \379 , \380 );
buf \U$5 ( \382 , RIc2274c0_3);
xor \U$6 ( \383 , \380 , \382 );
not \U$7 ( \384 , \383 );
and \U$8 ( \385 , \381 , \384 );
and \U$9 ( \386 , \378 , \385 );
not \U$10 ( \387 , \386 );
and \U$11 ( \388 , \380 , \382 );
not \U$12 ( \389 , \388 );
and \U$13 ( \390 , \379 , \389 );
xnor \U$14 ( \391 , \387 , \390 );
buf \U$15 ( \392 , RIc225738_66);
and \U$16 ( \393 , \392 , \379 );
or \U$17 ( \394 , \391 , \393 );
not \U$18 ( \395 , \390 );
xor \U$19 ( \396 , \394 , \395 );
and \U$20 ( \397 , \378 , \379 );
xor \U$21 ( \398 , \396 , \397 );
buf \U$22 ( \399 , RIc227448_4);
buf \U$23 ( \400 , RIc2273d0_5);
and \U$24 ( \401 , \399 , \400 );
not \U$25 ( \402 , \401 );
and \U$26 ( \403 , \382 , \402 );
not \U$27 ( \404 , \403 );
and \U$28 ( \405 , \392 , \385 );
and \U$29 ( \406 , \378 , \383 );
nor \U$30 ( \407 , \405 , \406 );
xnor \U$31 ( \408 , \407 , \390 );
and \U$32 ( \409 , \404 , \408 );
buf \U$33 ( \410 , RIc2256c0_67);
and \U$34 ( \411 , \410 , \379 );
and \U$35 ( \412 , \408 , \411 );
and \U$36 ( \413 , \404 , \411 );
or \U$37 ( \414 , \409 , \412 , \413 );
xnor \U$38 ( \415 , \391 , \393 );
and \U$39 ( \416 , \414 , \415 );
xor \U$40 ( \417 , \398 , \416 );
xor \U$41 ( \418 , \414 , \415 );
xor \U$42 ( \419 , \382 , \399 );
xor \U$43 ( \420 , \399 , \400 );
not \U$44 ( \421 , \420 );
and \U$45 ( \422 , \419 , \421 );
and \U$46 ( \423 , \378 , \422 );
not \U$47 ( \424 , \423 );
xnor \U$48 ( \425 , \424 , \403 );
and \U$49 ( \426 , \410 , \385 );
and \U$50 ( \427 , \392 , \383 );
nor \U$51 ( \428 , \426 , \427 );
xnor \U$52 ( \429 , \428 , \390 );
and \U$53 ( \430 , \425 , \429 );
buf \U$54 ( \431 , RIc225648_68);
and \U$55 ( \432 , \431 , \379 );
and \U$56 ( \433 , \429 , \432 );
and \U$57 ( \434 , \425 , \432 );
or \U$58 ( \435 , \430 , \433 , \434 );
buf \U$59 ( \436 , RIc227358_6);
buf \U$60 ( \437 , RIc2272e0_7);
and \U$61 ( \438 , \436 , \437 );
not \U$62 ( \439 , \438 );
and \U$63 ( \440 , \400 , \439 );
not \U$64 ( \441 , \440 );
and \U$65 ( \442 , \392 , \422 );
and \U$66 ( \443 , \378 , \420 );
nor \U$67 ( \444 , \442 , \443 );
xnor \U$68 ( \445 , \444 , \403 );
and \U$69 ( \446 , \441 , \445 );
and \U$70 ( \447 , \431 , \385 );
and \U$71 ( \448 , \410 , \383 );
nor \U$72 ( \449 , \447 , \448 );
xnor \U$73 ( \450 , \449 , \390 );
and \U$74 ( \451 , \445 , \450 );
and \U$75 ( \452 , \441 , \450 );
or \U$76 ( \453 , \446 , \451 , \452 );
xor \U$77 ( \454 , \425 , \429 );
xor \U$78 ( \455 , \454 , \432 );
or \U$79 ( \456 , \453 , \455 );
and \U$80 ( \457 , \435 , \456 );
xor \U$81 ( \458 , \404 , \408 );
xor \U$82 ( \459 , \458 , \411 );
and \U$83 ( \460 , \456 , \459 );
and \U$84 ( \461 , \435 , \459 );
or \U$85 ( \462 , \457 , \460 , \461 );
and \U$86 ( \463 , \418 , \462 );
xor \U$87 ( \464 , \418 , \462 );
xor \U$88 ( \465 , \435 , \456 );
xor \U$89 ( \466 , \465 , \459 );
xor \U$90 ( \467 , \400 , \436 );
xor \U$91 ( \468 , \436 , \437 );
not \U$92 ( \469 , \468 );
and \U$93 ( \470 , \467 , \469 );
and \U$94 ( \471 , \378 , \470 );
not \U$95 ( \472 , \471 );
xnor \U$96 ( \473 , \472 , \440 );
and \U$97 ( \474 , \410 , \422 );
and \U$98 ( \475 , \392 , \420 );
nor \U$99 ( \476 , \474 , \475 );
xnor \U$100 ( \477 , \476 , \403 );
and \U$101 ( \478 , \473 , \477 );
buf \U$102 ( \479 , RIc2255d0_69);
and \U$103 ( \480 , \479 , \385 );
and \U$104 ( \481 , \431 , \383 );
nor \U$105 ( \482 , \480 , \481 );
xnor \U$106 ( \483 , \482 , \390 );
and \U$107 ( \484 , \477 , \483 );
and \U$108 ( \485 , \473 , \483 );
or \U$109 ( \486 , \478 , \484 , \485 );
buf \U$110 ( \487 , RIc225558_70);
and \U$111 ( \488 , \487 , \379 );
buf \U$112 ( \489 , \488 );
and \U$113 ( \490 , \486 , \489 );
and \U$114 ( \491 , \479 , \379 );
and \U$115 ( \492 , \489 , \491 );
and \U$116 ( \493 , \486 , \491 );
or \U$117 ( \494 , \490 , \492 , \493 );
buf \U$118 ( \495 , RIc227268_8);
buf \U$119 ( \496 , RIc2271f0_9);
and \U$120 ( \497 , \495 , \496 );
not \U$121 ( \498 , \497 );
and \U$122 ( \499 , \437 , \498 );
not \U$123 ( \500 , \499 );
and \U$124 ( \501 , \392 , \470 );
and \U$125 ( \502 , \378 , \468 );
nor \U$126 ( \503 , \501 , \502 );
xnor \U$127 ( \504 , \503 , \440 );
and \U$128 ( \505 , \500 , \504 );
and \U$129 ( \506 , \431 , \422 );
and \U$130 ( \507 , \410 , \420 );
nor \U$131 ( \508 , \506 , \507 );
xnor \U$132 ( \509 , \508 , \403 );
and \U$133 ( \510 , \504 , \509 );
and \U$134 ( \511 , \500 , \509 );
or \U$135 ( \512 , \505 , \510 , \511 );
xor \U$136 ( \513 , \473 , \477 );
xor \U$137 ( \514 , \513 , \483 );
and \U$138 ( \515 , \512 , \514 );
not \U$139 ( \516 , \488 );
and \U$140 ( \517 , \514 , \516 );
and \U$141 ( \518 , \512 , \516 );
or \U$142 ( \519 , \515 , \517 , \518 );
xor \U$143 ( \520 , \441 , \445 );
xor \U$144 ( \521 , \520 , \450 );
and \U$145 ( \522 , \519 , \521 );
xor \U$146 ( \523 , \486 , \489 );
xor \U$147 ( \524 , \523 , \491 );
and \U$148 ( \525 , \521 , \524 );
and \U$149 ( \526 , \519 , \524 );
or \U$150 ( \527 , \522 , \525 , \526 );
and \U$151 ( \528 , \494 , \527 );
xnor \U$152 ( \529 , \453 , \455 );
and \U$153 ( \530 , \527 , \529 );
and \U$154 ( \531 , \494 , \529 );
or \U$155 ( \532 , \528 , \530 , \531 );
and \U$156 ( \533 , \466 , \532 );
xor \U$157 ( \534 , \466 , \532 );
xor \U$158 ( \535 , \494 , \527 );
xor \U$159 ( \536 , \535 , \529 );
xor \U$160 ( \537 , \437 , \495 );
xor \U$161 ( \538 , \495 , \496 );
not \U$162 ( \539 , \538 );
and \U$163 ( \540 , \537 , \539 );
and \U$164 ( \541 , \378 , \540 );
not \U$165 ( \542 , \541 );
xnor \U$166 ( \543 , \542 , \499 );
and \U$167 ( \544 , \410 , \470 );
and \U$168 ( \545 , \392 , \468 );
nor \U$169 ( \546 , \544 , \545 );
xnor \U$170 ( \547 , \546 , \440 );
and \U$171 ( \548 , \543 , \547 );
and \U$172 ( \549 , \479 , \422 );
and \U$173 ( \550 , \431 , \420 );
nor \U$174 ( \551 , \549 , \550 );
xnor \U$175 ( \552 , \551 , \403 );
and \U$176 ( \553 , \547 , \552 );
and \U$177 ( \554 , \543 , \552 );
or \U$178 ( \555 , \548 , \553 , \554 );
buf \U$179 ( \556 , RIc2254e0_71);
and \U$180 ( \557 , \556 , \385 );
and \U$181 ( \558 , \487 , \383 );
nor \U$182 ( \559 , \557 , \558 );
xnor \U$183 ( \560 , \559 , \390 );
buf \U$184 ( \561 , RIc225468_72);
and \U$185 ( \562 , \561 , \379 );
or \U$186 ( \563 , \560 , \562 );
and \U$187 ( \564 , \555 , \563 );
and \U$188 ( \565 , \487 , \385 );
and \U$189 ( \566 , \479 , \383 );
nor \U$190 ( \567 , \565 , \566 );
xnor \U$191 ( \568 , \567 , \390 );
and \U$192 ( \569 , \563 , \568 );
and \U$193 ( \570 , \555 , \568 );
or \U$194 ( \571 , \564 , \569 , \570 );
and \U$195 ( \572 , \556 , \379 );
xor \U$196 ( \573 , \500 , \504 );
xor \U$197 ( \574 , \573 , \509 );
and \U$198 ( \575 , \572 , \574 );
and \U$199 ( \576 , \571 , \575 );
xor \U$200 ( \577 , \512 , \514 );
xor \U$201 ( \578 , \577 , \516 );
and \U$202 ( \579 , \575 , \578 );
and \U$203 ( \580 , \571 , \578 );
or \U$204 ( \581 , \576 , \579 , \580 );
xor \U$205 ( \582 , \519 , \521 );
xor \U$206 ( \583 , \582 , \524 );
and \U$207 ( \584 , \581 , \583 );
and \U$208 ( \585 , \536 , \584 );
xor \U$209 ( \586 , \536 , \584 );
xor \U$210 ( \587 , \581 , \583 );
buf \U$211 ( \588 , RIc227178_10);
buf \U$212 ( \589 , RIc227100_11);
and \U$213 ( \590 , \588 , \589 );
not \U$214 ( \591 , \590 );
and \U$215 ( \592 , \496 , \591 );
not \U$216 ( \593 , \592 );
and \U$217 ( \594 , \392 , \540 );
and \U$218 ( \595 , \378 , \538 );
nor \U$219 ( \596 , \594 , \595 );
xnor \U$220 ( \597 , \596 , \499 );
and \U$221 ( \598 , \593 , \597 );
and \U$222 ( \599 , \431 , \470 );
and \U$223 ( \600 , \410 , \468 );
nor \U$224 ( \601 , \599 , \600 );
xnor \U$225 ( \602 , \601 , \440 );
and \U$226 ( \603 , \597 , \602 );
and \U$227 ( \604 , \593 , \602 );
or \U$228 ( \605 , \598 , \603 , \604 );
and \U$229 ( \606 , \487 , \422 );
and \U$230 ( \607 , \479 , \420 );
nor \U$231 ( \608 , \606 , \607 );
xnor \U$232 ( \609 , \608 , \403 );
and \U$233 ( \610 , \561 , \385 );
and \U$234 ( \611 , \556 , \383 );
nor \U$235 ( \612 , \610 , \611 );
xnor \U$236 ( \613 , \612 , \390 );
and \U$237 ( \614 , \609 , \613 );
buf \U$238 ( \615 , RIc2253f0_73);
and \U$239 ( \616 , \615 , \379 );
and \U$240 ( \617 , \613 , \616 );
and \U$241 ( \618 , \609 , \616 );
or \U$242 ( \619 , \614 , \617 , \618 );
and \U$243 ( \620 , \605 , \619 );
xnor \U$244 ( \621 , \560 , \562 );
and \U$245 ( \622 , \619 , \621 );
and \U$246 ( \623 , \605 , \621 );
or \U$247 ( \624 , \620 , \622 , \623 );
xor \U$248 ( \625 , \555 , \563 );
xor \U$249 ( \626 , \625 , \568 );
and \U$250 ( \627 , \624 , \626 );
xor \U$251 ( \628 , \572 , \574 );
and \U$252 ( \629 , \626 , \628 );
and \U$253 ( \630 , \624 , \628 );
or \U$254 ( \631 , \627 , \629 , \630 );
xor \U$255 ( \632 , \571 , \575 );
xor \U$256 ( \633 , \632 , \578 );
and \U$257 ( \634 , \631 , \633 );
and \U$258 ( \635 , \587 , \634 );
xor \U$259 ( \636 , \587 , \634 );
xor \U$260 ( \637 , \631 , \633 );
xor \U$261 ( \638 , \496 , \588 );
xor \U$262 ( \639 , \588 , \589 );
not \U$263 ( \640 , \639 );
and \U$264 ( \641 , \638 , \640 );
and \U$265 ( \642 , \378 , \641 );
not \U$266 ( \643 , \642 );
xnor \U$267 ( \644 , \643 , \592 );
and \U$268 ( \645 , \410 , \540 );
and \U$269 ( \646 , \392 , \538 );
nor \U$270 ( \647 , \645 , \646 );
xnor \U$271 ( \648 , \647 , \499 );
and \U$272 ( \649 , \644 , \648 );
and \U$273 ( \650 , \479 , \470 );
and \U$274 ( \651 , \431 , \468 );
nor \U$275 ( \652 , \650 , \651 );
xnor \U$276 ( \653 , \652 , \440 );
and \U$277 ( \654 , \648 , \653 );
and \U$278 ( \655 , \644 , \653 );
or \U$279 ( \656 , \649 , \654 , \655 );
and \U$280 ( \657 , \556 , \422 );
and \U$281 ( \658 , \487 , \420 );
nor \U$282 ( \659 , \657 , \658 );
xnor \U$283 ( \660 , \659 , \403 );
and \U$284 ( \661 , \615 , \385 );
and \U$285 ( \662 , \561 , \383 );
nor \U$286 ( \663 , \661 , \662 );
xnor \U$287 ( \664 , \663 , \390 );
and \U$288 ( \665 , \660 , \664 );
buf \U$289 ( \666 , RIc225378_74);
and \U$290 ( \667 , \666 , \379 );
and \U$291 ( \668 , \664 , \667 );
and \U$292 ( \669 , \660 , \667 );
or \U$293 ( \670 , \665 , \668 , \669 );
and \U$294 ( \671 , \656 , \670 );
xor \U$295 ( \672 , \609 , \613 );
xor \U$296 ( \673 , \672 , \616 );
and \U$297 ( \674 , \670 , \673 );
and \U$298 ( \675 , \656 , \673 );
or \U$299 ( \676 , \671 , \674 , \675 );
xor \U$300 ( \677 , \543 , \547 );
xor \U$301 ( \678 , \677 , \552 );
and \U$302 ( \679 , \676 , \678 );
xor \U$303 ( \680 , \605 , \619 );
xor \U$304 ( \681 , \680 , \621 );
and \U$305 ( \682 , \678 , \681 );
and \U$306 ( \683 , \676 , \681 );
or \U$307 ( \684 , \679 , \682 , \683 );
xor \U$308 ( \685 , \624 , \626 );
xor \U$309 ( \686 , \685 , \628 );
and \U$310 ( \687 , \684 , \686 );
and \U$311 ( \688 , \637 , \687 );
xor \U$312 ( \689 , \637 , \687 );
xor \U$313 ( \690 , \684 , \686 );
and \U$314 ( \691 , \487 , \470 );
and \U$315 ( \692 , \479 , \468 );
nor \U$316 ( \693 , \691 , \692 );
xnor \U$317 ( \694 , \693 , \440 );
and \U$318 ( \695 , \561 , \422 );
and \U$319 ( \696 , \556 , \420 );
nor \U$320 ( \697 , \695 , \696 );
xnor \U$321 ( \698 , \697 , \403 );
and \U$322 ( \699 , \694 , \698 );
and \U$323 ( \700 , \666 , \385 );
and \U$324 ( \701 , \615 , \383 );
nor \U$325 ( \702 , \700 , \701 );
xnor \U$326 ( \703 , \702 , \390 );
and \U$327 ( \704 , \698 , \703 );
and \U$328 ( \705 , \694 , \703 );
or \U$329 ( \706 , \699 , \704 , \705 );
buf \U$330 ( \707 , RIc227088_12);
buf \U$331 ( \708 , RIc227010_13);
and \U$332 ( \709 , \707 , \708 );
not \U$333 ( \710 , \709 );
and \U$334 ( \711 , \589 , \710 );
not \U$335 ( \712 , \711 );
and \U$336 ( \713 , \392 , \641 );
and \U$337 ( \714 , \378 , \639 );
nor \U$338 ( \715 , \713 , \714 );
xnor \U$339 ( \716 , \715 , \592 );
and \U$340 ( \717 , \712 , \716 );
and \U$341 ( \718 , \431 , \540 );
and \U$342 ( \719 , \410 , \538 );
nor \U$343 ( \720 , \718 , \719 );
xnor \U$344 ( \721 , \720 , \499 );
and \U$345 ( \722 , \716 , \721 );
and \U$346 ( \723 , \712 , \721 );
or \U$347 ( \724 , \717 , \722 , \723 );
or \U$348 ( \725 , \706 , \724 );
xor \U$349 ( \726 , \593 , \597 );
xor \U$350 ( \727 , \726 , \602 );
and \U$351 ( \728 , \725 , \727 );
xor \U$352 ( \729 , \656 , \670 );
xor \U$353 ( \730 , \729 , \673 );
and \U$354 ( \731 , \727 , \730 );
and \U$355 ( \732 , \725 , \730 );
or \U$356 ( \733 , \728 , \731 , \732 );
and \U$357 ( \734 , \556 , \470 );
and \U$358 ( \735 , \487 , \468 );
nor \U$359 ( \736 , \734 , \735 );
xnor \U$360 ( \737 , \736 , \440 );
and \U$361 ( \738 , \615 , \422 );
and \U$362 ( \739 , \561 , \420 );
nor \U$363 ( \740 , \738 , \739 );
xnor \U$364 ( \741 , \740 , \403 );
and \U$365 ( \742 , \737 , \741 );
buf \U$366 ( \743 , RIc225300_75);
and \U$367 ( \744 , \743 , \385 );
and \U$368 ( \745 , \666 , \383 );
nor \U$369 ( \746 , \744 , \745 );
xnor \U$370 ( \747 , \746 , \390 );
and \U$371 ( \748 , \741 , \747 );
and \U$372 ( \749 , \737 , \747 );
or \U$373 ( \750 , \742 , \748 , \749 );
xor \U$374 ( \751 , \589 , \707 );
xor \U$375 ( \752 , \707 , \708 );
not \U$376 ( \753 , \752 );
and \U$377 ( \754 , \751 , \753 );
and \U$378 ( \755 , \378 , \754 );
not \U$379 ( \756 , \755 );
xnor \U$380 ( \757 , \756 , \711 );
and \U$381 ( \758 , \410 , \641 );
and \U$382 ( \759 , \392 , \639 );
nor \U$383 ( \760 , \758 , \759 );
xnor \U$384 ( \761 , \760 , \592 );
and \U$385 ( \762 , \757 , \761 );
and \U$386 ( \763 , \479 , \540 );
and \U$387 ( \764 , \431 , \538 );
nor \U$388 ( \765 , \763 , \764 );
xnor \U$389 ( \766 , \765 , \499 );
and \U$390 ( \767 , \761 , \766 );
and \U$391 ( \768 , \757 , \766 );
or \U$392 ( \769 , \762 , \767 , \768 );
and \U$393 ( \770 , \750 , \769 );
buf \U$394 ( \771 , RIc225288_76);
and \U$395 ( \772 , \771 , \379 );
buf \U$396 ( \773 , \772 );
and \U$397 ( \774 , \769 , \773 );
and \U$398 ( \775 , \750 , \773 );
or \U$399 ( \776 , \770 , \774 , \775 );
and \U$400 ( \777 , \743 , \379 );
xor \U$401 ( \778 , \694 , \698 );
xor \U$402 ( \779 , \778 , \703 );
and \U$403 ( \780 , \777 , \779 );
xor \U$404 ( \781 , \712 , \716 );
xor \U$405 ( \782 , \781 , \721 );
and \U$406 ( \783 , \779 , \782 );
and \U$407 ( \784 , \777 , \782 );
or \U$408 ( \785 , \780 , \783 , \784 );
and \U$409 ( \786 , \776 , \785 );
xor \U$410 ( \787 , \660 , \664 );
xor \U$411 ( \788 , \787 , \667 );
and \U$412 ( \789 , \785 , \788 );
and \U$413 ( \790 , \776 , \788 );
or \U$414 ( \791 , \786 , \789 , \790 );
xor \U$415 ( \792 , \644 , \648 );
xor \U$416 ( \793 , \792 , \653 );
xnor \U$417 ( \794 , \706 , \724 );
and \U$418 ( \795 , \793 , \794 );
and \U$419 ( \796 , \791 , \795 );
xor \U$420 ( \797 , \725 , \727 );
xor \U$421 ( \798 , \797 , \730 );
and \U$422 ( \799 , \795 , \798 );
and \U$423 ( \800 , \791 , \798 );
or \U$424 ( \801 , \796 , \799 , \800 );
and \U$425 ( \802 , \733 , \801 );
xor \U$426 ( \803 , \676 , \678 );
xor \U$427 ( \804 , \803 , \681 );
and \U$428 ( \805 , \801 , \804 );
and \U$429 ( \806 , \733 , \804 );
or \U$430 ( \807 , \802 , \805 , \806 );
and \U$431 ( \808 , \690 , \807 );
xor \U$432 ( \809 , \690 , \807 );
xor \U$433 ( \810 , \733 , \801 );
xor \U$434 ( \811 , \810 , \804 );
buf \U$435 ( \812 , RIc226f98_14);
buf \U$436 ( \813 , RIc226f20_15);
and \U$437 ( \814 , \812 , \813 );
not \U$438 ( \815 , \814 );
and \U$439 ( \816 , \708 , \815 );
not \U$440 ( \817 , \816 );
and \U$441 ( \818 , \392 , \754 );
and \U$442 ( \819 , \378 , \752 );
nor \U$443 ( \820 , \818 , \819 );
xnor \U$444 ( \821 , \820 , \711 );
and \U$445 ( \822 , \817 , \821 );
and \U$446 ( \823 , \431 , \641 );
and \U$447 ( \824 , \410 , \639 );
nor \U$448 ( \825 , \823 , \824 );
xnor \U$449 ( \826 , \825 , \592 );
and \U$450 ( \827 , \821 , \826 );
and \U$451 ( \828 , \817 , \826 );
or \U$452 ( \829 , \822 , \827 , \828 );
and \U$453 ( \830 , \487 , \540 );
and \U$454 ( \831 , \479 , \538 );
nor \U$455 ( \832 , \830 , \831 );
xnor \U$456 ( \833 , \832 , \499 );
and \U$457 ( \834 , \561 , \470 );
and \U$458 ( \835 , \556 , \468 );
nor \U$459 ( \836 , \834 , \835 );
xnor \U$460 ( \837 , \836 , \440 );
and \U$461 ( \838 , \833 , \837 );
and \U$462 ( \839 , \666 , \422 );
and \U$463 ( \840 , \615 , \420 );
nor \U$464 ( \841 , \839 , \840 );
xnor \U$465 ( \842 , \841 , \403 );
and \U$466 ( \843 , \837 , \842 );
and \U$467 ( \844 , \833 , \842 );
or \U$468 ( \845 , \838 , \843 , \844 );
and \U$469 ( \846 , \829 , \845 );
and \U$470 ( \847 , \771 , \385 );
and \U$471 ( \848 , \743 , \383 );
nor \U$472 ( \849 , \847 , \848 );
xnor \U$473 ( \850 , \849 , \390 );
buf \U$474 ( \851 , RIc225210_77);
and \U$475 ( \852 , \851 , \379 );
and \U$476 ( \853 , \850 , \852 );
and \U$477 ( \854 , \845 , \853 );
and \U$478 ( \855 , \829 , \853 );
or \U$479 ( \856 , \846 , \854 , \855 );
xor \U$480 ( \857 , \737 , \741 );
xor \U$481 ( \858 , \857 , \747 );
xor \U$482 ( \859 , \757 , \761 );
xor \U$483 ( \860 , \859 , \766 );
and \U$484 ( \861 , \858 , \860 );
not \U$485 ( \862 , \772 );
and \U$486 ( \863 , \860 , \862 );
and \U$487 ( \864 , \858 , \862 );
or \U$488 ( \865 , \861 , \863 , \864 );
and \U$489 ( \866 , \856 , \865 );
xor \U$490 ( \867 , \777 , \779 );
xor \U$491 ( \868 , \867 , \782 );
and \U$492 ( \869 , \865 , \868 );
and \U$493 ( \870 , \856 , \868 );
or \U$494 ( \871 , \866 , \869 , \870 );
xor \U$495 ( \872 , \776 , \785 );
xor \U$496 ( \873 , \872 , \788 );
and \U$497 ( \874 , \871 , \873 );
xor \U$498 ( \875 , \793 , \794 );
and \U$499 ( \876 , \873 , \875 );
and \U$500 ( \877 , \871 , \875 );
or \U$501 ( \878 , \874 , \876 , \877 );
xor \U$502 ( \879 , \791 , \795 );
xor \U$503 ( \880 , \879 , \798 );
and \U$504 ( \881 , \878 , \880 );
and \U$505 ( \882 , \811 , \881 );
xor \U$506 ( \883 , \811 , \881 );
xor \U$507 ( \884 , \878 , \880 );
xor \U$508 ( \885 , \708 , \812 );
xor \U$509 ( \886 , \812 , \813 );
not \U$510 ( \887 , \886 );
and \U$511 ( \888 , \885 , \887 );
and \U$512 ( \889 , \378 , \888 );
not \U$513 ( \890 , \889 );
xnor \U$514 ( \891 , \890 , \816 );
and \U$515 ( \892 , \410 , \754 );
and \U$516 ( \893 , \392 , \752 );
nor \U$517 ( \894 , \892 , \893 );
xnor \U$518 ( \895 , \894 , \711 );
and \U$519 ( \896 , \891 , \895 );
and \U$520 ( \897 , \479 , \641 );
and \U$521 ( \898 , \431 , \639 );
nor \U$522 ( \899 , \897 , \898 );
xnor \U$523 ( \900 , \899 , \592 );
and \U$524 ( \901 , \895 , \900 );
and \U$525 ( \902 , \891 , \900 );
or \U$526 ( \903 , \896 , \901 , \902 );
and \U$527 ( \904 , \556 , \540 );
and \U$528 ( \905 , \487 , \538 );
nor \U$529 ( \906 , \904 , \905 );
xnor \U$530 ( \907 , \906 , \499 );
and \U$531 ( \908 , \615 , \470 );
and \U$532 ( \909 , \561 , \468 );
nor \U$533 ( \910 , \908 , \909 );
xnor \U$534 ( \911 , \910 , \440 );
and \U$535 ( \912 , \907 , \911 );
and \U$536 ( \913 , \743 , \422 );
and \U$537 ( \914 , \666 , \420 );
nor \U$538 ( \915 , \913 , \914 );
xnor \U$539 ( \916 , \915 , \403 );
and \U$540 ( \917 , \911 , \916 );
and \U$541 ( \918 , \907 , \916 );
or \U$542 ( \919 , \912 , \917 , \918 );
and \U$543 ( \920 , \903 , \919 );
and \U$544 ( \921 , \851 , \385 );
and \U$545 ( \922 , \771 , \383 );
nor \U$546 ( \923 , \921 , \922 );
xnor \U$547 ( \924 , \923 , \390 );
buf \U$548 ( \925 , RIc225198_78);
and \U$549 ( \926 , \925 , \379 );
or \U$550 ( \927 , \924 , \926 );
and \U$551 ( \928 , \919 , \927 );
and \U$552 ( \929 , \903 , \927 );
or \U$553 ( \930 , \920 , \928 , \929 );
xor \U$554 ( \931 , \817 , \821 );
xor \U$555 ( \932 , \931 , \826 );
xor \U$556 ( \933 , \833 , \837 );
xor \U$557 ( \934 , \933 , \842 );
and \U$558 ( \935 , \932 , \934 );
xor \U$559 ( \936 , \850 , \852 );
and \U$560 ( \937 , \934 , \936 );
and \U$561 ( \938 , \932 , \936 );
or \U$562 ( \939 , \935 , \937 , \938 );
and \U$563 ( \940 , \930 , \939 );
xor \U$564 ( \941 , \858 , \860 );
xor \U$565 ( \942 , \941 , \862 );
and \U$566 ( \943 , \939 , \942 );
and \U$567 ( \944 , \930 , \942 );
or \U$568 ( \945 , \940 , \943 , \944 );
xor \U$569 ( \946 , \750 , \769 );
xor \U$570 ( \947 , \946 , \773 );
and \U$571 ( \948 , \945 , \947 );
xor \U$572 ( \949 , \856 , \865 );
xor \U$573 ( \950 , \949 , \868 );
and \U$574 ( \951 , \947 , \950 );
and \U$575 ( \952 , \945 , \950 );
or \U$576 ( \953 , \948 , \951 , \952 );
xor \U$577 ( \954 , \871 , \873 );
xor \U$578 ( \955 , \954 , \875 );
and \U$579 ( \956 , \953 , \955 );
and \U$580 ( \957 , \884 , \956 );
xor \U$581 ( \958 , \884 , \956 );
xor \U$582 ( \959 , \953 , \955 );
buf \U$583 ( \960 , RIc226ea8_16);
buf \U$584 ( \961 , RIc226e30_17);
and \U$585 ( \962 , \960 , \961 );
not \U$586 ( \963 , \962 );
and \U$587 ( \964 , \813 , \963 );
not \U$588 ( \965 , \964 );
and \U$589 ( \966 , \392 , \888 );
and \U$590 ( \967 , \378 , \886 );
nor \U$591 ( \968 , \966 , \967 );
xnor \U$592 ( \969 , \968 , \816 );
and \U$593 ( \970 , \965 , \969 );
and \U$594 ( \971 , \431 , \754 );
and \U$595 ( \972 , \410 , \752 );
nor \U$596 ( \973 , \971 , \972 );
xnor \U$597 ( \974 , \973 , \711 );
and \U$598 ( \975 , \969 , \974 );
and \U$599 ( \976 , \965 , \974 );
or \U$600 ( \977 , \970 , \975 , \976 );
and \U$601 ( \978 , \771 , \422 );
and \U$602 ( \979 , \743 , \420 );
nor \U$603 ( \980 , \978 , \979 );
xnor \U$604 ( \981 , \980 , \403 );
and \U$605 ( \982 , \925 , \385 );
and \U$606 ( \983 , \851 , \383 );
nor \U$607 ( \984 , \982 , \983 );
xnor \U$608 ( \985 , \984 , \390 );
and \U$609 ( \986 , \981 , \985 );
buf \U$610 ( \987 , RIc225120_79);
and \U$611 ( \988 , \987 , \379 );
and \U$612 ( \989 , \985 , \988 );
and \U$613 ( \990 , \981 , \988 );
or \U$614 ( \991 , \986 , \989 , \990 );
and \U$615 ( \992 , \977 , \991 );
and \U$616 ( \993 , \487 , \641 );
and \U$617 ( \994 , \479 , \639 );
nor \U$618 ( \995 , \993 , \994 );
xnor \U$619 ( \996 , \995 , \592 );
and \U$620 ( \997 , \561 , \540 );
and \U$621 ( \998 , \556 , \538 );
nor \U$622 ( \999 , \997 , \998 );
xnor \U$623 ( \1000 , \999 , \499 );
and \U$624 ( \1001 , \996 , \1000 );
and \U$625 ( \1002 , \666 , \470 );
and \U$626 ( \1003 , \615 , \468 );
nor \U$627 ( \1004 , \1002 , \1003 );
xnor \U$628 ( \1005 , \1004 , \440 );
and \U$629 ( \1006 , \1000 , \1005 );
and \U$630 ( \1007 , \996 , \1005 );
or \U$631 ( \1008 , \1001 , \1006 , \1007 );
and \U$632 ( \1009 , \991 , \1008 );
and \U$633 ( \1010 , \977 , \1008 );
or \U$634 ( \1011 , \992 , \1009 , \1010 );
xor \U$635 ( \1012 , \891 , \895 );
xor \U$636 ( \1013 , \1012 , \900 );
xor \U$637 ( \1014 , \907 , \911 );
xor \U$638 ( \1015 , \1014 , \916 );
and \U$639 ( \1016 , \1013 , \1015 );
xnor \U$640 ( \1017 , \924 , \926 );
and \U$641 ( \1018 , \1015 , \1017 );
and \U$642 ( \1019 , \1013 , \1017 );
or \U$643 ( \1020 , \1016 , \1018 , \1019 );
and \U$644 ( \1021 , \1011 , \1020 );
xor \U$645 ( \1022 , \932 , \934 );
xor \U$646 ( \1023 , \1022 , \936 );
and \U$647 ( \1024 , \1020 , \1023 );
and \U$648 ( \1025 , \1011 , \1023 );
or \U$649 ( \1026 , \1021 , \1024 , \1025 );
xor \U$650 ( \1027 , \829 , \845 );
xor \U$651 ( \1028 , \1027 , \853 );
and \U$652 ( \1029 , \1026 , \1028 );
xor \U$653 ( \1030 , \930 , \939 );
xor \U$654 ( \1031 , \1030 , \942 );
and \U$655 ( \1032 , \1028 , \1031 );
and \U$656 ( \1033 , \1026 , \1031 );
or \U$657 ( \1034 , \1029 , \1032 , \1033 );
xor \U$658 ( \1035 , \945 , \947 );
xor \U$659 ( \1036 , \1035 , \950 );
and \U$660 ( \1037 , \1034 , \1036 );
and \U$661 ( \1038 , \959 , \1037 );
xor \U$662 ( \1039 , \959 , \1037 );
xor \U$663 ( \1040 , \1034 , \1036 );
and \U$664 ( \1041 , \851 , \422 );
and \U$665 ( \1042 , \771 , \420 );
nor \U$666 ( \1043 , \1041 , \1042 );
xnor \U$667 ( \1044 , \1043 , \403 );
and \U$668 ( \1045 , \987 , \385 );
and \U$669 ( \1046 , \925 , \383 );
nor \U$670 ( \1047 , \1045 , \1046 );
xnor \U$671 ( \1048 , \1047 , \390 );
and \U$672 ( \1049 , \1044 , \1048 );
buf \U$673 ( \1050 , RIc2250a8_80);
and \U$674 ( \1051 , \1050 , \379 );
and \U$675 ( \1052 , \1048 , \1051 );
and \U$676 ( \1053 , \1044 , \1051 );
or \U$677 ( \1054 , \1049 , \1052 , \1053 );
xor \U$678 ( \1055 , \813 , \960 );
xor \U$679 ( \1056 , \960 , \961 );
not \U$680 ( \1057 , \1056 );
and \U$681 ( \1058 , \1055 , \1057 );
and \U$682 ( \1059 , \378 , \1058 );
not \U$683 ( \1060 , \1059 );
xnor \U$684 ( \1061 , \1060 , \964 );
and \U$685 ( \1062 , \410 , \888 );
and \U$686 ( \1063 , \392 , \886 );
nor \U$687 ( \1064 , \1062 , \1063 );
xnor \U$688 ( \1065 , \1064 , \816 );
and \U$689 ( \1066 , \1061 , \1065 );
and \U$690 ( \1067 , \479 , \754 );
and \U$691 ( \1068 , \431 , \752 );
nor \U$692 ( \1069 , \1067 , \1068 );
xnor \U$693 ( \1070 , \1069 , \711 );
and \U$694 ( \1071 , \1065 , \1070 );
and \U$695 ( \1072 , \1061 , \1070 );
or \U$696 ( \1073 , \1066 , \1071 , \1072 );
and \U$697 ( \1074 , \1054 , \1073 );
and \U$698 ( \1075 , \556 , \641 );
and \U$699 ( \1076 , \487 , \639 );
nor \U$700 ( \1077 , \1075 , \1076 );
xnor \U$701 ( \1078 , \1077 , \592 );
and \U$702 ( \1079 , \615 , \540 );
and \U$703 ( \1080 , \561 , \538 );
nor \U$704 ( \1081 , \1079 , \1080 );
xnor \U$705 ( \1082 , \1081 , \499 );
and \U$706 ( \1083 , \1078 , \1082 );
and \U$707 ( \1084 , \743 , \470 );
and \U$708 ( \1085 , \666 , \468 );
nor \U$709 ( \1086 , \1084 , \1085 );
xnor \U$710 ( \1087 , \1086 , \440 );
and \U$711 ( \1088 , \1082 , \1087 );
and \U$712 ( \1089 , \1078 , \1087 );
or \U$713 ( \1090 , \1083 , \1088 , \1089 );
and \U$714 ( \1091 , \1073 , \1090 );
and \U$715 ( \1092 , \1054 , \1090 );
or \U$716 ( \1093 , \1074 , \1091 , \1092 );
xor \U$717 ( \1094 , \965 , \969 );
xor \U$718 ( \1095 , \1094 , \974 );
xor \U$719 ( \1096 , \981 , \985 );
xor \U$720 ( \1097 , \1096 , \988 );
and \U$721 ( \1098 , \1095 , \1097 );
xor \U$722 ( \1099 , \996 , \1000 );
xor \U$723 ( \1100 , \1099 , \1005 );
and \U$724 ( \1101 , \1097 , \1100 );
and \U$725 ( \1102 , \1095 , \1100 );
or \U$726 ( \1103 , \1098 , \1101 , \1102 );
and \U$727 ( \1104 , \1093 , \1103 );
xor \U$728 ( \1105 , \1013 , \1015 );
xor \U$729 ( \1106 , \1105 , \1017 );
and \U$730 ( \1107 , \1103 , \1106 );
and \U$731 ( \1108 , \1093 , \1106 );
or \U$732 ( \1109 , \1104 , \1107 , \1108 );
xor \U$733 ( \1110 , \903 , \919 );
xor \U$734 ( \1111 , \1110 , \927 );
and \U$735 ( \1112 , \1109 , \1111 );
xor \U$736 ( \1113 , \1011 , \1020 );
xor \U$737 ( \1114 , \1113 , \1023 );
and \U$738 ( \1115 , \1111 , \1114 );
and \U$739 ( \1116 , \1109 , \1114 );
or \U$740 ( \1117 , \1112 , \1115 , \1116 );
xor \U$741 ( \1118 , \1026 , \1028 );
xor \U$742 ( \1119 , \1118 , \1031 );
and \U$743 ( \1120 , \1117 , \1119 );
and \U$744 ( \1121 , \1040 , \1120 );
xor \U$745 ( \1122 , \1040 , \1120 );
xor \U$746 ( \1123 , \1117 , \1119 );
and \U$747 ( \1124 , \487 , \754 );
and \U$748 ( \1125 , \479 , \752 );
nor \U$749 ( \1126 , \1124 , \1125 );
xnor \U$750 ( \1127 , \1126 , \711 );
and \U$751 ( \1128 , \561 , \641 );
and \U$752 ( \1129 , \556 , \639 );
nor \U$753 ( \1130 , \1128 , \1129 );
xnor \U$754 ( \1131 , \1130 , \592 );
and \U$755 ( \1132 , \1127 , \1131 );
and \U$756 ( \1133 , \666 , \540 );
and \U$757 ( \1134 , \615 , \538 );
nor \U$758 ( \1135 , \1133 , \1134 );
xnor \U$759 ( \1136 , \1135 , \499 );
and \U$760 ( \1137 , \1131 , \1136 );
and \U$761 ( \1138 , \1127 , \1136 );
or \U$762 ( \1139 , \1132 , \1137 , \1138 );
buf \U$763 ( \1140 , RIc226db8_18);
buf \U$764 ( \1141 , RIc226d40_19);
and \U$765 ( \1142 , \1140 , \1141 );
not \U$766 ( \1143 , \1142 );
and \U$767 ( \1144 , \961 , \1143 );
not \U$768 ( \1145 , \1144 );
and \U$769 ( \1146 , \392 , \1058 );
and \U$770 ( \1147 , \378 , \1056 );
nor \U$771 ( \1148 , \1146 , \1147 );
xnor \U$772 ( \1149 , \1148 , \964 );
and \U$773 ( \1150 , \1145 , \1149 );
and \U$774 ( \1151 , \431 , \888 );
and \U$775 ( \1152 , \410 , \886 );
nor \U$776 ( \1153 , \1151 , \1152 );
xnor \U$777 ( \1154 , \1153 , \816 );
and \U$778 ( \1155 , \1149 , \1154 );
and \U$779 ( \1156 , \1145 , \1154 );
or \U$780 ( \1157 , \1150 , \1155 , \1156 );
and \U$781 ( \1158 , \1139 , \1157 );
and \U$782 ( \1159 , \771 , \470 );
and \U$783 ( \1160 , \743 , \468 );
nor \U$784 ( \1161 , \1159 , \1160 );
xnor \U$785 ( \1162 , \1161 , \440 );
and \U$786 ( \1163 , \925 , \422 );
and \U$787 ( \1164 , \851 , \420 );
nor \U$788 ( \1165 , \1163 , \1164 );
xnor \U$789 ( \1166 , \1165 , \403 );
and \U$790 ( \1167 , \1162 , \1166 );
and \U$791 ( \1168 , \1050 , \385 );
and \U$792 ( \1169 , \987 , \383 );
nor \U$793 ( \1170 , \1168 , \1169 );
xnor \U$794 ( \1171 , \1170 , \390 );
and \U$795 ( \1172 , \1166 , \1171 );
and \U$796 ( \1173 , \1162 , \1171 );
or \U$797 ( \1174 , \1167 , \1172 , \1173 );
and \U$798 ( \1175 , \1157 , \1174 );
and \U$799 ( \1176 , \1139 , \1174 );
or \U$800 ( \1177 , \1158 , \1175 , \1176 );
xor \U$801 ( \1178 , \1044 , \1048 );
xor \U$802 ( \1179 , \1178 , \1051 );
xor \U$803 ( \1180 , \1078 , \1082 );
xor \U$804 ( \1181 , \1180 , \1087 );
or \U$805 ( \1182 , \1179 , \1181 );
and \U$806 ( \1183 , \1177 , \1182 );
xor \U$807 ( \1184 , \1095 , \1097 );
xor \U$808 ( \1185 , \1184 , \1100 );
and \U$809 ( \1186 , \1182 , \1185 );
and \U$810 ( \1187 , \1177 , \1185 );
or \U$811 ( \1188 , \1183 , \1186 , \1187 );
xor \U$812 ( \1189 , \977 , \991 );
xor \U$813 ( \1190 , \1189 , \1008 );
and \U$814 ( \1191 , \1188 , \1190 );
xor \U$815 ( \1192 , \1093 , \1103 );
xor \U$816 ( \1193 , \1192 , \1106 );
and \U$817 ( \1194 , \1190 , \1193 );
and \U$818 ( \1195 , \1188 , \1193 );
or \U$819 ( \1196 , \1191 , \1194 , \1195 );
xor \U$820 ( \1197 , \1109 , \1111 );
xor \U$821 ( \1198 , \1197 , \1114 );
and \U$822 ( \1199 , \1196 , \1198 );
and \U$823 ( \1200 , \1123 , \1199 );
xor \U$824 ( \1201 , \1123 , \1199 );
xor \U$825 ( \1202 , \1196 , \1198 );
and \U$826 ( \1203 , \556 , \754 );
and \U$827 ( \1204 , \487 , \752 );
nor \U$828 ( \1205 , \1203 , \1204 );
xnor \U$829 ( \1206 , \1205 , \711 );
and \U$830 ( \1207 , \615 , \641 );
and \U$831 ( \1208 , \561 , \639 );
nor \U$832 ( \1209 , \1207 , \1208 );
xnor \U$833 ( \1210 , \1209 , \592 );
and \U$834 ( \1211 , \1206 , \1210 );
and \U$835 ( \1212 , \743 , \540 );
and \U$836 ( \1213 , \666 , \538 );
nor \U$837 ( \1214 , \1212 , \1213 );
xnor \U$838 ( \1215 , \1214 , \499 );
and \U$839 ( \1216 , \1210 , \1215 );
and \U$840 ( \1217 , \1206 , \1215 );
or \U$841 ( \1218 , \1211 , \1216 , \1217 );
xor \U$842 ( \1219 , \961 , \1140 );
xor \U$843 ( \1220 , \1140 , \1141 );
not \U$844 ( \1221 , \1220 );
and \U$845 ( \1222 , \1219 , \1221 );
and \U$846 ( \1223 , \378 , \1222 );
not \U$847 ( \1224 , \1223 );
xnor \U$848 ( \1225 , \1224 , \1144 );
and \U$849 ( \1226 , \410 , \1058 );
and \U$850 ( \1227 , \392 , \1056 );
nor \U$851 ( \1228 , \1226 , \1227 );
xnor \U$852 ( \1229 , \1228 , \964 );
and \U$853 ( \1230 , \1225 , \1229 );
and \U$854 ( \1231 , \479 , \888 );
and \U$855 ( \1232 , \431 , \886 );
nor \U$856 ( \1233 , \1231 , \1232 );
xnor \U$857 ( \1234 , \1233 , \816 );
and \U$858 ( \1235 , \1229 , \1234 );
and \U$859 ( \1236 , \1225 , \1234 );
or \U$860 ( \1237 , \1230 , \1235 , \1236 );
and \U$861 ( \1238 , \1218 , \1237 );
and \U$862 ( \1239 , \851 , \470 );
and \U$863 ( \1240 , \771 , \468 );
nor \U$864 ( \1241 , \1239 , \1240 );
xnor \U$865 ( \1242 , \1241 , \440 );
and \U$866 ( \1243 , \987 , \422 );
and \U$867 ( \1244 , \925 , \420 );
nor \U$868 ( \1245 , \1243 , \1244 );
xnor \U$869 ( \1246 , \1245 , \403 );
and \U$870 ( \1247 , \1242 , \1246 );
buf \U$871 ( \1248 , RIc225030_81);
and \U$872 ( \1249 , \1248 , \385 );
and \U$873 ( \1250 , \1050 , \383 );
nor \U$874 ( \1251 , \1249 , \1250 );
xnor \U$875 ( \1252 , \1251 , \390 );
and \U$876 ( \1253 , \1246 , \1252 );
and \U$877 ( \1254 , \1242 , \1252 );
or \U$878 ( \1255 , \1247 , \1253 , \1254 );
and \U$879 ( \1256 , \1237 , \1255 );
and \U$880 ( \1257 , \1218 , \1255 );
or \U$881 ( \1258 , \1238 , \1256 , \1257 );
and \U$882 ( \1259 , \1248 , \379 );
xor \U$883 ( \1260 , \1127 , \1131 );
xor \U$884 ( \1261 , \1260 , \1136 );
and \U$885 ( \1262 , \1259 , \1261 );
xor \U$886 ( \1263 , \1162 , \1166 );
xor \U$887 ( \1264 , \1263 , \1171 );
and \U$888 ( \1265 , \1261 , \1264 );
and \U$889 ( \1266 , \1259 , \1264 );
or \U$890 ( \1267 , \1262 , \1265 , \1266 );
and \U$891 ( \1268 , \1258 , \1267 );
xor \U$892 ( \1269 , \1061 , \1065 );
xor \U$893 ( \1270 , \1269 , \1070 );
and \U$894 ( \1271 , \1267 , \1270 );
and \U$895 ( \1272 , \1258 , \1270 );
or \U$896 ( \1273 , \1268 , \1271 , \1272 );
xor \U$897 ( \1274 , \1054 , \1073 );
xor \U$898 ( \1275 , \1274 , \1090 );
and \U$899 ( \1276 , \1273 , \1275 );
xor \U$900 ( \1277 , \1177 , \1182 );
xor \U$901 ( \1278 , \1277 , \1185 );
and \U$902 ( \1279 , \1275 , \1278 );
and \U$903 ( \1280 , \1273 , \1278 );
or \U$904 ( \1281 , \1276 , \1279 , \1280 );
buf \U$905 ( \1282 , RIc226cc8_20);
buf \U$906 ( \1283 , RIc226c50_21);
and \U$907 ( \1284 , \1282 , \1283 );
not \U$908 ( \1285 , \1284 );
and \U$909 ( \1286 , \1141 , \1285 );
not \U$910 ( \1287 , \1286 );
and \U$911 ( \1288 , \392 , \1222 );
and \U$912 ( \1289 , \378 , \1220 );
nor \U$913 ( \1290 , \1288 , \1289 );
xnor \U$914 ( \1291 , \1290 , \1144 );
and \U$915 ( \1292 , \1287 , \1291 );
and \U$916 ( \1293 , \431 , \1058 );
and \U$917 ( \1294 , \410 , \1056 );
nor \U$918 ( \1295 , \1293 , \1294 );
xnor \U$919 ( \1296 , \1295 , \964 );
and \U$920 ( \1297 , \1291 , \1296 );
and \U$921 ( \1298 , \1287 , \1296 );
or \U$922 ( \1299 , \1292 , \1297 , \1298 );
and \U$923 ( \1300 , \487 , \888 );
and \U$924 ( \1301 , \479 , \886 );
nor \U$925 ( \1302 , \1300 , \1301 );
xnor \U$926 ( \1303 , \1302 , \816 );
and \U$927 ( \1304 , \561 , \754 );
and \U$928 ( \1305 , \556 , \752 );
nor \U$929 ( \1306 , \1304 , \1305 );
xnor \U$930 ( \1307 , \1306 , \711 );
and \U$931 ( \1308 , \1303 , \1307 );
and \U$932 ( \1309 , \666 , \641 );
and \U$933 ( \1310 , \615 , \639 );
nor \U$934 ( \1311 , \1309 , \1310 );
xnor \U$935 ( \1312 , \1311 , \592 );
and \U$936 ( \1313 , \1307 , \1312 );
and \U$937 ( \1314 , \1303 , \1312 );
or \U$938 ( \1315 , \1308 , \1313 , \1314 );
and \U$939 ( \1316 , \1299 , \1315 );
and \U$940 ( \1317 , \771 , \540 );
and \U$941 ( \1318 , \743 , \538 );
nor \U$942 ( \1319 , \1317 , \1318 );
xnor \U$943 ( \1320 , \1319 , \499 );
and \U$944 ( \1321 , \925 , \470 );
and \U$945 ( \1322 , \851 , \468 );
nor \U$946 ( \1323 , \1321 , \1322 );
xnor \U$947 ( \1324 , \1323 , \440 );
and \U$948 ( \1325 , \1320 , \1324 );
and \U$949 ( \1326 , \1050 , \422 );
and \U$950 ( \1327 , \987 , \420 );
nor \U$951 ( \1328 , \1326 , \1327 );
xnor \U$952 ( \1329 , \1328 , \403 );
and \U$953 ( \1330 , \1324 , \1329 );
and \U$954 ( \1331 , \1320 , \1329 );
or \U$955 ( \1332 , \1325 , \1330 , \1331 );
and \U$956 ( \1333 , \1315 , \1332 );
and \U$957 ( \1334 , \1299 , \1332 );
or \U$958 ( \1335 , \1316 , \1333 , \1334 );
buf \U$959 ( \1336 , RIc224fb8_82);
and \U$960 ( \1337 , \1336 , \379 );
xor \U$961 ( \1338 , \1242 , \1246 );
xor \U$962 ( \1339 , \1338 , \1252 );
or \U$963 ( \1340 , \1337 , \1339 );
and \U$964 ( \1341 , \1335 , \1340 );
xor \U$965 ( \1342 , \1206 , \1210 );
xor \U$966 ( \1343 , \1342 , \1215 );
xor \U$967 ( \1344 , \1225 , \1229 );
xor \U$968 ( \1345 , \1344 , \1234 );
and \U$969 ( \1346 , \1343 , \1345 );
and \U$970 ( \1347 , \1340 , \1346 );
and \U$971 ( \1348 , \1335 , \1346 );
or \U$972 ( \1349 , \1341 , \1347 , \1348 );
xor \U$973 ( \1350 , \1145 , \1149 );
xor \U$974 ( \1351 , \1350 , \1154 );
xor \U$975 ( \1352 , \1218 , \1237 );
xor \U$976 ( \1353 , \1352 , \1255 );
and \U$977 ( \1354 , \1351 , \1353 );
xor \U$978 ( \1355 , \1259 , \1261 );
xor \U$979 ( \1356 , \1355 , \1264 );
and \U$980 ( \1357 , \1353 , \1356 );
and \U$981 ( \1358 , \1351 , \1356 );
or \U$982 ( \1359 , \1354 , \1357 , \1358 );
and \U$983 ( \1360 , \1349 , \1359 );
xnor \U$984 ( \1361 , \1179 , \1181 );
and \U$985 ( \1362 , \1359 , \1361 );
and \U$986 ( \1363 , \1349 , \1361 );
or \U$987 ( \1364 , \1360 , \1362 , \1363 );
xor \U$988 ( \1365 , \1139 , \1157 );
xor \U$989 ( \1366 , \1365 , \1174 );
xor \U$990 ( \1367 , \1258 , \1267 );
xor \U$991 ( \1368 , \1367 , \1270 );
and \U$992 ( \1369 , \1366 , \1368 );
and \U$993 ( \1370 , \1364 , \1369 );
xor \U$994 ( \1371 , \1273 , \1275 );
xor \U$995 ( \1372 , \1371 , \1278 );
and \U$996 ( \1373 , \1369 , \1372 );
and \U$997 ( \1374 , \1364 , \1372 );
or \U$998 ( \1375 , \1370 , \1373 , \1374 );
and \U$999 ( \1376 , \1281 , \1375 );
xor \U$1000 ( \1377 , \1188 , \1190 );
xor \U$1001 ( \1378 , \1377 , \1193 );
and \U$1002 ( \1379 , \1375 , \1378 );
and \U$1003 ( \1380 , \1281 , \1378 );
or \U$1004 ( \1381 , \1376 , \1379 , \1380 );
and \U$1005 ( \1382 , \1202 , \1381 );
xor \U$1006 ( \1383 , \1202 , \1381 );
xor \U$1007 ( \1384 , \1281 , \1375 );
xor \U$1008 ( \1385 , \1384 , \1378 );
and \U$1009 ( \1386 , \851 , \540 );
and \U$1010 ( \1387 , \771 , \538 );
nor \U$1011 ( \1388 , \1386 , \1387 );
xnor \U$1012 ( \1389 , \1388 , \499 );
and \U$1013 ( \1390 , \987 , \470 );
and \U$1014 ( \1391 , \925 , \468 );
nor \U$1015 ( \1392 , \1390 , \1391 );
xnor \U$1016 ( \1393 , \1392 , \440 );
and \U$1017 ( \1394 , \1389 , \1393 );
and \U$1018 ( \1395 , \1248 , \422 );
and \U$1019 ( \1396 , \1050 , \420 );
nor \U$1020 ( \1397 , \1395 , \1396 );
xnor \U$1021 ( \1398 , \1397 , \403 );
and \U$1022 ( \1399 , \1393 , \1398 );
and \U$1023 ( \1400 , \1389 , \1398 );
or \U$1024 ( \1401 , \1394 , \1399 , \1400 );
and \U$1025 ( \1402 , \556 , \888 );
and \U$1026 ( \1403 , \487 , \886 );
nor \U$1027 ( \1404 , \1402 , \1403 );
xnor \U$1028 ( \1405 , \1404 , \816 );
and \U$1029 ( \1406 , \615 , \754 );
and \U$1030 ( \1407 , \561 , \752 );
nor \U$1031 ( \1408 , \1406 , \1407 );
xnor \U$1032 ( \1409 , \1408 , \711 );
and \U$1033 ( \1410 , \1405 , \1409 );
and \U$1034 ( \1411 , \743 , \641 );
and \U$1035 ( \1412 , \666 , \639 );
nor \U$1036 ( \1413 , \1411 , \1412 );
xnor \U$1037 ( \1414 , \1413 , \592 );
and \U$1038 ( \1415 , \1409 , \1414 );
and \U$1039 ( \1416 , \1405 , \1414 );
or \U$1040 ( \1417 , \1410 , \1415 , \1416 );
and \U$1041 ( \1418 , \1401 , \1417 );
xor \U$1042 ( \1419 , \1141 , \1282 );
xor \U$1043 ( \1420 , \1282 , \1283 );
not \U$1044 ( \1421 , \1420 );
and \U$1045 ( \1422 , \1419 , \1421 );
and \U$1046 ( \1423 , \378 , \1422 );
not \U$1047 ( \1424 , \1423 );
xnor \U$1048 ( \1425 , \1424 , \1286 );
and \U$1049 ( \1426 , \410 , \1222 );
and \U$1050 ( \1427 , \392 , \1220 );
nor \U$1051 ( \1428 , \1426 , \1427 );
xnor \U$1052 ( \1429 , \1428 , \1144 );
and \U$1053 ( \1430 , \1425 , \1429 );
and \U$1054 ( \1431 , \479 , \1058 );
and \U$1055 ( \1432 , \431 , \1056 );
nor \U$1056 ( \1433 , \1431 , \1432 );
xnor \U$1057 ( \1434 , \1433 , \964 );
and \U$1058 ( \1435 , \1429 , \1434 );
and \U$1059 ( \1436 , \1425 , \1434 );
or \U$1060 ( \1437 , \1430 , \1435 , \1436 );
and \U$1061 ( \1438 , \1417 , \1437 );
and \U$1062 ( \1439 , \1401 , \1437 );
or \U$1063 ( \1440 , \1418 , \1438 , \1439 );
buf \U$1064 ( \1441 , RIc224f40_83);
and \U$1065 ( \1442 , \1441 , \385 );
and \U$1066 ( \1443 , \1336 , \383 );
nor \U$1067 ( \1444 , \1442 , \1443 );
xnor \U$1068 ( \1445 , \1444 , \390 );
buf \U$1069 ( \1446 , RIc224ec8_84);
and \U$1070 ( \1447 , \1446 , \379 );
or \U$1071 ( \1448 , \1445 , \1447 );
and \U$1072 ( \1449 , \1336 , \385 );
and \U$1073 ( \1450 , \1248 , \383 );
nor \U$1074 ( \1451 , \1449 , \1450 );
xnor \U$1075 ( \1452 , \1451 , \390 );
and \U$1076 ( \1453 , \1448 , \1452 );
and \U$1077 ( \1454 , \1441 , \379 );
and \U$1078 ( \1455 , \1452 , \1454 );
and \U$1079 ( \1456 , \1448 , \1454 );
or \U$1080 ( \1457 , \1453 , \1455 , \1456 );
and \U$1081 ( \1458 , \1440 , \1457 );
xor \U$1082 ( \1459 , \1287 , \1291 );
xor \U$1083 ( \1460 , \1459 , \1296 );
xor \U$1084 ( \1461 , \1303 , \1307 );
xor \U$1085 ( \1462 , \1461 , \1312 );
and \U$1086 ( \1463 , \1460 , \1462 );
xor \U$1087 ( \1464 , \1320 , \1324 );
xor \U$1088 ( \1465 , \1464 , \1329 );
and \U$1089 ( \1466 , \1462 , \1465 );
and \U$1090 ( \1467 , \1460 , \1465 );
or \U$1091 ( \1468 , \1463 , \1466 , \1467 );
and \U$1092 ( \1469 , \1457 , \1468 );
and \U$1093 ( \1470 , \1440 , \1468 );
or \U$1094 ( \1471 , \1458 , \1469 , \1470 );
xor \U$1095 ( \1472 , \1299 , \1315 );
xor \U$1096 ( \1473 , \1472 , \1332 );
xnor \U$1097 ( \1474 , \1337 , \1339 );
and \U$1098 ( \1475 , \1473 , \1474 );
xor \U$1099 ( \1476 , \1343 , \1345 );
and \U$1100 ( \1477 , \1474 , \1476 );
and \U$1101 ( \1478 , \1473 , \1476 );
or \U$1102 ( \1479 , \1475 , \1477 , \1478 );
and \U$1103 ( \1480 , \1471 , \1479 );
xor \U$1104 ( \1481 , \1351 , \1353 );
xor \U$1105 ( \1482 , \1481 , \1356 );
and \U$1106 ( \1483 , \1479 , \1482 );
and \U$1107 ( \1484 , \1471 , \1482 );
or \U$1108 ( \1485 , \1480 , \1483 , \1484 );
xor \U$1109 ( \1486 , \1349 , \1359 );
xor \U$1110 ( \1487 , \1486 , \1361 );
and \U$1111 ( \1488 , \1485 , \1487 );
xor \U$1112 ( \1489 , \1366 , \1368 );
and \U$1113 ( \1490 , \1487 , \1489 );
and \U$1114 ( \1491 , \1485 , \1489 );
or \U$1115 ( \1492 , \1488 , \1490 , \1491 );
xor \U$1116 ( \1493 , \1364 , \1369 );
xor \U$1117 ( \1494 , \1493 , \1372 );
and \U$1118 ( \1495 , \1492 , \1494 );
and \U$1119 ( \1496 , \1385 , \1495 );
xor \U$1120 ( \1497 , \1385 , \1495 );
xor \U$1121 ( \1498 , \1492 , \1494 );
buf \U$1122 ( \1499 , RIc226bd8_22);
buf \U$1123 ( \1500 , RIc226b60_23);
and \U$1124 ( \1501 , \1499 , \1500 );
not \U$1125 ( \1502 , \1501 );
and \U$1126 ( \1503 , \1283 , \1502 );
not \U$1127 ( \1504 , \1503 );
and \U$1128 ( \1505 , \392 , \1422 );
and \U$1129 ( \1506 , \378 , \1420 );
nor \U$1130 ( \1507 , \1505 , \1506 );
xnor \U$1131 ( \1508 , \1507 , \1286 );
and \U$1132 ( \1509 , \1504 , \1508 );
and \U$1133 ( \1510 , \431 , \1222 );
and \U$1134 ( \1511 , \410 , \1220 );
nor \U$1135 ( \1512 , \1510 , \1511 );
xnor \U$1136 ( \1513 , \1512 , \1144 );
and \U$1137 ( \1514 , \1508 , \1513 );
and \U$1138 ( \1515 , \1504 , \1513 );
or \U$1139 ( \1516 , \1509 , \1514 , \1515 );
and \U$1140 ( \1517 , \771 , \641 );
and \U$1141 ( \1518 , \743 , \639 );
nor \U$1142 ( \1519 , \1517 , \1518 );
xnor \U$1143 ( \1520 , \1519 , \592 );
and \U$1144 ( \1521 , \925 , \540 );
and \U$1145 ( \1522 , \851 , \538 );
nor \U$1146 ( \1523 , \1521 , \1522 );
xnor \U$1147 ( \1524 , \1523 , \499 );
and \U$1148 ( \1525 , \1520 , \1524 );
and \U$1149 ( \1526 , \1050 , \470 );
and \U$1150 ( \1527 , \987 , \468 );
nor \U$1151 ( \1528 , \1526 , \1527 );
xnor \U$1152 ( \1529 , \1528 , \440 );
and \U$1153 ( \1530 , \1524 , \1529 );
and \U$1154 ( \1531 , \1520 , \1529 );
or \U$1155 ( \1532 , \1525 , \1530 , \1531 );
and \U$1156 ( \1533 , \1516 , \1532 );
and \U$1157 ( \1534 , \487 , \1058 );
and \U$1158 ( \1535 , \479 , \1056 );
nor \U$1159 ( \1536 , \1534 , \1535 );
xnor \U$1160 ( \1537 , \1536 , \964 );
and \U$1161 ( \1538 , \561 , \888 );
and \U$1162 ( \1539 , \556 , \886 );
nor \U$1163 ( \1540 , \1538 , \1539 );
xnor \U$1164 ( \1541 , \1540 , \816 );
and \U$1165 ( \1542 , \1537 , \1541 );
and \U$1166 ( \1543 , \666 , \754 );
and \U$1167 ( \1544 , \615 , \752 );
nor \U$1168 ( \1545 , \1543 , \1544 );
xnor \U$1169 ( \1546 , \1545 , \711 );
and \U$1170 ( \1547 , \1541 , \1546 );
and \U$1171 ( \1548 , \1537 , \1546 );
or \U$1172 ( \1549 , \1542 , \1547 , \1548 );
and \U$1173 ( \1550 , \1532 , \1549 );
and \U$1174 ( \1551 , \1516 , \1549 );
or \U$1175 ( \1552 , \1533 , \1550 , \1551 );
and \U$1176 ( \1553 , \1336 , \422 );
and \U$1177 ( \1554 , \1248 , \420 );
nor \U$1178 ( \1555 , \1553 , \1554 );
xnor \U$1179 ( \1556 , \1555 , \403 );
and \U$1180 ( \1557 , \1446 , \385 );
and \U$1181 ( \1558 , \1441 , \383 );
nor \U$1182 ( \1559 , \1557 , \1558 );
xnor \U$1183 ( \1560 , \1559 , \390 );
and \U$1184 ( \1561 , \1556 , \1560 );
buf \U$1185 ( \1562 , RIc224e50_85);
and \U$1186 ( \1563 , \1562 , \379 );
and \U$1187 ( \1564 , \1560 , \1563 );
and \U$1188 ( \1565 , \1556 , \1563 );
or \U$1189 ( \1566 , \1561 , \1564 , \1565 );
xor \U$1190 ( \1567 , \1389 , \1393 );
xor \U$1191 ( \1568 , \1567 , \1398 );
and \U$1192 ( \1569 , \1566 , \1568 );
xnor \U$1193 ( \1570 , \1445 , \1447 );
and \U$1194 ( \1571 , \1568 , \1570 );
and \U$1195 ( \1572 , \1566 , \1570 );
or \U$1196 ( \1573 , \1569 , \1571 , \1572 );
and \U$1197 ( \1574 , \1552 , \1573 );
xor \U$1198 ( \1575 , \1405 , \1409 );
xor \U$1199 ( \1576 , \1575 , \1414 );
xor \U$1200 ( \1577 , \1425 , \1429 );
xor \U$1201 ( \1578 , \1577 , \1434 );
and \U$1202 ( \1579 , \1576 , \1578 );
and \U$1203 ( \1580 , \1573 , \1579 );
and \U$1204 ( \1581 , \1552 , \1579 );
or \U$1205 ( \1582 , \1574 , \1580 , \1581 );
xor \U$1206 ( \1583 , \1401 , \1417 );
xor \U$1207 ( \1584 , \1583 , \1437 );
xor \U$1208 ( \1585 , \1448 , \1452 );
xor \U$1209 ( \1586 , \1585 , \1454 );
and \U$1210 ( \1587 , \1584 , \1586 );
xor \U$1211 ( \1588 , \1460 , \1462 );
xor \U$1212 ( \1589 , \1588 , \1465 );
and \U$1213 ( \1590 , \1586 , \1589 );
and \U$1214 ( \1591 , \1584 , \1589 );
or \U$1215 ( \1592 , \1587 , \1590 , \1591 );
and \U$1216 ( \1593 , \1582 , \1592 );
xor \U$1217 ( \1594 , \1473 , \1474 );
xor \U$1218 ( \1595 , \1594 , \1476 );
and \U$1219 ( \1596 , \1592 , \1595 );
and \U$1220 ( \1597 , \1582 , \1595 );
or \U$1221 ( \1598 , \1593 , \1596 , \1597 );
xor \U$1222 ( \1599 , \1335 , \1340 );
xor \U$1223 ( \1600 , \1599 , \1346 );
and \U$1224 ( \1601 , \1598 , \1600 );
xor \U$1225 ( \1602 , \1471 , \1479 );
xor \U$1226 ( \1603 , \1602 , \1482 );
and \U$1227 ( \1604 , \1600 , \1603 );
and \U$1228 ( \1605 , \1598 , \1603 );
or \U$1229 ( \1606 , \1601 , \1604 , \1605 );
xor \U$1230 ( \1607 , \1485 , \1487 );
xor \U$1231 ( \1608 , \1607 , \1489 );
and \U$1232 ( \1609 , \1606 , \1608 );
and \U$1233 ( \1610 , \1498 , \1609 );
xor \U$1234 ( \1611 , \1498 , \1609 );
xor \U$1235 ( \1612 , \1606 , \1608 );
xor \U$1236 ( \1613 , \1283 , \1499 );
xor \U$1237 ( \1614 , \1499 , \1500 );
not \U$1238 ( \1615 , \1614 );
and \U$1239 ( \1616 , \1613 , \1615 );
and \U$1240 ( \1617 , \378 , \1616 );
not \U$1241 ( \1618 , \1617 );
xnor \U$1242 ( \1619 , \1618 , \1503 );
and \U$1243 ( \1620 , \410 , \1422 );
and \U$1244 ( \1621 , \392 , \1420 );
nor \U$1245 ( \1622 , \1620 , \1621 );
xnor \U$1246 ( \1623 , \1622 , \1286 );
and \U$1247 ( \1624 , \1619 , \1623 );
and \U$1248 ( \1625 , \479 , \1222 );
and \U$1249 ( \1626 , \431 , \1220 );
nor \U$1250 ( \1627 , \1625 , \1626 );
xnor \U$1251 ( \1628 , \1627 , \1144 );
and \U$1252 ( \1629 , \1623 , \1628 );
and \U$1253 ( \1630 , \1619 , \1628 );
or \U$1254 ( \1631 , \1624 , \1629 , \1630 );
and \U$1255 ( \1632 , \851 , \641 );
and \U$1256 ( \1633 , \771 , \639 );
nor \U$1257 ( \1634 , \1632 , \1633 );
xnor \U$1258 ( \1635 , \1634 , \592 );
and \U$1259 ( \1636 , \987 , \540 );
and \U$1260 ( \1637 , \925 , \538 );
nor \U$1261 ( \1638 , \1636 , \1637 );
xnor \U$1262 ( \1639 , \1638 , \499 );
and \U$1263 ( \1640 , \1635 , \1639 );
and \U$1264 ( \1641 , \1248 , \470 );
and \U$1265 ( \1642 , \1050 , \468 );
nor \U$1266 ( \1643 , \1641 , \1642 );
xnor \U$1267 ( \1644 , \1643 , \440 );
and \U$1268 ( \1645 , \1639 , \1644 );
and \U$1269 ( \1646 , \1635 , \1644 );
or \U$1270 ( \1647 , \1640 , \1645 , \1646 );
and \U$1271 ( \1648 , \1631 , \1647 );
and \U$1272 ( \1649 , \556 , \1058 );
and \U$1273 ( \1650 , \487 , \1056 );
nor \U$1274 ( \1651 , \1649 , \1650 );
xnor \U$1275 ( \1652 , \1651 , \964 );
and \U$1276 ( \1653 , \615 , \888 );
and \U$1277 ( \1654 , \561 , \886 );
nor \U$1278 ( \1655 , \1653 , \1654 );
xnor \U$1279 ( \1656 , \1655 , \816 );
and \U$1280 ( \1657 , \1652 , \1656 );
and \U$1281 ( \1658 , \743 , \754 );
and \U$1282 ( \1659 , \666 , \752 );
nor \U$1283 ( \1660 , \1658 , \1659 );
xnor \U$1284 ( \1661 , \1660 , \711 );
and \U$1285 ( \1662 , \1656 , \1661 );
and \U$1286 ( \1663 , \1652 , \1661 );
or \U$1287 ( \1664 , \1657 , \1662 , \1663 );
and \U$1288 ( \1665 , \1647 , \1664 );
and \U$1289 ( \1666 , \1631 , \1664 );
or \U$1290 ( \1667 , \1648 , \1665 , \1666 );
and \U$1291 ( \1668 , \1441 , \422 );
and \U$1292 ( \1669 , \1336 , \420 );
nor \U$1293 ( \1670 , \1668 , \1669 );
xnor \U$1294 ( \1671 , \1670 , \403 );
and \U$1295 ( \1672 , \1562 , \385 );
and \U$1296 ( \1673 , \1446 , \383 );
nor \U$1297 ( \1674 , \1672 , \1673 );
xnor \U$1298 ( \1675 , \1674 , \390 );
and \U$1299 ( \1676 , \1671 , \1675 );
buf \U$1300 ( \1677 , RIc224dd8_86);
and \U$1301 ( \1678 , \1677 , \379 );
and \U$1302 ( \1679 , \1675 , \1678 );
and \U$1303 ( \1680 , \1671 , \1678 );
or \U$1304 ( \1681 , \1676 , \1679 , \1680 );
xor \U$1305 ( \1682 , \1556 , \1560 );
xor \U$1306 ( \1683 , \1682 , \1563 );
and \U$1307 ( \1684 , \1681 , \1683 );
xor \U$1308 ( \1685 , \1520 , \1524 );
xor \U$1309 ( \1686 , \1685 , \1529 );
and \U$1310 ( \1687 , \1683 , \1686 );
and \U$1311 ( \1688 , \1681 , \1686 );
or \U$1312 ( \1689 , \1684 , \1687 , \1688 );
and \U$1313 ( \1690 , \1667 , \1689 );
xor \U$1314 ( \1691 , \1504 , \1508 );
xor \U$1315 ( \1692 , \1691 , \1513 );
xor \U$1316 ( \1693 , \1537 , \1541 );
xor \U$1317 ( \1694 , \1693 , \1546 );
and \U$1318 ( \1695 , \1692 , \1694 );
and \U$1319 ( \1696 , \1689 , \1695 );
and \U$1320 ( \1697 , \1667 , \1695 );
or \U$1321 ( \1698 , \1690 , \1696 , \1697 );
xor \U$1322 ( \1699 , \1516 , \1532 );
xor \U$1323 ( \1700 , \1699 , \1549 );
xor \U$1324 ( \1701 , \1566 , \1568 );
xor \U$1325 ( \1702 , \1701 , \1570 );
and \U$1326 ( \1703 , \1700 , \1702 );
xor \U$1327 ( \1704 , \1576 , \1578 );
and \U$1328 ( \1705 , \1702 , \1704 );
and \U$1329 ( \1706 , \1700 , \1704 );
or \U$1330 ( \1707 , \1703 , \1705 , \1706 );
and \U$1331 ( \1708 , \1698 , \1707 );
xor \U$1332 ( \1709 , \1584 , \1586 );
xor \U$1333 ( \1710 , \1709 , \1589 );
and \U$1334 ( \1711 , \1707 , \1710 );
and \U$1335 ( \1712 , \1698 , \1710 );
or \U$1336 ( \1713 , \1708 , \1711 , \1712 );
xor \U$1337 ( \1714 , \1440 , \1457 );
xor \U$1338 ( \1715 , \1714 , \1468 );
and \U$1339 ( \1716 , \1713 , \1715 );
xor \U$1340 ( \1717 , \1582 , \1592 );
xor \U$1341 ( \1718 , \1717 , \1595 );
and \U$1342 ( \1719 , \1715 , \1718 );
and \U$1343 ( \1720 , \1713 , \1718 );
or \U$1344 ( \1721 , \1716 , \1719 , \1720 );
xor \U$1345 ( \1722 , \1598 , \1600 );
xor \U$1346 ( \1723 , \1722 , \1603 );
and \U$1347 ( \1724 , \1721 , \1723 );
and \U$1348 ( \1725 , \1612 , \1724 );
xor \U$1349 ( \1726 , \1612 , \1724 );
xor \U$1350 ( \1727 , \1721 , \1723 );
buf \U$1351 ( \1728 , RIc226ae8_24);
buf \U$1352 ( \1729 , RIc226a70_25);
and \U$1353 ( \1730 , \1728 , \1729 );
not \U$1354 ( \1731 , \1730 );
and \U$1355 ( \1732 , \1500 , \1731 );
not \U$1356 ( \1733 , \1732 );
and \U$1357 ( \1734 , \392 , \1616 );
and \U$1358 ( \1735 , \378 , \1614 );
nor \U$1359 ( \1736 , \1734 , \1735 );
xnor \U$1360 ( \1737 , \1736 , \1503 );
and \U$1361 ( \1738 , \1733 , \1737 );
and \U$1362 ( \1739 , \431 , \1422 );
and \U$1363 ( \1740 , \410 , \1420 );
nor \U$1364 ( \1741 , \1739 , \1740 );
xnor \U$1365 ( \1742 , \1741 , \1286 );
and \U$1366 ( \1743 , \1737 , \1742 );
and \U$1367 ( \1744 , \1733 , \1742 );
or \U$1368 ( \1745 , \1738 , \1743 , \1744 );
and \U$1369 ( \1746 , \487 , \1222 );
and \U$1370 ( \1747 , \479 , \1220 );
nor \U$1371 ( \1748 , \1746 , \1747 );
xnor \U$1372 ( \1749 , \1748 , \1144 );
and \U$1373 ( \1750 , \561 , \1058 );
and \U$1374 ( \1751 , \556 , \1056 );
nor \U$1375 ( \1752 , \1750 , \1751 );
xnor \U$1376 ( \1753 , \1752 , \964 );
and \U$1377 ( \1754 , \1749 , \1753 );
and \U$1378 ( \1755 , \666 , \888 );
and \U$1379 ( \1756 , \615 , \886 );
nor \U$1380 ( \1757 , \1755 , \1756 );
xnor \U$1381 ( \1758 , \1757 , \816 );
and \U$1382 ( \1759 , \1753 , \1758 );
and \U$1383 ( \1760 , \1749 , \1758 );
or \U$1384 ( \1761 , \1754 , \1759 , \1760 );
and \U$1385 ( \1762 , \1745 , \1761 );
and \U$1386 ( \1763 , \771 , \754 );
and \U$1387 ( \1764 , \743 , \752 );
nor \U$1388 ( \1765 , \1763 , \1764 );
xnor \U$1389 ( \1766 , \1765 , \711 );
and \U$1390 ( \1767 , \925 , \641 );
and \U$1391 ( \1768 , \851 , \639 );
nor \U$1392 ( \1769 , \1767 , \1768 );
xnor \U$1393 ( \1770 , \1769 , \592 );
and \U$1394 ( \1771 , \1766 , \1770 );
and \U$1395 ( \1772 , \1050 , \540 );
and \U$1396 ( \1773 , \987 , \538 );
nor \U$1397 ( \1774 , \1772 , \1773 );
xnor \U$1398 ( \1775 , \1774 , \499 );
and \U$1399 ( \1776 , \1770 , \1775 );
and \U$1400 ( \1777 , \1766 , \1775 );
or \U$1401 ( \1778 , \1771 , \1776 , \1777 );
and \U$1402 ( \1779 , \1761 , \1778 );
and \U$1403 ( \1780 , \1745 , \1778 );
or \U$1404 ( \1781 , \1762 , \1779 , \1780 );
xor \U$1405 ( \1782 , \1619 , \1623 );
xor \U$1406 ( \1783 , \1782 , \1628 );
xor \U$1407 ( \1784 , \1635 , \1639 );
xor \U$1408 ( \1785 , \1784 , \1644 );
and \U$1409 ( \1786 , \1783 , \1785 );
xor \U$1410 ( \1787 , \1652 , \1656 );
xor \U$1411 ( \1788 , \1787 , \1661 );
and \U$1412 ( \1789 , \1785 , \1788 );
and \U$1413 ( \1790 , \1783 , \1788 );
or \U$1414 ( \1791 , \1786 , \1789 , \1790 );
and \U$1415 ( \1792 , \1781 , \1791 );
and \U$1416 ( \1793 , \1336 , \470 );
and \U$1417 ( \1794 , \1248 , \468 );
nor \U$1418 ( \1795 , \1793 , \1794 );
xnor \U$1419 ( \1796 , \1795 , \440 );
and \U$1420 ( \1797 , \1446 , \422 );
and \U$1421 ( \1798 , \1441 , \420 );
nor \U$1422 ( \1799 , \1797 , \1798 );
xnor \U$1423 ( \1800 , \1799 , \403 );
and \U$1424 ( \1801 , \1796 , \1800 );
and \U$1425 ( \1802 , \1677 , \385 );
and \U$1426 ( \1803 , \1562 , \383 );
nor \U$1427 ( \1804 , \1802 , \1803 );
xnor \U$1428 ( \1805 , \1804 , \390 );
and \U$1429 ( \1806 , \1800 , \1805 );
and \U$1430 ( \1807 , \1796 , \1805 );
or \U$1431 ( \1808 , \1801 , \1806 , \1807 );
xor \U$1432 ( \1809 , \1671 , \1675 );
xor \U$1433 ( \1810 , \1809 , \1678 );
or \U$1434 ( \1811 , \1808 , \1810 );
and \U$1435 ( \1812 , \1791 , \1811 );
and \U$1436 ( \1813 , \1781 , \1811 );
or \U$1437 ( \1814 , \1792 , \1812 , \1813 );
xor \U$1438 ( \1815 , \1631 , \1647 );
xor \U$1439 ( \1816 , \1815 , \1664 );
xor \U$1440 ( \1817 , \1681 , \1683 );
xor \U$1441 ( \1818 , \1817 , \1686 );
and \U$1442 ( \1819 , \1816 , \1818 );
xor \U$1443 ( \1820 , \1692 , \1694 );
and \U$1444 ( \1821 , \1818 , \1820 );
and \U$1445 ( \1822 , \1816 , \1820 );
or \U$1446 ( \1823 , \1819 , \1821 , \1822 );
and \U$1447 ( \1824 , \1814 , \1823 );
xor \U$1448 ( \1825 , \1700 , \1702 );
xor \U$1449 ( \1826 , \1825 , \1704 );
and \U$1450 ( \1827 , \1823 , \1826 );
and \U$1451 ( \1828 , \1814 , \1826 );
or \U$1452 ( \1829 , \1824 , \1827 , \1828 );
xor \U$1453 ( \1830 , \1552 , \1573 );
xor \U$1454 ( \1831 , \1830 , \1579 );
and \U$1455 ( \1832 , \1829 , \1831 );
xor \U$1456 ( \1833 , \1698 , \1707 );
xor \U$1457 ( \1834 , \1833 , \1710 );
and \U$1458 ( \1835 , \1831 , \1834 );
and \U$1459 ( \1836 , \1829 , \1834 );
or \U$1460 ( \1837 , \1832 , \1835 , \1836 );
xor \U$1461 ( \1838 , \1713 , \1715 );
xor \U$1462 ( \1839 , \1838 , \1718 );
and \U$1463 ( \1840 , \1837 , \1839 );
and \U$1464 ( \1841 , \1727 , \1840 );
xor \U$1465 ( \1842 , \1727 , \1840 );
xor \U$1466 ( \1843 , \1837 , \1839 );
and \U$1467 ( \1844 , \1441 , \470 );
and \U$1468 ( \1845 , \1336 , \468 );
nor \U$1469 ( \1846 , \1844 , \1845 );
xnor \U$1470 ( \1847 , \1846 , \440 );
and \U$1471 ( \1848 , \1562 , \422 );
and \U$1472 ( \1849 , \1446 , \420 );
nor \U$1473 ( \1850 , \1848 , \1849 );
xnor \U$1474 ( \1851 , \1850 , \403 );
and \U$1475 ( \1852 , \1847 , \1851 );
buf \U$1476 ( \1853 , RIc224d60_87);
and \U$1477 ( \1854 , \1853 , \385 );
and \U$1478 ( \1855 , \1677 , \383 );
nor \U$1479 ( \1856 , \1854 , \1855 );
xnor \U$1480 ( \1857 , \1856 , \390 );
and \U$1481 ( \1858 , \1851 , \1857 );
and \U$1482 ( \1859 , \1847 , \1857 );
or \U$1483 ( \1860 , \1852 , \1858 , \1859 );
buf \U$1484 ( \1861 , RIc224ce8_88);
and \U$1485 ( \1862 , \1861 , \379 );
buf \U$1486 ( \1863 , \1862 );
and \U$1487 ( \1864 , \1860 , \1863 );
and \U$1488 ( \1865 , \1853 , \379 );
and \U$1489 ( \1866 , \1863 , \1865 );
and \U$1490 ( \1867 , \1860 , \1865 );
or \U$1491 ( \1868 , \1864 , \1866 , \1867 );
and \U$1492 ( \1869 , \556 , \1222 );
and \U$1493 ( \1870 , \487 , \1220 );
nor \U$1494 ( \1871 , \1869 , \1870 );
xnor \U$1495 ( \1872 , \1871 , \1144 );
and \U$1496 ( \1873 , \615 , \1058 );
and \U$1497 ( \1874 , \561 , \1056 );
nor \U$1498 ( \1875 , \1873 , \1874 );
xnor \U$1499 ( \1876 , \1875 , \964 );
and \U$1500 ( \1877 , \1872 , \1876 );
and \U$1501 ( \1878 , \743 , \888 );
and \U$1502 ( \1879 , \666 , \886 );
nor \U$1503 ( \1880 , \1878 , \1879 );
xnor \U$1504 ( \1881 , \1880 , \816 );
and \U$1505 ( \1882 , \1876 , \1881 );
and \U$1506 ( \1883 , \1872 , \1881 );
or \U$1507 ( \1884 , \1877 , \1882 , \1883 );
xor \U$1508 ( \1885 , \1500 , \1728 );
xor \U$1509 ( \1886 , \1728 , \1729 );
not \U$1510 ( \1887 , \1886 );
and \U$1511 ( \1888 , \1885 , \1887 );
and \U$1512 ( \1889 , \378 , \1888 );
not \U$1513 ( \1890 , \1889 );
xnor \U$1514 ( \1891 , \1890 , \1732 );
and \U$1515 ( \1892 , \410 , \1616 );
and \U$1516 ( \1893 , \392 , \1614 );
nor \U$1517 ( \1894 , \1892 , \1893 );
xnor \U$1518 ( \1895 , \1894 , \1503 );
and \U$1519 ( \1896 , \1891 , \1895 );
and \U$1520 ( \1897 , \479 , \1422 );
and \U$1521 ( \1898 , \431 , \1420 );
nor \U$1522 ( \1899 , \1897 , \1898 );
xnor \U$1523 ( \1900 , \1899 , \1286 );
and \U$1524 ( \1901 , \1895 , \1900 );
and \U$1525 ( \1902 , \1891 , \1900 );
or \U$1526 ( \1903 , \1896 , \1901 , \1902 );
and \U$1527 ( \1904 , \1884 , \1903 );
and \U$1528 ( \1905 , \851 , \754 );
and \U$1529 ( \1906 , \771 , \752 );
nor \U$1530 ( \1907 , \1905 , \1906 );
xnor \U$1531 ( \1908 , \1907 , \711 );
and \U$1532 ( \1909 , \987 , \641 );
and \U$1533 ( \1910 , \925 , \639 );
nor \U$1534 ( \1911 , \1909 , \1910 );
xnor \U$1535 ( \1912 , \1911 , \592 );
and \U$1536 ( \1913 , \1908 , \1912 );
and \U$1537 ( \1914 , \1248 , \540 );
and \U$1538 ( \1915 , \1050 , \538 );
nor \U$1539 ( \1916 , \1914 , \1915 );
xnor \U$1540 ( \1917 , \1916 , \499 );
and \U$1541 ( \1918 , \1912 , \1917 );
and \U$1542 ( \1919 , \1908 , \1917 );
or \U$1543 ( \1920 , \1913 , \1918 , \1919 );
and \U$1544 ( \1921 , \1903 , \1920 );
and \U$1545 ( \1922 , \1884 , \1920 );
or \U$1546 ( \1923 , \1904 , \1921 , \1922 );
and \U$1547 ( \1924 , \1868 , \1923 );
xor \U$1548 ( \1925 , \1749 , \1753 );
xor \U$1549 ( \1926 , \1925 , \1758 );
xor \U$1550 ( \1927 , \1796 , \1800 );
xor \U$1551 ( \1928 , \1927 , \1805 );
and \U$1552 ( \1929 , \1926 , \1928 );
xor \U$1553 ( \1930 , \1766 , \1770 );
xor \U$1554 ( \1931 , \1930 , \1775 );
and \U$1555 ( \1932 , \1928 , \1931 );
and \U$1556 ( \1933 , \1926 , \1931 );
or \U$1557 ( \1934 , \1929 , \1932 , \1933 );
and \U$1558 ( \1935 , \1923 , \1934 );
and \U$1559 ( \1936 , \1868 , \1934 );
or \U$1560 ( \1937 , \1924 , \1935 , \1936 );
xor \U$1561 ( \1938 , \1745 , \1761 );
xor \U$1562 ( \1939 , \1938 , \1778 );
xor \U$1563 ( \1940 , \1783 , \1785 );
xor \U$1564 ( \1941 , \1940 , \1788 );
and \U$1565 ( \1942 , \1939 , \1941 );
xnor \U$1566 ( \1943 , \1808 , \1810 );
and \U$1567 ( \1944 , \1941 , \1943 );
and \U$1568 ( \1945 , \1939 , \1943 );
or \U$1569 ( \1946 , \1942 , \1944 , \1945 );
and \U$1570 ( \1947 , \1937 , \1946 );
xor \U$1571 ( \1948 , \1816 , \1818 );
xor \U$1572 ( \1949 , \1948 , \1820 );
and \U$1573 ( \1950 , \1946 , \1949 );
and \U$1574 ( \1951 , \1937 , \1949 );
or \U$1575 ( \1952 , \1947 , \1950 , \1951 );
xor \U$1576 ( \1953 , \1667 , \1689 );
xor \U$1577 ( \1954 , \1953 , \1695 );
and \U$1578 ( \1955 , \1952 , \1954 );
xor \U$1579 ( \1956 , \1814 , \1823 );
xor \U$1580 ( \1957 , \1956 , \1826 );
and \U$1581 ( \1958 , \1954 , \1957 );
and \U$1582 ( \1959 , \1952 , \1957 );
or \U$1583 ( \1960 , \1955 , \1958 , \1959 );
xor \U$1584 ( \1961 , \1829 , \1831 );
xor \U$1585 ( \1962 , \1961 , \1834 );
and \U$1586 ( \1963 , \1960 , \1962 );
and \U$1587 ( \1964 , \1843 , \1963 );
xor \U$1588 ( \1965 , \1843 , \1963 );
xor \U$1589 ( \1966 , \1960 , \1962 );
and \U$1590 ( \1967 , \771 , \888 );
and \U$1591 ( \1968 , \743 , \886 );
nor \U$1592 ( \1969 , \1967 , \1968 );
xnor \U$1593 ( \1970 , \1969 , \816 );
and \U$1594 ( \1971 , \925 , \754 );
and \U$1595 ( \1972 , \851 , \752 );
nor \U$1596 ( \1973 , \1971 , \1972 );
xnor \U$1597 ( \1974 , \1973 , \711 );
and \U$1598 ( \1975 , \1970 , \1974 );
and \U$1599 ( \1976 , \1050 , \641 );
and \U$1600 ( \1977 , \987 , \639 );
nor \U$1601 ( \1978 , \1976 , \1977 );
xnor \U$1602 ( \1979 , \1978 , \592 );
and \U$1603 ( \1980 , \1974 , \1979 );
and \U$1604 ( \1981 , \1970 , \1979 );
or \U$1605 ( \1982 , \1975 , \1980 , \1981 );
and \U$1606 ( \1983 , \487 , \1422 );
and \U$1607 ( \1984 , \479 , \1420 );
nor \U$1608 ( \1985 , \1983 , \1984 );
xnor \U$1609 ( \1986 , \1985 , \1286 );
and \U$1610 ( \1987 , \561 , \1222 );
and \U$1611 ( \1988 , \556 , \1220 );
nor \U$1612 ( \1989 , \1987 , \1988 );
xnor \U$1613 ( \1990 , \1989 , \1144 );
and \U$1614 ( \1991 , \1986 , \1990 );
and \U$1615 ( \1992 , \666 , \1058 );
and \U$1616 ( \1993 , \615 , \1056 );
nor \U$1617 ( \1994 , \1992 , \1993 );
xnor \U$1618 ( \1995 , \1994 , \964 );
and \U$1619 ( \1996 , \1990 , \1995 );
and \U$1620 ( \1997 , \1986 , \1995 );
or \U$1621 ( \1998 , \1991 , \1996 , \1997 );
and \U$1622 ( \1999 , \1982 , \1998 );
buf \U$1623 ( \2000 , RIc2269f8_26);
buf \U$1624 ( \2001 , RIc226980_27);
and \U$1625 ( \2002 , \2000 , \2001 );
not \U$1626 ( \2003 , \2002 );
and \U$1627 ( \2004 , \1729 , \2003 );
not \U$1628 ( \2005 , \2004 );
and \U$1629 ( \2006 , \392 , \1888 );
and \U$1630 ( \2007 , \378 , \1886 );
nor \U$1631 ( \2008 , \2006 , \2007 );
xnor \U$1632 ( \2009 , \2008 , \1732 );
and \U$1633 ( \2010 , \2005 , \2009 );
and \U$1634 ( \2011 , \431 , \1616 );
and \U$1635 ( \2012 , \410 , \1614 );
nor \U$1636 ( \2013 , \2011 , \2012 );
xnor \U$1637 ( \2014 , \2013 , \1503 );
and \U$1638 ( \2015 , \2009 , \2014 );
and \U$1639 ( \2016 , \2005 , \2014 );
or \U$1640 ( \2017 , \2010 , \2015 , \2016 );
and \U$1641 ( \2018 , \1998 , \2017 );
and \U$1642 ( \2019 , \1982 , \2017 );
or \U$1643 ( \2020 , \1999 , \2018 , \2019 );
xor \U$1644 ( \2021 , \1872 , \1876 );
xor \U$1645 ( \2022 , \2021 , \1881 );
xor \U$1646 ( \2023 , \1891 , \1895 );
xor \U$1647 ( \2024 , \2023 , \1900 );
and \U$1648 ( \2025 , \2022 , \2024 );
xor \U$1649 ( \2026 , \1908 , \1912 );
xor \U$1650 ( \2027 , \2026 , \1917 );
and \U$1651 ( \2028 , \2024 , \2027 );
and \U$1652 ( \2029 , \2022 , \2027 );
or \U$1653 ( \2030 , \2025 , \2028 , \2029 );
and \U$1654 ( \2031 , \2020 , \2030 );
and \U$1655 ( \2032 , \1336 , \540 );
and \U$1656 ( \2033 , \1248 , \538 );
nor \U$1657 ( \2034 , \2032 , \2033 );
xnor \U$1658 ( \2035 , \2034 , \499 );
and \U$1659 ( \2036 , \1446 , \470 );
and \U$1660 ( \2037 , \1441 , \468 );
nor \U$1661 ( \2038 , \2036 , \2037 );
xnor \U$1662 ( \2039 , \2038 , \440 );
and \U$1663 ( \2040 , \2035 , \2039 );
and \U$1664 ( \2041 , \1677 , \422 );
and \U$1665 ( \2042 , \1562 , \420 );
nor \U$1666 ( \2043 , \2041 , \2042 );
xnor \U$1667 ( \2044 , \2043 , \403 );
and \U$1668 ( \2045 , \2039 , \2044 );
and \U$1669 ( \2046 , \2035 , \2044 );
or \U$1670 ( \2047 , \2040 , \2045 , \2046 );
xor \U$1671 ( \2048 , \1847 , \1851 );
xor \U$1672 ( \2049 , \2048 , \1857 );
and \U$1673 ( \2050 , \2047 , \2049 );
not \U$1674 ( \2051 , \1862 );
and \U$1675 ( \2052 , \2049 , \2051 );
and \U$1676 ( \2053 , \2047 , \2051 );
or \U$1677 ( \2054 , \2050 , \2052 , \2053 );
and \U$1678 ( \2055 , \2030 , \2054 );
and \U$1679 ( \2056 , \2020 , \2054 );
or \U$1680 ( \2057 , \2031 , \2055 , \2056 );
xor \U$1681 ( \2058 , \1733 , \1737 );
xor \U$1682 ( \2059 , \2058 , \1742 );
xor \U$1683 ( \2060 , \1860 , \1863 );
xor \U$1684 ( \2061 , \2060 , \1865 );
and \U$1685 ( \2062 , \2059 , \2061 );
xor \U$1686 ( \2063 , \1926 , \1928 );
xor \U$1687 ( \2064 , \2063 , \1931 );
and \U$1688 ( \2065 , \2061 , \2064 );
and \U$1689 ( \2066 , \2059 , \2064 );
or \U$1690 ( \2067 , \2062 , \2065 , \2066 );
and \U$1691 ( \2068 , \2057 , \2067 );
xor \U$1692 ( \2069 , \1939 , \1941 );
xor \U$1693 ( \2070 , \2069 , \1943 );
and \U$1694 ( \2071 , \2067 , \2070 );
and \U$1695 ( \2072 , \2057 , \2070 );
or \U$1696 ( \2073 , \2068 , \2071 , \2072 );
xor \U$1697 ( \2074 , \1781 , \1791 );
xor \U$1698 ( \2075 , \2074 , \1811 );
and \U$1699 ( \2076 , \2073 , \2075 );
xor \U$1700 ( \2077 , \1937 , \1946 );
xor \U$1701 ( \2078 , \2077 , \1949 );
and \U$1702 ( \2079 , \2075 , \2078 );
and \U$1703 ( \2080 , \2073 , \2078 );
or \U$1704 ( \2081 , \2076 , \2079 , \2080 );
xor \U$1705 ( \2082 , \1952 , \1954 );
xor \U$1706 ( \2083 , \2082 , \1957 );
and \U$1707 ( \2084 , \2081 , \2083 );
and \U$1708 ( \2085 , \1966 , \2084 );
xor \U$1709 ( \2086 , \1966 , \2084 );
xor \U$1710 ( \2087 , \2081 , \2083 );
and \U$1711 ( \2088 , \1441 , \540 );
and \U$1712 ( \2089 , \1336 , \538 );
nor \U$1713 ( \2090 , \2088 , \2089 );
xnor \U$1714 ( \2091 , \2090 , \499 );
and \U$1715 ( \2092 , \1562 , \470 );
and \U$1716 ( \2093 , \1446 , \468 );
nor \U$1717 ( \2094 , \2092 , \2093 );
xnor \U$1718 ( \2095 , \2094 , \440 );
and \U$1719 ( \2096 , \2091 , \2095 );
and \U$1720 ( \2097 , \1853 , \422 );
and \U$1721 ( \2098 , \1677 , \420 );
nor \U$1722 ( \2099 , \2097 , \2098 );
xnor \U$1723 ( \2100 , \2099 , \403 );
and \U$1724 ( \2101 , \2095 , \2100 );
and \U$1725 ( \2102 , \2091 , \2100 );
or \U$1726 ( \2103 , \2096 , \2101 , \2102 );
buf \U$1727 ( \2104 , RIc224c70_89);
and \U$1728 ( \2105 , \2104 , \385 );
and \U$1729 ( \2106 , \1861 , \383 );
nor \U$1730 ( \2107 , \2105 , \2106 );
xnor \U$1731 ( \2108 , \2107 , \390 );
buf \U$1732 ( \2109 , RIc224bf8_90);
and \U$1733 ( \2110 , \2109 , \379 );
or \U$1734 ( \2111 , \2108 , \2110 );
and \U$1735 ( \2112 , \2103 , \2111 );
and \U$1736 ( \2113 , \1861 , \385 );
and \U$1737 ( \2114 , \1853 , \383 );
nor \U$1738 ( \2115 , \2113 , \2114 );
xnor \U$1739 ( \2116 , \2115 , \390 );
and \U$1740 ( \2117 , \2111 , \2116 );
and \U$1741 ( \2118 , \2103 , \2116 );
or \U$1742 ( \2119 , \2112 , \2117 , \2118 );
and \U$1743 ( \2120 , \851 , \888 );
and \U$1744 ( \2121 , \771 , \886 );
nor \U$1745 ( \2122 , \2120 , \2121 );
xnor \U$1746 ( \2123 , \2122 , \816 );
and \U$1747 ( \2124 , \987 , \754 );
and \U$1748 ( \2125 , \925 , \752 );
nor \U$1749 ( \2126 , \2124 , \2125 );
xnor \U$1750 ( \2127 , \2126 , \711 );
and \U$1751 ( \2128 , \2123 , \2127 );
and \U$1752 ( \2129 , \1248 , \641 );
and \U$1753 ( \2130 , \1050 , \639 );
nor \U$1754 ( \2131 , \2129 , \2130 );
xnor \U$1755 ( \2132 , \2131 , \592 );
and \U$1756 ( \2133 , \2127 , \2132 );
and \U$1757 ( \2134 , \2123 , \2132 );
or \U$1758 ( \2135 , \2128 , \2133 , \2134 );
and \U$1759 ( \2136 , \556 , \1422 );
and \U$1760 ( \2137 , \487 , \1420 );
nor \U$1761 ( \2138 , \2136 , \2137 );
xnor \U$1762 ( \2139 , \2138 , \1286 );
and \U$1763 ( \2140 , \615 , \1222 );
and \U$1764 ( \2141 , \561 , \1220 );
nor \U$1765 ( \2142 , \2140 , \2141 );
xnor \U$1766 ( \2143 , \2142 , \1144 );
and \U$1767 ( \2144 , \2139 , \2143 );
and \U$1768 ( \2145 , \743 , \1058 );
and \U$1769 ( \2146 , \666 , \1056 );
nor \U$1770 ( \2147 , \2145 , \2146 );
xnor \U$1771 ( \2148 , \2147 , \964 );
and \U$1772 ( \2149 , \2143 , \2148 );
and \U$1773 ( \2150 , \2139 , \2148 );
or \U$1774 ( \2151 , \2144 , \2149 , \2150 );
and \U$1775 ( \2152 , \2135 , \2151 );
xor \U$1776 ( \2153 , \1729 , \2000 );
xor \U$1777 ( \2154 , \2000 , \2001 );
not \U$1778 ( \2155 , \2154 );
and \U$1779 ( \2156 , \2153 , \2155 );
and \U$1780 ( \2157 , \378 , \2156 );
not \U$1781 ( \2158 , \2157 );
xnor \U$1782 ( \2159 , \2158 , \2004 );
and \U$1783 ( \2160 , \410 , \1888 );
and \U$1784 ( \2161 , \392 , \1886 );
nor \U$1785 ( \2162 , \2160 , \2161 );
xnor \U$1786 ( \2163 , \2162 , \1732 );
and \U$1787 ( \2164 , \2159 , \2163 );
and \U$1788 ( \2165 , \479 , \1616 );
and \U$1789 ( \2166 , \431 , \1614 );
nor \U$1790 ( \2167 , \2165 , \2166 );
xnor \U$1791 ( \2168 , \2167 , \1503 );
and \U$1792 ( \2169 , \2163 , \2168 );
and \U$1793 ( \2170 , \2159 , \2168 );
or \U$1794 ( \2171 , \2164 , \2169 , \2170 );
and \U$1795 ( \2172 , \2151 , \2171 );
and \U$1796 ( \2173 , \2135 , \2171 );
or \U$1797 ( \2174 , \2152 , \2172 , \2173 );
and \U$1798 ( \2175 , \2119 , \2174 );
and \U$1799 ( \2176 , \2104 , \379 );
xor \U$1800 ( \2177 , \1970 , \1974 );
xor \U$1801 ( \2178 , \2177 , \1979 );
and \U$1802 ( \2179 , \2176 , \2178 );
xor \U$1803 ( \2180 , \2035 , \2039 );
xor \U$1804 ( \2181 , \2180 , \2044 );
and \U$1805 ( \2182 , \2178 , \2181 );
and \U$1806 ( \2183 , \2176 , \2181 );
or \U$1807 ( \2184 , \2179 , \2182 , \2183 );
and \U$1808 ( \2185 , \2174 , \2184 );
and \U$1809 ( \2186 , \2119 , \2184 );
or \U$1810 ( \2187 , \2175 , \2185 , \2186 );
xor \U$1811 ( \2188 , \1982 , \1998 );
xor \U$1812 ( \2189 , \2188 , \2017 );
xor \U$1813 ( \2190 , \2022 , \2024 );
xor \U$1814 ( \2191 , \2190 , \2027 );
and \U$1815 ( \2192 , \2189 , \2191 );
xor \U$1816 ( \2193 , \2047 , \2049 );
xor \U$1817 ( \2194 , \2193 , \2051 );
and \U$1818 ( \2195 , \2191 , \2194 );
and \U$1819 ( \2196 , \2189 , \2194 );
or \U$1820 ( \2197 , \2192 , \2195 , \2196 );
and \U$1821 ( \2198 , \2187 , \2197 );
xor \U$1822 ( \2199 , \1884 , \1903 );
xor \U$1823 ( \2200 , \2199 , \1920 );
and \U$1824 ( \2201 , \2197 , \2200 );
and \U$1825 ( \2202 , \2187 , \2200 );
or \U$1826 ( \2203 , \2198 , \2201 , \2202 );
xor \U$1827 ( \2204 , \2020 , \2030 );
xor \U$1828 ( \2205 , \2204 , \2054 );
xor \U$1829 ( \2206 , \2059 , \2061 );
xor \U$1830 ( \2207 , \2206 , \2064 );
and \U$1831 ( \2208 , \2205 , \2207 );
and \U$1832 ( \2209 , \2203 , \2208 );
xor \U$1833 ( \2210 , \1868 , \1923 );
xor \U$1834 ( \2211 , \2210 , \1934 );
and \U$1835 ( \2212 , \2208 , \2211 );
and \U$1836 ( \2213 , \2203 , \2211 );
or \U$1837 ( \2214 , \2209 , \2212 , \2213 );
xor \U$1838 ( \2215 , \2073 , \2075 );
xor \U$1839 ( \2216 , \2215 , \2078 );
and \U$1840 ( \2217 , \2214 , \2216 );
and \U$1841 ( \2218 , \2087 , \2217 );
xor \U$1842 ( \2219 , \2087 , \2217 );
xor \U$1843 ( \2220 , \2214 , \2216 );
buf \U$1844 ( \2221 , RIc226908_28);
buf \U$1845 ( \2222 , RIc226890_29);
and \U$1846 ( \2223 , \2221 , \2222 );
not \U$1847 ( \2224 , \2223 );
and \U$1848 ( \2225 , \2001 , \2224 );
not \U$1849 ( \2226 , \2225 );
and \U$1850 ( \2227 , \392 , \2156 );
and \U$1851 ( \2228 , \378 , \2154 );
nor \U$1852 ( \2229 , \2227 , \2228 );
xnor \U$1853 ( \2230 , \2229 , \2004 );
and \U$1854 ( \2231 , \2226 , \2230 );
and \U$1855 ( \2232 , \431 , \1888 );
and \U$1856 ( \2233 , \410 , \1886 );
nor \U$1857 ( \2234 , \2232 , \2233 );
xnor \U$1858 ( \2235 , \2234 , \1732 );
and \U$1859 ( \2236 , \2230 , \2235 );
and \U$1860 ( \2237 , \2226 , \2235 );
or \U$1861 ( \2238 , \2231 , \2236 , \2237 );
and \U$1862 ( \2239 , \487 , \1616 );
and \U$1863 ( \2240 , \479 , \1614 );
nor \U$1864 ( \2241 , \2239 , \2240 );
xnor \U$1865 ( \2242 , \2241 , \1503 );
and \U$1866 ( \2243 , \561 , \1422 );
and \U$1867 ( \2244 , \556 , \1420 );
nor \U$1868 ( \2245 , \2243 , \2244 );
xnor \U$1869 ( \2246 , \2245 , \1286 );
and \U$1870 ( \2247 , \2242 , \2246 );
and \U$1871 ( \2248 , \666 , \1222 );
and \U$1872 ( \2249 , \615 , \1220 );
nor \U$1873 ( \2250 , \2248 , \2249 );
xnor \U$1874 ( \2251 , \2250 , \1144 );
and \U$1875 ( \2252 , \2246 , \2251 );
and \U$1876 ( \2253 , \2242 , \2251 );
or \U$1877 ( \2254 , \2247 , \2252 , \2253 );
and \U$1878 ( \2255 , \2238 , \2254 );
and \U$1879 ( \2256 , \771 , \1058 );
and \U$1880 ( \2257 , \743 , \1056 );
nor \U$1881 ( \2258 , \2256 , \2257 );
xnor \U$1882 ( \2259 , \2258 , \964 );
and \U$1883 ( \2260 , \925 , \888 );
and \U$1884 ( \2261 , \851 , \886 );
nor \U$1885 ( \2262 , \2260 , \2261 );
xnor \U$1886 ( \2263 , \2262 , \816 );
and \U$1887 ( \2264 , \2259 , \2263 );
and \U$1888 ( \2265 , \1050 , \754 );
and \U$1889 ( \2266 , \987 , \752 );
nor \U$1890 ( \2267 , \2265 , \2266 );
xnor \U$1891 ( \2268 , \2267 , \711 );
and \U$1892 ( \2269 , \2263 , \2268 );
and \U$1893 ( \2270 , \2259 , \2268 );
or \U$1894 ( \2271 , \2264 , \2269 , \2270 );
and \U$1895 ( \2272 , \2254 , \2271 );
and \U$1896 ( \2273 , \2238 , \2271 );
or \U$1897 ( \2274 , \2255 , \2272 , \2273 );
xor \U$1898 ( \2275 , \2123 , \2127 );
xor \U$1899 ( \2276 , \2275 , \2132 );
xor \U$1900 ( \2277 , \2139 , \2143 );
xor \U$1901 ( \2278 , \2277 , \2148 );
and \U$1902 ( \2279 , \2276 , \2278 );
xor \U$1903 ( \2280 , \2091 , \2095 );
xor \U$1904 ( \2281 , \2280 , \2100 );
and \U$1905 ( \2282 , \2278 , \2281 );
and \U$1906 ( \2283 , \2276 , \2281 );
or \U$1907 ( \2284 , \2279 , \2282 , \2283 );
and \U$1908 ( \2285 , \2274 , \2284 );
and \U$1909 ( \2286 , \1861 , \422 );
and \U$1910 ( \2287 , \1853 , \420 );
nor \U$1911 ( \2288 , \2286 , \2287 );
xnor \U$1912 ( \2289 , \2288 , \403 );
and \U$1913 ( \2290 , \2109 , \385 );
and \U$1914 ( \2291 , \2104 , \383 );
nor \U$1915 ( \2292 , \2290 , \2291 );
xnor \U$1916 ( \2293 , \2292 , \390 );
and \U$1917 ( \2294 , \2289 , \2293 );
buf \U$1918 ( \2295 , RIc224b80_91);
and \U$1919 ( \2296 , \2295 , \379 );
and \U$1920 ( \2297 , \2293 , \2296 );
and \U$1921 ( \2298 , \2289 , \2296 );
or \U$1922 ( \2299 , \2294 , \2297 , \2298 );
and \U$1923 ( \2300 , \1336 , \641 );
and \U$1924 ( \2301 , \1248 , \639 );
nor \U$1925 ( \2302 , \2300 , \2301 );
xnor \U$1926 ( \2303 , \2302 , \592 );
and \U$1927 ( \2304 , \1446 , \540 );
and \U$1928 ( \2305 , \1441 , \538 );
nor \U$1929 ( \2306 , \2304 , \2305 );
xnor \U$1930 ( \2307 , \2306 , \499 );
and \U$1931 ( \2308 , \2303 , \2307 );
and \U$1932 ( \2309 , \1677 , \470 );
and \U$1933 ( \2310 , \1562 , \468 );
nor \U$1934 ( \2311 , \2309 , \2310 );
xnor \U$1935 ( \2312 , \2311 , \440 );
and \U$1936 ( \2313 , \2307 , \2312 );
and \U$1937 ( \2314 , \2303 , \2312 );
or \U$1938 ( \2315 , \2308 , \2313 , \2314 );
and \U$1939 ( \2316 , \2299 , \2315 );
xnor \U$1940 ( \2317 , \2108 , \2110 );
and \U$1941 ( \2318 , \2315 , \2317 );
and \U$1942 ( \2319 , \2299 , \2317 );
or \U$1943 ( \2320 , \2316 , \2318 , \2319 );
and \U$1944 ( \2321 , \2284 , \2320 );
and \U$1945 ( \2322 , \2274 , \2320 );
or \U$1946 ( \2323 , \2285 , \2321 , \2322 );
xor \U$1947 ( \2324 , \1986 , \1990 );
xor \U$1948 ( \2325 , \2324 , \1995 );
xor \U$1949 ( \2326 , \2005 , \2009 );
xor \U$1950 ( \2327 , \2326 , \2014 );
and \U$1951 ( \2328 , \2325 , \2327 );
xor \U$1952 ( \2329 , \2176 , \2178 );
xor \U$1953 ( \2330 , \2329 , \2181 );
and \U$1954 ( \2331 , \2327 , \2330 );
and \U$1955 ( \2332 , \2325 , \2330 );
or \U$1956 ( \2333 , \2328 , \2331 , \2332 );
and \U$1957 ( \2334 , \2323 , \2333 );
xor \U$1958 ( \2335 , \2189 , \2191 );
xor \U$1959 ( \2336 , \2335 , \2194 );
and \U$1960 ( \2337 , \2333 , \2336 );
and \U$1961 ( \2338 , \2323 , \2336 );
or \U$1962 ( \2339 , \2334 , \2337 , \2338 );
xor \U$1963 ( \2340 , \2187 , \2197 );
xor \U$1964 ( \2341 , \2340 , \2200 );
and \U$1965 ( \2342 , \2339 , \2341 );
xor \U$1966 ( \2343 , \2205 , \2207 );
and \U$1967 ( \2344 , \2341 , \2343 );
and \U$1968 ( \2345 , \2339 , \2343 );
or \U$1969 ( \2346 , \2342 , \2344 , \2345 );
xor \U$1970 ( \2347 , \2203 , \2208 );
xor \U$1971 ( \2348 , \2347 , \2211 );
and \U$1972 ( \2349 , \2346 , \2348 );
xor \U$1973 ( \2350 , \2057 , \2067 );
xor \U$1974 ( \2351 , \2350 , \2070 );
and \U$1975 ( \2352 , \2348 , \2351 );
and \U$1976 ( \2353 , \2346 , \2351 );
or \U$1977 ( \2354 , \2349 , \2352 , \2353 );
and \U$1978 ( \2355 , \2220 , \2354 );
xor \U$1979 ( \2356 , \2220 , \2354 );
xor \U$1980 ( \2357 , \2346 , \2348 );
xor \U$1981 ( \2358 , \2357 , \2351 );
xor \U$1982 ( \2359 , \2001 , \2221 );
xor \U$1983 ( \2360 , \2221 , \2222 );
not \U$1984 ( \2361 , \2360 );
and \U$1985 ( \2362 , \2359 , \2361 );
and \U$1986 ( \2363 , \378 , \2362 );
not \U$1987 ( \2364 , \2363 );
xnor \U$1988 ( \2365 , \2364 , \2225 );
and \U$1989 ( \2366 , \410 , \2156 );
and \U$1990 ( \2367 , \392 , \2154 );
nor \U$1991 ( \2368 , \2366 , \2367 );
xnor \U$1992 ( \2369 , \2368 , \2004 );
and \U$1993 ( \2370 , \2365 , \2369 );
and \U$1994 ( \2371 , \479 , \1888 );
and \U$1995 ( \2372 , \431 , \1886 );
nor \U$1996 ( \2373 , \2371 , \2372 );
xnor \U$1997 ( \2374 , \2373 , \1732 );
and \U$1998 ( \2375 , \2369 , \2374 );
and \U$1999 ( \2376 , \2365 , \2374 );
or \U$2000 ( \2377 , \2370 , \2375 , \2376 );
and \U$2001 ( \2378 , \556 , \1616 );
and \U$2002 ( \2379 , \487 , \1614 );
nor \U$2003 ( \2380 , \2378 , \2379 );
xnor \U$2004 ( \2381 , \2380 , \1503 );
and \U$2005 ( \2382 , \615 , \1422 );
and \U$2006 ( \2383 , \561 , \1420 );
nor \U$2007 ( \2384 , \2382 , \2383 );
xnor \U$2008 ( \2385 , \2384 , \1286 );
and \U$2009 ( \2386 , \2381 , \2385 );
and \U$2010 ( \2387 , \743 , \1222 );
and \U$2011 ( \2388 , \666 , \1220 );
nor \U$2012 ( \2389 , \2387 , \2388 );
xnor \U$2013 ( \2390 , \2389 , \1144 );
and \U$2014 ( \2391 , \2385 , \2390 );
and \U$2015 ( \2392 , \2381 , \2390 );
or \U$2016 ( \2393 , \2386 , \2391 , \2392 );
and \U$2017 ( \2394 , \2377 , \2393 );
and \U$2018 ( \2395 , \851 , \1058 );
and \U$2019 ( \2396 , \771 , \1056 );
nor \U$2020 ( \2397 , \2395 , \2396 );
xnor \U$2021 ( \2398 , \2397 , \964 );
and \U$2022 ( \2399 , \987 , \888 );
and \U$2023 ( \2400 , \925 , \886 );
nor \U$2024 ( \2401 , \2399 , \2400 );
xnor \U$2025 ( \2402 , \2401 , \816 );
and \U$2026 ( \2403 , \2398 , \2402 );
and \U$2027 ( \2404 , \1248 , \754 );
and \U$2028 ( \2405 , \1050 , \752 );
nor \U$2029 ( \2406 , \2404 , \2405 );
xnor \U$2030 ( \2407 , \2406 , \711 );
and \U$2031 ( \2408 , \2402 , \2407 );
and \U$2032 ( \2409 , \2398 , \2407 );
or \U$2033 ( \2410 , \2403 , \2408 , \2409 );
and \U$2034 ( \2411 , \2393 , \2410 );
and \U$2035 ( \2412 , \2377 , \2410 );
or \U$2036 ( \2413 , \2394 , \2411 , \2412 );
and \U$2037 ( \2414 , \1441 , \641 );
and \U$2038 ( \2415 , \1336 , \639 );
nor \U$2039 ( \2416 , \2414 , \2415 );
xnor \U$2040 ( \2417 , \2416 , \592 );
and \U$2041 ( \2418 , \1562 , \540 );
and \U$2042 ( \2419 , \1446 , \538 );
nor \U$2043 ( \2420 , \2418 , \2419 );
xnor \U$2044 ( \2421 , \2420 , \499 );
and \U$2045 ( \2422 , \2417 , \2421 );
and \U$2046 ( \2423 , \1853 , \470 );
and \U$2047 ( \2424 , \1677 , \468 );
nor \U$2048 ( \2425 , \2423 , \2424 );
xnor \U$2049 ( \2426 , \2425 , \440 );
and \U$2050 ( \2427 , \2421 , \2426 );
and \U$2051 ( \2428 , \2417 , \2426 );
or \U$2052 ( \2429 , \2422 , \2427 , \2428 );
and \U$2053 ( \2430 , \2104 , \422 );
and \U$2054 ( \2431 , \1861 , \420 );
nor \U$2055 ( \2432 , \2430 , \2431 );
xnor \U$2056 ( \2433 , \2432 , \403 );
and \U$2057 ( \2434 , \2295 , \385 );
and \U$2058 ( \2435 , \2109 , \383 );
nor \U$2059 ( \2436 , \2434 , \2435 );
xnor \U$2060 ( \2437 , \2436 , \390 );
and \U$2061 ( \2438 , \2433 , \2437 );
buf \U$2062 ( \2439 , RIc224b08_92);
and \U$2063 ( \2440 , \2439 , \379 );
and \U$2064 ( \2441 , \2437 , \2440 );
and \U$2065 ( \2442 , \2433 , \2440 );
or \U$2066 ( \2443 , \2438 , \2441 , \2442 );
and \U$2067 ( \2444 , \2429 , \2443 );
xor \U$2068 ( \2445 , \2289 , \2293 );
xor \U$2069 ( \2446 , \2445 , \2296 );
and \U$2070 ( \2447 , \2443 , \2446 );
and \U$2071 ( \2448 , \2429 , \2446 );
or \U$2072 ( \2449 , \2444 , \2447 , \2448 );
and \U$2073 ( \2450 , \2413 , \2449 );
xor \U$2074 ( \2451 , \2242 , \2246 );
xor \U$2075 ( \2452 , \2451 , \2251 );
xor \U$2076 ( \2453 , \2303 , \2307 );
xor \U$2077 ( \2454 , \2453 , \2312 );
and \U$2078 ( \2455 , \2452 , \2454 );
xor \U$2079 ( \2456 , \2259 , \2263 );
xor \U$2080 ( \2457 , \2456 , \2268 );
and \U$2081 ( \2458 , \2454 , \2457 );
and \U$2082 ( \2459 , \2452 , \2457 );
or \U$2083 ( \2460 , \2455 , \2458 , \2459 );
and \U$2084 ( \2461 , \2449 , \2460 );
and \U$2085 ( \2462 , \2413 , \2460 );
or \U$2086 ( \2463 , \2450 , \2461 , \2462 );
xor \U$2087 ( \2464 , \2159 , \2163 );
xor \U$2088 ( \2465 , \2464 , \2168 );
xor \U$2089 ( \2466 , \2276 , \2278 );
xor \U$2090 ( \2467 , \2466 , \2281 );
and \U$2091 ( \2468 , \2465 , \2467 );
xor \U$2092 ( \2469 , \2299 , \2315 );
xor \U$2093 ( \2470 , \2469 , \2317 );
and \U$2094 ( \2471 , \2467 , \2470 );
and \U$2095 ( \2472 , \2465 , \2470 );
or \U$2096 ( \2473 , \2468 , \2471 , \2472 );
and \U$2097 ( \2474 , \2463 , \2473 );
xor \U$2098 ( \2475 , \2103 , \2111 );
xor \U$2099 ( \2476 , \2475 , \2116 );
and \U$2100 ( \2477 , \2473 , \2476 );
and \U$2101 ( \2478 , \2463 , \2476 );
or \U$2102 ( \2479 , \2474 , \2477 , \2478 );
xor \U$2103 ( \2480 , \2135 , \2151 );
xor \U$2104 ( \2481 , \2480 , \2171 );
xor \U$2105 ( \2482 , \2274 , \2284 );
xor \U$2106 ( \2483 , \2482 , \2320 );
and \U$2107 ( \2484 , \2481 , \2483 );
xor \U$2108 ( \2485 , \2325 , \2327 );
xor \U$2109 ( \2486 , \2485 , \2330 );
and \U$2110 ( \2487 , \2483 , \2486 );
and \U$2111 ( \2488 , \2481 , \2486 );
or \U$2112 ( \2489 , \2484 , \2487 , \2488 );
and \U$2113 ( \2490 , \2479 , \2489 );
xor \U$2114 ( \2491 , \2119 , \2174 );
xor \U$2115 ( \2492 , \2491 , \2184 );
and \U$2116 ( \2493 , \2489 , \2492 );
and \U$2117 ( \2494 , \2479 , \2492 );
or \U$2118 ( \2495 , \2490 , \2493 , \2494 );
and \U$2119 ( \2496 , \487 , \1888 );
and \U$2120 ( \2497 , \479 , \1886 );
nor \U$2121 ( \2498 , \2496 , \2497 );
xnor \U$2122 ( \2499 , \2498 , \1732 );
and \U$2123 ( \2500 , \561 , \1616 );
and \U$2124 ( \2501 , \556 , \1614 );
nor \U$2125 ( \2502 , \2500 , \2501 );
xnor \U$2126 ( \2503 , \2502 , \1503 );
and \U$2127 ( \2504 , \2499 , \2503 );
and \U$2128 ( \2505 , \666 , \1422 );
and \U$2129 ( \2506 , \615 , \1420 );
nor \U$2130 ( \2507 , \2505 , \2506 );
xnor \U$2131 ( \2508 , \2507 , \1286 );
and \U$2132 ( \2509 , \2503 , \2508 );
and \U$2133 ( \2510 , \2499 , \2508 );
or \U$2134 ( \2511 , \2504 , \2509 , \2510 );
buf \U$2135 ( \2512 , RIc226818_30);
buf \U$2136 ( \2513 , RIc2267a0_31);
and \U$2137 ( \2514 , \2512 , \2513 );
not \U$2138 ( \2515 , \2514 );
and \U$2139 ( \2516 , \2222 , \2515 );
not \U$2140 ( \2517 , \2516 );
and \U$2141 ( \2518 , \392 , \2362 );
and \U$2142 ( \2519 , \378 , \2360 );
nor \U$2143 ( \2520 , \2518 , \2519 );
xnor \U$2144 ( \2521 , \2520 , \2225 );
and \U$2145 ( \2522 , \2517 , \2521 );
and \U$2146 ( \2523 , \431 , \2156 );
and \U$2147 ( \2524 , \410 , \2154 );
nor \U$2148 ( \2525 , \2523 , \2524 );
xnor \U$2149 ( \2526 , \2525 , \2004 );
and \U$2150 ( \2527 , \2521 , \2526 );
and \U$2151 ( \2528 , \2517 , \2526 );
or \U$2152 ( \2529 , \2522 , \2527 , \2528 );
and \U$2153 ( \2530 , \2511 , \2529 );
and \U$2154 ( \2531 , \771 , \1222 );
and \U$2155 ( \2532 , \743 , \1220 );
nor \U$2156 ( \2533 , \2531 , \2532 );
xnor \U$2157 ( \2534 , \2533 , \1144 );
and \U$2158 ( \2535 , \925 , \1058 );
and \U$2159 ( \2536 , \851 , \1056 );
nor \U$2160 ( \2537 , \2535 , \2536 );
xnor \U$2161 ( \2538 , \2537 , \964 );
and \U$2162 ( \2539 , \2534 , \2538 );
and \U$2163 ( \2540 , \1050 , \888 );
and \U$2164 ( \2541 , \987 , \886 );
nor \U$2165 ( \2542 , \2540 , \2541 );
xnor \U$2166 ( \2543 , \2542 , \816 );
and \U$2167 ( \2544 , \2538 , \2543 );
and \U$2168 ( \2545 , \2534 , \2543 );
or \U$2169 ( \2546 , \2539 , \2544 , \2545 );
and \U$2170 ( \2547 , \2529 , \2546 );
and \U$2171 ( \2548 , \2511 , \2546 );
or \U$2172 ( \2549 , \2530 , \2547 , \2548 );
xor \U$2173 ( \2550 , \2417 , \2421 );
xor \U$2174 ( \2551 , \2550 , \2426 );
xor \U$2175 ( \2552 , \2433 , \2437 );
xor \U$2176 ( \2553 , \2552 , \2440 );
and \U$2177 ( \2554 , \2551 , \2553 );
xor \U$2178 ( \2555 , \2398 , \2402 );
xor \U$2179 ( \2556 , \2555 , \2407 );
and \U$2180 ( \2557 , \2553 , \2556 );
and \U$2181 ( \2558 , \2551 , \2556 );
or \U$2182 ( \2559 , \2554 , \2557 , \2558 );
and \U$2183 ( \2560 , \2549 , \2559 );
and \U$2184 ( \2561 , \1861 , \470 );
and \U$2185 ( \2562 , \1853 , \468 );
nor \U$2186 ( \2563 , \2561 , \2562 );
xnor \U$2187 ( \2564 , \2563 , \440 );
and \U$2188 ( \2565 , \2109 , \422 );
and \U$2189 ( \2566 , \2104 , \420 );
nor \U$2190 ( \2567 , \2565 , \2566 );
xnor \U$2191 ( \2568 , \2567 , \403 );
and \U$2192 ( \2569 , \2564 , \2568 );
and \U$2193 ( \2570 , \2439 , \385 );
and \U$2194 ( \2571 , \2295 , \383 );
nor \U$2195 ( \2572 , \2570 , \2571 );
xnor \U$2196 ( \2573 , \2572 , \390 );
and \U$2197 ( \2574 , \2568 , \2573 );
and \U$2198 ( \2575 , \2564 , \2573 );
or \U$2199 ( \2576 , \2569 , \2574 , \2575 );
and \U$2200 ( \2577 , \1336 , \754 );
and \U$2201 ( \2578 , \1248 , \752 );
nor \U$2202 ( \2579 , \2577 , \2578 );
xnor \U$2203 ( \2580 , \2579 , \711 );
and \U$2204 ( \2581 , \1446 , \641 );
and \U$2205 ( \2582 , \1441 , \639 );
nor \U$2206 ( \2583 , \2581 , \2582 );
xnor \U$2207 ( \2584 , \2583 , \592 );
and \U$2208 ( \2585 , \2580 , \2584 );
and \U$2209 ( \2586 , \1677 , \540 );
and \U$2210 ( \2587 , \1562 , \538 );
nor \U$2211 ( \2588 , \2586 , \2587 );
xnor \U$2212 ( \2589 , \2588 , \499 );
and \U$2213 ( \2590 , \2584 , \2589 );
and \U$2214 ( \2591 , \2580 , \2589 );
or \U$2215 ( \2592 , \2585 , \2590 , \2591 );
or \U$2216 ( \2593 , \2576 , \2592 );
and \U$2217 ( \2594 , \2559 , \2593 );
and \U$2218 ( \2595 , \2549 , \2593 );
or \U$2219 ( \2596 , \2560 , \2594 , \2595 );
xor \U$2220 ( \2597 , \2226 , \2230 );
xor \U$2221 ( \2598 , \2597 , \2235 );
xor \U$2222 ( \2599 , \2429 , \2443 );
xor \U$2223 ( \2600 , \2599 , \2446 );
and \U$2224 ( \2601 , \2598 , \2600 );
xor \U$2225 ( \2602 , \2452 , \2454 );
xor \U$2226 ( \2603 , \2602 , \2457 );
and \U$2227 ( \2604 , \2600 , \2603 );
and \U$2228 ( \2605 , \2598 , \2603 );
or \U$2229 ( \2606 , \2601 , \2604 , \2605 );
and \U$2230 ( \2607 , \2596 , \2606 );
xor \U$2231 ( \2608 , \2238 , \2254 );
xor \U$2232 ( \2609 , \2608 , \2271 );
and \U$2233 ( \2610 , \2606 , \2609 );
and \U$2234 ( \2611 , \2596 , \2609 );
or \U$2235 ( \2612 , \2607 , \2610 , \2611 );
xor \U$2236 ( \2613 , \2463 , \2473 );
xor \U$2237 ( \2614 , \2613 , \2476 );
and \U$2238 ( \2615 , \2612 , \2614 );
xor \U$2239 ( \2616 , \2481 , \2483 );
xor \U$2240 ( \2617 , \2616 , \2486 );
and \U$2241 ( \2618 , \2614 , \2617 );
and \U$2242 ( \2619 , \2612 , \2617 );
or \U$2243 ( \2620 , \2615 , \2618 , \2619 );
xor \U$2244 ( \2621 , \2479 , \2489 );
xor \U$2245 ( \2622 , \2621 , \2492 );
and \U$2246 ( \2623 , \2620 , \2622 );
xor \U$2247 ( \2624 , \2323 , \2333 );
xor \U$2248 ( \2625 , \2624 , \2336 );
and \U$2249 ( \2626 , \2622 , \2625 );
and \U$2250 ( \2627 , \2620 , \2625 );
or \U$2251 ( \2628 , \2623 , \2626 , \2627 );
and \U$2252 ( \2629 , \2495 , \2628 );
xor \U$2253 ( \2630 , \2339 , \2341 );
xor \U$2254 ( \2631 , \2630 , \2343 );
and \U$2255 ( \2632 , \2628 , \2631 );
and \U$2256 ( \2633 , \2495 , \2631 );
or \U$2257 ( \2634 , \2629 , \2632 , \2633 );
and \U$2258 ( \2635 , \2358 , \2634 );
xor \U$2259 ( \2636 , \2358 , \2634 );
xor \U$2260 ( \2637 , \2495 , \2628 );
xor \U$2261 ( \2638 , \2637 , \2631 );
and \U$2262 ( \2639 , \556 , \1888 );
and \U$2263 ( \2640 , \487 , \1886 );
nor \U$2264 ( \2641 , \2639 , \2640 );
xnor \U$2265 ( \2642 , \2641 , \1732 );
and \U$2266 ( \2643 , \615 , \1616 );
and \U$2267 ( \2644 , \561 , \1614 );
nor \U$2268 ( \2645 , \2643 , \2644 );
xnor \U$2269 ( \2646 , \2645 , \1503 );
and \U$2270 ( \2647 , \2642 , \2646 );
and \U$2271 ( \2648 , \743 , \1422 );
and \U$2272 ( \2649 , \666 , \1420 );
nor \U$2273 ( \2650 , \2648 , \2649 );
xnor \U$2274 ( \2651 , \2650 , \1286 );
and \U$2275 ( \2652 , \2646 , \2651 );
and \U$2276 ( \2653 , \2642 , \2651 );
or \U$2277 ( \2654 , \2647 , \2652 , \2653 );
xor \U$2278 ( \2655 , \2222 , \2512 );
xor \U$2279 ( \2656 , \2512 , \2513 );
not \U$2280 ( \2657 , \2656 );
and \U$2281 ( \2658 , \2655 , \2657 );
and \U$2282 ( \2659 , \378 , \2658 );
not \U$2283 ( \2660 , \2659 );
xnor \U$2284 ( \2661 , \2660 , \2516 );
and \U$2285 ( \2662 , \410 , \2362 );
and \U$2286 ( \2663 , \392 , \2360 );
nor \U$2287 ( \2664 , \2662 , \2663 );
xnor \U$2288 ( \2665 , \2664 , \2225 );
and \U$2289 ( \2666 , \2661 , \2665 );
and \U$2290 ( \2667 , \479 , \2156 );
and \U$2291 ( \2668 , \431 , \2154 );
nor \U$2292 ( \2669 , \2667 , \2668 );
xnor \U$2293 ( \2670 , \2669 , \2004 );
and \U$2294 ( \2671 , \2665 , \2670 );
and \U$2295 ( \2672 , \2661 , \2670 );
or \U$2296 ( \2673 , \2666 , \2671 , \2672 );
and \U$2297 ( \2674 , \2654 , \2673 );
and \U$2298 ( \2675 , \851 , \1222 );
and \U$2299 ( \2676 , \771 , \1220 );
nor \U$2300 ( \2677 , \2675 , \2676 );
xnor \U$2301 ( \2678 , \2677 , \1144 );
and \U$2302 ( \2679 , \987 , \1058 );
and \U$2303 ( \2680 , \925 , \1056 );
nor \U$2304 ( \2681 , \2679 , \2680 );
xnor \U$2305 ( \2682 , \2681 , \964 );
and \U$2306 ( \2683 , \2678 , \2682 );
and \U$2307 ( \2684 , \1248 , \888 );
and \U$2308 ( \2685 , \1050 , \886 );
nor \U$2309 ( \2686 , \2684 , \2685 );
xnor \U$2310 ( \2687 , \2686 , \816 );
and \U$2311 ( \2688 , \2682 , \2687 );
and \U$2312 ( \2689 , \2678 , \2687 );
or \U$2313 ( \2690 , \2683 , \2688 , \2689 );
and \U$2314 ( \2691 , \2673 , \2690 );
and \U$2315 ( \2692 , \2654 , \2690 );
or \U$2316 ( \2693 , \2674 , \2691 , \2692 );
and \U$2317 ( \2694 , \2104 , \470 );
and \U$2318 ( \2695 , \1861 , \468 );
nor \U$2319 ( \2696 , \2694 , \2695 );
xnor \U$2320 ( \2697 , \2696 , \440 );
and \U$2321 ( \2698 , \2295 , \422 );
and \U$2322 ( \2699 , \2109 , \420 );
nor \U$2323 ( \2700 , \2698 , \2699 );
xnor \U$2324 ( \2701 , \2700 , \403 );
and \U$2325 ( \2702 , \2697 , \2701 );
buf \U$2326 ( \2703 , RIc224a90_93);
and \U$2327 ( \2704 , \2703 , \385 );
and \U$2328 ( \2705 , \2439 , \383 );
nor \U$2329 ( \2706 , \2704 , \2705 );
xnor \U$2330 ( \2707 , \2706 , \390 );
and \U$2331 ( \2708 , \2701 , \2707 );
and \U$2332 ( \2709 , \2697 , \2707 );
or \U$2333 ( \2710 , \2702 , \2708 , \2709 );
and \U$2334 ( \2711 , \1441 , \754 );
and \U$2335 ( \2712 , \1336 , \752 );
nor \U$2336 ( \2713 , \2711 , \2712 );
xnor \U$2337 ( \2714 , \2713 , \711 );
and \U$2338 ( \2715 , \1562 , \641 );
and \U$2339 ( \2716 , \1446 , \639 );
nor \U$2340 ( \2717 , \2715 , \2716 );
xnor \U$2341 ( \2718 , \2717 , \592 );
and \U$2342 ( \2719 , \2714 , \2718 );
and \U$2343 ( \2720 , \1853 , \540 );
and \U$2344 ( \2721 , \1677 , \538 );
nor \U$2345 ( \2722 , \2720 , \2721 );
xnor \U$2346 ( \2723 , \2722 , \499 );
and \U$2347 ( \2724 , \2718 , \2723 );
and \U$2348 ( \2725 , \2714 , \2723 );
or \U$2349 ( \2726 , \2719 , \2724 , \2725 );
and \U$2350 ( \2727 , \2710 , \2726 );
buf \U$2351 ( \2728 , RIc224a18_94);
and \U$2352 ( \2729 , \2728 , \379 );
buf \U$2353 ( \2730 , \2729 );
and \U$2354 ( \2731 , \2726 , \2730 );
and \U$2355 ( \2732 , \2710 , \2730 );
or \U$2356 ( \2733 , \2727 , \2731 , \2732 );
and \U$2357 ( \2734 , \2693 , \2733 );
and \U$2358 ( \2735 , \2703 , \379 );
xor \U$2359 ( \2736 , \2564 , \2568 );
xor \U$2360 ( \2737 , \2736 , \2573 );
and \U$2361 ( \2738 , \2735 , \2737 );
xor \U$2362 ( \2739 , \2580 , \2584 );
xor \U$2363 ( \2740 , \2739 , \2589 );
and \U$2364 ( \2741 , \2737 , \2740 );
and \U$2365 ( \2742 , \2735 , \2740 );
or \U$2366 ( \2743 , \2738 , \2741 , \2742 );
and \U$2367 ( \2744 , \2733 , \2743 );
and \U$2368 ( \2745 , \2693 , \2743 );
or \U$2369 ( \2746 , \2734 , \2744 , \2745 );
xor \U$2370 ( \2747 , \2499 , \2503 );
xor \U$2371 ( \2748 , \2747 , \2508 );
xor \U$2372 ( \2749 , \2517 , \2521 );
xor \U$2373 ( \2750 , \2749 , \2526 );
and \U$2374 ( \2751 , \2748 , \2750 );
xor \U$2375 ( \2752 , \2534 , \2538 );
xor \U$2376 ( \2753 , \2752 , \2543 );
and \U$2377 ( \2754 , \2750 , \2753 );
and \U$2378 ( \2755 , \2748 , \2753 );
or \U$2379 ( \2756 , \2751 , \2754 , \2755 );
xor \U$2380 ( \2757 , \2365 , \2369 );
xor \U$2381 ( \2758 , \2757 , \2374 );
and \U$2382 ( \2759 , \2756 , \2758 );
xor \U$2383 ( \2760 , \2381 , \2385 );
xor \U$2384 ( \2761 , \2760 , \2390 );
and \U$2385 ( \2762 , \2758 , \2761 );
and \U$2386 ( \2763 , \2756 , \2761 );
or \U$2387 ( \2764 , \2759 , \2762 , \2763 );
and \U$2388 ( \2765 , \2746 , \2764 );
xor \U$2389 ( \2766 , \2511 , \2529 );
xor \U$2390 ( \2767 , \2766 , \2546 );
xor \U$2391 ( \2768 , \2551 , \2553 );
xor \U$2392 ( \2769 , \2768 , \2556 );
and \U$2393 ( \2770 , \2767 , \2769 );
xnor \U$2394 ( \2771 , \2576 , \2592 );
and \U$2395 ( \2772 , \2769 , \2771 );
and \U$2396 ( \2773 , \2767 , \2771 );
or \U$2397 ( \2774 , \2770 , \2772 , \2773 );
and \U$2398 ( \2775 , \2764 , \2774 );
and \U$2399 ( \2776 , \2746 , \2774 );
or \U$2400 ( \2777 , \2765 , \2775 , \2776 );
xor \U$2401 ( \2778 , \2377 , \2393 );
xor \U$2402 ( \2779 , \2778 , \2410 );
xor \U$2403 ( \2780 , \2549 , \2559 );
xor \U$2404 ( \2781 , \2780 , \2593 );
and \U$2405 ( \2782 , \2779 , \2781 );
xor \U$2406 ( \2783 , \2598 , \2600 );
xor \U$2407 ( \2784 , \2783 , \2603 );
and \U$2408 ( \2785 , \2781 , \2784 );
and \U$2409 ( \2786 , \2779 , \2784 );
or \U$2410 ( \2787 , \2782 , \2785 , \2786 );
and \U$2411 ( \2788 , \2777 , \2787 );
xor \U$2412 ( \2789 , \2465 , \2467 );
xor \U$2413 ( \2790 , \2789 , \2470 );
and \U$2414 ( \2791 , \2787 , \2790 );
and \U$2415 ( \2792 , \2777 , \2790 );
or \U$2416 ( \2793 , \2788 , \2791 , \2792 );
xor \U$2417 ( \2794 , \2413 , \2449 );
xor \U$2418 ( \2795 , \2794 , \2460 );
xor \U$2419 ( \2796 , \2596 , \2606 );
xor \U$2420 ( \2797 , \2796 , \2609 );
and \U$2421 ( \2798 , \2795 , \2797 );
and \U$2422 ( \2799 , \2793 , \2798 );
xor \U$2423 ( \2800 , \2612 , \2614 );
xor \U$2424 ( \2801 , \2800 , \2617 );
and \U$2425 ( \2802 , \2798 , \2801 );
and \U$2426 ( \2803 , \2793 , \2801 );
or \U$2427 ( \2804 , \2799 , \2802 , \2803 );
xor \U$2428 ( \2805 , \2620 , \2622 );
xor \U$2429 ( \2806 , \2805 , \2625 );
and \U$2430 ( \2807 , \2804 , \2806 );
and \U$2431 ( \2808 , \2638 , \2807 );
xor \U$2432 ( \2809 , \2638 , \2807 );
xor \U$2433 ( \2810 , \2804 , \2806 );
and \U$2434 ( \2811 , \771 , \1422 );
and \U$2435 ( \2812 , \743 , \1420 );
nor \U$2436 ( \2813 , \2811 , \2812 );
xnor \U$2437 ( \2814 , \2813 , \1286 );
and \U$2438 ( \2815 , \925 , \1222 );
and \U$2439 ( \2816 , \851 , \1220 );
nor \U$2440 ( \2817 , \2815 , \2816 );
xnor \U$2441 ( \2818 , \2817 , \1144 );
and \U$2442 ( \2819 , \2814 , \2818 );
and \U$2443 ( \2820 , \1050 , \1058 );
and \U$2444 ( \2821 , \987 , \1056 );
nor \U$2445 ( \2822 , \2820 , \2821 );
xnor \U$2446 ( \2823 , \2822 , \964 );
and \U$2447 ( \2824 , \2818 , \2823 );
and \U$2448 ( \2825 , \2814 , \2823 );
or \U$2449 ( \2826 , \2819 , \2824 , \2825 );
buf \U$2450 ( \2827 , RIc226728_32);
buf \U$2451 ( \2828 , RIc2266b0_33);
and \U$2452 ( \2829 , \2827 , \2828 );
not \U$2453 ( \2830 , \2829 );
and \U$2454 ( \2831 , \2513 , \2830 );
not \U$2455 ( \2832 , \2831 );
and \U$2456 ( \2833 , \392 , \2658 );
and \U$2457 ( \2834 , \378 , \2656 );
nor \U$2458 ( \2835 , \2833 , \2834 );
xnor \U$2459 ( \2836 , \2835 , \2516 );
and \U$2460 ( \2837 , \2832 , \2836 );
and \U$2461 ( \2838 , \431 , \2362 );
and \U$2462 ( \2839 , \410 , \2360 );
nor \U$2463 ( \2840 , \2838 , \2839 );
xnor \U$2464 ( \2841 , \2840 , \2225 );
and \U$2465 ( \2842 , \2836 , \2841 );
and \U$2466 ( \2843 , \2832 , \2841 );
or \U$2467 ( \2844 , \2837 , \2842 , \2843 );
and \U$2468 ( \2845 , \2826 , \2844 );
and \U$2469 ( \2846 , \487 , \2156 );
and \U$2470 ( \2847 , \479 , \2154 );
nor \U$2471 ( \2848 , \2846 , \2847 );
xnor \U$2472 ( \2849 , \2848 , \2004 );
and \U$2473 ( \2850 , \561 , \1888 );
and \U$2474 ( \2851 , \556 , \1886 );
nor \U$2475 ( \2852 , \2850 , \2851 );
xnor \U$2476 ( \2853 , \2852 , \1732 );
and \U$2477 ( \2854 , \2849 , \2853 );
and \U$2478 ( \2855 , \666 , \1616 );
and \U$2479 ( \2856 , \615 , \1614 );
nor \U$2480 ( \2857 , \2855 , \2856 );
xnor \U$2481 ( \2858 , \2857 , \1503 );
and \U$2482 ( \2859 , \2853 , \2858 );
and \U$2483 ( \2860 , \2849 , \2858 );
or \U$2484 ( \2861 , \2854 , \2859 , \2860 );
and \U$2485 ( \2862 , \2844 , \2861 );
and \U$2486 ( \2863 , \2826 , \2861 );
or \U$2487 ( \2864 , \2845 , \2862 , \2863 );
and \U$2488 ( \2865 , \1861 , \540 );
and \U$2489 ( \2866 , \1853 , \538 );
nor \U$2490 ( \2867 , \2865 , \2866 );
xnor \U$2491 ( \2868 , \2867 , \499 );
and \U$2492 ( \2869 , \2109 , \470 );
and \U$2493 ( \2870 , \2104 , \468 );
nor \U$2494 ( \2871 , \2869 , \2870 );
xnor \U$2495 ( \2872 , \2871 , \440 );
and \U$2496 ( \2873 , \2868 , \2872 );
and \U$2497 ( \2874 , \2439 , \422 );
and \U$2498 ( \2875 , \2295 , \420 );
nor \U$2499 ( \2876 , \2874 , \2875 );
xnor \U$2500 ( \2877 , \2876 , \403 );
and \U$2501 ( \2878 , \2872 , \2877 );
and \U$2502 ( \2879 , \2868 , \2877 );
or \U$2503 ( \2880 , \2873 , \2878 , \2879 );
and \U$2504 ( \2881 , \1336 , \888 );
and \U$2505 ( \2882 , \1248 , \886 );
nor \U$2506 ( \2883 , \2881 , \2882 );
xnor \U$2507 ( \2884 , \2883 , \816 );
and \U$2508 ( \2885 , \1446 , \754 );
and \U$2509 ( \2886 , \1441 , \752 );
nor \U$2510 ( \2887 , \2885 , \2886 );
xnor \U$2511 ( \2888 , \2887 , \711 );
and \U$2512 ( \2889 , \2884 , \2888 );
and \U$2513 ( \2890 , \1677 , \641 );
and \U$2514 ( \2891 , \1562 , \639 );
nor \U$2515 ( \2892 , \2890 , \2891 );
xnor \U$2516 ( \2893 , \2892 , \592 );
and \U$2517 ( \2894 , \2888 , \2893 );
and \U$2518 ( \2895 , \2884 , \2893 );
or \U$2519 ( \2896 , \2889 , \2894 , \2895 );
and \U$2520 ( \2897 , \2880 , \2896 );
and \U$2521 ( \2898 , \2728 , \385 );
and \U$2522 ( \2899 , \2703 , \383 );
nor \U$2523 ( \2900 , \2898 , \2899 );
xnor \U$2524 ( \2901 , \2900 , \390 );
buf \U$2525 ( \2902 , RIc2249a0_95);
and \U$2526 ( \2903 , \2902 , \379 );
and \U$2527 ( \2904 , \2901 , \2903 );
and \U$2528 ( \2905 , \2896 , \2904 );
and \U$2529 ( \2906 , \2880 , \2904 );
or \U$2530 ( \2907 , \2897 , \2905 , \2906 );
and \U$2531 ( \2908 , \2864 , \2907 );
xor \U$2532 ( \2909 , \2697 , \2701 );
xor \U$2533 ( \2910 , \2909 , \2707 );
xor \U$2534 ( \2911 , \2714 , \2718 );
xor \U$2535 ( \2912 , \2911 , \2723 );
and \U$2536 ( \2913 , \2910 , \2912 );
not \U$2537 ( \2914 , \2729 );
and \U$2538 ( \2915 , \2912 , \2914 );
and \U$2539 ( \2916 , \2910 , \2914 );
or \U$2540 ( \2917 , \2913 , \2915 , \2916 );
and \U$2541 ( \2918 , \2907 , \2917 );
and \U$2542 ( \2919 , \2864 , \2917 );
or \U$2543 ( \2920 , \2908 , \2918 , \2919 );
xor \U$2544 ( \2921 , \2642 , \2646 );
xor \U$2545 ( \2922 , \2921 , \2651 );
xor \U$2546 ( \2923 , \2661 , \2665 );
xor \U$2547 ( \2924 , \2923 , \2670 );
and \U$2548 ( \2925 , \2922 , \2924 );
xor \U$2549 ( \2926 , \2678 , \2682 );
xor \U$2550 ( \2927 , \2926 , \2687 );
and \U$2551 ( \2928 , \2924 , \2927 );
and \U$2552 ( \2929 , \2922 , \2927 );
or \U$2553 ( \2930 , \2925 , \2928 , \2929 );
xor \U$2554 ( \2931 , \2748 , \2750 );
xor \U$2555 ( \2932 , \2931 , \2753 );
and \U$2556 ( \2933 , \2930 , \2932 );
xor \U$2557 ( \2934 , \2735 , \2737 );
xor \U$2558 ( \2935 , \2934 , \2740 );
and \U$2559 ( \2936 , \2932 , \2935 );
and \U$2560 ( \2937 , \2930 , \2935 );
or \U$2561 ( \2938 , \2933 , \2936 , \2937 );
and \U$2562 ( \2939 , \2920 , \2938 );
xor \U$2563 ( \2940 , \2654 , \2673 );
xor \U$2564 ( \2941 , \2940 , \2690 );
xor \U$2565 ( \2942 , \2710 , \2726 );
xor \U$2566 ( \2943 , \2942 , \2730 );
and \U$2567 ( \2944 , \2941 , \2943 );
and \U$2568 ( \2945 , \2938 , \2944 );
and \U$2569 ( \2946 , \2920 , \2944 );
or \U$2570 ( \2947 , \2939 , \2945 , \2946 );
xor \U$2571 ( \2948 , \2693 , \2733 );
xor \U$2572 ( \2949 , \2948 , \2743 );
xor \U$2573 ( \2950 , \2756 , \2758 );
xor \U$2574 ( \2951 , \2950 , \2761 );
and \U$2575 ( \2952 , \2949 , \2951 );
xor \U$2576 ( \2953 , \2767 , \2769 );
xor \U$2577 ( \2954 , \2953 , \2771 );
and \U$2578 ( \2955 , \2951 , \2954 );
and \U$2579 ( \2956 , \2949 , \2954 );
or \U$2580 ( \2957 , \2952 , \2955 , \2956 );
and \U$2581 ( \2958 , \2947 , \2957 );
xor \U$2582 ( \2959 , \2779 , \2781 );
xor \U$2583 ( \2960 , \2959 , \2784 );
and \U$2584 ( \2961 , \2957 , \2960 );
and \U$2585 ( \2962 , \2947 , \2960 );
or \U$2586 ( \2963 , \2958 , \2961 , \2962 );
xor \U$2587 ( \2964 , \2777 , \2787 );
xor \U$2588 ( \2965 , \2964 , \2790 );
and \U$2589 ( \2966 , \2963 , \2965 );
xor \U$2590 ( \2967 , \2795 , \2797 );
and \U$2591 ( \2968 , \2965 , \2967 );
and \U$2592 ( \2969 , \2963 , \2967 );
or \U$2593 ( \2970 , \2966 , \2968 , \2969 );
xor \U$2594 ( \2971 , \2793 , \2798 );
xor \U$2595 ( \2972 , \2971 , \2801 );
and \U$2596 ( \2973 , \2970 , \2972 );
and \U$2597 ( \2974 , \2810 , \2973 );
xor \U$2598 ( \2975 , \2810 , \2973 );
xor \U$2599 ( \2976 , \2970 , \2972 );
xor \U$2600 ( \2977 , \2513 , \2827 );
xor \U$2601 ( \2978 , \2827 , \2828 );
not \U$2602 ( \2979 , \2978 );
and \U$2603 ( \2980 , \2977 , \2979 );
and \U$2604 ( \2981 , \378 , \2980 );
not \U$2605 ( \2982 , \2981 );
xnor \U$2606 ( \2983 , \2982 , \2831 );
and \U$2607 ( \2984 , \410 , \2658 );
and \U$2608 ( \2985 , \392 , \2656 );
nor \U$2609 ( \2986 , \2984 , \2985 );
xnor \U$2610 ( \2987 , \2986 , \2516 );
and \U$2611 ( \2988 , \2983 , \2987 );
and \U$2612 ( \2989 , \479 , \2362 );
and \U$2613 ( \2990 , \431 , \2360 );
nor \U$2614 ( \2991 , \2989 , \2990 );
xnor \U$2615 ( \2992 , \2991 , \2225 );
and \U$2616 ( \2993 , \2987 , \2992 );
and \U$2617 ( \2994 , \2983 , \2992 );
or \U$2618 ( \2995 , \2988 , \2993 , \2994 );
and \U$2619 ( \2996 , \851 , \1422 );
and \U$2620 ( \2997 , \771 , \1420 );
nor \U$2621 ( \2998 , \2996 , \2997 );
xnor \U$2622 ( \2999 , \2998 , \1286 );
and \U$2623 ( \3000 , \987 , \1222 );
and \U$2624 ( \3001 , \925 , \1220 );
nor \U$2625 ( \3002 , \3000 , \3001 );
xnor \U$2626 ( \3003 , \3002 , \1144 );
and \U$2627 ( \3004 , \2999 , \3003 );
and \U$2628 ( \3005 , \1248 , \1058 );
and \U$2629 ( \3006 , \1050 , \1056 );
nor \U$2630 ( \3007 , \3005 , \3006 );
xnor \U$2631 ( \3008 , \3007 , \964 );
and \U$2632 ( \3009 , \3003 , \3008 );
and \U$2633 ( \3010 , \2999 , \3008 );
or \U$2634 ( \3011 , \3004 , \3009 , \3010 );
and \U$2635 ( \3012 , \2995 , \3011 );
and \U$2636 ( \3013 , \556 , \2156 );
and \U$2637 ( \3014 , \487 , \2154 );
nor \U$2638 ( \3015 , \3013 , \3014 );
xnor \U$2639 ( \3016 , \3015 , \2004 );
and \U$2640 ( \3017 , \615 , \1888 );
and \U$2641 ( \3018 , \561 , \1886 );
nor \U$2642 ( \3019 , \3017 , \3018 );
xnor \U$2643 ( \3020 , \3019 , \1732 );
and \U$2644 ( \3021 , \3016 , \3020 );
and \U$2645 ( \3022 , \743 , \1616 );
and \U$2646 ( \3023 , \666 , \1614 );
nor \U$2647 ( \3024 , \3022 , \3023 );
xnor \U$2648 ( \3025 , \3024 , \1503 );
and \U$2649 ( \3026 , \3020 , \3025 );
and \U$2650 ( \3027 , \3016 , \3025 );
or \U$2651 ( \3028 , \3021 , \3026 , \3027 );
and \U$2652 ( \3029 , \3011 , \3028 );
and \U$2653 ( \3030 , \2995 , \3028 );
or \U$2654 ( \3031 , \3012 , \3029 , \3030 );
and \U$2655 ( \3032 , \2104 , \540 );
and \U$2656 ( \3033 , \1861 , \538 );
nor \U$2657 ( \3034 , \3032 , \3033 );
xnor \U$2658 ( \3035 , \3034 , \499 );
and \U$2659 ( \3036 , \2295 , \470 );
and \U$2660 ( \3037 , \2109 , \468 );
nor \U$2661 ( \3038 , \3036 , \3037 );
xnor \U$2662 ( \3039 , \3038 , \440 );
and \U$2663 ( \3040 , \3035 , \3039 );
and \U$2664 ( \3041 , \2703 , \422 );
and \U$2665 ( \3042 , \2439 , \420 );
nor \U$2666 ( \3043 , \3041 , \3042 );
xnor \U$2667 ( \3044 , \3043 , \403 );
and \U$2668 ( \3045 , \3039 , \3044 );
and \U$2669 ( \3046 , \3035 , \3044 );
or \U$2670 ( \3047 , \3040 , \3045 , \3046 );
and \U$2671 ( \3048 , \1441 , \888 );
and \U$2672 ( \3049 , \1336 , \886 );
nor \U$2673 ( \3050 , \3048 , \3049 );
xnor \U$2674 ( \3051 , \3050 , \816 );
and \U$2675 ( \3052 , \1562 , \754 );
and \U$2676 ( \3053 , \1446 , \752 );
nor \U$2677 ( \3054 , \3052 , \3053 );
xnor \U$2678 ( \3055 , \3054 , \711 );
and \U$2679 ( \3056 , \3051 , \3055 );
and \U$2680 ( \3057 , \1853 , \641 );
and \U$2681 ( \3058 , \1677 , \639 );
nor \U$2682 ( \3059 , \3057 , \3058 );
xnor \U$2683 ( \3060 , \3059 , \592 );
and \U$2684 ( \3061 , \3055 , \3060 );
and \U$2685 ( \3062 , \3051 , \3060 );
or \U$2686 ( \3063 , \3056 , \3061 , \3062 );
and \U$2687 ( \3064 , \3047 , \3063 );
and \U$2688 ( \3065 , \2902 , \385 );
and \U$2689 ( \3066 , \2728 , \383 );
nor \U$2690 ( \3067 , \3065 , \3066 );
xnor \U$2691 ( \3068 , \3067 , \390 );
buf \U$2692 ( \3069 , RIc224928_96);
and \U$2693 ( \3070 , \3069 , \379 );
or \U$2694 ( \3071 , \3068 , \3070 );
and \U$2695 ( \3072 , \3063 , \3071 );
and \U$2696 ( \3073 , \3047 , \3071 );
or \U$2697 ( \3074 , \3064 , \3072 , \3073 );
and \U$2698 ( \3075 , \3031 , \3074 );
xor \U$2699 ( \3076 , \2868 , \2872 );
xor \U$2700 ( \3077 , \3076 , \2877 );
xor \U$2701 ( \3078 , \2884 , \2888 );
xor \U$2702 ( \3079 , \3078 , \2893 );
and \U$2703 ( \3080 , \3077 , \3079 );
xor \U$2704 ( \3081 , \2901 , \2903 );
and \U$2705 ( \3082 , \3079 , \3081 );
and \U$2706 ( \3083 , \3077 , \3081 );
or \U$2707 ( \3084 , \3080 , \3082 , \3083 );
and \U$2708 ( \3085 , \3074 , \3084 );
and \U$2709 ( \3086 , \3031 , \3084 );
or \U$2710 ( \3087 , \3075 , \3085 , \3086 );
xor \U$2711 ( \3088 , \2814 , \2818 );
xor \U$2712 ( \3089 , \3088 , \2823 );
xor \U$2713 ( \3090 , \2832 , \2836 );
xor \U$2714 ( \3091 , \3090 , \2841 );
and \U$2715 ( \3092 , \3089 , \3091 );
xor \U$2716 ( \3093 , \2849 , \2853 );
xor \U$2717 ( \3094 , \3093 , \2858 );
and \U$2718 ( \3095 , \3091 , \3094 );
and \U$2719 ( \3096 , \3089 , \3094 );
or \U$2720 ( \3097 , \3092 , \3095 , \3096 );
xor \U$2721 ( \3098 , \2922 , \2924 );
xor \U$2722 ( \3099 , \3098 , \2927 );
and \U$2723 ( \3100 , \3097 , \3099 );
xor \U$2724 ( \3101 , \2910 , \2912 );
xor \U$2725 ( \3102 , \3101 , \2914 );
and \U$2726 ( \3103 , \3099 , \3102 );
and \U$2727 ( \3104 , \3097 , \3102 );
or \U$2728 ( \3105 , \3100 , \3103 , \3104 );
and \U$2729 ( \3106 , \3087 , \3105 );
xor \U$2730 ( \3107 , \2826 , \2844 );
xor \U$2731 ( \3108 , \3107 , \2861 );
xor \U$2732 ( \3109 , \2880 , \2896 );
xor \U$2733 ( \3110 , \3109 , \2904 );
and \U$2734 ( \3111 , \3108 , \3110 );
and \U$2735 ( \3112 , \3105 , \3111 );
and \U$2736 ( \3113 , \3087 , \3111 );
or \U$2737 ( \3114 , \3106 , \3112 , \3113 );
xor \U$2738 ( \3115 , \2864 , \2907 );
xor \U$2739 ( \3116 , \3115 , \2917 );
xor \U$2740 ( \3117 , \2930 , \2932 );
xor \U$2741 ( \3118 , \3117 , \2935 );
and \U$2742 ( \3119 , \3116 , \3118 );
xor \U$2743 ( \3120 , \2941 , \2943 );
and \U$2744 ( \3121 , \3118 , \3120 );
and \U$2745 ( \3122 , \3116 , \3120 );
or \U$2746 ( \3123 , \3119 , \3121 , \3122 );
and \U$2747 ( \3124 , \3114 , \3123 );
xor \U$2748 ( \3125 , \2949 , \2951 );
xor \U$2749 ( \3126 , \3125 , \2954 );
and \U$2750 ( \3127 , \3123 , \3126 );
and \U$2751 ( \3128 , \3114 , \3126 );
or \U$2752 ( \3129 , \3124 , \3127 , \3128 );
xor \U$2753 ( \3130 , \2746 , \2764 );
xor \U$2754 ( \3131 , \3130 , \2774 );
and \U$2755 ( \3132 , \3129 , \3131 );
xor \U$2756 ( \3133 , \2947 , \2957 );
xor \U$2757 ( \3134 , \3133 , \2960 );
and \U$2758 ( \3135 , \3131 , \3134 );
and \U$2759 ( \3136 , \3129 , \3134 );
or \U$2760 ( \3137 , \3132 , \3135 , \3136 );
xor \U$2761 ( \3138 , \2963 , \2965 );
xor \U$2762 ( \3139 , \3138 , \2967 );
and \U$2763 ( \3140 , \3137 , \3139 );
and \U$2764 ( \3141 , \2976 , \3140 );
xor \U$2765 ( \3142 , \2976 , \3140 );
xor \U$2766 ( \3143 , \3137 , \3139 );
and \U$2767 ( \3144 , \487 , \2362 );
and \U$2768 ( \3145 , \479 , \2360 );
nor \U$2769 ( \3146 , \3144 , \3145 );
xnor \U$2770 ( \3147 , \3146 , \2225 );
and \U$2771 ( \3148 , \561 , \2156 );
and \U$2772 ( \3149 , \556 , \2154 );
nor \U$2773 ( \3150 , \3148 , \3149 );
xnor \U$2774 ( \3151 , \3150 , \2004 );
and \U$2775 ( \3152 , \3147 , \3151 );
and \U$2776 ( \3153 , \666 , \1888 );
and \U$2777 ( \3154 , \615 , \1886 );
nor \U$2778 ( \3155 , \3153 , \3154 );
xnor \U$2779 ( \3156 , \3155 , \1732 );
and \U$2780 ( \3157 , \3151 , \3156 );
and \U$2781 ( \3158 , \3147 , \3156 );
or \U$2782 ( \3159 , \3152 , \3157 , \3158 );
and \U$2783 ( \3160 , \771 , \1616 );
and \U$2784 ( \3161 , \743 , \1614 );
nor \U$2785 ( \3162 , \3160 , \3161 );
xnor \U$2786 ( \3163 , \3162 , \1503 );
and \U$2787 ( \3164 , \925 , \1422 );
and \U$2788 ( \3165 , \851 , \1420 );
nor \U$2789 ( \3166 , \3164 , \3165 );
xnor \U$2790 ( \3167 , \3166 , \1286 );
and \U$2791 ( \3168 , \3163 , \3167 );
and \U$2792 ( \3169 , \1050 , \1222 );
and \U$2793 ( \3170 , \987 , \1220 );
nor \U$2794 ( \3171 , \3169 , \3170 );
xnor \U$2795 ( \3172 , \3171 , \1144 );
and \U$2796 ( \3173 , \3167 , \3172 );
and \U$2797 ( \3174 , \3163 , \3172 );
or \U$2798 ( \3175 , \3168 , \3173 , \3174 );
and \U$2799 ( \3176 , \3159 , \3175 );
buf \U$2800 ( \3177 , RIc226638_34);
buf \U$2801 ( \3178 , RIc2265c0_35);
and \U$2802 ( \3179 , \3177 , \3178 );
not \U$2803 ( \3180 , \3179 );
and \U$2804 ( \3181 , \2828 , \3180 );
not \U$2805 ( \3182 , \3181 );
and \U$2806 ( \3183 , \392 , \2980 );
and \U$2807 ( \3184 , \378 , \2978 );
nor \U$2808 ( \3185 , \3183 , \3184 );
xnor \U$2809 ( \3186 , \3185 , \2831 );
and \U$2810 ( \3187 , \3182 , \3186 );
and \U$2811 ( \3188 , \431 , \2658 );
and \U$2812 ( \3189 , \410 , \2656 );
nor \U$2813 ( \3190 , \3188 , \3189 );
xnor \U$2814 ( \3191 , \3190 , \2516 );
and \U$2815 ( \3192 , \3186 , \3191 );
and \U$2816 ( \3193 , \3182 , \3191 );
or \U$2817 ( \3194 , \3187 , \3192 , \3193 );
and \U$2818 ( \3195 , \3175 , \3194 );
and \U$2819 ( \3196 , \3159 , \3194 );
or \U$2820 ( \3197 , \3176 , \3195 , \3196 );
and \U$2821 ( \3198 , \2728 , \422 );
and \U$2822 ( \3199 , \2703 , \420 );
nor \U$2823 ( \3200 , \3198 , \3199 );
xnor \U$2824 ( \3201 , \3200 , \403 );
and \U$2825 ( \3202 , \3069 , \385 );
and \U$2826 ( \3203 , \2902 , \383 );
nor \U$2827 ( \3204 , \3202 , \3203 );
xnor \U$2828 ( \3205 , \3204 , \390 );
and \U$2829 ( \3206 , \3201 , \3205 );
buf \U$2830 ( \3207 , RIc2248b0_97);
and \U$2831 ( \3208 , \3207 , \379 );
and \U$2832 ( \3209 , \3205 , \3208 );
and \U$2833 ( \3210 , \3201 , \3208 );
or \U$2834 ( \3211 , \3206 , \3209 , \3210 );
and \U$2835 ( \3212 , \1861 , \641 );
and \U$2836 ( \3213 , \1853 , \639 );
nor \U$2837 ( \3214 , \3212 , \3213 );
xnor \U$2838 ( \3215 , \3214 , \592 );
and \U$2839 ( \3216 , \2109 , \540 );
and \U$2840 ( \3217 , \2104 , \538 );
nor \U$2841 ( \3218 , \3216 , \3217 );
xnor \U$2842 ( \3219 , \3218 , \499 );
and \U$2843 ( \3220 , \3215 , \3219 );
and \U$2844 ( \3221 , \2439 , \470 );
and \U$2845 ( \3222 , \2295 , \468 );
nor \U$2846 ( \3223 , \3221 , \3222 );
xnor \U$2847 ( \3224 , \3223 , \440 );
and \U$2848 ( \3225 , \3219 , \3224 );
and \U$2849 ( \3226 , \3215 , \3224 );
or \U$2850 ( \3227 , \3220 , \3225 , \3226 );
and \U$2851 ( \3228 , \3211 , \3227 );
and \U$2852 ( \3229 , \1336 , \1058 );
and \U$2853 ( \3230 , \1248 , \1056 );
nor \U$2854 ( \3231 , \3229 , \3230 );
xnor \U$2855 ( \3232 , \3231 , \964 );
and \U$2856 ( \3233 , \1446 , \888 );
and \U$2857 ( \3234 , \1441 , \886 );
nor \U$2858 ( \3235 , \3233 , \3234 );
xnor \U$2859 ( \3236 , \3235 , \816 );
and \U$2860 ( \3237 , \3232 , \3236 );
and \U$2861 ( \3238 , \1677 , \754 );
and \U$2862 ( \3239 , \1562 , \752 );
nor \U$2863 ( \3240 , \3238 , \3239 );
xnor \U$2864 ( \3241 , \3240 , \711 );
and \U$2865 ( \3242 , \3236 , \3241 );
and \U$2866 ( \3243 , \3232 , \3241 );
or \U$2867 ( \3244 , \3237 , \3242 , \3243 );
and \U$2868 ( \3245 , \3227 , \3244 );
and \U$2869 ( \3246 , \3211 , \3244 );
or \U$2870 ( \3247 , \3228 , \3245 , \3246 );
and \U$2871 ( \3248 , \3197 , \3247 );
xor \U$2872 ( \3249 , \3035 , \3039 );
xor \U$2873 ( \3250 , \3249 , \3044 );
xor \U$2874 ( \3251 , \3051 , \3055 );
xor \U$2875 ( \3252 , \3251 , \3060 );
and \U$2876 ( \3253 , \3250 , \3252 );
xnor \U$2877 ( \3254 , \3068 , \3070 );
and \U$2878 ( \3255 , \3252 , \3254 );
and \U$2879 ( \3256 , \3250 , \3254 );
or \U$2880 ( \3257 , \3253 , \3255 , \3256 );
and \U$2881 ( \3258 , \3247 , \3257 );
and \U$2882 ( \3259 , \3197 , \3257 );
or \U$2883 ( \3260 , \3248 , \3258 , \3259 );
xor \U$2884 ( \3261 , \2983 , \2987 );
xor \U$2885 ( \3262 , \3261 , \2992 );
xor \U$2886 ( \3263 , \2999 , \3003 );
xor \U$2887 ( \3264 , \3263 , \3008 );
and \U$2888 ( \3265 , \3262 , \3264 );
xor \U$2889 ( \3266 , \3016 , \3020 );
xor \U$2890 ( \3267 , \3266 , \3025 );
and \U$2891 ( \3268 , \3264 , \3267 );
and \U$2892 ( \3269 , \3262 , \3267 );
or \U$2893 ( \3270 , \3265 , \3268 , \3269 );
xor \U$2894 ( \3271 , \3089 , \3091 );
xor \U$2895 ( \3272 , \3271 , \3094 );
and \U$2896 ( \3273 , \3270 , \3272 );
xor \U$2897 ( \3274 , \3077 , \3079 );
xor \U$2898 ( \3275 , \3274 , \3081 );
and \U$2899 ( \3276 , \3272 , \3275 );
and \U$2900 ( \3277 , \3270 , \3275 );
or \U$2901 ( \3278 , \3273 , \3276 , \3277 );
and \U$2902 ( \3279 , \3260 , \3278 );
xor \U$2903 ( \3280 , \2995 , \3011 );
xor \U$2904 ( \3281 , \3280 , \3028 );
xor \U$2905 ( \3282 , \3047 , \3063 );
xor \U$2906 ( \3283 , \3282 , \3071 );
and \U$2907 ( \3284 , \3281 , \3283 );
and \U$2908 ( \3285 , \3278 , \3284 );
and \U$2909 ( \3286 , \3260 , \3284 );
or \U$2910 ( \3287 , \3279 , \3285 , \3286 );
xor \U$2911 ( \3288 , \3031 , \3074 );
xor \U$2912 ( \3289 , \3288 , \3084 );
xor \U$2913 ( \3290 , \3097 , \3099 );
xor \U$2914 ( \3291 , \3290 , \3102 );
and \U$2915 ( \3292 , \3289 , \3291 );
xor \U$2916 ( \3293 , \3108 , \3110 );
and \U$2917 ( \3294 , \3291 , \3293 );
and \U$2918 ( \3295 , \3289 , \3293 );
or \U$2919 ( \3296 , \3292 , \3294 , \3295 );
and \U$2920 ( \3297 , \3287 , \3296 );
xor \U$2921 ( \3298 , \3116 , \3118 );
xor \U$2922 ( \3299 , \3298 , \3120 );
and \U$2923 ( \3300 , \3296 , \3299 );
and \U$2924 ( \3301 , \3287 , \3299 );
or \U$2925 ( \3302 , \3297 , \3300 , \3301 );
xor \U$2926 ( \3303 , \2920 , \2938 );
xor \U$2927 ( \3304 , \3303 , \2944 );
and \U$2928 ( \3305 , \3302 , \3304 );
xor \U$2929 ( \3306 , \3114 , \3123 );
xor \U$2930 ( \3307 , \3306 , \3126 );
and \U$2931 ( \3308 , \3304 , \3307 );
and \U$2932 ( \3309 , \3302 , \3307 );
or \U$2933 ( \3310 , \3305 , \3308 , \3309 );
xor \U$2934 ( \3311 , \3129 , \3131 );
xor \U$2935 ( \3312 , \3311 , \3134 );
and \U$2936 ( \3313 , \3310 , \3312 );
and \U$2937 ( \3314 , \3143 , \3313 );
xor \U$2938 ( \3315 , \3143 , \3313 );
xor \U$2939 ( \3316 , \3310 , \3312 );
and \U$2940 ( \3317 , \2902 , \422 );
and \U$2941 ( \3318 , \2728 , \420 );
nor \U$2942 ( \3319 , \3317 , \3318 );
xnor \U$2943 ( \3320 , \3319 , \403 );
and \U$2944 ( \3321 , \3207 , \385 );
and \U$2945 ( \3322 , \3069 , \383 );
nor \U$2946 ( \3323 , \3321 , \3322 );
xnor \U$2947 ( \3324 , \3323 , \390 );
and \U$2948 ( \3325 , \3320 , \3324 );
buf \U$2949 ( \3326 , RIc224838_98);
and \U$2950 ( \3327 , \3326 , \379 );
and \U$2951 ( \3328 , \3324 , \3327 );
and \U$2952 ( \3329 , \3320 , \3327 );
or \U$2953 ( \3330 , \3325 , \3328 , \3329 );
and \U$2954 ( \3331 , \2104 , \641 );
and \U$2955 ( \3332 , \1861 , \639 );
nor \U$2956 ( \3333 , \3331 , \3332 );
xnor \U$2957 ( \3334 , \3333 , \592 );
and \U$2958 ( \3335 , \2295 , \540 );
and \U$2959 ( \3336 , \2109 , \538 );
nor \U$2960 ( \3337 , \3335 , \3336 );
xnor \U$2961 ( \3338 , \3337 , \499 );
and \U$2962 ( \3339 , \3334 , \3338 );
and \U$2963 ( \3340 , \2703 , \470 );
and \U$2964 ( \3341 , \2439 , \468 );
nor \U$2965 ( \3342 , \3340 , \3341 );
xnor \U$2966 ( \3343 , \3342 , \440 );
and \U$2967 ( \3344 , \3338 , \3343 );
and \U$2968 ( \3345 , \3334 , \3343 );
or \U$2969 ( \3346 , \3339 , \3344 , \3345 );
and \U$2970 ( \3347 , \3330 , \3346 );
and \U$2971 ( \3348 , \1441 , \1058 );
and \U$2972 ( \3349 , \1336 , \1056 );
nor \U$2973 ( \3350 , \3348 , \3349 );
xnor \U$2974 ( \3351 , \3350 , \964 );
and \U$2975 ( \3352 , \1562 , \888 );
and \U$2976 ( \3353 , \1446 , \886 );
nor \U$2977 ( \3354 , \3352 , \3353 );
xnor \U$2978 ( \3355 , \3354 , \816 );
and \U$2979 ( \3356 , \3351 , \3355 );
and \U$2980 ( \3357 , \1853 , \754 );
and \U$2981 ( \3358 , \1677 , \752 );
nor \U$2982 ( \3359 , \3357 , \3358 );
xnor \U$2983 ( \3360 , \3359 , \711 );
and \U$2984 ( \3361 , \3355 , \3360 );
and \U$2985 ( \3362 , \3351 , \3360 );
or \U$2986 ( \3363 , \3356 , \3361 , \3362 );
and \U$2987 ( \3364 , \3346 , \3363 );
and \U$2988 ( \3365 , \3330 , \3363 );
or \U$2989 ( \3366 , \3347 , \3364 , \3365 );
and \U$2990 ( \3367 , \556 , \2362 );
and \U$2991 ( \3368 , \487 , \2360 );
nor \U$2992 ( \3369 , \3367 , \3368 );
xnor \U$2993 ( \3370 , \3369 , \2225 );
and \U$2994 ( \3371 , \615 , \2156 );
and \U$2995 ( \3372 , \561 , \2154 );
nor \U$2996 ( \3373 , \3371 , \3372 );
xnor \U$2997 ( \3374 , \3373 , \2004 );
and \U$2998 ( \3375 , \3370 , \3374 );
and \U$2999 ( \3376 , \743 , \1888 );
and \U$3000 ( \3377 , \666 , \1886 );
nor \U$3001 ( \3378 , \3376 , \3377 );
xnor \U$3002 ( \3379 , \3378 , \1732 );
and \U$3003 ( \3380 , \3374 , \3379 );
and \U$3004 ( \3381 , \3370 , \3379 );
or \U$3005 ( \3382 , \3375 , \3380 , \3381 );
xor \U$3006 ( \3383 , \2828 , \3177 );
xor \U$3007 ( \3384 , \3177 , \3178 );
not \U$3008 ( \3385 , \3384 );
and \U$3009 ( \3386 , \3383 , \3385 );
and \U$3010 ( \3387 , \378 , \3386 );
not \U$3011 ( \3388 , \3387 );
xnor \U$3012 ( \3389 , \3388 , \3181 );
and \U$3013 ( \3390 , \410 , \2980 );
and \U$3014 ( \3391 , \392 , \2978 );
nor \U$3015 ( \3392 , \3390 , \3391 );
xnor \U$3016 ( \3393 , \3392 , \2831 );
and \U$3017 ( \3394 , \3389 , \3393 );
and \U$3018 ( \3395 , \479 , \2658 );
and \U$3019 ( \3396 , \431 , \2656 );
nor \U$3020 ( \3397 , \3395 , \3396 );
xnor \U$3021 ( \3398 , \3397 , \2516 );
and \U$3022 ( \3399 , \3393 , \3398 );
and \U$3023 ( \3400 , \3389 , \3398 );
or \U$3024 ( \3401 , \3394 , \3399 , \3400 );
and \U$3025 ( \3402 , \3382 , \3401 );
and \U$3026 ( \3403 , \851 , \1616 );
and \U$3027 ( \3404 , \771 , \1614 );
nor \U$3028 ( \3405 , \3403 , \3404 );
xnor \U$3029 ( \3406 , \3405 , \1503 );
and \U$3030 ( \3407 , \987 , \1422 );
and \U$3031 ( \3408 , \925 , \1420 );
nor \U$3032 ( \3409 , \3407 , \3408 );
xnor \U$3033 ( \3410 , \3409 , \1286 );
and \U$3034 ( \3411 , \3406 , \3410 );
and \U$3035 ( \3412 , \1248 , \1222 );
and \U$3036 ( \3413 , \1050 , \1220 );
nor \U$3037 ( \3414 , \3412 , \3413 );
xnor \U$3038 ( \3415 , \3414 , \1144 );
and \U$3039 ( \3416 , \3410 , \3415 );
and \U$3040 ( \3417 , \3406 , \3415 );
or \U$3041 ( \3418 , \3411 , \3416 , \3417 );
and \U$3042 ( \3419 , \3401 , \3418 );
and \U$3043 ( \3420 , \3382 , \3418 );
or \U$3044 ( \3421 , \3402 , \3419 , \3420 );
and \U$3045 ( \3422 , \3366 , \3421 );
xor \U$3046 ( \3423 , \3201 , \3205 );
xor \U$3047 ( \3424 , \3423 , \3208 );
xor \U$3048 ( \3425 , \3215 , \3219 );
xor \U$3049 ( \3426 , \3425 , \3224 );
and \U$3050 ( \3427 , \3424 , \3426 );
xor \U$3051 ( \3428 , \3232 , \3236 );
xor \U$3052 ( \3429 , \3428 , \3241 );
and \U$3053 ( \3430 , \3426 , \3429 );
and \U$3054 ( \3431 , \3424 , \3429 );
or \U$3055 ( \3432 , \3427 , \3430 , \3431 );
and \U$3056 ( \3433 , \3421 , \3432 );
and \U$3057 ( \3434 , \3366 , \3432 );
or \U$3058 ( \3435 , \3422 , \3433 , \3434 );
xor \U$3059 ( \3436 , \3147 , \3151 );
xor \U$3060 ( \3437 , \3436 , \3156 );
xor \U$3061 ( \3438 , \3163 , \3167 );
xor \U$3062 ( \3439 , \3438 , \3172 );
and \U$3063 ( \3440 , \3437 , \3439 );
xor \U$3064 ( \3441 , \3182 , \3186 );
xor \U$3065 ( \3442 , \3441 , \3191 );
and \U$3066 ( \3443 , \3439 , \3442 );
and \U$3067 ( \3444 , \3437 , \3442 );
or \U$3068 ( \3445 , \3440 , \3443 , \3444 );
xor \U$3069 ( \3446 , \3262 , \3264 );
xor \U$3070 ( \3447 , \3446 , \3267 );
and \U$3071 ( \3448 , \3445 , \3447 );
xor \U$3072 ( \3449 , \3250 , \3252 );
xor \U$3073 ( \3450 , \3449 , \3254 );
and \U$3074 ( \3451 , \3447 , \3450 );
and \U$3075 ( \3452 , \3445 , \3450 );
or \U$3076 ( \3453 , \3448 , \3451 , \3452 );
and \U$3077 ( \3454 , \3435 , \3453 );
xor \U$3078 ( \3455 , \3159 , \3175 );
xor \U$3079 ( \3456 , \3455 , \3194 );
xor \U$3080 ( \3457 , \3211 , \3227 );
xor \U$3081 ( \3458 , \3457 , \3244 );
and \U$3082 ( \3459 , \3456 , \3458 );
and \U$3083 ( \3460 , \3453 , \3459 );
and \U$3084 ( \3461 , \3435 , \3459 );
or \U$3085 ( \3462 , \3454 , \3460 , \3461 );
xor \U$3086 ( \3463 , \3197 , \3247 );
xor \U$3087 ( \3464 , \3463 , \3257 );
xor \U$3088 ( \3465 , \3270 , \3272 );
xor \U$3089 ( \3466 , \3465 , \3275 );
and \U$3090 ( \3467 , \3464 , \3466 );
xor \U$3091 ( \3468 , \3281 , \3283 );
and \U$3092 ( \3469 , \3466 , \3468 );
and \U$3093 ( \3470 , \3464 , \3468 );
or \U$3094 ( \3471 , \3467 , \3469 , \3470 );
and \U$3095 ( \3472 , \3462 , \3471 );
xor \U$3096 ( \3473 , \3289 , \3291 );
xor \U$3097 ( \3474 , \3473 , \3293 );
and \U$3098 ( \3475 , \3471 , \3474 );
and \U$3099 ( \3476 , \3462 , \3474 );
or \U$3100 ( \3477 , \3472 , \3475 , \3476 );
xor \U$3101 ( \3478 , \3087 , \3105 );
xor \U$3102 ( \3479 , \3478 , \3111 );
and \U$3103 ( \3480 , \3477 , \3479 );
xor \U$3104 ( \3481 , \3287 , \3296 );
xor \U$3105 ( \3482 , \3481 , \3299 );
and \U$3106 ( \3483 , \3479 , \3482 );
and \U$3107 ( \3484 , \3477 , \3482 );
or \U$3108 ( \3485 , \3480 , \3483 , \3484 );
xor \U$3109 ( \3486 , \3302 , \3304 );
xor \U$3110 ( \3487 , \3486 , \3307 );
and \U$3111 ( \3488 , \3485 , \3487 );
and \U$3112 ( \3489 , \3316 , \3488 );
xor \U$3113 ( \3490 , \3316 , \3488 );
xor \U$3114 ( \3491 , \3485 , \3487 );
and \U$3115 ( \3492 , \771 , \1888 );
and \U$3116 ( \3493 , \743 , \1886 );
nor \U$3117 ( \3494 , \3492 , \3493 );
xnor \U$3118 ( \3495 , \3494 , \1732 );
and \U$3119 ( \3496 , \925 , \1616 );
and \U$3120 ( \3497 , \851 , \1614 );
nor \U$3121 ( \3498 , \3496 , \3497 );
xnor \U$3122 ( \3499 , \3498 , \1503 );
and \U$3123 ( \3500 , \3495 , \3499 );
and \U$3124 ( \3501 , \1050 , \1422 );
and \U$3125 ( \3502 , \987 , \1420 );
nor \U$3126 ( \3503 , \3501 , \3502 );
xnor \U$3127 ( \3504 , \3503 , \1286 );
and \U$3128 ( \3505 , \3499 , \3504 );
and \U$3129 ( \3506 , \3495 , \3504 );
or \U$3130 ( \3507 , \3500 , \3505 , \3506 );
buf \U$3131 ( \3508 , RIc226548_36);
buf \U$3132 ( \3509 , RIc2264d0_37);
and \U$3133 ( \3510 , \3508 , \3509 );
not \U$3134 ( \3511 , \3510 );
and \U$3135 ( \3512 , \3178 , \3511 );
not \U$3136 ( \3513 , \3512 );
and \U$3137 ( \3514 , \392 , \3386 );
and \U$3138 ( \3515 , \378 , \3384 );
nor \U$3139 ( \3516 , \3514 , \3515 );
xnor \U$3140 ( \3517 , \3516 , \3181 );
and \U$3141 ( \3518 , \3513 , \3517 );
and \U$3142 ( \3519 , \431 , \2980 );
and \U$3143 ( \3520 , \410 , \2978 );
nor \U$3144 ( \3521 , \3519 , \3520 );
xnor \U$3145 ( \3522 , \3521 , \2831 );
and \U$3146 ( \3523 , \3517 , \3522 );
and \U$3147 ( \3524 , \3513 , \3522 );
or \U$3148 ( \3525 , \3518 , \3523 , \3524 );
and \U$3149 ( \3526 , \3507 , \3525 );
and \U$3150 ( \3527 , \487 , \2658 );
and \U$3151 ( \3528 , \479 , \2656 );
nor \U$3152 ( \3529 , \3527 , \3528 );
xnor \U$3153 ( \3530 , \3529 , \2516 );
and \U$3154 ( \3531 , \561 , \2362 );
and \U$3155 ( \3532 , \556 , \2360 );
nor \U$3156 ( \3533 , \3531 , \3532 );
xnor \U$3157 ( \3534 , \3533 , \2225 );
and \U$3158 ( \3535 , \3530 , \3534 );
and \U$3159 ( \3536 , \666 , \2156 );
and \U$3160 ( \3537 , \615 , \2154 );
nor \U$3161 ( \3538 , \3536 , \3537 );
xnor \U$3162 ( \3539 , \3538 , \2004 );
and \U$3163 ( \3540 , \3534 , \3539 );
and \U$3164 ( \3541 , \3530 , \3539 );
or \U$3165 ( \3542 , \3535 , \3540 , \3541 );
and \U$3166 ( \3543 , \3525 , \3542 );
and \U$3167 ( \3544 , \3507 , \3542 );
or \U$3168 ( \3545 , \3526 , \3543 , \3544 );
and \U$3169 ( \3546 , \2728 , \470 );
and \U$3170 ( \3547 , \2703 , \468 );
nor \U$3171 ( \3548 , \3546 , \3547 );
xnor \U$3172 ( \3549 , \3548 , \440 );
and \U$3173 ( \3550 , \3069 , \422 );
and \U$3174 ( \3551 , \2902 , \420 );
nor \U$3175 ( \3552 , \3550 , \3551 );
xnor \U$3176 ( \3553 , \3552 , \403 );
and \U$3177 ( \3554 , \3549 , \3553 );
and \U$3178 ( \3555 , \3326 , \385 );
and \U$3179 ( \3556 , \3207 , \383 );
nor \U$3180 ( \3557 , \3555 , \3556 );
xnor \U$3181 ( \3558 , \3557 , \390 );
and \U$3182 ( \3559 , \3553 , \3558 );
and \U$3183 ( \3560 , \3549 , \3558 );
or \U$3184 ( \3561 , \3554 , \3559 , \3560 );
and \U$3185 ( \3562 , \1336 , \1222 );
and \U$3186 ( \3563 , \1248 , \1220 );
nor \U$3187 ( \3564 , \3562 , \3563 );
xnor \U$3188 ( \3565 , \3564 , \1144 );
and \U$3189 ( \3566 , \1446 , \1058 );
and \U$3190 ( \3567 , \1441 , \1056 );
nor \U$3191 ( \3568 , \3566 , \3567 );
xnor \U$3192 ( \3569 , \3568 , \964 );
and \U$3193 ( \3570 , \3565 , \3569 );
and \U$3194 ( \3571 , \1677 , \888 );
and \U$3195 ( \3572 , \1562 , \886 );
nor \U$3196 ( \3573 , \3571 , \3572 );
xnor \U$3197 ( \3574 , \3573 , \816 );
and \U$3198 ( \3575 , \3569 , \3574 );
and \U$3199 ( \3576 , \3565 , \3574 );
or \U$3200 ( \3577 , \3570 , \3575 , \3576 );
and \U$3201 ( \3578 , \3561 , \3577 );
and \U$3202 ( \3579 , \1861 , \754 );
and \U$3203 ( \3580 , \1853 , \752 );
nor \U$3204 ( \3581 , \3579 , \3580 );
xnor \U$3205 ( \3582 , \3581 , \711 );
and \U$3206 ( \3583 , \2109 , \641 );
and \U$3207 ( \3584 , \2104 , \639 );
nor \U$3208 ( \3585 , \3583 , \3584 );
xnor \U$3209 ( \3586 , \3585 , \592 );
and \U$3210 ( \3587 , \3582 , \3586 );
and \U$3211 ( \3588 , \2439 , \540 );
and \U$3212 ( \3589 , \2295 , \538 );
nor \U$3213 ( \3590 , \3588 , \3589 );
xnor \U$3214 ( \3591 , \3590 , \499 );
and \U$3215 ( \3592 , \3586 , \3591 );
and \U$3216 ( \3593 , \3582 , \3591 );
or \U$3217 ( \3594 , \3587 , \3592 , \3593 );
and \U$3218 ( \3595 , \3577 , \3594 );
and \U$3219 ( \3596 , \3561 , \3594 );
or \U$3220 ( \3597 , \3578 , \3595 , \3596 );
and \U$3221 ( \3598 , \3545 , \3597 );
xor \U$3222 ( \3599 , \3320 , \3324 );
xor \U$3223 ( \3600 , \3599 , \3327 );
xor \U$3224 ( \3601 , \3334 , \3338 );
xor \U$3225 ( \3602 , \3601 , \3343 );
or \U$3226 ( \3603 , \3600 , \3602 );
and \U$3227 ( \3604 , \3597 , \3603 );
and \U$3228 ( \3605 , \3545 , \3603 );
or \U$3229 ( \3606 , \3598 , \3604 , \3605 );
xor \U$3230 ( \3607 , \3370 , \3374 );
xor \U$3231 ( \3608 , \3607 , \3379 );
xor \U$3232 ( \3609 , \3406 , \3410 );
xor \U$3233 ( \3610 , \3609 , \3415 );
and \U$3234 ( \3611 , \3608 , \3610 );
xor \U$3235 ( \3612 , \3351 , \3355 );
xor \U$3236 ( \3613 , \3612 , \3360 );
and \U$3237 ( \3614 , \3610 , \3613 );
and \U$3238 ( \3615 , \3608 , \3613 );
or \U$3239 ( \3616 , \3611 , \3614 , \3615 );
xor \U$3240 ( \3617 , \3424 , \3426 );
xor \U$3241 ( \3618 , \3617 , \3429 );
and \U$3242 ( \3619 , \3616 , \3618 );
xor \U$3243 ( \3620 , \3437 , \3439 );
xor \U$3244 ( \3621 , \3620 , \3442 );
and \U$3245 ( \3622 , \3618 , \3621 );
and \U$3246 ( \3623 , \3616 , \3621 );
or \U$3247 ( \3624 , \3619 , \3622 , \3623 );
and \U$3248 ( \3625 , \3606 , \3624 );
xor \U$3249 ( \3626 , \3330 , \3346 );
xor \U$3250 ( \3627 , \3626 , \3363 );
xor \U$3251 ( \3628 , \3382 , \3401 );
xor \U$3252 ( \3629 , \3628 , \3418 );
and \U$3253 ( \3630 , \3627 , \3629 );
and \U$3254 ( \3631 , \3624 , \3630 );
and \U$3255 ( \3632 , \3606 , \3630 );
or \U$3256 ( \3633 , \3625 , \3631 , \3632 );
xor \U$3257 ( \3634 , \3366 , \3421 );
xor \U$3258 ( \3635 , \3634 , \3432 );
xor \U$3259 ( \3636 , \3445 , \3447 );
xor \U$3260 ( \3637 , \3636 , \3450 );
and \U$3261 ( \3638 , \3635 , \3637 );
xor \U$3262 ( \3639 , \3456 , \3458 );
and \U$3263 ( \3640 , \3637 , \3639 );
and \U$3264 ( \3641 , \3635 , \3639 );
or \U$3265 ( \3642 , \3638 , \3640 , \3641 );
and \U$3266 ( \3643 , \3633 , \3642 );
xor \U$3267 ( \3644 , \3464 , \3466 );
xor \U$3268 ( \3645 , \3644 , \3468 );
and \U$3269 ( \3646 , \3642 , \3645 );
and \U$3270 ( \3647 , \3633 , \3645 );
or \U$3271 ( \3648 , \3643 , \3646 , \3647 );
xor \U$3272 ( \3649 , \3260 , \3278 );
xor \U$3273 ( \3650 , \3649 , \3284 );
and \U$3274 ( \3651 , \3648 , \3650 );
xor \U$3275 ( \3652 , \3462 , \3471 );
xor \U$3276 ( \3653 , \3652 , \3474 );
and \U$3277 ( \3654 , \3650 , \3653 );
and \U$3278 ( \3655 , \3648 , \3653 );
or \U$3279 ( \3656 , \3651 , \3654 , \3655 );
xor \U$3280 ( \3657 , \3477 , \3479 );
xor \U$3281 ( \3658 , \3657 , \3482 );
and \U$3282 ( \3659 , \3656 , \3658 );
and \U$3283 ( \3660 , \3491 , \3659 );
xor \U$3284 ( \3661 , \3491 , \3659 );
xor \U$3285 ( \3662 , \3656 , \3658 );
and \U$3286 ( \3663 , \851 , \1888 );
and \U$3287 ( \3664 , \771 , \1886 );
nor \U$3288 ( \3665 , \3663 , \3664 );
xnor \U$3289 ( \3666 , \3665 , \1732 );
and \U$3290 ( \3667 , \987 , \1616 );
and \U$3291 ( \3668 , \925 , \1614 );
nor \U$3292 ( \3669 , \3667 , \3668 );
xnor \U$3293 ( \3670 , \3669 , \1503 );
and \U$3294 ( \3671 , \3666 , \3670 );
and \U$3295 ( \3672 , \1248 , \1422 );
and \U$3296 ( \3673 , \1050 , \1420 );
nor \U$3297 ( \3674 , \3672 , \3673 );
xnor \U$3298 ( \3675 , \3674 , \1286 );
and \U$3299 ( \3676 , \3670 , \3675 );
and \U$3300 ( \3677 , \3666 , \3675 );
or \U$3301 ( \3678 , \3671 , \3676 , \3677 );
and \U$3302 ( \3679 , \556 , \2658 );
and \U$3303 ( \3680 , \487 , \2656 );
nor \U$3304 ( \3681 , \3679 , \3680 );
xnor \U$3305 ( \3682 , \3681 , \2516 );
and \U$3306 ( \3683 , \615 , \2362 );
and \U$3307 ( \3684 , \561 , \2360 );
nor \U$3308 ( \3685 , \3683 , \3684 );
xnor \U$3309 ( \3686 , \3685 , \2225 );
and \U$3310 ( \3687 , \3682 , \3686 );
and \U$3311 ( \3688 , \743 , \2156 );
and \U$3312 ( \3689 , \666 , \2154 );
nor \U$3313 ( \3690 , \3688 , \3689 );
xnor \U$3314 ( \3691 , \3690 , \2004 );
and \U$3315 ( \3692 , \3686 , \3691 );
and \U$3316 ( \3693 , \3682 , \3691 );
or \U$3317 ( \3694 , \3687 , \3692 , \3693 );
and \U$3318 ( \3695 , \3678 , \3694 );
xor \U$3319 ( \3696 , \3178 , \3508 );
xor \U$3320 ( \3697 , \3508 , \3509 );
not \U$3321 ( \3698 , \3697 );
and \U$3322 ( \3699 , \3696 , \3698 );
and \U$3323 ( \3700 , \378 , \3699 );
not \U$3324 ( \3701 , \3700 );
xnor \U$3325 ( \3702 , \3701 , \3512 );
and \U$3326 ( \3703 , \410 , \3386 );
and \U$3327 ( \3704 , \392 , \3384 );
nor \U$3328 ( \3705 , \3703 , \3704 );
xnor \U$3329 ( \3706 , \3705 , \3181 );
and \U$3330 ( \3707 , \3702 , \3706 );
and \U$3331 ( \3708 , \479 , \2980 );
and \U$3332 ( \3709 , \431 , \2978 );
nor \U$3333 ( \3710 , \3708 , \3709 );
xnor \U$3334 ( \3711 , \3710 , \2831 );
and \U$3335 ( \3712 , \3706 , \3711 );
and \U$3336 ( \3713 , \3702 , \3711 );
or \U$3337 ( \3714 , \3707 , \3712 , \3713 );
and \U$3338 ( \3715 , \3694 , \3714 );
and \U$3339 ( \3716 , \3678 , \3714 );
or \U$3340 ( \3717 , \3695 , \3715 , \3716 );
and \U$3341 ( \3718 , \1441 , \1222 );
and \U$3342 ( \3719 , \1336 , \1220 );
nor \U$3343 ( \3720 , \3718 , \3719 );
xnor \U$3344 ( \3721 , \3720 , \1144 );
and \U$3345 ( \3722 , \1562 , \1058 );
and \U$3346 ( \3723 , \1446 , \1056 );
nor \U$3347 ( \3724 , \3722 , \3723 );
xnor \U$3348 ( \3725 , \3724 , \964 );
and \U$3349 ( \3726 , \3721 , \3725 );
and \U$3350 ( \3727 , \1853 , \888 );
and \U$3351 ( \3728 , \1677 , \886 );
nor \U$3352 ( \3729 , \3727 , \3728 );
xnor \U$3353 ( \3730 , \3729 , \816 );
and \U$3354 ( \3731 , \3725 , \3730 );
and \U$3355 ( \3732 , \3721 , \3730 );
or \U$3356 ( \3733 , \3726 , \3731 , \3732 );
and \U$3357 ( \3734 , \2902 , \470 );
and \U$3358 ( \3735 , \2728 , \468 );
nor \U$3359 ( \3736 , \3734 , \3735 );
xnor \U$3360 ( \3737 , \3736 , \440 );
and \U$3361 ( \3738 , \3207 , \422 );
and \U$3362 ( \3739 , \3069 , \420 );
nor \U$3363 ( \3740 , \3738 , \3739 );
xnor \U$3364 ( \3741 , \3740 , \403 );
and \U$3365 ( \3742 , \3737 , \3741 );
buf \U$3366 ( \3743 , RIc2247c0_99);
and \U$3367 ( \3744 , \3743 , \385 );
and \U$3368 ( \3745 , \3326 , \383 );
nor \U$3369 ( \3746 , \3744 , \3745 );
xnor \U$3370 ( \3747 , \3746 , \390 );
and \U$3371 ( \3748 , \3741 , \3747 );
and \U$3372 ( \3749 , \3737 , \3747 );
or \U$3373 ( \3750 , \3742 , \3748 , \3749 );
and \U$3374 ( \3751 , \3733 , \3750 );
and \U$3375 ( \3752 , \2104 , \754 );
and \U$3376 ( \3753 , \1861 , \752 );
nor \U$3377 ( \3754 , \3752 , \3753 );
xnor \U$3378 ( \3755 , \3754 , \711 );
and \U$3379 ( \3756 , \2295 , \641 );
and \U$3380 ( \3757 , \2109 , \639 );
nor \U$3381 ( \3758 , \3756 , \3757 );
xnor \U$3382 ( \3759 , \3758 , \592 );
and \U$3383 ( \3760 , \3755 , \3759 );
and \U$3384 ( \3761 , \2703 , \540 );
and \U$3385 ( \3762 , \2439 , \538 );
nor \U$3386 ( \3763 , \3761 , \3762 );
xnor \U$3387 ( \3764 , \3763 , \499 );
and \U$3388 ( \3765 , \3759 , \3764 );
and \U$3389 ( \3766 , \3755 , \3764 );
or \U$3390 ( \3767 , \3760 , \3765 , \3766 );
and \U$3391 ( \3768 , \3750 , \3767 );
and \U$3392 ( \3769 , \3733 , \3767 );
or \U$3393 ( \3770 , \3751 , \3768 , \3769 );
and \U$3394 ( \3771 , \3717 , \3770 );
and \U$3395 ( \3772 , \3743 , \379 );
xor \U$3396 ( \3773 , \3549 , \3553 );
xor \U$3397 ( \3774 , \3773 , \3558 );
and \U$3398 ( \3775 , \3772 , \3774 );
xor \U$3399 ( \3776 , \3582 , \3586 );
xor \U$3400 ( \3777 , \3776 , \3591 );
and \U$3401 ( \3778 , \3774 , \3777 );
and \U$3402 ( \3779 , \3772 , \3777 );
or \U$3403 ( \3780 , \3775 , \3778 , \3779 );
and \U$3404 ( \3781 , \3770 , \3780 );
and \U$3405 ( \3782 , \3717 , \3780 );
or \U$3406 ( \3783 , \3771 , \3781 , \3782 );
xor \U$3407 ( \3784 , \3495 , \3499 );
xor \U$3408 ( \3785 , \3784 , \3504 );
xor \U$3409 ( \3786 , \3565 , \3569 );
xor \U$3410 ( \3787 , \3786 , \3574 );
and \U$3411 ( \3788 , \3785 , \3787 );
xor \U$3412 ( \3789 , \3530 , \3534 );
xor \U$3413 ( \3790 , \3789 , \3539 );
and \U$3414 ( \3791 , \3787 , \3790 );
and \U$3415 ( \3792 , \3785 , \3790 );
or \U$3416 ( \3793 , \3788 , \3791 , \3792 );
xor \U$3417 ( \3794 , \3389 , \3393 );
xor \U$3418 ( \3795 , \3794 , \3398 );
and \U$3419 ( \3796 , \3793 , \3795 );
xor \U$3420 ( \3797 , \3608 , \3610 );
xor \U$3421 ( \3798 , \3797 , \3613 );
and \U$3422 ( \3799 , \3795 , \3798 );
and \U$3423 ( \3800 , \3793 , \3798 );
or \U$3424 ( \3801 , \3796 , \3799 , \3800 );
and \U$3425 ( \3802 , \3783 , \3801 );
xor \U$3426 ( \3803 , \3507 , \3525 );
xor \U$3427 ( \3804 , \3803 , \3542 );
xor \U$3428 ( \3805 , \3561 , \3577 );
xor \U$3429 ( \3806 , \3805 , \3594 );
and \U$3430 ( \3807 , \3804 , \3806 );
xnor \U$3431 ( \3808 , \3600 , \3602 );
and \U$3432 ( \3809 , \3806 , \3808 );
and \U$3433 ( \3810 , \3804 , \3808 );
or \U$3434 ( \3811 , \3807 , \3809 , \3810 );
and \U$3435 ( \3812 , \3801 , \3811 );
and \U$3436 ( \3813 , \3783 , \3811 );
or \U$3437 ( \3814 , \3802 , \3812 , \3813 );
xor \U$3438 ( \3815 , \3545 , \3597 );
xor \U$3439 ( \3816 , \3815 , \3603 );
xor \U$3440 ( \3817 , \3616 , \3618 );
xor \U$3441 ( \3818 , \3817 , \3621 );
and \U$3442 ( \3819 , \3816 , \3818 );
xor \U$3443 ( \3820 , \3627 , \3629 );
and \U$3444 ( \3821 , \3818 , \3820 );
and \U$3445 ( \3822 , \3816 , \3820 );
or \U$3446 ( \3823 , \3819 , \3821 , \3822 );
and \U$3447 ( \3824 , \3814 , \3823 );
xor \U$3448 ( \3825 , \3635 , \3637 );
xor \U$3449 ( \3826 , \3825 , \3639 );
and \U$3450 ( \3827 , \3823 , \3826 );
and \U$3451 ( \3828 , \3814 , \3826 );
or \U$3452 ( \3829 , \3824 , \3827 , \3828 );
xor \U$3453 ( \3830 , \3435 , \3453 );
xor \U$3454 ( \3831 , \3830 , \3459 );
and \U$3455 ( \3832 , \3829 , \3831 );
xor \U$3456 ( \3833 , \3633 , \3642 );
xor \U$3457 ( \3834 , \3833 , \3645 );
and \U$3458 ( \3835 , \3831 , \3834 );
and \U$3459 ( \3836 , \3829 , \3834 );
or \U$3460 ( \3837 , \3832 , \3835 , \3836 );
xor \U$3461 ( \3838 , \3648 , \3650 );
xor \U$3462 ( \3839 , \3838 , \3653 );
and \U$3463 ( \3840 , \3837 , \3839 );
and \U$3464 ( \3841 , \3662 , \3840 );
xor \U$3465 ( \3842 , \3662 , \3840 );
xor \U$3466 ( \3843 , \3837 , \3839 );
buf \U$3467 ( \3844 , RIc226458_38);
buf \U$3468 ( \3845 , RIc2263e0_39);
and \U$3469 ( \3846 , \3844 , \3845 );
not \U$3470 ( \3847 , \3846 );
and \U$3471 ( \3848 , \3509 , \3847 );
not \U$3472 ( \3849 , \3848 );
and \U$3473 ( \3850 , \392 , \3699 );
and \U$3474 ( \3851 , \378 , \3697 );
nor \U$3475 ( \3852 , \3850 , \3851 );
xnor \U$3476 ( \3853 , \3852 , \3512 );
and \U$3477 ( \3854 , \3849 , \3853 );
and \U$3478 ( \3855 , \431 , \3386 );
and \U$3479 ( \3856 , \410 , \3384 );
nor \U$3480 ( \3857 , \3855 , \3856 );
xnor \U$3481 ( \3858 , \3857 , \3181 );
and \U$3482 ( \3859 , \3853 , \3858 );
and \U$3483 ( \3860 , \3849 , \3858 );
or \U$3484 ( \3861 , \3854 , \3859 , \3860 );
and \U$3485 ( \3862 , \487 , \2980 );
and \U$3486 ( \3863 , \479 , \2978 );
nor \U$3487 ( \3864 , \3862 , \3863 );
xnor \U$3488 ( \3865 , \3864 , \2831 );
and \U$3489 ( \3866 , \561 , \2658 );
and \U$3490 ( \3867 , \556 , \2656 );
nor \U$3491 ( \3868 , \3866 , \3867 );
xnor \U$3492 ( \3869 , \3868 , \2516 );
and \U$3493 ( \3870 , \3865 , \3869 );
and \U$3494 ( \3871 , \666 , \2362 );
and \U$3495 ( \3872 , \615 , \2360 );
nor \U$3496 ( \3873 , \3871 , \3872 );
xnor \U$3497 ( \3874 , \3873 , \2225 );
and \U$3498 ( \3875 , \3869 , \3874 );
and \U$3499 ( \3876 , \3865 , \3874 );
or \U$3500 ( \3877 , \3870 , \3875 , \3876 );
and \U$3501 ( \3878 , \3861 , \3877 );
and \U$3502 ( \3879 , \771 , \2156 );
and \U$3503 ( \3880 , \743 , \2154 );
nor \U$3504 ( \3881 , \3879 , \3880 );
xnor \U$3505 ( \3882 , \3881 , \2004 );
and \U$3506 ( \3883 , \925 , \1888 );
and \U$3507 ( \3884 , \851 , \1886 );
nor \U$3508 ( \3885 , \3883 , \3884 );
xnor \U$3509 ( \3886 , \3885 , \1732 );
and \U$3510 ( \3887 , \3882 , \3886 );
and \U$3511 ( \3888 , \1050 , \1616 );
and \U$3512 ( \3889 , \987 , \1614 );
nor \U$3513 ( \3890 , \3888 , \3889 );
xnor \U$3514 ( \3891 , \3890 , \1503 );
and \U$3515 ( \3892 , \3886 , \3891 );
and \U$3516 ( \3893 , \3882 , \3891 );
or \U$3517 ( \3894 , \3887 , \3892 , \3893 );
and \U$3518 ( \3895 , \3877 , \3894 );
and \U$3519 ( \3896 , \3861 , \3894 );
or \U$3520 ( \3897 , \3878 , \3895 , \3896 );
and \U$3521 ( \3898 , \1861 , \888 );
and \U$3522 ( \3899 , \1853 , \886 );
nor \U$3523 ( \3900 , \3898 , \3899 );
xnor \U$3524 ( \3901 , \3900 , \816 );
and \U$3525 ( \3902 , \2109 , \754 );
and \U$3526 ( \3903 , \2104 , \752 );
nor \U$3527 ( \3904 , \3902 , \3903 );
xnor \U$3528 ( \3905 , \3904 , \711 );
and \U$3529 ( \3906 , \3901 , \3905 );
and \U$3530 ( \3907 , \2439 , \641 );
and \U$3531 ( \3908 , \2295 , \639 );
nor \U$3532 ( \3909 , \3907 , \3908 );
xnor \U$3533 ( \3910 , \3909 , \592 );
and \U$3534 ( \3911 , \3905 , \3910 );
and \U$3535 ( \3912 , \3901 , \3910 );
or \U$3536 ( \3913 , \3906 , \3911 , \3912 );
and \U$3537 ( \3914 , \1336 , \1422 );
and \U$3538 ( \3915 , \1248 , \1420 );
nor \U$3539 ( \3916 , \3914 , \3915 );
xnor \U$3540 ( \3917 , \3916 , \1286 );
and \U$3541 ( \3918 , \1446 , \1222 );
and \U$3542 ( \3919 , \1441 , \1220 );
nor \U$3543 ( \3920 , \3918 , \3919 );
xnor \U$3544 ( \3921 , \3920 , \1144 );
and \U$3545 ( \3922 , \3917 , \3921 );
and \U$3546 ( \3923 , \1677 , \1058 );
and \U$3547 ( \3924 , \1562 , \1056 );
nor \U$3548 ( \3925 , \3923 , \3924 );
xnor \U$3549 ( \3926 , \3925 , \964 );
and \U$3550 ( \3927 , \3921 , \3926 );
and \U$3551 ( \3928 , \3917 , \3926 );
or \U$3552 ( \3929 , \3922 , \3927 , \3928 );
and \U$3553 ( \3930 , \3913 , \3929 );
and \U$3554 ( \3931 , \2728 , \540 );
and \U$3555 ( \3932 , \2703 , \538 );
nor \U$3556 ( \3933 , \3931 , \3932 );
xnor \U$3557 ( \3934 , \3933 , \499 );
and \U$3558 ( \3935 , \3069 , \470 );
and \U$3559 ( \3936 , \2902 , \468 );
nor \U$3560 ( \3937 , \3935 , \3936 );
xnor \U$3561 ( \3938 , \3937 , \440 );
and \U$3562 ( \3939 , \3934 , \3938 );
and \U$3563 ( \3940 , \3326 , \422 );
and \U$3564 ( \3941 , \3207 , \420 );
nor \U$3565 ( \3942 , \3940 , \3941 );
xnor \U$3566 ( \3943 , \3942 , \403 );
and \U$3567 ( \3944 , \3938 , \3943 );
and \U$3568 ( \3945 , \3934 , \3943 );
or \U$3569 ( \3946 , \3939 , \3944 , \3945 );
and \U$3570 ( \3947 , \3929 , \3946 );
and \U$3571 ( \3948 , \3913 , \3946 );
or \U$3572 ( \3949 , \3930 , \3947 , \3948 );
and \U$3573 ( \3950 , \3897 , \3949 );
buf \U$3574 ( \3951 , RIc224748_100);
and \U$3575 ( \3952 , \3951 , \379 );
xor \U$3576 ( \3953 , \3737 , \3741 );
xor \U$3577 ( \3954 , \3953 , \3747 );
or \U$3578 ( \3955 , \3952 , \3954 );
and \U$3579 ( \3956 , \3949 , \3955 );
and \U$3580 ( \3957 , \3897 , \3955 );
or \U$3581 ( \3958 , \3950 , \3956 , \3957 );
xor \U$3582 ( \3959 , \3666 , \3670 );
xor \U$3583 ( \3960 , \3959 , \3675 );
xor \U$3584 ( \3961 , \3721 , \3725 );
xor \U$3585 ( \3962 , \3961 , \3730 );
and \U$3586 ( \3963 , \3960 , \3962 );
xor \U$3587 ( \3964 , \3755 , \3759 );
xor \U$3588 ( \3965 , \3964 , \3764 );
and \U$3589 ( \3966 , \3962 , \3965 );
and \U$3590 ( \3967 , \3960 , \3965 );
or \U$3591 ( \3968 , \3963 , \3966 , \3967 );
xor \U$3592 ( \3969 , \3513 , \3517 );
xor \U$3593 ( \3970 , \3969 , \3522 );
and \U$3594 ( \3971 , \3968 , \3970 );
xor \U$3595 ( \3972 , \3785 , \3787 );
xor \U$3596 ( \3973 , \3972 , \3790 );
and \U$3597 ( \3974 , \3970 , \3973 );
and \U$3598 ( \3975 , \3968 , \3973 );
or \U$3599 ( \3976 , \3971 , \3974 , \3975 );
and \U$3600 ( \3977 , \3958 , \3976 );
xor \U$3601 ( \3978 , \3678 , \3694 );
xor \U$3602 ( \3979 , \3978 , \3714 );
xor \U$3603 ( \3980 , \3733 , \3750 );
xor \U$3604 ( \3981 , \3980 , \3767 );
and \U$3605 ( \3982 , \3979 , \3981 );
xor \U$3606 ( \3983 , \3772 , \3774 );
xor \U$3607 ( \3984 , \3983 , \3777 );
and \U$3608 ( \3985 , \3981 , \3984 );
and \U$3609 ( \3986 , \3979 , \3984 );
or \U$3610 ( \3987 , \3982 , \3985 , \3986 );
and \U$3611 ( \3988 , \3976 , \3987 );
and \U$3612 ( \3989 , \3958 , \3987 );
or \U$3613 ( \3990 , \3977 , \3988 , \3989 );
xor \U$3614 ( \3991 , \3717 , \3770 );
xor \U$3615 ( \3992 , \3991 , \3780 );
xor \U$3616 ( \3993 , \3793 , \3795 );
xor \U$3617 ( \3994 , \3993 , \3798 );
and \U$3618 ( \3995 , \3992 , \3994 );
xor \U$3619 ( \3996 , \3804 , \3806 );
xor \U$3620 ( \3997 , \3996 , \3808 );
and \U$3621 ( \3998 , \3994 , \3997 );
and \U$3622 ( \3999 , \3992 , \3997 );
or \U$3623 ( \4000 , \3995 , \3998 , \3999 );
and \U$3624 ( \4001 , \3990 , \4000 );
xor \U$3625 ( \4002 , \3816 , \3818 );
xor \U$3626 ( \4003 , \4002 , \3820 );
and \U$3627 ( \4004 , \4000 , \4003 );
and \U$3628 ( \4005 , \3990 , \4003 );
or \U$3629 ( \4006 , \4001 , \4004 , \4005 );
xor \U$3630 ( \4007 , \3606 , \3624 );
xor \U$3631 ( \4008 , \4007 , \3630 );
and \U$3632 ( \4009 , \4006 , \4008 );
xor \U$3633 ( \4010 , \3814 , \3823 );
xor \U$3634 ( \4011 , \4010 , \3826 );
and \U$3635 ( \4012 , \4008 , \4011 );
and \U$3636 ( \4013 , \4006 , \4011 );
or \U$3637 ( \4014 , \4009 , \4012 , \4013 );
xor \U$3638 ( \4015 , \3829 , \3831 );
xor \U$3639 ( \4016 , \4015 , \3834 );
and \U$3640 ( \4017 , \4014 , \4016 );
and \U$3641 ( \4018 , \3843 , \4017 );
xor \U$3642 ( \4019 , \3843 , \4017 );
xor \U$3643 ( \4020 , \4014 , \4016 );
and \U$3644 ( \4021 , \1441 , \1422 );
and \U$3645 ( \4022 , \1336 , \1420 );
nor \U$3646 ( \4023 , \4021 , \4022 );
xnor \U$3647 ( \4024 , \4023 , \1286 );
and \U$3648 ( \4025 , \1562 , \1222 );
and \U$3649 ( \4026 , \1446 , \1220 );
nor \U$3650 ( \4027 , \4025 , \4026 );
xnor \U$3651 ( \4028 , \4027 , \1144 );
and \U$3652 ( \4029 , \4024 , \4028 );
and \U$3653 ( \4030 , \1853 , \1058 );
and \U$3654 ( \4031 , \1677 , \1056 );
nor \U$3655 ( \4032 , \4030 , \4031 );
xnor \U$3656 ( \4033 , \4032 , \964 );
and \U$3657 ( \4034 , \4028 , \4033 );
and \U$3658 ( \4035 , \4024 , \4033 );
or \U$3659 ( \4036 , \4029 , \4034 , \4035 );
and \U$3660 ( \4037 , \2104 , \888 );
and \U$3661 ( \4038 , \1861 , \886 );
nor \U$3662 ( \4039 , \4037 , \4038 );
xnor \U$3663 ( \4040 , \4039 , \816 );
and \U$3664 ( \4041 , \2295 , \754 );
and \U$3665 ( \4042 , \2109 , \752 );
nor \U$3666 ( \4043 , \4041 , \4042 );
xnor \U$3667 ( \4044 , \4043 , \711 );
and \U$3668 ( \4045 , \4040 , \4044 );
and \U$3669 ( \4046 , \2703 , \641 );
and \U$3670 ( \4047 , \2439 , \639 );
nor \U$3671 ( \4048 , \4046 , \4047 );
xnor \U$3672 ( \4049 , \4048 , \592 );
and \U$3673 ( \4050 , \4044 , \4049 );
and \U$3674 ( \4051 , \4040 , \4049 );
or \U$3675 ( \4052 , \4045 , \4050 , \4051 );
and \U$3676 ( \4053 , \4036 , \4052 );
and \U$3677 ( \4054 , \2902 , \540 );
and \U$3678 ( \4055 , \2728 , \538 );
nor \U$3679 ( \4056 , \4054 , \4055 );
xnor \U$3680 ( \4057 , \4056 , \499 );
and \U$3681 ( \4058 , \3207 , \470 );
and \U$3682 ( \4059 , \3069 , \468 );
nor \U$3683 ( \4060 , \4058 , \4059 );
xnor \U$3684 ( \4061 , \4060 , \440 );
and \U$3685 ( \4062 , \4057 , \4061 );
and \U$3686 ( \4063 , \3743 , \422 );
and \U$3687 ( \4064 , \3326 , \420 );
nor \U$3688 ( \4065 , \4063 , \4064 );
xnor \U$3689 ( \4066 , \4065 , \403 );
and \U$3690 ( \4067 , \4061 , \4066 );
and \U$3691 ( \4068 , \4057 , \4066 );
or \U$3692 ( \4069 , \4062 , \4067 , \4068 );
and \U$3693 ( \4070 , \4052 , \4069 );
and \U$3694 ( \4071 , \4036 , \4069 );
or \U$3695 ( \4072 , \4053 , \4070 , \4071 );
buf \U$3696 ( \4073 , RIc2246d0_101);
and \U$3697 ( \4074 , \4073 , \385 );
and \U$3698 ( \4075 , \3951 , \383 );
nor \U$3699 ( \4076 , \4074 , \4075 );
xnor \U$3700 ( \4077 , \4076 , \390 );
buf \U$3701 ( \4078 , RIc224658_102);
and \U$3702 ( \4079 , \4078 , \379 );
or \U$3703 ( \4080 , \4077 , \4079 );
and \U$3704 ( \4081 , \3951 , \385 );
and \U$3705 ( \4082 , \3743 , \383 );
nor \U$3706 ( \4083 , \4081 , \4082 );
xnor \U$3707 ( \4084 , \4083 , \390 );
and \U$3708 ( \4085 , \4080 , \4084 );
and \U$3709 ( \4086 , \4073 , \379 );
and \U$3710 ( \4087 , \4084 , \4086 );
and \U$3711 ( \4088 , \4080 , \4086 );
or \U$3712 ( \4089 , \4085 , \4087 , \4088 );
and \U$3713 ( \4090 , \4072 , \4089 );
xor \U$3714 ( \4091 , \3509 , \3844 );
xor \U$3715 ( \4092 , \3844 , \3845 );
not \U$3716 ( \4093 , \4092 );
and \U$3717 ( \4094 , \4091 , \4093 );
and \U$3718 ( \4095 , \378 , \4094 );
not \U$3719 ( \4096 , \4095 );
xnor \U$3720 ( \4097 , \4096 , \3848 );
and \U$3721 ( \4098 , \410 , \3699 );
and \U$3722 ( \4099 , \392 , \3697 );
nor \U$3723 ( \4100 , \4098 , \4099 );
xnor \U$3724 ( \4101 , \4100 , \3512 );
and \U$3725 ( \4102 , \4097 , \4101 );
and \U$3726 ( \4103 , \479 , \3386 );
and \U$3727 ( \4104 , \431 , \3384 );
nor \U$3728 ( \4105 , \4103 , \4104 );
xnor \U$3729 ( \4106 , \4105 , \3181 );
and \U$3730 ( \4107 , \4101 , \4106 );
and \U$3731 ( \4108 , \4097 , \4106 );
or \U$3732 ( \4109 , \4102 , \4107 , \4108 );
and \U$3733 ( \4110 , \556 , \2980 );
and \U$3734 ( \4111 , \487 , \2978 );
nor \U$3735 ( \4112 , \4110 , \4111 );
xnor \U$3736 ( \4113 , \4112 , \2831 );
and \U$3737 ( \4114 , \615 , \2658 );
and \U$3738 ( \4115 , \561 , \2656 );
nor \U$3739 ( \4116 , \4114 , \4115 );
xnor \U$3740 ( \4117 , \4116 , \2516 );
and \U$3741 ( \4118 , \4113 , \4117 );
and \U$3742 ( \4119 , \743 , \2362 );
and \U$3743 ( \4120 , \666 , \2360 );
nor \U$3744 ( \4121 , \4119 , \4120 );
xnor \U$3745 ( \4122 , \4121 , \2225 );
and \U$3746 ( \4123 , \4117 , \4122 );
and \U$3747 ( \4124 , \4113 , \4122 );
or \U$3748 ( \4125 , \4118 , \4123 , \4124 );
and \U$3749 ( \4126 , \4109 , \4125 );
and \U$3750 ( \4127 , \851 , \2156 );
and \U$3751 ( \4128 , \771 , \2154 );
nor \U$3752 ( \4129 , \4127 , \4128 );
xnor \U$3753 ( \4130 , \4129 , \2004 );
and \U$3754 ( \4131 , \987 , \1888 );
and \U$3755 ( \4132 , \925 , \1886 );
nor \U$3756 ( \4133 , \4131 , \4132 );
xnor \U$3757 ( \4134 , \4133 , \1732 );
and \U$3758 ( \4135 , \4130 , \4134 );
and \U$3759 ( \4136 , \1248 , \1616 );
and \U$3760 ( \4137 , \1050 , \1614 );
nor \U$3761 ( \4138 , \4136 , \4137 );
xnor \U$3762 ( \4139 , \4138 , \1503 );
and \U$3763 ( \4140 , \4134 , \4139 );
and \U$3764 ( \4141 , \4130 , \4139 );
or \U$3765 ( \4142 , \4135 , \4140 , \4141 );
and \U$3766 ( \4143 , \4125 , \4142 );
and \U$3767 ( \4144 , \4109 , \4142 );
or \U$3768 ( \4145 , \4126 , \4143 , \4144 );
and \U$3769 ( \4146 , \4089 , \4145 );
and \U$3770 ( \4147 , \4072 , \4145 );
or \U$3771 ( \4148 , \4090 , \4146 , \4147 );
xor \U$3772 ( \4149 , \3901 , \3905 );
xor \U$3773 ( \4150 , \4149 , \3910 );
xor \U$3774 ( \4151 , \3917 , \3921 );
xor \U$3775 ( \4152 , \4151 , \3926 );
and \U$3776 ( \4153 , \4150 , \4152 );
xor \U$3777 ( \4154 , \3934 , \3938 );
xor \U$3778 ( \4155 , \4154 , \3943 );
and \U$3779 ( \4156 , \4152 , \4155 );
and \U$3780 ( \4157 , \4150 , \4155 );
or \U$3781 ( \4158 , \4153 , \4156 , \4157 );
xor \U$3782 ( \4159 , \3849 , \3853 );
xor \U$3783 ( \4160 , \4159 , \3858 );
xor \U$3784 ( \4161 , \3865 , \3869 );
xor \U$3785 ( \4162 , \4161 , \3874 );
and \U$3786 ( \4163 , \4160 , \4162 );
xor \U$3787 ( \4164 , \3882 , \3886 );
xor \U$3788 ( \4165 , \4164 , \3891 );
and \U$3789 ( \4166 , \4162 , \4165 );
and \U$3790 ( \4167 , \4160 , \4165 );
or \U$3791 ( \4168 , \4163 , \4166 , \4167 );
and \U$3792 ( \4169 , \4158 , \4168 );
xor \U$3793 ( \4170 , \3682 , \3686 );
xor \U$3794 ( \4171 , \4170 , \3691 );
and \U$3795 ( \4172 , \4168 , \4171 );
and \U$3796 ( \4173 , \4158 , \4171 );
or \U$3797 ( \4174 , \4169 , \4172 , \4173 );
and \U$3798 ( \4175 , \4148 , \4174 );
xor \U$3799 ( \4176 , \3702 , \3706 );
xor \U$3800 ( \4177 , \4176 , \3711 );
xor \U$3801 ( \4178 , \3960 , \3962 );
xor \U$3802 ( \4179 , \4178 , \3965 );
and \U$3803 ( \4180 , \4177 , \4179 );
xnor \U$3804 ( \4181 , \3952 , \3954 );
and \U$3805 ( \4182 , \4179 , \4181 );
and \U$3806 ( \4183 , \4177 , \4181 );
or \U$3807 ( \4184 , \4180 , \4182 , \4183 );
and \U$3808 ( \4185 , \4174 , \4184 );
and \U$3809 ( \4186 , \4148 , \4184 );
or \U$3810 ( \4187 , \4175 , \4185 , \4186 );
xor \U$3811 ( \4188 , \3897 , \3949 );
xor \U$3812 ( \4189 , \4188 , \3955 );
xor \U$3813 ( \4190 , \3968 , \3970 );
xor \U$3814 ( \4191 , \4190 , \3973 );
and \U$3815 ( \4192 , \4189 , \4191 );
xor \U$3816 ( \4193 , \3979 , \3981 );
xor \U$3817 ( \4194 , \4193 , \3984 );
and \U$3818 ( \4195 , \4191 , \4194 );
and \U$3819 ( \4196 , \4189 , \4194 );
or \U$3820 ( \4197 , \4192 , \4195 , \4196 );
and \U$3821 ( \4198 , \4187 , \4197 );
xor \U$3822 ( \4199 , \3992 , \3994 );
xor \U$3823 ( \4200 , \4199 , \3997 );
and \U$3824 ( \4201 , \4197 , \4200 );
and \U$3825 ( \4202 , \4187 , \4200 );
or \U$3826 ( \4203 , \4198 , \4201 , \4202 );
xor \U$3827 ( \4204 , \3783 , \3801 );
xor \U$3828 ( \4205 , \4204 , \3811 );
and \U$3829 ( \4206 , \4203 , \4205 );
xor \U$3830 ( \4207 , \3990 , \4000 );
xor \U$3831 ( \4208 , \4207 , \4003 );
and \U$3832 ( \4209 , \4205 , \4208 );
and \U$3833 ( \4210 , \4203 , \4208 );
or \U$3834 ( \4211 , \4206 , \4209 , \4210 );
xor \U$3835 ( \4212 , \4006 , \4008 );
xor \U$3836 ( \4213 , \4212 , \4011 );
and \U$3837 ( \4214 , \4211 , \4213 );
and \U$3838 ( \4215 , \4020 , \4214 );
xor \U$3839 ( \4216 , \4020 , \4214 );
xor \U$3840 ( \4217 , \4211 , \4213 );
and \U$3841 ( \4218 , \1861 , \1058 );
and \U$3842 ( \4219 , \1853 , \1056 );
nor \U$3843 ( \4220 , \4218 , \4219 );
xnor \U$3844 ( \4221 , \4220 , \964 );
and \U$3845 ( \4222 , \2109 , \888 );
and \U$3846 ( \4223 , \2104 , \886 );
nor \U$3847 ( \4224 , \4222 , \4223 );
xnor \U$3848 ( \4225 , \4224 , \816 );
and \U$3849 ( \4226 , \4221 , \4225 );
and \U$3850 ( \4227 , \2439 , \754 );
and \U$3851 ( \4228 , \2295 , \752 );
nor \U$3852 ( \4229 , \4227 , \4228 );
xnor \U$3853 ( \4230 , \4229 , \711 );
and \U$3854 ( \4231 , \4225 , \4230 );
and \U$3855 ( \4232 , \4221 , \4230 );
or \U$3856 ( \4233 , \4226 , \4231 , \4232 );
and \U$3857 ( \4234 , \1336 , \1616 );
and \U$3858 ( \4235 , \1248 , \1614 );
nor \U$3859 ( \4236 , \4234 , \4235 );
xnor \U$3860 ( \4237 , \4236 , \1503 );
and \U$3861 ( \4238 , \1446 , \1422 );
and \U$3862 ( \4239 , \1441 , \1420 );
nor \U$3863 ( \4240 , \4238 , \4239 );
xnor \U$3864 ( \4241 , \4240 , \1286 );
and \U$3865 ( \4242 , \4237 , \4241 );
and \U$3866 ( \4243 , \1677 , \1222 );
and \U$3867 ( \4244 , \1562 , \1220 );
nor \U$3868 ( \4245 , \4243 , \4244 );
xnor \U$3869 ( \4246 , \4245 , \1144 );
and \U$3870 ( \4247 , \4241 , \4246 );
and \U$3871 ( \4248 , \4237 , \4246 );
or \U$3872 ( \4249 , \4242 , \4247 , \4248 );
and \U$3873 ( \4250 , \4233 , \4249 );
and \U$3874 ( \4251 , \2728 , \641 );
and \U$3875 ( \4252 , \2703 , \639 );
nor \U$3876 ( \4253 , \4251 , \4252 );
xnor \U$3877 ( \4254 , \4253 , \592 );
and \U$3878 ( \4255 , \3069 , \540 );
and \U$3879 ( \4256 , \2902 , \538 );
nor \U$3880 ( \4257 , \4255 , \4256 );
xnor \U$3881 ( \4258 , \4257 , \499 );
and \U$3882 ( \4259 , \4254 , \4258 );
and \U$3883 ( \4260 , \3326 , \470 );
and \U$3884 ( \4261 , \3207 , \468 );
nor \U$3885 ( \4262 , \4260 , \4261 );
xnor \U$3886 ( \4263 , \4262 , \440 );
and \U$3887 ( \4264 , \4258 , \4263 );
and \U$3888 ( \4265 , \4254 , \4263 );
or \U$3889 ( \4266 , \4259 , \4264 , \4265 );
and \U$3890 ( \4267 , \4249 , \4266 );
and \U$3891 ( \4268 , \4233 , \4266 );
or \U$3892 ( \4269 , \4250 , \4267 , \4268 );
buf \U$3893 ( \4270 , RIc226368_40);
buf \U$3894 ( \4271 , RIc2262f0_41);
and \U$3895 ( \4272 , \4270 , \4271 );
not \U$3896 ( \4273 , \4272 );
and \U$3897 ( \4274 , \3845 , \4273 );
not \U$3898 ( \4275 , \4274 );
and \U$3899 ( \4276 , \392 , \4094 );
and \U$3900 ( \4277 , \378 , \4092 );
nor \U$3901 ( \4278 , \4276 , \4277 );
xnor \U$3902 ( \4279 , \4278 , \3848 );
and \U$3903 ( \4280 , \4275 , \4279 );
and \U$3904 ( \4281 , \431 , \3699 );
and \U$3905 ( \4282 , \410 , \3697 );
nor \U$3906 ( \4283 , \4281 , \4282 );
xnor \U$3907 ( \4284 , \4283 , \3512 );
and \U$3908 ( \4285 , \4279 , \4284 );
and \U$3909 ( \4286 , \4275 , \4284 );
or \U$3910 ( \4287 , \4280 , \4285 , \4286 );
and \U$3911 ( \4288 , \487 , \3386 );
and \U$3912 ( \4289 , \479 , \3384 );
nor \U$3913 ( \4290 , \4288 , \4289 );
xnor \U$3914 ( \4291 , \4290 , \3181 );
and \U$3915 ( \4292 , \561 , \2980 );
and \U$3916 ( \4293 , \556 , \2978 );
nor \U$3917 ( \4294 , \4292 , \4293 );
xnor \U$3918 ( \4295 , \4294 , \2831 );
and \U$3919 ( \4296 , \4291 , \4295 );
and \U$3920 ( \4297 , \666 , \2658 );
and \U$3921 ( \4298 , \615 , \2656 );
nor \U$3922 ( \4299 , \4297 , \4298 );
xnor \U$3923 ( \4300 , \4299 , \2516 );
and \U$3924 ( \4301 , \4295 , \4300 );
and \U$3925 ( \4302 , \4291 , \4300 );
or \U$3926 ( \4303 , \4296 , \4301 , \4302 );
and \U$3927 ( \4304 , \4287 , \4303 );
and \U$3928 ( \4305 , \771 , \2362 );
and \U$3929 ( \4306 , \743 , \2360 );
nor \U$3930 ( \4307 , \4305 , \4306 );
xnor \U$3931 ( \4308 , \4307 , \2225 );
and \U$3932 ( \4309 , \925 , \2156 );
and \U$3933 ( \4310 , \851 , \2154 );
nor \U$3934 ( \4311 , \4309 , \4310 );
xnor \U$3935 ( \4312 , \4311 , \2004 );
and \U$3936 ( \4313 , \4308 , \4312 );
and \U$3937 ( \4314 , \1050 , \1888 );
and \U$3938 ( \4315 , \987 , \1886 );
nor \U$3939 ( \4316 , \4314 , \4315 );
xnor \U$3940 ( \4317 , \4316 , \1732 );
and \U$3941 ( \4318 , \4312 , \4317 );
and \U$3942 ( \4319 , \4308 , \4317 );
or \U$3943 ( \4320 , \4313 , \4318 , \4319 );
and \U$3944 ( \4321 , \4303 , \4320 );
and \U$3945 ( \4322 , \4287 , \4320 );
or \U$3946 ( \4323 , \4304 , \4321 , \4322 );
and \U$3947 ( \4324 , \4269 , \4323 );
and \U$3948 ( \4325 , \3951 , \422 );
and \U$3949 ( \4326 , \3743 , \420 );
nor \U$3950 ( \4327 , \4325 , \4326 );
xnor \U$3951 ( \4328 , \4327 , \403 );
and \U$3952 ( \4329 , \4078 , \385 );
and \U$3953 ( \4330 , \4073 , \383 );
nor \U$3954 ( \4331 , \4329 , \4330 );
xnor \U$3955 ( \4332 , \4331 , \390 );
and \U$3956 ( \4333 , \4328 , \4332 );
buf \U$3957 ( \4334 , RIc2245e0_103);
and \U$3958 ( \4335 , \4334 , \379 );
and \U$3959 ( \4336 , \4332 , \4335 );
and \U$3960 ( \4337 , \4328 , \4335 );
or \U$3961 ( \4338 , \4333 , \4336 , \4337 );
xor \U$3962 ( \4339 , \4057 , \4061 );
xor \U$3963 ( \4340 , \4339 , \4066 );
and \U$3964 ( \4341 , \4338 , \4340 );
xnor \U$3965 ( \4342 , \4077 , \4079 );
and \U$3966 ( \4343 , \4340 , \4342 );
and \U$3967 ( \4344 , \4338 , \4342 );
or \U$3968 ( \4345 , \4341 , \4343 , \4344 );
and \U$3969 ( \4346 , \4323 , \4345 );
and \U$3970 ( \4347 , \4269 , \4345 );
or \U$3971 ( \4348 , \4324 , \4346 , \4347 );
xor \U$3972 ( \4349 , \4024 , \4028 );
xor \U$3973 ( \4350 , \4349 , \4033 );
xor \U$3974 ( \4351 , \4040 , \4044 );
xor \U$3975 ( \4352 , \4351 , \4049 );
and \U$3976 ( \4353 , \4350 , \4352 );
xor \U$3977 ( \4354 , \4130 , \4134 );
xor \U$3978 ( \4355 , \4354 , \4139 );
and \U$3979 ( \4356 , \4352 , \4355 );
and \U$3980 ( \4357 , \4350 , \4355 );
or \U$3981 ( \4358 , \4353 , \4356 , \4357 );
xor \U$3982 ( \4359 , \4097 , \4101 );
xor \U$3983 ( \4360 , \4359 , \4106 );
xor \U$3984 ( \4361 , \4113 , \4117 );
xor \U$3985 ( \4362 , \4361 , \4122 );
and \U$3986 ( \4363 , \4360 , \4362 );
and \U$3987 ( \4364 , \4358 , \4363 );
xor \U$3988 ( \4365 , \4160 , \4162 );
xor \U$3989 ( \4366 , \4365 , \4165 );
and \U$3990 ( \4367 , \4363 , \4366 );
and \U$3991 ( \4368 , \4358 , \4366 );
or \U$3992 ( \4369 , \4364 , \4367 , \4368 );
and \U$3993 ( \4370 , \4348 , \4369 );
xor \U$3994 ( \4371 , \4036 , \4052 );
xor \U$3995 ( \4372 , \4371 , \4069 );
xor \U$3996 ( \4373 , \4080 , \4084 );
xor \U$3997 ( \4374 , \4373 , \4086 );
and \U$3998 ( \4375 , \4372 , \4374 );
xor \U$3999 ( \4376 , \4150 , \4152 );
xor \U$4000 ( \4377 , \4376 , \4155 );
and \U$4001 ( \4378 , \4374 , \4377 );
and \U$4002 ( \4379 , \4372 , \4377 );
or \U$4003 ( \4380 , \4375 , \4378 , \4379 );
and \U$4004 ( \4381 , \4369 , \4380 );
and \U$4005 ( \4382 , \4348 , \4380 );
or \U$4006 ( \4383 , \4370 , \4381 , \4382 );
xor \U$4007 ( \4384 , \3861 , \3877 );
xor \U$4008 ( \4385 , \4384 , \3894 );
xor \U$4009 ( \4386 , \3913 , \3929 );
xor \U$4010 ( \4387 , \4386 , \3946 );
and \U$4011 ( \4388 , \4385 , \4387 );
xor \U$4012 ( \4389 , \4177 , \4179 );
xor \U$4013 ( \4390 , \4389 , \4181 );
and \U$4014 ( \4391 , \4387 , \4390 );
and \U$4015 ( \4392 , \4385 , \4390 );
or \U$4016 ( \4393 , \4388 , \4391 , \4392 );
and \U$4017 ( \4394 , \4383 , \4393 );
xor \U$4018 ( \4395 , \4189 , \4191 );
xor \U$4019 ( \4396 , \4395 , \4194 );
and \U$4020 ( \4397 , \4393 , \4396 );
and \U$4021 ( \4398 , \4383 , \4396 );
or \U$4022 ( \4399 , \4394 , \4397 , \4398 );
xor \U$4023 ( \4400 , \3958 , \3976 );
xor \U$4024 ( \4401 , \4400 , \3987 );
and \U$4025 ( \4402 , \4399 , \4401 );
xor \U$4026 ( \4403 , \4187 , \4197 );
xor \U$4027 ( \4404 , \4403 , \4200 );
and \U$4028 ( \4405 , \4401 , \4404 );
and \U$4029 ( \4406 , \4399 , \4404 );
or \U$4030 ( \4407 , \4402 , \4405 , \4406 );
xor \U$4031 ( \4408 , \4203 , \4205 );
xor \U$4032 ( \4409 , \4408 , \4208 );
and \U$4033 ( \4410 , \4407 , \4409 );
and \U$4034 ( \4411 , \4217 , \4410 );
xor \U$4035 ( \4412 , \4217 , \4410 );
xor \U$4036 ( \4413 , \4407 , \4409 );
xor \U$4037 ( \4414 , \3845 , \4270 );
xor \U$4038 ( \4415 , \4270 , \4271 );
not \U$4039 ( \4416 , \4415 );
and \U$4040 ( \4417 , \4414 , \4416 );
and \U$4041 ( \4418 , \378 , \4417 );
not \U$4042 ( \4419 , \4418 );
xnor \U$4043 ( \4420 , \4419 , \4274 );
and \U$4044 ( \4421 , \410 , \4094 );
and \U$4045 ( \4422 , \392 , \4092 );
nor \U$4046 ( \4423 , \4421 , \4422 );
xnor \U$4047 ( \4424 , \4423 , \3848 );
and \U$4048 ( \4425 , \4420 , \4424 );
and \U$4049 ( \4426 , \479 , \3699 );
and \U$4050 ( \4427 , \431 , \3697 );
nor \U$4051 ( \4428 , \4426 , \4427 );
xnor \U$4052 ( \4429 , \4428 , \3512 );
and \U$4053 ( \4430 , \4424 , \4429 );
and \U$4054 ( \4431 , \4420 , \4429 );
or \U$4055 ( \4432 , \4425 , \4430 , \4431 );
and \U$4056 ( \4433 , \556 , \3386 );
and \U$4057 ( \4434 , \487 , \3384 );
nor \U$4058 ( \4435 , \4433 , \4434 );
xnor \U$4059 ( \4436 , \4435 , \3181 );
and \U$4060 ( \4437 , \615 , \2980 );
and \U$4061 ( \4438 , \561 , \2978 );
nor \U$4062 ( \4439 , \4437 , \4438 );
xnor \U$4063 ( \4440 , \4439 , \2831 );
and \U$4064 ( \4441 , \4436 , \4440 );
and \U$4065 ( \4442 , \743 , \2658 );
and \U$4066 ( \4443 , \666 , \2656 );
nor \U$4067 ( \4444 , \4442 , \4443 );
xnor \U$4068 ( \4445 , \4444 , \2516 );
and \U$4069 ( \4446 , \4440 , \4445 );
and \U$4070 ( \4447 , \4436 , \4445 );
or \U$4071 ( \4448 , \4441 , \4446 , \4447 );
and \U$4072 ( \4449 , \4432 , \4448 );
and \U$4073 ( \4450 , \851 , \2362 );
and \U$4074 ( \4451 , \771 , \2360 );
nor \U$4075 ( \4452 , \4450 , \4451 );
xnor \U$4076 ( \4453 , \4452 , \2225 );
and \U$4077 ( \4454 , \987 , \2156 );
and \U$4078 ( \4455 , \925 , \2154 );
nor \U$4079 ( \4456 , \4454 , \4455 );
xnor \U$4080 ( \4457 , \4456 , \2004 );
and \U$4081 ( \4458 , \4453 , \4457 );
and \U$4082 ( \4459 , \1248 , \1888 );
and \U$4083 ( \4460 , \1050 , \1886 );
nor \U$4084 ( \4461 , \4459 , \4460 );
xnor \U$4085 ( \4462 , \4461 , \1732 );
and \U$4086 ( \4463 , \4457 , \4462 );
and \U$4087 ( \4464 , \4453 , \4462 );
or \U$4088 ( \4465 , \4458 , \4463 , \4464 );
and \U$4089 ( \4466 , \4448 , \4465 );
and \U$4090 ( \4467 , \4432 , \4465 );
or \U$4091 ( \4468 , \4449 , \4466 , \4467 );
and \U$4092 ( \4469 , \2902 , \641 );
and \U$4093 ( \4470 , \2728 , \639 );
nor \U$4094 ( \4471 , \4469 , \4470 );
xnor \U$4095 ( \4472 , \4471 , \592 );
and \U$4096 ( \4473 , \3207 , \540 );
and \U$4097 ( \4474 , \3069 , \538 );
nor \U$4098 ( \4475 , \4473 , \4474 );
xnor \U$4099 ( \4476 , \4475 , \499 );
and \U$4100 ( \4477 , \4472 , \4476 );
and \U$4101 ( \4478 , \3743 , \470 );
and \U$4102 ( \4479 , \3326 , \468 );
nor \U$4103 ( \4480 , \4478 , \4479 );
xnor \U$4104 ( \4481 , \4480 , \440 );
and \U$4105 ( \4482 , \4476 , \4481 );
and \U$4106 ( \4483 , \4472 , \4481 );
or \U$4107 ( \4484 , \4477 , \4482 , \4483 );
and \U$4108 ( \4485 , \1441 , \1616 );
and \U$4109 ( \4486 , \1336 , \1614 );
nor \U$4110 ( \4487 , \4485 , \4486 );
xnor \U$4111 ( \4488 , \4487 , \1503 );
and \U$4112 ( \4489 , \1562 , \1422 );
and \U$4113 ( \4490 , \1446 , \1420 );
nor \U$4114 ( \4491 , \4489 , \4490 );
xnor \U$4115 ( \4492 , \4491 , \1286 );
and \U$4116 ( \4493 , \4488 , \4492 );
and \U$4117 ( \4494 , \1853 , \1222 );
and \U$4118 ( \4495 , \1677 , \1220 );
nor \U$4119 ( \4496 , \4494 , \4495 );
xnor \U$4120 ( \4497 , \4496 , \1144 );
and \U$4121 ( \4498 , \4492 , \4497 );
and \U$4122 ( \4499 , \4488 , \4497 );
or \U$4123 ( \4500 , \4493 , \4498 , \4499 );
and \U$4124 ( \4501 , \4484 , \4500 );
and \U$4125 ( \4502 , \2104 , \1058 );
and \U$4126 ( \4503 , \1861 , \1056 );
nor \U$4127 ( \4504 , \4502 , \4503 );
xnor \U$4128 ( \4505 , \4504 , \964 );
and \U$4129 ( \4506 , \2295 , \888 );
and \U$4130 ( \4507 , \2109 , \886 );
nor \U$4131 ( \4508 , \4506 , \4507 );
xnor \U$4132 ( \4509 , \4508 , \816 );
and \U$4133 ( \4510 , \4505 , \4509 );
and \U$4134 ( \4511 , \2703 , \754 );
and \U$4135 ( \4512 , \2439 , \752 );
nor \U$4136 ( \4513 , \4511 , \4512 );
xnor \U$4137 ( \4514 , \4513 , \711 );
and \U$4138 ( \4515 , \4509 , \4514 );
and \U$4139 ( \4516 , \4505 , \4514 );
or \U$4140 ( \4517 , \4510 , \4515 , \4516 );
and \U$4141 ( \4518 , \4500 , \4517 );
and \U$4142 ( \4519 , \4484 , \4517 );
or \U$4143 ( \4520 , \4501 , \4518 , \4519 );
and \U$4144 ( \4521 , \4468 , \4520 );
and \U$4145 ( \4522 , \4073 , \422 );
and \U$4146 ( \4523 , \3951 , \420 );
nor \U$4147 ( \4524 , \4522 , \4523 );
xnor \U$4148 ( \4525 , \4524 , \403 );
and \U$4149 ( \4526 , \4334 , \385 );
and \U$4150 ( \4527 , \4078 , \383 );
nor \U$4151 ( \4528 , \4526 , \4527 );
xnor \U$4152 ( \4529 , \4528 , \390 );
and \U$4153 ( \4530 , \4525 , \4529 );
buf \U$4154 ( \4531 , RIc224568_104);
and \U$4155 ( \4532 , \4531 , \379 );
and \U$4156 ( \4533 , \4529 , \4532 );
and \U$4157 ( \4534 , \4525 , \4532 );
or \U$4158 ( \4535 , \4530 , \4533 , \4534 );
xor \U$4159 ( \4536 , \4328 , \4332 );
xor \U$4160 ( \4537 , \4536 , \4335 );
and \U$4161 ( \4538 , \4535 , \4537 );
xor \U$4162 ( \4539 , \4254 , \4258 );
xor \U$4163 ( \4540 , \4539 , \4263 );
and \U$4164 ( \4541 , \4537 , \4540 );
and \U$4165 ( \4542 , \4535 , \4540 );
or \U$4166 ( \4543 , \4538 , \4541 , \4542 );
and \U$4167 ( \4544 , \4520 , \4543 );
and \U$4168 ( \4545 , \4468 , \4543 );
or \U$4169 ( \4546 , \4521 , \4544 , \4545 );
xor \U$4170 ( \4547 , \4233 , \4249 );
xor \U$4171 ( \4548 , \4547 , \4266 );
xor \U$4172 ( \4549 , \4287 , \4303 );
xor \U$4173 ( \4550 , \4549 , \4320 );
and \U$4174 ( \4551 , \4548 , \4550 );
xor \U$4175 ( \4552 , \4338 , \4340 );
xor \U$4176 ( \4553 , \4552 , \4342 );
and \U$4177 ( \4554 , \4550 , \4553 );
and \U$4178 ( \4555 , \4548 , \4553 );
or \U$4179 ( \4556 , \4551 , \4554 , \4555 );
and \U$4180 ( \4557 , \4546 , \4556 );
xor \U$4181 ( \4558 , \4221 , \4225 );
xor \U$4182 ( \4559 , \4558 , \4230 );
xor \U$4183 ( \4560 , \4237 , \4241 );
xor \U$4184 ( \4561 , \4560 , \4246 );
and \U$4185 ( \4562 , \4559 , \4561 );
xor \U$4186 ( \4563 , \4308 , \4312 );
xor \U$4187 ( \4564 , \4563 , \4317 );
and \U$4188 ( \4565 , \4561 , \4564 );
and \U$4189 ( \4566 , \4559 , \4564 );
or \U$4190 ( \4567 , \4562 , \4565 , \4566 );
xor \U$4191 ( \4568 , \4350 , \4352 );
xor \U$4192 ( \4569 , \4568 , \4355 );
and \U$4193 ( \4570 , \4567 , \4569 );
xor \U$4194 ( \4571 , \4360 , \4362 );
and \U$4195 ( \4572 , \4569 , \4571 );
and \U$4196 ( \4573 , \4567 , \4571 );
or \U$4197 ( \4574 , \4570 , \4572 , \4573 );
and \U$4198 ( \4575 , \4556 , \4574 );
and \U$4199 ( \4576 , \4546 , \4574 );
or \U$4200 ( \4577 , \4557 , \4575 , \4576 );
xor \U$4201 ( \4578 , \4109 , \4125 );
xor \U$4202 ( \4579 , \4578 , \4142 );
xor \U$4203 ( \4580 , \4358 , \4363 );
xor \U$4204 ( \4581 , \4580 , \4366 );
and \U$4205 ( \4582 , \4579 , \4581 );
xor \U$4206 ( \4583 , \4372 , \4374 );
xor \U$4207 ( \4584 , \4583 , \4377 );
and \U$4208 ( \4585 , \4581 , \4584 );
and \U$4209 ( \4586 , \4579 , \4584 );
or \U$4210 ( \4587 , \4582 , \4585 , \4586 );
and \U$4211 ( \4588 , \4577 , \4587 );
xor \U$4212 ( \4589 , \4158 , \4168 );
xor \U$4213 ( \4590 , \4589 , \4171 );
and \U$4214 ( \4591 , \4587 , \4590 );
and \U$4215 ( \4592 , \4577 , \4590 );
or \U$4216 ( \4593 , \4588 , \4591 , \4592 );
xor \U$4217 ( \4594 , \4072 , \4089 );
xor \U$4218 ( \4595 , \4594 , \4145 );
xor \U$4219 ( \4596 , \4348 , \4369 );
xor \U$4220 ( \4597 , \4596 , \4380 );
and \U$4221 ( \4598 , \4595 , \4597 );
xor \U$4222 ( \4599 , \4385 , \4387 );
xor \U$4223 ( \4600 , \4599 , \4390 );
and \U$4224 ( \4601 , \4597 , \4600 );
and \U$4225 ( \4602 , \4595 , \4600 );
or \U$4226 ( \4603 , \4598 , \4601 , \4602 );
and \U$4227 ( \4604 , \4593 , \4603 );
xor \U$4228 ( \4605 , \4148 , \4174 );
xor \U$4229 ( \4606 , \4605 , \4184 );
and \U$4230 ( \4607 , \4603 , \4606 );
and \U$4231 ( \4608 , \4593 , \4606 );
or \U$4232 ( \4609 , \4604 , \4607 , \4608 );
xor \U$4233 ( \4610 , \4399 , \4401 );
xor \U$4234 ( \4611 , \4610 , \4404 );
and \U$4235 ( \4612 , \4609 , \4611 );
and \U$4236 ( \4613 , \4413 , \4612 );
xor \U$4237 ( \4614 , \4413 , \4612 );
xor \U$4238 ( \4615 , \4609 , \4611 );
and \U$4239 ( \4616 , \771 , \2658 );
and \U$4240 ( \4617 , \743 , \2656 );
nor \U$4241 ( \4618 , \4616 , \4617 );
xnor \U$4242 ( \4619 , \4618 , \2516 );
and \U$4243 ( \4620 , \925 , \2362 );
and \U$4244 ( \4621 , \851 , \2360 );
nor \U$4245 ( \4622 , \4620 , \4621 );
xnor \U$4246 ( \4623 , \4622 , \2225 );
and \U$4247 ( \4624 , \4619 , \4623 );
and \U$4248 ( \4625 , \1050 , \2156 );
and \U$4249 ( \4626 , \987 , \2154 );
nor \U$4250 ( \4627 , \4625 , \4626 );
xnor \U$4251 ( \4628 , \4627 , \2004 );
and \U$4252 ( \4629 , \4623 , \4628 );
and \U$4253 ( \4630 , \4619 , \4628 );
or \U$4254 ( \4631 , \4624 , \4629 , \4630 );
buf \U$4255 ( \4632 , RIc226278_42);
buf \U$4256 ( \4633 , RIc226200_43);
and \U$4257 ( \4634 , \4632 , \4633 );
not \U$4258 ( \4635 , \4634 );
and \U$4259 ( \4636 , \4271 , \4635 );
not \U$4260 ( \4637 , \4636 );
and \U$4261 ( \4638 , \392 , \4417 );
and \U$4262 ( \4639 , \378 , \4415 );
nor \U$4263 ( \4640 , \4638 , \4639 );
xnor \U$4264 ( \4641 , \4640 , \4274 );
and \U$4265 ( \4642 , \4637 , \4641 );
and \U$4266 ( \4643 , \431 , \4094 );
and \U$4267 ( \4644 , \410 , \4092 );
nor \U$4268 ( \4645 , \4643 , \4644 );
xnor \U$4269 ( \4646 , \4645 , \3848 );
and \U$4270 ( \4647 , \4641 , \4646 );
and \U$4271 ( \4648 , \4637 , \4646 );
or \U$4272 ( \4649 , \4642 , \4647 , \4648 );
and \U$4273 ( \4650 , \4631 , \4649 );
and \U$4274 ( \4651 , \487 , \3699 );
and \U$4275 ( \4652 , \479 , \3697 );
nor \U$4276 ( \4653 , \4651 , \4652 );
xnor \U$4277 ( \4654 , \4653 , \3512 );
and \U$4278 ( \4655 , \561 , \3386 );
and \U$4279 ( \4656 , \556 , \3384 );
nor \U$4280 ( \4657 , \4655 , \4656 );
xnor \U$4281 ( \4658 , \4657 , \3181 );
and \U$4282 ( \4659 , \4654 , \4658 );
and \U$4283 ( \4660 , \666 , \2980 );
and \U$4284 ( \4661 , \615 , \2978 );
nor \U$4285 ( \4662 , \4660 , \4661 );
xnor \U$4286 ( \4663 , \4662 , \2831 );
and \U$4287 ( \4664 , \4658 , \4663 );
and \U$4288 ( \4665 , \4654 , \4663 );
or \U$4289 ( \4666 , \4659 , \4664 , \4665 );
and \U$4290 ( \4667 , \4649 , \4666 );
and \U$4291 ( \4668 , \4631 , \4666 );
or \U$4292 ( \4669 , \4650 , \4667 , \4668 );
and \U$4293 ( \4670 , \2728 , \754 );
and \U$4294 ( \4671 , \2703 , \752 );
nor \U$4295 ( \4672 , \4670 , \4671 );
xnor \U$4296 ( \4673 , \4672 , \711 );
and \U$4297 ( \4674 , \3069 , \641 );
and \U$4298 ( \4675 , \2902 , \639 );
nor \U$4299 ( \4676 , \4674 , \4675 );
xnor \U$4300 ( \4677 , \4676 , \592 );
and \U$4301 ( \4678 , \4673 , \4677 );
and \U$4302 ( \4679 , \3326 , \540 );
and \U$4303 ( \4680 , \3207 , \538 );
nor \U$4304 ( \4681 , \4679 , \4680 );
xnor \U$4305 ( \4682 , \4681 , \499 );
and \U$4306 ( \4683 , \4677 , \4682 );
and \U$4307 ( \4684 , \4673 , \4682 );
or \U$4308 ( \4685 , \4678 , \4683 , \4684 );
and \U$4309 ( \4686 , \1336 , \1888 );
and \U$4310 ( \4687 , \1248 , \1886 );
nor \U$4311 ( \4688 , \4686 , \4687 );
xnor \U$4312 ( \4689 , \4688 , \1732 );
and \U$4313 ( \4690 , \1446 , \1616 );
and \U$4314 ( \4691 , \1441 , \1614 );
nor \U$4315 ( \4692 , \4690 , \4691 );
xnor \U$4316 ( \4693 , \4692 , \1503 );
and \U$4317 ( \4694 , \4689 , \4693 );
and \U$4318 ( \4695 , \1677 , \1422 );
and \U$4319 ( \4696 , \1562 , \1420 );
nor \U$4320 ( \4697 , \4695 , \4696 );
xnor \U$4321 ( \4698 , \4697 , \1286 );
and \U$4322 ( \4699 , \4693 , \4698 );
and \U$4323 ( \4700 , \4689 , \4698 );
or \U$4324 ( \4701 , \4694 , \4699 , \4700 );
and \U$4325 ( \4702 , \4685 , \4701 );
and \U$4326 ( \4703 , \1861 , \1222 );
and \U$4327 ( \4704 , \1853 , \1220 );
nor \U$4328 ( \4705 , \4703 , \4704 );
xnor \U$4329 ( \4706 , \4705 , \1144 );
and \U$4330 ( \4707 , \2109 , \1058 );
and \U$4331 ( \4708 , \2104 , \1056 );
nor \U$4332 ( \4709 , \4707 , \4708 );
xnor \U$4333 ( \4710 , \4709 , \964 );
and \U$4334 ( \4711 , \4706 , \4710 );
and \U$4335 ( \4712 , \2439 , \888 );
and \U$4336 ( \4713 , \2295 , \886 );
nor \U$4337 ( \4714 , \4712 , \4713 );
xnor \U$4338 ( \4715 , \4714 , \816 );
and \U$4339 ( \4716 , \4710 , \4715 );
and \U$4340 ( \4717 , \4706 , \4715 );
or \U$4341 ( \4718 , \4711 , \4716 , \4717 );
and \U$4342 ( \4719 , \4701 , \4718 );
and \U$4343 ( \4720 , \4685 , \4718 );
or \U$4344 ( \4721 , \4702 , \4719 , \4720 );
and \U$4345 ( \4722 , \4669 , \4721 );
and \U$4346 ( \4723 , \3951 , \470 );
and \U$4347 ( \4724 , \3743 , \468 );
nor \U$4348 ( \4725 , \4723 , \4724 );
xnor \U$4349 ( \4726 , \4725 , \440 );
and \U$4350 ( \4727 , \4078 , \422 );
and \U$4351 ( \4728 , \4073 , \420 );
nor \U$4352 ( \4729 , \4727 , \4728 );
xnor \U$4353 ( \4730 , \4729 , \403 );
and \U$4354 ( \4731 , \4726 , \4730 );
and \U$4355 ( \4732 , \4531 , \385 );
and \U$4356 ( \4733 , \4334 , \383 );
nor \U$4357 ( \4734 , \4732 , \4733 );
xnor \U$4358 ( \4735 , \4734 , \390 );
and \U$4359 ( \4736 , \4730 , \4735 );
and \U$4360 ( \4737 , \4726 , \4735 );
or \U$4361 ( \4738 , \4731 , \4736 , \4737 );
xor \U$4362 ( \4739 , \4525 , \4529 );
xor \U$4363 ( \4740 , \4739 , \4532 );
or \U$4364 ( \4741 , \4738 , \4740 );
and \U$4365 ( \4742 , \4721 , \4741 );
and \U$4366 ( \4743 , \4669 , \4741 );
or \U$4367 ( \4744 , \4722 , \4742 , \4743 );
xor \U$4368 ( \4745 , \4472 , \4476 );
xor \U$4369 ( \4746 , \4745 , \4481 );
xor \U$4370 ( \4747 , \4488 , \4492 );
xor \U$4371 ( \4748 , \4747 , \4497 );
and \U$4372 ( \4749 , \4746 , \4748 );
xor \U$4373 ( \4750 , \4505 , \4509 );
xor \U$4374 ( \4751 , \4750 , \4514 );
and \U$4375 ( \4752 , \4748 , \4751 );
and \U$4376 ( \4753 , \4746 , \4751 );
or \U$4377 ( \4754 , \4749 , \4752 , \4753 );
xor \U$4378 ( \4755 , \4420 , \4424 );
xor \U$4379 ( \4756 , \4755 , \4429 );
xor \U$4380 ( \4757 , \4436 , \4440 );
xor \U$4381 ( \4758 , \4757 , \4445 );
and \U$4382 ( \4759 , \4756 , \4758 );
xor \U$4383 ( \4760 , \4453 , \4457 );
xor \U$4384 ( \4761 , \4760 , \4462 );
and \U$4385 ( \4762 , \4758 , \4761 );
and \U$4386 ( \4763 , \4756 , \4761 );
or \U$4387 ( \4764 , \4759 , \4762 , \4763 );
and \U$4388 ( \4765 , \4754 , \4764 );
xor \U$4389 ( \4766 , \4291 , \4295 );
xor \U$4390 ( \4767 , \4766 , \4300 );
and \U$4391 ( \4768 , \4764 , \4767 );
and \U$4392 ( \4769 , \4754 , \4767 );
or \U$4393 ( \4770 , \4765 , \4768 , \4769 );
and \U$4394 ( \4771 , \4744 , \4770 );
xor \U$4395 ( \4772 , \4275 , \4279 );
xor \U$4396 ( \4773 , \4772 , \4284 );
xor \U$4397 ( \4774 , \4559 , \4561 );
xor \U$4398 ( \4775 , \4774 , \4564 );
and \U$4399 ( \4776 , \4773 , \4775 );
xor \U$4400 ( \4777 , \4535 , \4537 );
xor \U$4401 ( \4778 , \4777 , \4540 );
and \U$4402 ( \4779 , \4775 , \4778 );
and \U$4403 ( \4780 , \4773 , \4778 );
or \U$4404 ( \4781 , \4776 , \4779 , \4780 );
and \U$4405 ( \4782 , \4770 , \4781 );
and \U$4406 ( \4783 , \4744 , \4781 );
or \U$4407 ( \4784 , \4771 , \4782 , \4783 );
xor \U$4408 ( \4785 , \4468 , \4520 );
xor \U$4409 ( \4786 , \4785 , \4543 );
xor \U$4410 ( \4787 , \4548 , \4550 );
xor \U$4411 ( \4788 , \4787 , \4553 );
and \U$4412 ( \4789 , \4786 , \4788 );
xor \U$4413 ( \4790 , \4567 , \4569 );
xor \U$4414 ( \4791 , \4790 , \4571 );
and \U$4415 ( \4792 , \4788 , \4791 );
and \U$4416 ( \4793 , \4786 , \4791 );
or \U$4417 ( \4794 , \4789 , \4792 , \4793 );
and \U$4418 ( \4795 , \4784 , \4794 );
xor \U$4419 ( \4796 , \4269 , \4323 );
xor \U$4420 ( \4797 , \4796 , \4345 );
and \U$4421 ( \4798 , \4794 , \4797 );
and \U$4422 ( \4799 , \4784 , \4797 );
or \U$4423 ( \4800 , \4795 , \4798 , \4799 );
xor \U$4424 ( \4801 , \4546 , \4556 );
xor \U$4425 ( \4802 , \4801 , \4574 );
xor \U$4426 ( \4803 , \4579 , \4581 );
xor \U$4427 ( \4804 , \4803 , \4584 );
and \U$4428 ( \4805 , \4802 , \4804 );
and \U$4429 ( \4806 , \4800 , \4805 );
xor \U$4430 ( \4807 , \4595 , \4597 );
xor \U$4431 ( \4808 , \4807 , \4600 );
and \U$4432 ( \4809 , \4805 , \4808 );
and \U$4433 ( \4810 , \4800 , \4808 );
or \U$4434 ( \4811 , \4806 , \4809 , \4810 );
xor \U$4435 ( \4812 , \4593 , \4603 );
xor \U$4436 ( \4813 , \4812 , \4606 );
and \U$4437 ( \4814 , \4811 , \4813 );
xor \U$4438 ( \4815 , \4383 , \4393 );
xor \U$4439 ( \4816 , \4815 , \4396 );
and \U$4440 ( \4817 , \4813 , \4816 );
and \U$4441 ( \4818 , \4811 , \4816 );
or \U$4442 ( \4819 , \4814 , \4817 , \4818 );
and \U$4443 ( \4820 , \4615 , \4819 );
xor \U$4444 ( \4821 , \4615 , \4819 );
xor \U$4445 ( \4822 , \4811 , \4813 );
xor \U$4446 ( \4823 , \4822 , \4816 );
and \U$4447 ( \4824 , \4073 , \470 );
and \U$4448 ( \4825 , \3951 , \468 );
nor \U$4449 ( \4826 , \4824 , \4825 );
xnor \U$4450 ( \4827 , \4826 , \440 );
and \U$4451 ( \4828 , \4334 , \422 );
and \U$4452 ( \4829 , \4078 , \420 );
nor \U$4453 ( \4830 , \4828 , \4829 );
xnor \U$4454 ( \4831 , \4830 , \403 );
and \U$4455 ( \4832 , \4827 , \4831 );
buf \U$4456 ( \4833 , RIc2244f0_105);
and \U$4457 ( \4834 , \4833 , \385 );
and \U$4458 ( \4835 , \4531 , \383 );
nor \U$4459 ( \4836 , \4834 , \4835 );
xnor \U$4460 ( \4837 , \4836 , \390 );
and \U$4461 ( \4838 , \4831 , \4837 );
and \U$4462 ( \4839 , \4827 , \4837 );
or \U$4463 ( \4840 , \4832 , \4838 , \4839 );
buf \U$4464 ( \4841 , RIc224478_106);
and \U$4465 ( \4842 , \4841 , \379 );
buf \U$4466 ( \4843 , \4842 );
and \U$4467 ( \4844 , \4840 , \4843 );
and \U$4468 ( \4845 , \4833 , \379 );
and \U$4469 ( \4846 , \4843 , \4845 );
and \U$4470 ( \4847 , \4840 , \4845 );
or \U$4471 ( \4848 , \4844 , \4846 , \4847 );
and \U$4472 ( \4849 , \851 , \2658 );
and \U$4473 ( \4850 , \771 , \2656 );
nor \U$4474 ( \4851 , \4849 , \4850 );
xnor \U$4475 ( \4852 , \4851 , \2516 );
and \U$4476 ( \4853 , \987 , \2362 );
and \U$4477 ( \4854 , \925 , \2360 );
nor \U$4478 ( \4855 , \4853 , \4854 );
xnor \U$4479 ( \4856 , \4855 , \2225 );
and \U$4480 ( \4857 , \4852 , \4856 );
and \U$4481 ( \4858 , \1248 , \2156 );
and \U$4482 ( \4859 , \1050 , \2154 );
nor \U$4483 ( \4860 , \4858 , \4859 );
xnor \U$4484 ( \4861 , \4860 , \2004 );
and \U$4485 ( \4862 , \4856 , \4861 );
and \U$4486 ( \4863 , \4852 , \4861 );
or \U$4487 ( \4864 , \4857 , \4862 , \4863 );
xor \U$4488 ( \4865 , \4271 , \4632 );
xor \U$4489 ( \4866 , \4632 , \4633 );
not \U$4490 ( \4867 , \4866 );
and \U$4491 ( \4868 , \4865 , \4867 );
and \U$4492 ( \4869 , \378 , \4868 );
not \U$4493 ( \4870 , \4869 );
xnor \U$4494 ( \4871 , \4870 , \4636 );
and \U$4495 ( \4872 , \410 , \4417 );
and \U$4496 ( \4873 , \392 , \4415 );
nor \U$4497 ( \4874 , \4872 , \4873 );
xnor \U$4498 ( \4875 , \4874 , \4274 );
and \U$4499 ( \4876 , \4871 , \4875 );
and \U$4500 ( \4877 , \479 , \4094 );
and \U$4501 ( \4878 , \431 , \4092 );
nor \U$4502 ( \4879 , \4877 , \4878 );
xnor \U$4503 ( \4880 , \4879 , \3848 );
and \U$4504 ( \4881 , \4875 , \4880 );
and \U$4505 ( \4882 , \4871 , \4880 );
or \U$4506 ( \4883 , \4876 , \4881 , \4882 );
and \U$4507 ( \4884 , \4864 , \4883 );
and \U$4508 ( \4885 , \556 , \3699 );
and \U$4509 ( \4886 , \487 , \3697 );
nor \U$4510 ( \4887 , \4885 , \4886 );
xnor \U$4511 ( \4888 , \4887 , \3512 );
and \U$4512 ( \4889 , \615 , \3386 );
and \U$4513 ( \4890 , \561 , \3384 );
nor \U$4514 ( \4891 , \4889 , \4890 );
xnor \U$4515 ( \4892 , \4891 , \3181 );
and \U$4516 ( \4893 , \4888 , \4892 );
and \U$4517 ( \4894 , \743 , \2980 );
and \U$4518 ( \4895 , \666 , \2978 );
nor \U$4519 ( \4896 , \4894 , \4895 );
xnor \U$4520 ( \4897 , \4896 , \2831 );
and \U$4521 ( \4898 , \4892 , \4897 );
and \U$4522 ( \4899 , \4888 , \4897 );
or \U$4523 ( \4900 , \4893 , \4898 , \4899 );
and \U$4524 ( \4901 , \4883 , \4900 );
and \U$4525 ( \4902 , \4864 , \4900 );
or \U$4526 ( \4903 , \4884 , \4901 , \4902 );
and \U$4527 ( \4904 , \4848 , \4903 );
and \U$4528 ( \4905 , \2902 , \754 );
and \U$4529 ( \4906 , \2728 , \752 );
nor \U$4530 ( \4907 , \4905 , \4906 );
xnor \U$4531 ( \4908 , \4907 , \711 );
and \U$4532 ( \4909 , \3207 , \641 );
and \U$4533 ( \4910 , \3069 , \639 );
nor \U$4534 ( \4911 , \4909 , \4910 );
xnor \U$4535 ( \4912 , \4911 , \592 );
and \U$4536 ( \4913 , \4908 , \4912 );
and \U$4537 ( \4914 , \3743 , \540 );
and \U$4538 ( \4915 , \3326 , \538 );
nor \U$4539 ( \4916 , \4914 , \4915 );
xnor \U$4540 ( \4917 , \4916 , \499 );
and \U$4541 ( \4918 , \4912 , \4917 );
and \U$4542 ( \4919 , \4908 , \4917 );
or \U$4543 ( \4920 , \4913 , \4918 , \4919 );
and \U$4544 ( \4921 , \2104 , \1222 );
and \U$4545 ( \4922 , \1861 , \1220 );
nor \U$4546 ( \4923 , \4921 , \4922 );
xnor \U$4547 ( \4924 , \4923 , \1144 );
and \U$4548 ( \4925 , \2295 , \1058 );
and \U$4549 ( \4926 , \2109 , \1056 );
nor \U$4550 ( \4927 , \4925 , \4926 );
xnor \U$4551 ( \4928 , \4927 , \964 );
and \U$4552 ( \4929 , \4924 , \4928 );
and \U$4553 ( \4930 , \2703 , \888 );
and \U$4554 ( \4931 , \2439 , \886 );
nor \U$4555 ( \4932 , \4930 , \4931 );
xnor \U$4556 ( \4933 , \4932 , \816 );
and \U$4557 ( \4934 , \4928 , \4933 );
and \U$4558 ( \4935 , \4924 , \4933 );
or \U$4559 ( \4936 , \4929 , \4934 , \4935 );
and \U$4560 ( \4937 , \4920 , \4936 );
and \U$4561 ( \4938 , \1441 , \1888 );
and \U$4562 ( \4939 , \1336 , \1886 );
nor \U$4563 ( \4940 , \4938 , \4939 );
xnor \U$4564 ( \4941 , \4940 , \1732 );
and \U$4565 ( \4942 , \1562 , \1616 );
and \U$4566 ( \4943 , \1446 , \1614 );
nor \U$4567 ( \4944 , \4942 , \4943 );
xnor \U$4568 ( \4945 , \4944 , \1503 );
and \U$4569 ( \4946 , \4941 , \4945 );
and \U$4570 ( \4947 , \1853 , \1422 );
and \U$4571 ( \4948 , \1677 , \1420 );
nor \U$4572 ( \4949 , \4947 , \4948 );
xnor \U$4573 ( \4950 , \4949 , \1286 );
and \U$4574 ( \4951 , \4945 , \4950 );
and \U$4575 ( \4952 , \4941 , \4950 );
or \U$4576 ( \4953 , \4946 , \4951 , \4952 );
and \U$4577 ( \4954 , \4936 , \4953 );
and \U$4578 ( \4955 , \4920 , \4953 );
or \U$4579 ( \4956 , \4937 , \4954 , \4955 );
and \U$4580 ( \4957 , \4903 , \4956 );
and \U$4581 ( \4958 , \4848 , \4956 );
or \U$4582 ( \4959 , \4904 , \4957 , \4958 );
xor \U$4583 ( \4960 , \4673 , \4677 );
xor \U$4584 ( \4961 , \4960 , \4682 );
xor \U$4585 ( \4962 , \4706 , \4710 );
xor \U$4586 ( \4963 , \4962 , \4715 );
and \U$4587 ( \4964 , \4961 , \4963 );
xor \U$4588 ( \4965 , \4726 , \4730 );
xor \U$4589 ( \4966 , \4965 , \4735 );
and \U$4590 ( \4967 , \4963 , \4966 );
and \U$4591 ( \4968 , \4961 , \4966 );
or \U$4592 ( \4969 , \4964 , \4967 , \4968 );
xor \U$4593 ( \4970 , \4619 , \4623 );
xor \U$4594 ( \4971 , \4970 , \4628 );
xor \U$4595 ( \4972 , \4689 , \4693 );
xor \U$4596 ( \4973 , \4972 , \4698 );
and \U$4597 ( \4974 , \4971 , \4973 );
xor \U$4598 ( \4975 , \4654 , \4658 );
xor \U$4599 ( \4976 , \4975 , \4663 );
and \U$4600 ( \4977 , \4973 , \4976 );
and \U$4601 ( \4978 , \4971 , \4976 );
or \U$4602 ( \4979 , \4974 , \4977 , \4978 );
and \U$4603 ( \4980 , \4969 , \4979 );
xor \U$4604 ( \4981 , \4756 , \4758 );
xor \U$4605 ( \4982 , \4981 , \4761 );
and \U$4606 ( \4983 , \4979 , \4982 );
and \U$4607 ( \4984 , \4969 , \4982 );
or \U$4608 ( \4985 , \4980 , \4983 , \4984 );
and \U$4609 ( \4986 , \4959 , \4985 );
xor \U$4610 ( \4987 , \4685 , \4701 );
xor \U$4611 ( \4988 , \4987 , \4718 );
xor \U$4612 ( \4989 , \4746 , \4748 );
xor \U$4613 ( \4990 , \4989 , \4751 );
and \U$4614 ( \4991 , \4988 , \4990 );
xnor \U$4615 ( \4992 , \4738 , \4740 );
and \U$4616 ( \4993 , \4990 , \4992 );
and \U$4617 ( \4994 , \4988 , \4992 );
or \U$4618 ( \4995 , \4991 , \4993 , \4994 );
and \U$4619 ( \4996 , \4985 , \4995 );
and \U$4620 ( \4997 , \4959 , \4995 );
or \U$4621 ( \4998 , \4986 , \4996 , \4997 );
xor \U$4622 ( \4999 , \4432 , \4448 );
xor \U$4623 ( \5000 , \4999 , \4465 );
xor \U$4624 ( \5001 , \4484 , \4500 );
xor \U$4625 ( \5002 , \5001 , \4517 );
and \U$4626 ( \5003 , \5000 , \5002 );
xor \U$4627 ( \5004 , \4773 , \4775 );
xor \U$4628 ( \5005 , \5004 , \4778 );
and \U$4629 ( \5006 , \5002 , \5005 );
and \U$4630 ( \5007 , \5000 , \5005 );
or \U$4631 ( \5008 , \5003 , \5006 , \5007 );
and \U$4632 ( \5009 , \4998 , \5008 );
xor \U$4633 ( \5010 , \4786 , \4788 );
xor \U$4634 ( \5011 , \5010 , \4791 );
and \U$4635 ( \5012 , \5008 , \5011 );
and \U$4636 ( \5013 , \4998 , \5011 );
or \U$4637 ( \5014 , \5009 , \5012 , \5013 );
xor \U$4638 ( \5015 , \4784 , \4794 );
xor \U$4639 ( \5016 , \5015 , \4797 );
and \U$4640 ( \5017 , \5014 , \5016 );
xor \U$4641 ( \5018 , \4802 , \4804 );
and \U$4642 ( \5019 , \5016 , \5018 );
and \U$4643 ( \5020 , \5014 , \5018 );
or \U$4644 ( \5021 , \5017 , \5019 , \5020 );
xor \U$4645 ( \5022 , \4577 , \4587 );
xor \U$4646 ( \5023 , \5022 , \4590 );
and \U$4647 ( \5024 , \5021 , \5023 );
xor \U$4648 ( \5025 , \4800 , \4805 );
xor \U$4649 ( \5026 , \5025 , \4808 );
and \U$4650 ( \5027 , \5023 , \5026 );
and \U$4651 ( \5028 , \5021 , \5026 );
or \U$4652 ( \5029 , \5024 , \5027 , \5028 );
and \U$4653 ( \5030 , \4823 , \5029 );
xor \U$4654 ( \5031 , \4823 , \5029 );
xor \U$4655 ( \5032 , \5021 , \5023 );
xor \U$4656 ( \5033 , \5032 , \5026 );
and \U$4657 ( \5034 , \771 , \2980 );
and \U$4658 ( \5035 , \743 , \2978 );
nor \U$4659 ( \5036 , \5034 , \5035 );
xnor \U$4660 ( \5037 , \5036 , \2831 );
and \U$4661 ( \5038 , \925 , \2658 );
and \U$4662 ( \5039 , \851 , \2656 );
nor \U$4663 ( \5040 , \5038 , \5039 );
xnor \U$4664 ( \5041 , \5040 , \2516 );
and \U$4665 ( \5042 , \5037 , \5041 );
and \U$4666 ( \5043 , \1050 , \2362 );
and \U$4667 ( \5044 , \987 , \2360 );
nor \U$4668 ( \5045 , \5043 , \5044 );
xnor \U$4669 ( \5046 , \5045 , \2225 );
and \U$4670 ( \5047 , \5041 , \5046 );
and \U$4671 ( \5048 , \5037 , \5046 );
or \U$4672 ( \5049 , \5042 , \5047 , \5048 );
buf \U$4673 ( \5050 , RIc226188_44);
buf \U$4674 ( \5051 , RIc226110_45);
and \U$4675 ( \5052 , \5050 , \5051 );
not \U$4676 ( \5053 , \5052 );
and \U$4677 ( \5054 , \4633 , \5053 );
not \U$4678 ( \5055 , \5054 );
and \U$4679 ( \5056 , \392 , \4868 );
and \U$4680 ( \5057 , \378 , \4866 );
nor \U$4681 ( \5058 , \5056 , \5057 );
xnor \U$4682 ( \5059 , \5058 , \4636 );
and \U$4683 ( \5060 , \5055 , \5059 );
and \U$4684 ( \5061 , \431 , \4417 );
and \U$4685 ( \5062 , \410 , \4415 );
nor \U$4686 ( \5063 , \5061 , \5062 );
xnor \U$4687 ( \5064 , \5063 , \4274 );
and \U$4688 ( \5065 , \5059 , \5064 );
and \U$4689 ( \5066 , \5055 , \5064 );
or \U$4690 ( \5067 , \5060 , \5065 , \5066 );
and \U$4691 ( \5068 , \5049 , \5067 );
and \U$4692 ( \5069 , \487 , \4094 );
and \U$4693 ( \5070 , \479 , \4092 );
nor \U$4694 ( \5071 , \5069 , \5070 );
xnor \U$4695 ( \5072 , \5071 , \3848 );
and \U$4696 ( \5073 , \561 , \3699 );
and \U$4697 ( \5074 , \556 , \3697 );
nor \U$4698 ( \5075 , \5073 , \5074 );
xnor \U$4699 ( \5076 , \5075 , \3512 );
and \U$4700 ( \5077 , \5072 , \5076 );
and \U$4701 ( \5078 , \666 , \3386 );
and \U$4702 ( \5079 , \615 , \3384 );
nor \U$4703 ( \5080 , \5078 , \5079 );
xnor \U$4704 ( \5081 , \5080 , \3181 );
and \U$4705 ( \5082 , \5076 , \5081 );
and \U$4706 ( \5083 , \5072 , \5081 );
or \U$4707 ( \5084 , \5077 , \5082 , \5083 );
and \U$4708 ( \5085 , \5067 , \5084 );
and \U$4709 ( \5086 , \5049 , \5084 );
or \U$4710 ( \5087 , \5068 , \5085 , \5086 );
and \U$4711 ( \5088 , \1336 , \2156 );
and \U$4712 ( \5089 , \1248 , \2154 );
nor \U$4713 ( \5090 , \5088 , \5089 );
xnor \U$4714 ( \5091 , \5090 , \2004 );
and \U$4715 ( \5092 , \1446 , \1888 );
and \U$4716 ( \5093 , \1441 , \1886 );
nor \U$4717 ( \5094 , \5092 , \5093 );
xnor \U$4718 ( \5095 , \5094 , \1732 );
and \U$4719 ( \5096 , \5091 , \5095 );
and \U$4720 ( \5097 , \1677 , \1616 );
and \U$4721 ( \5098 , \1562 , \1614 );
nor \U$4722 ( \5099 , \5097 , \5098 );
xnor \U$4723 ( \5100 , \5099 , \1503 );
and \U$4724 ( \5101 , \5095 , \5100 );
and \U$4725 ( \5102 , \5091 , \5100 );
or \U$4726 ( \5103 , \5096 , \5101 , \5102 );
and \U$4727 ( \5104 , \2728 , \888 );
and \U$4728 ( \5105 , \2703 , \886 );
nor \U$4729 ( \5106 , \5104 , \5105 );
xnor \U$4730 ( \5107 , \5106 , \816 );
and \U$4731 ( \5108 , \3069 , \754 );
and \U$4732 ( \5109 , \2902 , \752 );
nor \U$4733 ( \5110 , \5108 , \5109 );
xnor \U$4734 ( \5111 , \5110 , \711 );
and \U$4735 ( \5112 , \5107 , \5111 );
and \U$4736 ( \5113 , \3326 , \641 );
and \U$4737 ( \5114 , \3207 , \639 );
nor \U$4738 ( \5115 , \5113 , \5114 );
xnor \U$4739 ( \5116 , \5115 , \592 );
and \U$4740 ( \5117 , \5111 , \5116 );
and \U$4741 ( \5118 , \5107 , \5116 );
or \U$4742 ( \5119 , \5112 , \5117 , \5118 );
and \U$4743 ( \5120 , \5103 , \5119 );
and \U$4744 ( \5121 , \1861 , \1422 );
and \U$4745 ( \5122 , \1853 , \1420 );
nor \U$4746 ( \5123 , \5121 , \5122 );
xnor \U$4747 ( \5124 , \5123 , \1286 );
and \U$4748 ( \5125 , \2109 , \1222 );
and \U$4749 ( \5126 , \2104 , \1220 );
nor \U$4750 ( \5127 , \5125 , \5126 );
xnor \U$4751 ( \5128 , \5127 , \1144 );
and \U$4752 ( \5129 , \5124 , \5128 );
and \U$4753 ( \5130 , \2439 , \1058 );
and \U$4754 ( \5131 , \2295 , \1056 );
nor \U$4755 ( \5132 , \5130 , \5131 );
xnor \U$4756 ( \5133 , \5132 , \964 );
and \U$4757 ( \5134 , \5128 , \5133 );
and \U$4758 ( \5135 , \5124 , \5133 );
or \U$4759 ( \5136 , \5129 , \5134 , \5135 );
and \U$4760 ( \5137 , \5119 , \5136 );
and \U$4761 ( \5138 , \5103 , \5136 );
or \U$4762 ( \5139 , \5120 , \5137 , \5138 );
and \U$4763 ( \5140 , \5087 , \5139 );
and \U$4764 ( \5141 , \3951 , \540 );
and \U$4765 ( \5142 , \3743 , \538 );
nor \U$4766 ( \5143 , \5141 , \5142 );
xnor \U$4767 ( \5144 , \5143 , \499 );
and \U$4768 ( \5145 , \4078 , \470 );
and \U$4769 ( \5146 , \4073 , \468 );
nor \U$4770 ( \5147 , \5145 , \5146 );
xnor \U$4771 ( \5148 , \5147 , \440 );
and \U$4772 ( \5149 , \5144 , \5148 );
and \U$4773 ( \5150 , \4531 , \422 );
and \U$4774 ( \5151 , \4334 , \420 );
nor \U$4775 ( \5152 , \5150 , \5151 );
xnor \U$4776 ( \5153 , \5152 , \403 );
and \U$4777 ( \5154 , \5148 , \5153 );
and \U$4778 ( \5155 , \5144 , \5153 );
or \U$4779 ( \5156 , \5149 , \5154 , \5155 );
xor \U$4780 ( \5157 , \4827 , \4831 );
xor \U$4781 ( \5158 , \5157 , \4837 );
and \U$4782 ( \5159 , \5156 , \5158 );
not \U$4783 ( \5160 , \4842 );
and \U$4784 ( \5161 , \5158 , \5160 );
and \U$4785 ( \5162 , \5156 , \5160 );
or \U$4786 ( \5163 , \5159 , \5161 , \5162 );
and \U$4787 ( \5164 , \5139 , \5163 );
and \U$4788 ( \5165 , \5087 , \5163 );
or \U$4789 ( \5166 , \5140 , \5164 , \5165 );
xor \U$4790 ( \5167 , \4908 , \4912 );
xor \U$4791 ( \5168 , \5167 , \4917 );
xor \U$4792 ( \5169 , \4924 , \4928 );
xor \U$4793 ( \5170 , \5169 , \4933 );
and \U$4794 ( \5171 , \5168 , \5170 );
xor \U$4795 ( \5172 , \4941 , \4945 );
xor \U$4796 ( \5173 , \5172 , \4950 );
and \U$4797 ( \5174 , \5170 , \5173 );
and \U$4798 ( \5175 , \5168 , \5173 );
or \U$4799 ( \5176 , \5171 , \5174 , \5175 );
xor \U$4800 ( \5177 , \4852 , \4856 );
xor \U$4801 ( \5178 , \5177 , \4861 );
xor \U$4802 ( \5179 , \4871 , \4875 );
xor \U$4803 ( \5180 , \5179 , \4880 );
and \U$4804 ( \5181 , \5178 , \5180 );
xor \U$4805 ( \5182 , \4888 , \4892 );
xor \U$4806 ( \5183 , \5182 , \4897 );
and \U$4807 ( \5184 , \5180 , \5183 );
and \U$4808 ( \5185 , \5178 , \5183 );
or \U$4809 ( \5186 , \5181 , \5184 , \5185 );
and \U$4810 ( \5187 , \5176 , \5186 );
xor \U$4811 ( \5188 , \4637 , \4641 );
xor \U$4812 ( \5189 , \5188 , \4646 );
and \U$4813 ( \5190 , \5186 , \5189 );
and \U$4814 ( \5191 , \5176 , \5189 );
or \U$4815 ( \5192 , \5187 , \5190 , \5191 );
and \U$4816 ( \5193 , \5166 , \5192 );
xor \U$4817 ( \5194 , \4840 , \4843 );
xor \U$4818 ( \5195 , \5194 , \4845 );
xor \U$4819 ( \5196 , \4961 , \4963 );
xor \U$4820 ( \5197 , \5196 , \4966 );
and \U$4821 ( \5198 , \5195 , \5197 );
xor \U$4822 ( \5199 , \4971 , \4973 );
xor \U$4823 ( \5200 , \5199 , \4976 );
and \U$4824 ( \5201 , \5197 , \5200 );
and \U$4825 ( \5202 , \5195 , \5200 );
or \U$4826 ( \5203 , \5198 , \5201 , \5202 );
and \U$4827 ( \5204 , \5192 , \5203 );
and \U$4828 ( \5205 , \5166 , \5203 );
or \U$4829 ( \5206 , \5193 , \5204 , \5205 );
xor \U$4830 ( \5207 , \4631 , \4649 );
xor \U$4831 ( \5208 , \5207 , \4666 );
xor \U$4832 ( \5209 , \4969 , \4979 );
xor \U$4833 ( \5210 , \5209 , \4982 );
and \U$4834 ( \5211 , \5208 , \5210 );
xor \U$4835 ( \5212 , \4988 , \4990 );
xor \U$4836 ( \5213 , \5212 , \4992 );
and \U$4837 ( \5214 , \5210 , \5213 );
and \U$4838 ( \5215 , \5208 , \5213 );
or \U$4839 ( \5216 , \5211 , \5214 , \5215 );
and \U$4840 ( \5217 , \5206 , \5216 );
xor \U$4841 ( \5218 , \4754 , \4764 );
xor \U$4842 ( \5219 , \5218 , \4767 );
and \U$4843 ( \5220 , \5216 , \5219 );
and \U$4844 ( \5221 , \5206 , \5219 );
or \U$4845 ( \5222 , \5217 , \5220 , \5221 );
xor \U$4846 ( \5223 , \4669 , \4721 );
xor \U$4847 ( \5224 , \5223 , \4741 );
xor \U$4848 ( \5225 , \4959 , \4985 );
xor \U$4849 ( \5226 , \5225 , \4995 );
and \U$4850 ( \5227 , \5224 , \5226 );
xor \U$4851 ( \5228 , \5000 , \5002 );
xor \U$4852 ( \5229 , \5228 , \5005 );
and \U$4853 ( \5230 , \5226 , \5229 );
and \U$4854 ( \5231 , \5224 , \5229 );
or \U$4855 ( \5232 , \5227 , \5230 , \5231 );
and \U$4856 ( \5233 , \5222 , \5232 );
xor \U$4857 ( \5234 , \4744 , \4770 );
xor \U$4858 ( \5235 , \5234 , \4781 );
and \U$4859 ( \5236 , \5232 , \5235 );
and \U$4860 ( \5237 , \5222 , \5235 );
or \U$4861 ( \5238 , \5233 , \5236 , \5237 );
xor \U$4862 ( \5239 , \4633 , \5050 );
xor \U$4863 ( \5240 , \5050 , \5051 );
not \U$4864 ( \5241 , \5240 );
and \U$4865 ( \5242 , \5239 , \5241 );
and \U$4866 ( \5243 , \378 , \5242 );
not \U$4867 ( \5244 , \5243 );
xnor \U$4868 ( \5245 , \5244 , \5054 );
and \U$4869 ( \5246 , \410 , \4868 );
and \U$4870 ( \5247 , \392 , \4866 );
nor \U$4871 ( \5248 , \5246 , \5247 );
xnor \U$4872 ( \5249 , \5248 , \4636 );
and \U$4873 ( \5250 , \5245 , \5249 );
and \U$4874 ( \5251 , \479 , \4417 );
and \U$4875 ( \5252 , \431 , \4415 );
nor \U$4876 ( \5253 , \5251 , \5252 );
xnor \U$4877 ( \5254 , \5253 , \4274 );
and \U$4878 ( \5255 , \5249 , \5254 );
and \U$4879 ( \5256 , \5245 , \5254 );
or \U$4880 ( \5257 , \5250 , \5255 , \5256 );
and \U$4881 ( \5258 , \851 , \2980 );
and \U$4882 ( \5259 , \771 , \2978 );
nor \U$4883 ( \5260 , \5258 , \5259 );
xnor \U$4884 ( \5261 , \5260 , \2831 );
and \U$4885 ( \5262 , \987 , \2658 );
and \U$4886 ( \5263 , \925 , \2656 );
nor \U$4887 ( \5264 , \5262 , \5263 );
xnor \U$4888 ( \5265 , \5264 , \2516 );
and \U$4889 ( \5266 , \5261 , \5265 );
and \U$4890 ( \5267 , \1248 , \2362 );
and \U$4891 ( \5268 , \1050 , \2360 );
nor \U$4892 ( \5269 , \5267 , \5268 );
xnor \U$4893 ( \5270 , \5269 , \2225 );
and \U$4894 ( \5271 , \5265 , \5270 );
and \U$4895 ( \5272 , \5261 , \5270 );
or \U$4896 ( \5273 , \5266 , \5271 , \5272 );
and \U$4897 ( \5274 , \5257 , \5273 );
and \U$4898 ( \5275 , \556 , \4094 );
and \U$4899 ( \5276 , \487 , \4092 );
nor \U$4900 ( \5277 , \5275 , \5276 );
xnor \U$4901 ( \5278 , \5277 , \3848 );
and \U$4902 ( \5279 , \615 , \3699 );
and \U$4903 ( \5280 , \561 , \3697 );
nor \U$4904 ( \5281 , \5279 , \5280 );
xnor \U$4905 ( \5282 , \5281 , \3512 );
and \U$4906 ( \5283 , \5278 , \5282 );
and \U$4907 ( \5284 , \743 , \3386 );
and \U$4908 ( \5285 , \666 , \3384 );
nor \U$4909 ( \5286 , \5284 , \5285 );
xnor \U$4910 ( \5287 , \5286 , \3181 );
and \U$4911 ( \5288 , \5282 , \5287 );
and \U$4912 ( \5289 , \5278 , \5287 );
or \U$4913 ( \5290 , \5283 , \5288 , \5289 );
and \U$4914 ( \5291 , \5273 , \5290 );
and \U$4915 ( \5292 , \5257 , \5290 );
or \U$4916 ( \5293 , \5274 , \5291 , \5292 );
and \U$4917 ( \5294 , \4073 , \540 );
and \U$4918 ( \5295 , \3951 , \538 );
nor \U$4919 ( \5296 , \5294 , \5295 );
xnor \U$4920 ( \5297 , \5296 , \499 );
and \U$4921 ( \5298 , \4334 , \470 );
and \U$4922 ( \5299 , \4078 , \468 );
nor \U$4923 ( \5300 , \5298 , \5299 );
xnor \U$4924 ( \5301 , \5300 , \440 );
and \U$4925 ( \5302 , \5297 , \5301 );
and \U$4926 ( \5303 , \4833 , \422 );
and \U$4927 ( \5304 , \4531 , \420 );
nor \U$4928 ( \5305 , \5303 , \5304 );
xnor \U$4929 ( \5306 , \5305 , \403 );
and \U$4930 ( \5307 , \5301 , \5306 );
and \U$4931 ( \5308 , \5297 , \5306 );
or \U$4932 ( \5309 , \5302 , \5307 , \5308 );
buf \U$4933 ( \5310 , RIc224400_107);
and \U$4934 ( \5311 , \5310 , \385 );
and \U$4935 ( \5312 , \4841 , \383 );
nor \U$4936 ( \5313 , \5311 , \5312 );
xnor \U$4937 ( \5314 , \5313 , \390 );
buf \U$4938 ( \5315 , RIc224388_108);
and \U$4939 ( \5316 , \5315 , \379 );
or \U$4940 ( \5317 , \5314 , \5316 );
and \U$4941 ( \5318 , \5309 , \5317 );
and \U$4942 ( \5319 , \4841 , \385 );
and \U$4943 ( \5320 , \4833 , \383 );
nor \U$4944 ( \5321 , \5319 , \5320 );
xnor \U$4945 ( \5322 , \5321 , \390 );
and \U$4946 ( \5323 , \5317 , \5322 );
and \U$4947 ( \5324 , \5309 , \5322 );
or \U$4948 ( \5325 , \5318 , \5323 , \5324 );
and \U$4949 ( \5326 , \5293 , \5325 );
and \U$4950 ( \5327 , \1441 , \2156 );
and \U$4951 ( \5328 , \1336 , \2154 );
nor \U$4952 ( \5329 , \5327 , \5328 );
xnor \U$4953 ( \5330 , \5329 , \2004 );
and \U$4954 ( \5331 , \1562 , \1888 );
and \U$4955 ( \5332 , \1446 , \1886 );
nor \U$4956 ( \5333 , \5331 , \5332 );
xnor \U$4957 ( \5334 , \5333 , \1732 );
and \U$4958 ( \5335 , \5330 , \5334 );
and \U$4959 ( \5336 , \1853 , \1616 );
and \U$4960 ( \5337 , \1677 , \1614 );
nor \U$4961 ( \5338 , \5336 , \5337 );
xnor \U$4962 ( \5339 , \5338 , \1503 );
and \U$4963 ( \5340 , \5334 , \5339 );
and \U$4964 ( \5341 , \5330 , \5339 );
or \U$4965 ( \5342 , \5335 , \5340 , \5341 );
and \U$4966 ( \5343 , \2104 , \1422 );
and \U$4967 ( \5344 , \1861 , \1420 );
nor \U$4968 ( \5345 , \5343 , \5344 );
xnor \U$4969 ( \5346 , \5345 , \1286 );
and \U$4970 ( \5347 , \2295 , \1222 );
and \U$4971 ( \5348 , \2109 , \1220 );
nor \U$4972 ( \5349 , \5347 , \5348 );
xnor \U$4973 ( \5350 , \5349 , \1144 );
and \U$4974 ( \5351 , \5346 , \5350 );
and \U$4975 ( \5352 , \2703 , \1058 );
and \U$4976 ( \5353 , \2439 , \1056 );
nor \U$4977 ( \5354 , \5352 , \5353 );
xnor \U$4978 ( \5355 , \5354 , \964 );
and \U$4979 ( \5356 , \5350 , \5355 );
and \U$4980 ( \5357 , \5346 , \5355 );
or \U$4981 ( \5358 , \5351 , \5356 , \5357 );
and \U$4982 ( \5359 , \5342 , \5358 );
and \U$4983 ( \5360 , \2902 , \888 );
and \U$4984 ( \5361 , \2728 , \886 );
nor \U$4985 ( \5362 , \5360 , \5361 );
xnor \U$4986 ( \5363 , \5362 , \816 );
and \U$4987 ( \5364 , \3207 , \754 );
and \U$4988 ( \5365 , \3069 , \752 );
nor \U$4989 ( \5366 , \5364 , \5365 );
xnor \U$4990 ( \5367 , \5366 , \711 );
and \U$4991 ( \5368 , \5363 , \5367 );
and \U$4992 ( \5369 , \3743 , \641 );
and \U$4993 ( \5370 , \3326 , \639 );
nor \U$4994 ( \5371 , \5369 , \5370 );
xnor \U$4995 ( \5372 , \5371 , \592 );
and \U$4996 ( \5373 , \5367 , \5372 );
and \U$4997 ( \5374 , \5363 , \5372 );
or \U$4998 ( \5375 , \5368 , \5373 , \5374 );
and \U$4999 ( \5376 , \5358 , \5375 );
and \U$5000 ( \5377 , \5342 , \5375 );
or \U$5001 ( \5378 , \5359 , \5376 , \5377 );
and \U$5002 ( \5379 , \5325 , \5378 );
and \U$5003 ( \5380 , \5293 , \5378 );
or \U$5004 ( \5381 , \5326 , \5379 , \5380 );
and \U$5005 ( \5382 , \5310 , \379 );
xor \U$5006 ( \5383 , \5144 , \5148 );
xor \U$5007 ( \5384 , \5383 , \5153 );
and \U$5008 ( \5385 , \5382 , \5384 );
xor \U$5009 ( \5386 , \5107 , \5111 );
xor \U$5010 ( \5387 , \5386 , \5116 );
and \U$5011 ( \5388 , \5384 , \5387 );
and \U$5012 ( \5389 , \5382 , \5387 );
or \U$5013 ( \5390 , \5385 , \5388 , \5389 );
xor \U$5014 ( \5391 , \5091 , \5095 );
xor \U$5015 ( \5392 , \5391 , \5100 );
xor \U$5016 ( \5393 , \5037 , \5041 );
xor \U$5017 ( \5394 , \5393 , \5046 );
and \U$5018 ( \5395 , \5392 , \5394 );
xor \U$5019 ( \5396 , \5124 , \5128 );
xor \U$5020 ( \5397 , \5396 , \5133 );
and \U$5021 ( \5398 , \5394 , \5397 );
and \U$5022 ( \5399 , \5392 , \5397 );
or \U$5023 ( \5400 , \5395 , \5398 , \5399 );
and \U$5024 ( \5401 , \5390 , \5400 );
xor \U$5025 ( \5402 , \5178 , \5180 );
xor \U$5026 ( \5403 , \5402 , \5183 );
and \U$5027 ( \5404 , \5400 , \5403 );
and \U$5028 ( \5405 , \5390 , \5403 );
or \U$5029 ( \5406 , \5401 , \5404 , \5405 );
and \U$5030 ( \5407 , \5381 , \5406 );
xor \U$5031 ( \5408 , \5103 , \5119 );
xor \U$5032 ( \5409 , \5408 , \5136 );
xor \U$5033 ( \5410 , \5168 , \5170 );
xor \U$5034 ( \5411 , \5410 , \5173 );
and \U$5035 ( \5412 , \5409 , \5411 );
xor \U$5036 ( \5413 , \5156 , \5158 );
xor \U$5037 ( \5414 , \5413 , \5160 );
and \U$5038 ( \5415 , \5411 , \5414 );
and \U$5039 ( \5416 , \5409 , \5414 );
or \U$5040 ( \5417 , \5412 , \5415 , \5416 );
and \U$5041 ( \5418 , \5406 , \5417 );
and \U$5042 ( \5419 , \5381 , \5417 );
or \U$5043 ( \5420 , \5407 , \5418 , \5419 );
xor \U$5044 ( \5421 , \4864 , \4883 );
xor \U$5045 ( \5422 , \5421 , \4900 );
xor \U$5046 ( \5423 , \4920 , \4936 );
xor \U$5047 ( \5424 , \5423 , \4953 );
and \U$5048 ( \5425 , \5422 , \5424 );
xor \U$5049 ( \5426 , \5195 , \5197 );
xor \U$5050 ( \5427 , \5426 , \5200 );
and \U$5051 ( \5428 , \5424 , \5427 );
and \U$5052 ( \5429 , \5422 , \5427 );
or \U$5053 ( \5430 , \5425 , \5428 , \5429 );
and \U$5054 ( \5431 , \5420 , \5430 );
xor \U$5055 ( \5432 , \4848 , \4903 );
xor \U$5056 ( \5433 , \5432 , \4956 );
and \U$5057 ( \5434 , \5430 , \5433 );
and \U$5058 ( \5435 , \5420 , \5433 );
or \U$5059 ( \5436 , \5431 , \5434 , \5435 );
xor \U$5060 ( \5437 , \5206 , \5216 );
xor \U$5061 ( \5438 , \5437 , \5219 );
and \U$5062 ( \5439 , \5436 , \5438 );
xor \U$5063 ( \5440 , \5224 , \5226 );
xor \U$5064 ( \5441 , \5440 , \5229 );
and \U$5065 ( \5442 , \5438 , \5441 );
and \U$5066 ( \5443 , \5436 , \5441 );
or \U$5067 ( \5444 , \5439 , \5442 , \5443 );
xor \U$5068 ( \5445 , \5222 , \5232 );
xor \U$5069 ( \5446 , \5445 , \5235 );
and \U$5070 ( \5447 , \5444 , \5446 );
xor \U$5071 ( \5448 , \4998 , \5008 );
xor \U$5072 ( \5449 , \5448 , \5011 );
and \U$5073 ( \5450 , \5446 , \5449 );
and \U$5074 ( \5451 , \5444 , \5449 );
or \U$5075 ( \5452 , \5447 , \5450 , \5451 );
and \U$5076 ( \5453 , \5238 , \5452 );
xor \U$5077 ( \5454 , \5014 , \5016 );
xor \U$5078 ( \5455 , \5454 , \5018 );
and \U$5079 ( \5456 , \5452 , \5455 );
and \U$5080 ( \5457 , \5238 , \5455 );
or \U$5081 ( \5458 , \5453 , \5456 , \5457 );
and \U$5082 ( \5459 , \5033 , \5458 );
xor \U$5083 ( \5460 , \5033 , \5458 );
xor \U$5084 ( \5461 , \5238 , \5452 );
xor \U$5085 ( \5462 , \5461 , \5455 );
buf \U$5086 ( \5463 , RIc226098_46);
buf \U$5087 ( \5464 , RIc226020_47);
and \U$5088 ( \5465 , \5463 , \5464 );
not \U$5089 ( \5466 , \5465 );
and \U$5090 ( \5467 , \5051 , \5466 );
not \U$5091 ( \5468 , \5467 );
and \U$5092 ( \5469 , \392 , \5242 );
and \U$5093 ( \5470 , \378 , \5240 );
nor \U$5094 ( \5471 , \5469 , \5470 );
xnor \U$5095 ( \5472 , \5471 , \5054 );
and \U$5096 ( \5473 , \5468 , \5472 );
and \U$5097 ( \5474 , \431 , \4868 );
and \U$5098 ( \5475 , \410 , \4866 );
nor \U$5099 ( \5476 , \5474 , \5475 );
xnor \U$5100 ( \5477 , \5476 , \4636 );
and \U$5101 ( \5478 , \5472 , \5477 );
and \U$5102 ( \5479 , \5468 , \5477 );
or \U$5103 ( \5480 , \5473 , \5478 , \5479 );
and \U$5104 ( \5481 , \487 , \4417 );
and \U$5105 ( \5482 , \479 , \4415 );
nor \U$5106 ( \5483 , \5481 , \5482 );
xnor \U$5107 ( \5484 , \5483 , \4274 );
and \U$5108 ( \5485 , \561 , \4094 );
and \U$5109 ( \5486 , \556 , \4092 );
nor \U$5110 ( \5487 , \5485 , \5486 );
xnor \U$5111 ( \5488 , \5487 , \3848 );
and \U$5112 ( \5489 , \5484 , \5488 );
and \U$5113 ( \5490 , \666 , \3699 );
and \U$5114 ( \5491 , \615 , \3697 );
nor \U$5115 ( \5492 , \5490 , \5491 );
xnor \U$5116 ( \5493 , \5492 , \3512 );
and \U$5117 ( \5494 , \5488 , \5493 );
and \U$5118 ( \5495 , \5484 , \5493 );
or \U$5119 ( \5496 , \5489 , \5494 , \5495 );
and \U$5120 ( \5497 , \5480 , \5496 );
and \U$5121 ( \5498 , \771 , \3386 );
and \U$5122 ( \5499 , \743 , \3384 );
nor \U$5123 ( \5500 , \5498 , \5499 );
xnor \U$5124 ( \5501 , \5500 , \3181 );
and \U$5125 ( \5502 , \925 , \2980 );
and \U$5126 ( \5503 , \851 , \2978 );
nor \U$5127 ( \5504 , \5502 , \5503 );
xnor \U$5128 ( \5505 , \5504 , \2831 );
and \U$5129 ( \5506 , \5501 , \5505 );
and \U$5130 ( \5507 , \1050 , \2658 );
and \U$5131 ( \5508 , \987 , \2656 );
nor \U$5132 ( \5509 , \5507 , \5508 );
xnor \U$5133 ( \5510 , \5509 , \2516 );
and \U$5134 ( \5511 , \5505 , \5510 );
and \U$5135 ( \5512 , \5501 , \5510 );
or \U$5136 ( \5513 , \5506 , \5511 , \5512 );
and \U$5137 ( \5514 , \5496 , \5513 );
and \U$5138 ( \5515 , \5480 , \5513 );
or \U$5139 ( \5516 , \5497 , \5514 , \5515 );
and \U$5140 ( \5517 , \1336 , \2362 );
and \U$5141 ( \5518 , \1248 , \2360 );
nor \U$5142 ( \5519 , \5517 , \5518 );
xnor \U$5143 ( \5520 , \5519 , \2225 );
and \U$5144 ( \5521 , \1446 , \2156 );
and \U$5145 ( \5522 , \1441 , \2154 );
nor \U$5146 ( \5523 , \5521 , \5522 );
xnor \U$5147 ( \5524 , \5523 , \2004 );
and \U$5148 ( \5525 , \5520 , \5524 );
and \U$5149 ( \5526 , \1677 , \1888 );
and \U$5150 ( \5527 , \1562 , \1886 );
nor \U$5151 ( \5528 , \5526 , \5527 );
xnor \U$5152 ( \5529 , \5528 , \1732 );
and \U$5153 ( \5530 , \5524 , \5529 );
and \U$5154 ( \5531 , \5520 , \5529 );
or \U$5155 ( \5532 , \5525 , \5530 , \5531 );
and \U$5156 ( \5533 , \1861 , \1616 );
and \U$5157 ( \5534 , \1853 , \1614 );
nor \U$5158 ( \5535 , \5533 , \5534 );
xnor \U$5159 ( \5536 , \5535 , \1503 );
and \U$5160 ( \5537 , \2109 , \1422 );
and \U$5161 ( \5538 , \2104 , \1420 );
nor \U$5162 ( \5539 , \5537 , \5538 );
xnor \U$5163 ( \5540 , \5539 , \1286 );
and \U$5164 ( \5541 , \5536 , \5540 );
and \U$5165 ( \5542 , \2439 , \1222 );
and \U$5166 ( \5543 , \2295 , \1220 );
nor \U$5167 ( \5544 , \5542 , \5543 );
xnor \U$5168 ( \5545 , \5544 , \1144 );
and \U$5169 ( \5546 , \5540 , \5545 );
and \U$5170 ( \5547 , \5536 , \5545 );
or \U$5171 ( \5548 , \5541 , \5546 , \5547 );
and \U$5172 ( \5549 , \5532 , \5548 );
and \U$5173 ( \5550 , \2728 , \1058 );
and \U$5174 ( \5551 , \2703 , \1056 );
nor \U$5175 ( \5552 , \5550 , \5551 );
xnor \U$5176 ( \5553 , \5552 , \964 );
and \U$5177 ( \5554 , \3069 , \888 );
and \U$5178 ( \5555 , \2902 , \886 );
nor \U$5179 ( \5556 , \5554 , \5555 );
xnor \U$5180 ( \5557 , \5556 , \816 );
and \U$5181 ( \5558 , \5553 , \5557 );
and \U$5182 ( \5559 , \3326 , \754 );
and \U$5183 ( \5560 , \3207 , \752 );
nor \U$5184 ( \5561 , \5559 , \5560 );
xnor \U$5185 ( \5562 , \5561 , \711 );
and \U$5186 ( \5563 , \5557 , \5562 );
and \U$5187 ( \5564 , \5553 , \5562 );
or \U$5188 ( \5565 , \5558 , \5563 , \5564 );
and \U$5189 ( \5566 , \5548 , \5565 );
and \U$5190 ( \5567 , \5532 , \5565 );
or \U$5191 ( \5568 , \5549 , \5566 , \5567 );
and \U$5192 ( \5569 , \5516 , \5568 );
and \U$5193 ( \5570 , \4841 , \422 );
and \U$5194 ( \5571 , \4833 , \420 );
nor \U$5195 ( \5572 , \5570 , \5571 );
xnor \U$5196 ( \5573 , \5572 , \403 );
and \U$5197 ( \5574 , \5315 , \385 );
and \U$5198 ( \5575 , \5310 , \383 );
nor \U$5199 ( \5576 , \5574 , \5575 );
xnor \U$5200 ( \5577 , \5576 , \390 );
and \U$5201 ( \5578 , \5573 , \5577 );
buf \U$5202 ( \5579 , RIc224310_109);
and \U$5203 ( \5580 , \5579 , \379 );
and \U$5204 ( \5581 , \5577 , \5580 );
and \U$5205 ( \5582 , \5573 , \5580 );
or \U$5206 ( \5583 , \5578 , \5581 , \5582 );
and \U$5207 ( \5584 , \3951 , \641 );
and \U$5208 ( \5585 , \3743 , \639 );
nor \U$5209 ( \5586 , \5584 , \5585 );
xnor \U$5210 ( \5587 , \5586 , \592 );
and \U$5211 ( \5588 , \4078 , \540 );
and \U$5212 ( \5589 , \4073 , \538 );
nor \U$5213 ( \5590 , \5588 , \5589 );
xnor \U$5214 ( \5591 , \5590 , \499 );
and \U$5215 ( \5592 , \5587 , \5591 );
and \U$5216 ( \5593 , \4531 , \470 );
and \U$5217 ( \5594 , \4334 , \468 );
nor \U$5218 ( \5595 , \5593 , \5594 );
xnor \U$5219 ( \5596 , \5595 , \440 );
and \U$5220 ( \5597 , \5591 , \5596 );
and \U$5221 ( \5598 , \5587 , \5596 );
or \U$5222 ( \5599 , \5592 , \5597 , \5598 );
and \U$5223 ( \5600 , \5583 , \5599 );
xnor \U$5224 ( \5601 , \5314 , \5316 );
and \U$5225 ( \5602 , \5599 , \5601 );
and \U$5226 ( \5603 , \5583 , \5601 );
or \U$5227 ( \5604 , \5600 , \5602 , \5603 );
and \U$5228 ( \5605 , \5568 , \5604 );
and \U$5229 ( \5606 , \5516 , \5604 );
or \U$5230 ( \5607 , \5569 , \5605 , \5606 );
xor \U$5231 ( \5608 , \5297 , \5301 );
xor \U$5232 ( \5609 , \5608 , \5306 );
xor \U$5233 ( \5610 , \5346 , \5350 );
xor \U$5234 ( \5611 , \5610 , \5355 );
and \U$5235 ( \5612 , \5609 , \5611 );
xor \U$5236 ( \5613 , \5363 , \5367 );
xor \U$5237 ( \5614 , \5613 , \5372 );
and \U$5238 ( \5615 , \5611 , \5614 );
and \U$5239 ( \5616 , \5609 , \5614 );
or \U$5240 ( \5617 , \5612 , \5615 , \5616 );
xor \U$5241 ( \5618 , \5330 , \5334 );
xor \U$5242 ( \5619 , \5618 , \5339 );
xor \U$5243 ( \5620 , \5261 , \5265 );
xor \U$5244 ( \5621 , \5620 , \5270 );
and \U$5245 ( \5622 , \5619 , \5621 );
xor \U$5246 ( \5623 , \5278 , \5282 );
xor \U$5247 ( \5624 , \5623 , \5287 );
and \U$5248 ( \5625 , \5621 , \5624 );
and \U$5249 ( \5626 , \5619 , \5624 );
or \U$5250 ( \5627 , \5622 , \5625 , \5626 );
and \U$5251 ( \5628 , \5617 , \5627 );
xor \U$5252 ( \5629 , \5072 , \5076 );
xor \U$5253 ( \5630 , \5629 , \5081 );
and \U$5254 ( \5631 , \5627 , \5630 );
and \U$5255 ( \5632 , \5617 , \5630 );
or \U$5256 ( \5633 , \5628 , \5631 , \5632 );
and \U$5257 ( \5634 , \5607 , \5633 );
xor \U$5258 ( \5635 , \5055 , \5059 );
xor \U$5259 ( \5636 , \5635 , \5064 );
xor \U$5260 ( \5637 , \5382 , \5384 );
xor \U$5261 ( \5638 , \5637 , \5387 );
and \U$5262 ( \5639 , \5636 , \5638 );
xor \U$5263 ( \5640 , \5392 , \5394 );
xor \U$5264 ( \5641 , \5640 , \5397 );
and \U$5265 ( \5642 , \5638 , \5641 );
and \U$5266 ( \5643 , \5636 , \5641 );
or \U$5267 ( \5644 , \5639 , \5642 , \5643 );
and \U$5268 ( \5645 , \5633 , \5644 );
and \U$5269 ( \5646 , \5607 , \5644 );
or \U$5270 ( \5647 , \5634 , \5645 , \5646 );
xor \U$5271 ( \5648 , \5257 , \5273 );
xor \U$5272 ( \5649 , \5648 , \5290 );
xor \U$5273 ( \5650 , \5309 , \5317 );
xor \U$5274 ( \5651 , \5650 , \5322 );
and \U$5275 ( \5652 , \5649 , \5651 );
xor \U$5276 ( \5653 , \5342 , \5358 );
xor \U$5277 ( \5654 , \5653 , \5375 );
and \U$5278 ( \5655 , \5651 , \5654 );
and \U$5279 ( \5656 , \5649 , \5654 );
or \U$5280 ( \5657 , \5652 , \5655 , \5656 );
xor \U$5281 ( \5658 , \5049 , \5067 );
xor \U$5282 ( \5659 , \5658 , \5084 );
and \U$5283 ( \5660 , \5657 , \5659 );
xor \U$5284 ( \5661 , \5409 , \5411 );
xor \U$5285 ( \5662 , \5661 , \5414 );
and \U$5286 ( \5663 , \5659 , \5662 );
and \U$5287 ( \5664 , \5657 , \5662 );
or \U$5288 ( \5665 , \5660 , \5663 , \5664 );
and \U$5289 ( \5666 , \5647 , \5665 );
xor \U$5290 ( \5667 , \5176 , \5186 );
xor \U$5291 ( \5668 , \5667 , \5189 );
and \U$5292 ( \5669 , \5665 , \5668 );
and \U$5293 ( \5670 , \5647 , \5668 );
or \U$5294 ( \5671 , \5666 , \5669 , \5670 );
xor \U$5295 ( \5672 , \5087 , \5139 );
xor \U$5296 ( \5673 , \5672 , \5163 );
xor \U$5297 ( \5674 , \5381 , \5406 );
xor \U$5298 ( \5675 , \5674 , \5417 );
and \U$5299 ( \5676 , \5673 , \5675 );
xor \U$5300 ( \5677 , \5422 , \5424 );
xor \U$5301 ( \5678 , \5677 , \5427 );
and \U$5302 ( \5679 , \5675 , \5678 );
and \U$5303 ( \5680 , \5673 , \5678 );
or \U$5304 ( \5681 , \5676 , \5679 , \5680 );
and \U$5305 ( \5682 , \5671 , \5681 );
xor \U$5306 ( \5683 , \5208 , \5210 );
xor \U$5307 ( \5684 , \5683 , \5213 );
and \U$5308 ( \5685 , \5681 , \5684 );
and \U$5309 ( \5686 , \5671 , \5684 );
or \U$5310 ( \5687 , \5682 , \5685 , \5686 );
xor \U$5311 ( \5688 , \5166 , \5192 );
xor \U$5312 ( \5689 , \5688 , \5203 );
xor \U$5313 ( \5690 , \5420 , \5430 );
xor \U$5314 ( \5691 , \5690 , \5433 );
and \U$5315 ( \5692 , \5689 , \5691 );
and \U$5316 ( \5693 , \5687 , \5692 );
xor \U$5317 ( \5694 , \5436 , \5438 );
xor \U$5318 ( \5695 , \5694 , \5441 );
and \U$5319 ( \5696 , \5692 , \5695 );
and \U$5320 ( \5697 , \5687 , \5695 );
or \U$5321 ( \5698 , \5693 , \5696 , \5697 );
xor \U$5322 ( \5699 , \5444 , \5446 );
xor \U$5323 ( \5700 , \5699 , \5449 );
and \U$5324 ( \5701 , \5698 , \5700 );
and \U$5325 ( \5702 , \5462 , \5701 );
xor \U$5326 ( \5703 , \5462 , \5701 );
xor \U$5327 ( \5704 , \5698 , \5700 );
xor \U$5328 ( \5705 , \5051 , \5463 );
xor \U$5329 ( \5706 , \5463 , \5464 );
not \U$5330 ( \5707 , \5706 );
and \U$5331 ( \5708 , \5705 , \5707 );
and \U$5332 ( \5709 , \378 , \5708 );
not \U$5333 ( \5710 , \5709 );
xnor \U$5334 ( \5711 , \5710 , \5467 );
and \U$5335 ( \5712 , \410 , \5242 );
and \U$5336 ( \5713 , \392 , \5240 );
nor \U$5337 ( \5714 , \5712 , \5713 );
xnor \U$5338 ( \5715 , \5714 , \5054 );
and \U$5339 ( \5716 , \5711 , \5715 );
and \U$5340 ( \5717 , \479 , \4868 );
and \U$5341 ( \5718 , \431 , \4866 );
nor \U$5342 ( \5719 , \5717 , \5718 );
xnor \U$5343 ( \5720 , \5719 , \4636 );
and \U$5344 ( \5721 , \5715 , \5720 );
and \U$5345 ( \5722 , \5711 , \5720 );
or \U$5346 ( \5723 , \5716 , \5721 , \5722 );
and \U$5347 ( \5724 , \556 , \4417 );
and \U$5348 ( \5725 , \487 , \4415 );
nor \U$5349 ( \5726 , \5724 , \5725 );
xnor \U$5350 ( \5727 , \5726 , \4274 );
and \U$5351 ( \5728 , \615 , \4094 );
and \U$5352 ( \5729 , \561 , \4092 );
nor \U$5353 ( \5730 , \5728 , \5729 );
xnor \U$5354 ( \5731 , \5730 , \3848 );
and \U$5355 ( \5732 , \5727 , \5731 );
and \U$5356 ( \5733 , \743 , \3699 );
and \U$5357 ( \5734 , \666 , \3697 );
nor \U$5358 ( \5735 , \5733 , \5734 );
xnor \U$5359 ( \5736 , \5735 , \3512 );
and \U$5360 ( \5737 , \5731 , \5736 );
and \U$5361 ( \5738 , \5727 , \5736 );
or \U$5362 ( \5739 , \5732 , \5737 , \5738 );
and \U$5363 ( \5740 , \5723 , \5739 );
and \U$5364 ( \5741 , \851 , \3386 );
and \U$5365 ( \5742 , \771 , \3384 );
nor \U$5366 ( \5743 , \5741 , \5742 );
xnor \U$5367 ( \5744 , \5743 , \3181 );
and \U$5368 ( \5745 , \987 , \2980 );
and \U$5369 ( \5746 , \925 , \2978 );
nor \U$5370 ( \5747 , \5745 , \5746 );
xnor \U$5371 ( \5748 , \5747 , \2831 );
and \U$5372 ( \5749 , \5744 , \5748 );
and \U$5373 ( \5750 , \1248 , \2658 );
and \U$5374 ( \5751 , \1050 , \2656 );
nor \U$5375 ( \5752 , \5750 , \5751 );
xnor \U$5376 ( \5753 , \5752 , \2516 );
and \U$5377 ( \5754 , \5748 , \5753 );
and \U$5378 ( \5755 , \5744 , \5753 );
or \U$5379 ( \5756 , \5749 , \5754 , \5755 );
and \U$5380 ( \5757 , \5739 , \5756 );
and \U$5381 ( \5758 , \5723 , \5756 );
or \U$5382 ( \5759 , \5740 , \5757 , \5758 );
and \U$5383 ( \5760 , \1441 , \2362 );
and \U$5384 ( \5761 , \1336 , \2360 );
nor \U$5385 ( \5762 , \5760 , \5761 );
xnor \U$5386 ( \5763 , \5762 , \2225 );
and \U$5387 ( \5764 , \1562 , \2156 );
and \U$5388 ( \5765 , \1446 , \2154 );
nor \U$5389 ( \5766 , \5764 , \5765 );
xnor \U$5390 ( \5767 , \5766 , \2004 );
and \U$5391 ( \5768 , \5763 , \5767 );
and \U$5392 ( \5769 , \1853 , \1888 );
and \U$5393 ( \5770 , \1677 , \1886 );
nor \U$5394 ( \5771 , \5769 , \5770 );
xnor \U$5395 ( \5772 , \5771 , \1732 );
and \U$5396 ( \5773 , \5767 , \5772 );
and \U$5397 ( \5774 , \5763 , \5772 );
or \U$5398 ( \5775 , \5768 , \5773 , \5774 );
and \U$5399 ( \5776 , \2104 , \1616 );
and \U$5400 ( \5777 , \1861 , \1614 );
nor \U$5401 ( \5778 , \5776 , \5777 );
xnor \U$5402 ( \5779 , \5778 , \1503 );
and \U$5403 ( \5780 , \2295 , \1422 );
and \U$5404 ( \5781 , \2109 , \1420 );
nor \U$5405 ( \5782 , \5780 , \5781 );
xnor \U$5406 ( \5783 , \5782 , \1286 );
and \U$5407 ( \5784 , \5779 , \5783 );
and \U$5408 ( \5785 , \2703 , \1222 );
and \U$5409 ( \5786 , \2439 , \1220 );
nor \U$5410 ( \5787 , \5785 , \5786 );
xnor \U$5411 ( \5788 , \5787 , \1144 );
and \U$5412 ( \5789 , \5783 , \5788 );
and \U$5413 ( \5790 , \5779 , \5788 );
or \U$5414 ( \5791 , \5784 , \5789 , \5790 );
and \U$5415 ( \5792 , \5775 , \5791 );
and \U$5416 ( \5793 , \2902 , \1058 );
and \U$5417 ( \5794 , \2728 , \1056 );
nor \U$5418 ( \5795 , \5793 , \5794 );
xnor \U$5419 ( \5796 , \5795 , \964 );
and \U$5420 ( \5797 , \3207 , \888 );
and \U$5421 ( \5798 , \3069 , \886 );
nor \U$5422 ( \5799 , \5797 , \5798 );
xnor \U$5423 ( \5800 , \5799 , \816 );
and \U$5424 ( \5801 , \5796 , \5800 );
and \U$5425 ( \5802 , \3743 , \754 );
and \U$5426 ( \5803 , \3326 , \752 );
nor \U$5427 ( \5804 , \5802 , \5803 );
xnor \U$5428 ( \5805 , \5804 , \711 );
and \U$5429 ( \5806 , \5800 , \5805 );
and \U$5430 ( \5807 , \5796 , \5805 );
or \U$5431 ( \5808 , \5801 , \5806 , \5807 );
and \U$5432 ( \5809 , \5791 , \5808 );
and \U$5433 ( \5810 , \5775 , \5808 );
or \U$5434 ( \5811 , \5792 , \5809 , \5810 );
and \U$5435 ( \5812 , \5759 , \5811 );
and \U$5436 ( \5813 , \4073 , \641 );
and \U$5437 ( \5814 , \3951 , \639 );
nor \U$5438 ( \5815 , \5813 , \5814 );
xnor \U$5439 ( \5816 , \5815 , \592 );
and \U$5440 ( \5817 , \4334 , \540 );
and \U$5441 ( \5818 , \4078 , \538 );
nor \U$5442 ( \5819 , \5817 , \5818 );
xnor \U$5443 ( \5820 , \5819 , \499 );
and \U$5444 ( \5821 , \5816 , \5820 );
and \U$5445 ( \5822 , \4833 , \470 );
and \U$5446 ( \5823 , \4531 , \468 );
nor \U$5447 ( \5824 , \5822 , \5823 );
xnor \U$5448 ( \5825 , \5824 , \440 );
and \U$5449 ( \5826 , \5820 , \5825 );
and \U$5450 ( \5827 , \5816 , \5825 );
or \U$5451 ( \5828 , \5821 , \5826 , \5827 );
and \U$5452 ( \5829 , \5310 , \422 );
and \U$5453 ( \5830 , \4841 , \420 );
nor \U$5454 ( \5831 , \5829 , \5830 );
xnor \U$5455 ( \5832 , \5831 , \403 );
and \U$5456 ( \5833 , \5579 , \385 );
and \U$5457 ( \5834 , \5315 , \383 );
nor \U$5458 ( \5835 , \5833 , \5834 );
xnor \U$5459 ( \5836 , \5835 , \390 );
and \U$5460 ( \5837 , \5832 , \5836 );
buf \U$5461 ( \5838 , RIc224298_110);
and \U$5462 ( \5839 , \5838 , \379 );
and \U$5463 ( \5840 , \5836 , \5839 );
and \U$5464 ( \5841 , \5832 , \5839 );
or \U$5465 ( \5842 , \5837 , \5840 , \5841 );
and \U$5466 ( \5843 , \5828 , \5842 );
xor \U$5467 ( \5844 , \5573 , \5577 );
xor \U$5468 ( \5845 , \5844 , \5580 );
and \U$5469 ( \5846 , \5842 , \5845 );
and \U$5470 ( \5847 , \5828 , \5845 );
or \U$5471 ( \5848 , \5843 , \5846 , \5847 );
and \U$5472 ( \5849 , \5811 , \5848 );
and \U$5473 ( \5850 , \5759 , \5848 );
or \U$5474 ( \5851 , \5812 , \5849 , \5850 );
xor \U$5475 ( \5852 , \5520 , \5524 );
xor \U$5476 ( \5853 , \5852 , \5529 );
xor \U$5477 ( \5854 , \5484 , \5488 );
xor \U$5478 ( \5855 , \5854 , \5493 );
and \U$5479 ( \5856 , \5853 , \5855 );
xor \U$5480 ( \5857 , \5501 , \5505 );
xor \U$5481 ( \5858 , \5857 , \5510 );
and \U$5482 ( \5859 , \5855 , \5858 );
and \U$5483 ( \5860 , \5853 , \5858 );
or \U$5484 ( \5861 , \5856 , \5859 , \5860 );
xor \U$5485 ( \5862 , \5536 , \5540 );
xor \U$5486 ( \5863 , \5862 , \5545 );
xor \U$5487 ( \5864 , \5553 , \5557 );
xor \U$5488 ( \5865 , \5864 , \5562 );
and \U$5489 ( \5866 , \5863 , \5865 );
xor \U$5490 ( \5867 , \5587 , \5591 );
xor \U$5491 ( \5868 , \5867 , \5596 );
and \U$5492 ( \5869 , \5865 , \5868 );
and \U$5493 ( \5870 , \5863 , \5868 );
or \U$5494 ( \5871 , \5866 , \5869 , \5870 );
and \U$5495 ( \5872 , \5861 , \5871 );
xor \U$5496 ( \5873 , \5245 , \5249 );
xor \U$5497 ( \5874 , \5873 , \5254 );
and \U$5498 ( \5875 , \5871 , \5874 );
and \U$5499 ( \5876 , \5861 , \5874 );
or \U$5500 ( \5877 , \5872 , \5875 , \5876 );
and \U$5501 ( \5878 , \5851 , \5877 );
xor \U$5502 ( \5879 , \5609 , \5611 );
xor \U$5503 ( \5880 , \5879 , \5614 );
xor \U$5504 ( \5881 , \5619 , \5621 );
xor \U$5505 ( \5882 , \5881 , \5624 );
and \U$5506 ( \5883 , \5880 , \5882 );
xor \U$5507 ( \5884 , \5583 , \5599 );
xor \U$5508 ( \5885 , \5884 , \5601 );
and \U$5509 ( \5886 , \5882 , \5885 );
and \U$5510 ( \5887 , \5880 , \5885 );
or \U$5511 ( \5888 , \5883 , \5886 , \5887 );
and \U$5512 ( \5889 , \5877 , \5888 );
and \U$5513 ( \5890 , \5851 , \5888 );
or \U$5514 ( \5891 , \5878 , \5889 , \5890 );
xor \U$5515 ( \5892 , \5617 , \5627 );
xor \U$5516 ( \5893 , \5892 , \5630 );
xor \U$5517 ( \5894 , \5649 , \5651 );
xor \U$5518 ( \5895 , \5894 , \5654 );
and \U$5519 ( \5896 , \5893 , \5895 );
xor \U$5520 ( \5897 , \5636 , \5638 );
xor \U$5521 ( \5898 , \5897 , \5641 );
and \U$5522 ( \5899 , \5895 , \5898 );
and \U$5523 ( \5900 , \5893 , \5898 );
or \U$5524 ( \5901 , \5896 , \5899 , \5900 );
and \U$5525 ( \5902 , \5891 , \5901 );
xor \U$5526 ( \5903 , \5390 , \5400 );
xor \U$5527 ( \5904 , \5903 , \5403 );
and \U$5528 ( \5905 , \5901 , \5904 );
and \U$5529 ( \5906 , \5891 , \5904 );
or \U$5530 ( \5907 , \5902 , \5905 , \5906 );
xor \U$5531 ( \5908 , \5293 , \5325 );
xor \U$5532 ( \5909 , \5908 , \5378 );
xor \U$5533 ( \5910 , \5607 , \5633 );
xor \U$5534 ( \5911 , \5910 , \5644 );
and \U$5535 ( \5912 , \5909 , \5911 );
xor \U$5536 ( \5913 , \5657 , \5659 );
xor \U$5537 ( \5914 , \5913 , \5662 );
and \U$5538 ( \5915 , \5911 , \5914 );
and \U$5539 ( \5916 , \5909 , \5914 );
or \U$5540 ( \5917 , \5912 , \5915 , \5916 );
and \U$5541 ( \5918 , \5907 , \5917 );
xor \U$5542 ( \5919 , \5673 , \5675 );
xor \U$5543 ( \5920 , \5919 , \5678 );
and \U$5544 ( \5921 , \5917 , \5920 );
and \U$5545 ( \5922 , \5907 , \5920 );
or \U$5546 ( \5923 , \5918 , \5921 , \5922 );
xor \U$5547 ( \5924 , \5671 , \5681 );
xor \U$5548 ( \5925 , \5924 , \5684 );
and \U$5549 ( \5926 , \5923 , \5925 );
xor \U$5550 ( \5927 , \5689 , \5691 );
and \U$5551 ( \5928 , \5925 , \5927 );
and \U$5552 ( \5929 , \5923 , \5927 );
or \U$5553 ( \5930 , \5926 , \5928 , \5929 );
xor \U$5554 ( \5931 , \5687 , \5692 );
xor \U$5555 ( \5932 , \5931 , \5695 );
and \U$5556 ( \5933 , \5930 , \5932 );
and \U$5557 ( \5934 , \5704 , \5933 );
xor \U$5558 ( \5935 , \5704 , \5933 );
xor \U$5559 ( \5936 , \5930 , \5932 );
and \U$5560 ( \5937 , \487 , \4868 );
and \U$5561 ( \5938 , \479 , \4866 );
nor \U$5562 ( \5939 , \5937 , \5938 );
xnor \U$5563 ( \5940 , \5939 , \4636 );
and \U$5564 ( \5941 , \561 , \4417 );
and \U$5565 ( \5942 , \556 , \4415 );
nor \U$5566 ( \5943 , \5941 , \5942 );
xnor \U$5567 ( \5944 , \5943 , \4274 );
and \U$5568 ( \5945 , \5940 , \5944 );
and \U$5569 ( \5946 , \666 , \4094 );
and \U$5570 ( \5947 , \615 , \4092 );
nor \U$5571 ( \5948 , \5946 , \5947 );
xnor \U$5572 ( \5949 , \5948 , \3848 );
and \U$5573 ( \5950 , \5944 , \5949 );
and \U$5574 ( \5951 , \5940 , \5949 );
or \U$5575 ( \5952 , \5945 , \5950 , \5951 );
buf \U$5576 ( \5953 , RIc225fa8_48);
buf \U$5577 ( \5954 , RIc225f30_49);
and \U$5578 ( \5955 , \5953 , \5954 );
not \U$5579 ( \5956 , \5955 );
and \U$5580 ( \5957 , \5464 , \5956 );
not \U$5581 ( \5958 , \5957 );
and \U$5582 ( \5959 , \392 , \5708 );
and \U$5583 ( \5960 , \378 , \5706 );
nor \U$5584 ( \5961 , \5959 , \5960 );
xnor \U$5585 ( \5962 , \5961 , \5467 );
and \U$5586 ( \5963 , \5958 , \5962 );
and \U$5587 ( \5964 , \431 , \5242 );
and \U$5588 ( \5965 , \410 , \5240 );
nor \U$5589 ( \5966 , \5964 , \5965 );
xnor \U$5590 ( \5967 , \5966 , \5054 );
and \U$5591 ( \5968 , \5962 , \5967 );
and \U$5592 ( \5969 , \5958 , \5967 );
or \U$5593 ( \5970 , \5963 , \5968 , \5969 );
and \U$5594 ( \5971 , \5952 , \5970 );
and \U$5595 ( \5972 , \771 , \3699 );
and \U$5596 ( \5973 , \743 , \3697 );
nor \U$5597 ( \5974 , \5972 , \5973 );
xnor \U$5598 ( \5975 , \5974 , \3512 );
and \U$5599 ( \5976 , \925 , \3386 );
and \U$5600 ( \5977 , \851 , \3384 );
nor \U$5601 ( \5978 , \5976 , \5977 );
xnor \U$5602 ( \5979 , \5978 , \3181 );
and \U$5603 ( \5980 , \5975 , \5979 );
and \U$5604 ( \5981 , \1050 , \2980 );
and \U$5605 ( \5982 , \987 , \2978 );
nor \U$5606 ( \5983 , \5981 , \5982 );
xnor \U$5607 ( \5984 , \5983 , \2831 );
and \U$5608 ( \5985 , \5979 , \5984 );
and \U$5609 ( \5986 , \5975 , \5984 );
or \U$5610 ( \5987 , \5980 , \5985 , \5986 );
and \U$5611 ( \5988 , \5970 , \5987 );
and \U$5612 ( \5989 , \5952 , \5987 );
or \U$5613 ( \5990 , \5971 , \5988 , \5989 );
and \U$5614 ( \5991 , \2728 , \1222 );
and \U$5615 ( \5992 , \2703 , \1220 );
nor \U$5616 ( \5993 , \5991 , \5992 );
xnor \U$5617 ( \5994 , \5993 , \1144 );
and \U$5618 ( \5995 , \3069 , \1058 );
and \U$5619 ( \5996 , \2902 , \1056 );
nor \U$5620 ( \5997 , \5995 , \5996 );
xnor \U$5621 ( \5998 , \5997 , \964 );
and \U$5622 ( \5999 , \5994 , \5998 );
and \U$5623 ( \6000 , \3326 , \888 );
and \U$5624 ( \6001 , \3207 , \886 );
nor \U$5625 ( \6002 , \6000 , \6001 );
xnor \U$5626 ( \6003 , \6002 , \816 );
and \U$5627 ( \6004 , \5998 , \6003 );
and \U$5628 ( \6005 , \5994 , \6003 );
or \U$5629 ( \6006 , \5999 , \6004 , \6005 );
and \U$5630 ( \6007 , \1861 , \1888 );
and \U$5631 ( \6008 , \1853 , \1886 );
nor \U$5632 ( \6009 , \6007 , \6008 );
xnor \U$5633 ( \6010 , \6009 , \1732 );
and \U$5634 ( \6011 , \2109 , \1616 );
and \U$5635 ( \6012 , \2104 , \1614 );
nor \U$5636 ( \6013 , \6011 , \6012 );
xnor \U$5637 ( \6014 , \6013 , \1503 );
and \U$5638 ( \6015 , \6010 , \6014 );
and \U$5639 ( \6016 , \2439 , \1422 );
and \U$5640 ( \6017 , \2295 , \1420 );
nor \U$5641 ( \6018 , \6016 , \6017 );
xnor \U$5642 ( \6019 , \6018 , \1286 );
and \U$5643 ( \6020 , \6014 , \6019 );
and \U$5644 ( \6021 , \6010 , \6019 );
or \U$5645 ( \6022 , \6015 , \6020 , \6021 );
and \U$5646 ( \6023 , \6006 , \6022 );
and \U$5647 ( \6024 , \1336 , \2658 );
and \U$5648 ( \6025 , \1248 , \2656 );
nor \U$5649 ( \6026 , \6024 , \6025 );
xnor \U$5650 ( \6027 , \6026 , \2516 );
and \U$5651 ( \6028 , \1446 , \2362 );
and \U$5652 ( \6029 , \1441 , \2360 );
nor \U$5653 ( \6030 , \6028 , \6029 );
xnor \U$5654 ( \6031 , \6030 , \2225 );
and \U$5655 ( \6032 , \6027 , \6031 );
and \U$5656 ( \6033 , \1677 , \2156 );
and \U$5657 ( \6034 , \1562 , \2154 );
nor \U$5658 ( \6035 , \6033 , \6034 );
xnor \U$5659 ( \6036 , \6035 , \2004 );
and \U$5660 ( \6037 , \6031 , \6036 );
and \U$5661 ( \6038 , \6027 , \6036 );
or \U$5662 ( \6039 , \6032 , \6037 , \6038 );
and \U$5663 ( \6040 , \6022 , \6039 );
and \U$5664 ( \6041 , \6006 , \6039 );
or \U$5665 ( \6042 , \6023 , \6040 , \6041 );
and \U$5666 ( \6043 , \5990 , \6042 );
and \U$5667 ( \6044 , \3951 , \754 );
and \U$5668 ( \6045 , \3743 , \752 );
nor \U$5669 ( \6046 , \6044 , \6045 );
xnor \U$5670 ( \6047 , \6046 , \711 );
and \U$5671 ( \6048 , \4078 , \641 );
and \U$5672 ( \6049 , \4073 , \639 );
nor \U$5673 ( \6050 , \6048 , \6049 );
xnor \U$5674 ( \6051 , \6050 , \592 );
and \U$5675 ( \6052 , \6047 , \6051 );
and \U$5676 ( \6053 , \4531 , \540 );
and \U$5677 ( \6054 , \4334 , \538 );
nor \U$5678 ( \6055 , \6053 , \6054 );
xnor \U$5679 ( \6056 , \6055 , \499 );
and \U$5680 ( \6057 , \6051 , \6056 );
and \U$5681 ( \6058 , \6047 , \6056 );
or \U$5682 ( \6059 , \6052 , \6057 , \6058 );
and \U$5683 ( \6060 , \4841 , \470 );
and \U$5684 ( \6061 , \4833 , \468 );
nor \U$5685 ( \6062 , \6060 , \6061 );
xnor \U$5686 ( \6063 , \6062 , \440 );
and \U$5687 ( \6064 , \5315 , \422 );
and \U$5688 ( \6065 , \5310 , \420 );
nor \U$5689 ( \6066 , \6064 , \6065 );
xnor \U$5690 ( \6067 , \6066 , \403 );
and \U$5691 ( \6068 , \6063 , \6067 );
and \U$5692 ( \6069 , \5838 , \385 );
and \U$5693 ( \6070 , \5579 , \383 );
nor \U$5694 ( \6071 , \6069 , \6070 );
xnor \U$5695 ( \6072 , \6071 , \390 );
and \U$5696 ( \6073 , \6067 , \6072 );
and \U$5697 ( \6074 , \6063 , \6072 );
or \U$5698 ( \6075 , \6068 , \6073 , \6074 );
or \U$5699 ( \6076 , \6059 , \6075 );
and \U$5700 ( \6077 , \6042 , \6076 );
and \U$5701 ( \6078 , \5990 , \6076 );
or \U$5702 ( \6079 , \6043 , \6077 , \6078 );
xor \U$5703 ( \6080 , \5763 , \5767 );
xor \U$5704 ( \6081 , \6080 , \5772 );
xor \U$5705 ( \6082 , \5779 , \5783 );
xor \U$5706 ( \6083 , \6082 , \5788 );
and \U$5707 ( \6084 , \6081 , \6083 );
xor \U$5708 ( \6085 , \5744 , \5748 );
xor \U$5709 ( \6086 , \6085 , \5753 );
and \U$5710 ( \6087 , \6083 , \6086 );
and \U$5711 ( \6088 , \6081 , \6086 );
or \U$5712 ( \6089 , \6084 , \6087 , \6088 );
xor \U$5713 ( \6090 , \5796 , \5800 );
xor \U$5714 ( \6091 , \6090 , \5805 );
xor \U$5715 ( \6092 , \5816 , \5820 );
xor \U$5716 ( \6093 , \6092 , \5825 );
and \U$5717 ( \6094 , \6091 , \6093 );
xor \U$5718 ( \6095 , \5832 , \5836 );
xor \U$5719 ( \6096 , \6095 , \5839 );
and \U$5720 ( \6097 , \6093 , \6096 );
and \U$5721 ( \6098 , \6091 , \6096 );
or \U$5722 ( \6099 , \6094 , \6097 , \6098 );
and \U$5723 ( \6100 , \6089 , \6099 );
xor \U$5724 ( \6101 , \5711 , \5715 );
xor \U$5725 ( \6102 , \6101 , \5720 );
xor \U$5726 ( \6103 , \5727 , \5731 );
xor \U$5727 ( \6104 , \6103 , \5736 );
and \U$5728 ( \6105 , \6102 , \6104 );
and \U$5729 ( \6106 , \6099 , \6105 );
and \U$5730 ( \6107 , \6089 , \6105 );
or \U$5731 ( \6108 , \6100 , \6106 , \6107 );
and \U$5732 ( \6109 , \6079 , \6108 );
xor \U$5733 ( \6110 , \5468 , \5472 );
xor \U$5734 ( \6111 , \6110 , \5477 );
xor \U$5735 ( \6112 , \5853 , \5855 );
xor \U$5736 ( \6113 , \6112 , \5858 );
and \U$5737 ( \6114 , \6111 , \6113 );
xor \U$5738 ( \6115 , \5863 , \5865 );
xor \U$5739 ( \6116 , \6115 , \5868 );
and \U$5740 ( \6117 , \6113 , \6116 );
and \U$5741 ( \6118 , \6111 , \6116 );
or \U$5742 ( \6119 , \6114 , \6117 , \6118 );
and \U$5743 ( \6120 , \6108 , \6119 );
and \U$5744 ( \6121 , \6079 , \6119 );
or \U$5745 ( \6122 , \6109 , \6120 , \6121 );
xor \U$5746 ( \6123 , \5723 , \5739 );
xor \U$5747 ( \6124 , \6123 , \5756 );
xor \U$5748 ( \6125 , \5775 , \5791 );
xor \U$5749 ( \6126 , \6125 , \5808 );
and \U$5750 ( \6127 , \6124 , \6126 );
xor \U$5751 ( \6128 , \5828 , \5842 );
xor \U$5752 ( \6129 , \6128 , \5845 );
and \U$5753 ( \6130 , \6126 , \6129 );
and \U$5754 ( \6131 , \6124 , \6129 );
or \U$5755 ( \6132 , \6127 , \6130 , \6131 );
xor \U$5756 ( \6133 , \5480 , \5496 );
xor \U$5757 ( \6134 , \6133 , \5513 );
and \U$5758 ( \6135 , \6132 , \6134 );
xor \U$5759 ( \6136 , \5532 , \5548 );
xor \U$5760 ( \6137 , \6136 , \5565 );
and \U$5761 ( \6138 , \6134 , \6137 );
and \U$5762 ( \6139 , \6132 , \6137 );
or \U$5763 ( \6140 , \6135 , \6138 , \6139 );
and \U$5764 ( \6141 , \6122 , \6140 );
xor \U$5765 ( \6142 , \5759 , \5811 );
xor \U$5766 ( \6143 , \6142 , \5848 );
xor \U$5767 ( \6144 , \5861 , \5871 );
xor \U$5768 ( \6145 , \6144 , \5874 );
and \U$5769 ( \6146 , \6143 , \6145 );
xor \U$5770 ( \6147 , \5880 , \5882 );
xor \U$5771 ( \6148 , \6147 , \5885 );
and \U$5772 ( \6149 , \6145 , \6148 );
and \U$5773 ( \6150 , \6143 , \6148 );
or \U$5774 ( \6151 , \6146 , \6149 , \6150 );
and \U$5775 ( \6152 , \6140 , \6151 );
and \U$5776 ( \6153 , \6122 , \6151 );
or \U$5777 ( \6154 , \6141 , \6152 , \6153 );
xor \U$5778 ( \6155 , \5516 , \5568 );
xor \U$5779 ( \6156 , \6155 , \5604 );
xor \U$5780 ( \6157 , \5851 , \5877 );
xor \U$5781 ( \6158 , \6157 , \5888 );
and \U$5782 ( \6159 , \6156 , \6158 );
xor \U$5783 ( \6160 , \5893 , \5895 );
xor \U$5784 ( \6161 , \6160 , \5898 );
and \U$5785 ( \6162 , \6158 , \6161 );
and \U$5786 ( \6163 , \6156 , \6161 );
or \U$5787 ( \6164 , \6159 , \6162 , \6163 );
and \U$5788 ( \6165 , \6154 , \6164 );
xor \U$5789 ( \6166 , \5909 , \5911 );
xor \U$5790 ( \6167 , \6166 , \5914 );
and \U$5791 ( \6168 , \6164 , \6167 );
and \U$5792 ( \6169 , \6154 , \6167 );
or \U$5793 ( \6170 , \6165 , \6168 , \6169 );
xor \U$5794 ( \6171 , \5647 , \5665 );
xor \U$5795 ( \6172 , \6171 , \5668 );
and \U$5796 ( \6173 , \6170 , \6172 );
xor \U$5797 ( \6174 , \5907 , \5917 );
xor \U$5798 ( \6175 , \6174 , \5920 );
and \U$5799 ( \6176 , \6172 , \6175 );
and \U$5800 ( \6177 , \6170 , \6175 );
or \U$5801 ( \6178 , \6173 , \6176 , \6177 );
xor \U$5802 ( \6179 , \5923 , \5925 );
xor \U$5803 ( \6180 , \6179 , \5927 );
and \U$5804 ( \6181 , \6178 , \6180 );
and \U$5805 ( \6182 , \5936 , \6181 );
xor \U$5806 ( \6183 , \5936 , \6181 );
xor \U$5807 ( \6184 , \6178 , \6180 );
and \U$5808 ( \6185 , \4073 , \754 );
and \U$5809 ( \6186 , \3951 , \752 );
nor \U$5810 ( \6187 , \6185 , \6186 );
xnor \U$5811 ( \6188 , \6187 , \711 );
and \U$5812 ( \6189 , \4334 , \641 );
and \U$5813 ( \6190 , \4078 , \639 );
nor \U$5814 ( \6191 , \6189 , \6190 );
xnor \U$5815 ( \6192 , \6191 , \592 );
and \U$5816 ( \6193 , \6188 , \6192 );
and \U$5817 ( \6194 , \4833 , \540 );
and \U$5818 ( \6195 , \4531 , \538 );
nor \U$5819 ( \6196 , \6194 , \6195 );
xnor \U$5820 ( \6197 , \6196 , \499 );
and \U$5821 ( \6198 , \6192 , \6197 );
and \U$5822 ( \6199 , \6188 , \6197 );
or \U$5823 ( \6200 , \6193 , \6198 , \6199 );
and \U$5824 ( \6201 , \5310 , \470 );
and \U$5825 ( \6202 , \4841 , \468 );
nor \U$5826 ( \6203 , \6201 , \6202 );
xnor \U$5827 ( \6204 , \6203 , \440 );
and \U$5828 ( \6205 , \5579 , \422 );
and \U$5829 ( \6206 , \5315 , \420 );
nor \U$5830 ( \6207 , \6205 , \6206 );
xnor \U$5831 ( \6208 , \6207 , \403 );
and \U$5832 ( \6209 , \6204 , \6208 );
buf \U$5833 ( \6210 , RIc224220_111);
and \U$5834 ( \6211 , \6210 , \385 );
and \U$5835 ( \6212 , \5838 , \383 );
nor \U$5836 ( \6213 , \6211 , \6212 );
xnor \U$5837 ( \6214 , \6213 , \390 );
and \U$5838 ( \6215 , \6208 , \6214 );
and \U$5839 ( \6216 , \6204 , \6214 );
or \U$5840 ( \6217 , \6209 , \6215 , \6216 );
and \U$5841 ( \6218 , \6200 , \6217 );
buf \U$5842 ( \6219 , RIc2241a8_112);
and \U$5843 ( \6220 , \6219 , \379 );
buf \U$5844 ( \6221 , \6220 );
and \U$5845 ( \6222 , \6217 , \6221 );
and \U$5846 ( \6223 , \6200 , \6221 );
or \U$5847 ( \6224 , \6218 , \6222 , \6223 );
and \U$5848 ( \6225 , \2104 , \1888 );
and \U$5849 ( \6226 , \1861 , \1886 );
nor \U$5850 ( \6227 , \6225 , \6226 );
xnor \U$5851 ( \6228 , \6227 , \1732 );
and \U$5852 ( \6229 , \2295 , \1616 );
and \U$5853 ( \6230 , \2109 , \1614 );
nor \U$5854 ( \6231 , \6229 , \6230 );
xnor \U$5855 ( \6232 , \6231 , \1503 );
and \U$5856 ( \6233 , \6228 , \6232 );
and \U$5857 ( \6234 , \2703 , \1422 );
and \U$5858 ( \6235 , \2439 , \1420 );
nor \U$5859 ( \6236 , \6234 , \6235 );
xnor \U$5860 ( \6237 , \6236 , \1286 );
and \U$5861 ( \6238 , \6232 , \6237 );
and \U$5862 ( \6239 , \6228 , \6237 );
or \U$5863 ( \6240 , \6233 , \6238 , \6239 );
and \U$5864 ( \6241 , \1441 , \2658 );
and \U$5865 ( \6242 , \1336 , \2656 );
nor \U$5866 ( \6243 , \6241 , \6242 );
xnor \U$5867 ( \6244 , \6243 , \2516 );
and \U$5868 ( \6245 , \1562 , \2362 );
and \U$5869 ( \6246 , \1446 , \2360 );
nor \U$5870 ( \6247 , \6245 , \6246 );
xnor \U$5871 ( \6248 , \6247 , \2225 );
and \U$5872 ( \6249 , \6244 , \6248 );
and \U$5873 ( \6250 , \1853 , \2156 );
and \U$5874 ( \6251 , \1677 , \2154 );
nor \U$5875 ( \6252 , \6250 , \6251 );
xnor \U$5876 ( \6253 , \6252 , \2004 );
and \U$5877 ( \6254 , \6248 , \6253 );
and \U$5878 ( \6255 , \6244 , \6253 );
or \U$5879 ( \6256 , \6249 , \6254 , \6255 );
and \U$5880 ( \6257 , \6240 , \6256 );
and \U$5881 ( \6258 , \2902 , \1222 );
and \U$5882 ( \6259 , \2728 , \1220 );
nor \U$5883 ( \6260 , \6258 , \6259 );
xnor \U$5884 ( \6261 , \6260 , \1144 );
and \U$5885 ( \6262 , \3207 , \1058 );
and \U$5886 ( \6263 , \3069 , \1056 );
nor \U$5887 ( \6264 , \6262 , \6263 );
xnor \U$5888 ( \6265 , \6264 , \964 );
and \U$5889 ( \6266 , \6261 , \6265 );
and \U$5890 ( \6267 , \3743 , \888 );
and \U$5891 ( \6268 , \3326 , \886 );
nor \U$5892 ( \6269 , \6267 , \6268 );
xnor \U$5893 ( \6270 , \6269 , \816 );
and \U$5894 ( \6271 , \6265 , \6270 );
and \U$5895 ( \6272 , \6261 , \6270 );
or \U$5896 ( \6273 , \6266 , \6271 , \6272 );
and \U$5897 ( \6274 , \6256 , \6273 );
and \U$5898 ( \6275 , \6240 , \6273 );
or \U$5899 ( \6276 , \6257 , \6274 , \6275 );
and \U$5900 ( \6277 , \6224 , \6276 );
and \U$5901 ( \6278 , \556 , \4868 );
and \U$5902 ( \6279 , \487 , \4866 );
nor \U$5903 ( \6280 , \6278 , \6279 );
xnor \U$5904 ( \6281 , \6280 , \4636 );
and \U$5905 ( \6282 , \615 , \4417 );
and \U$5906 ( \6283 , \561 , \4415 );
nor \U$5907 ( \6284 , \6282 , \6283 );
xnor \U$5908 ( \6285 , \6284 , \4274 );
and \U$5909 ( \6286 , \6281 , \6285 );
and \U$5910 ( \6287 , \743 , \4094 );
and \U$5911 ( \6288 , \666 , \4092 );
nor \U$5912 ( \6289 , \6287 , \6288 );
xnor \U$5913 ( \6290 , \6289 , \3848 );
and \U$5914 ( \6291 , \6285 , \6290 );
and \U$5915 ( \6292 , \6281 , \6290 );
or \U$5916 ( \6293 , \6286 , \6291 , \6292 );
xor \U$5917 ( \6294 , \5464 , \5953 );
xor \U$5918 ( \6295 , \5953 , \5954 );
not \U$5919 ( \6296 , \6295 );
and \U$5920 ( \6297 , \6294 , \6296 );
and \U$5921 ( \6298 , \378 , \6297 );
not \U$5922 ( \6299 , \6298 );
xnor \U$5923 ( \6300 , \6299 , \5957 );
and \U$5924 ( \6301 , \410 , \5708 );
and \U$5925 ( \6302 , \392 , \5706 );
nor \U$5926 ( \6303 , \6301 , \6302 );
xnor \U$5927 ( \6304 , \6303 , \5467 );
and \U$5928 ( \6305 , \6300 , \6304 );
and \U$5929 ( \6306 , \479 , \5242 );
and \U$5930 ( \6307 , \431 , \5240 );
nor \U$5931 ( \6308 , \6306 , \6307 );
xnor \U$5932 ( \6309 , \6308 , \5054 );
and \U$5933 ( \6310 , \6304 , \6309 );
and \U$5934 ( \6311 , \6300 , \6309 );
or \U$5935 ( \6312 , \6305 , \6310 , \6311 );
and \U$5936 ( \6313 , \6293 , \6312 );
and \U$5937 ( \6314 , \851 , \3699 );
and \U$5938 ( \6315 , \771 , \3697 );
nor \U$5939 ( \6316 , \6314 , \6315 );
xnor \U$5940 ( \6317 , \6316 , \3512 );
and \U$5941 ( \6318 , \987 , \3386 );
and \U$5942 ( \6319 , \925 , \3384 );
nor \U$5943 ( \6320 , \6318 , \6319 );
xnor \U$5944 ( \6321 , \6320 , \3181 );
and \U$5945 ( \6322 , \6317 , \6321 );
and \U$5946 ( \6323 , \1248 , \2980 );
and \U$5947 ( \6324 , \1050 , \2978 );
nor \U$5948 ( \6325 , \6323 , \6324 );
xnor \U$5949 ( \6326 , \6325 , \2831 );
and \U$5950 ( \6327 , \6321 , \6326 );
and \U$5951 ( \6328 , \6317 , \6326 );
or \U$5952 ( \6329 , \6322 , \6327 , \6328 );
and \U$5953 ( \6330 , \6312 , \6329 );
and \U$5954 ( \6331 , \6293 , \6329 );
or \U$5955 ( \6332 , \6313 , \6330 , \6331 );
and \U$5956 ( \6333 , \6276 , \6332 );
and \U$5957 ( \6334 , \6224 , \6332 );
or \U$5958 ( \6335 , \6277 , \6333 , \6334 );
xor \U$5959 ( \6336 , \5940 , \5944 );
xor \U$5960 ( \6337 , \6336 , \5949 );
xor \U$5961 ( \6338 , \5958 , \5962 );
xor \U$5962 ( \6339 , \6338 , \5967 );
and \U$5963 ( \6340 , \6337 , \6339 );
xor \U$5964 ( \6341 , \5975 , \5979 );
xor \U$5965 ( \6342 , \6341 , \5984 );
and \U$5966 ( \6343 , \6339 , \6342 );
and \U$5967 ( \6344 , \6337 , \6342 );
or \U$5968 ( \6345 , \6340 , \6343 , \6344 );
xor \U$5969 ( \6346 , \5994 , \5998 );
xor \U$5970 ( \6347 , \6346 , \6003 );
xor \U$5971 ( \6348 , \6010 , \6014 );
xor \U$5972 ( \6349 , \6348 , \6019 );
and \U$5973 ( \6350 , \6347 , \6349 );
xor \U$5974 ( \6351 , \6027 , \6031 );
xor \U$5975 ( \6352 , \6351 , \6036 );
and \U$5976 ( \6353 , \6349 , \6352 );
and \U$5977 ( \6354 , \6347 , \6352 );
or \U$5978 ( \6355 , \6350 , \6353 , \6354 );
and \U$5979 ( \6356 , \6345 , \6355 );
and \U$5980 ( \6357 , \6210 , \379 );
xor \U$5981 ( \6358 , \6047 , \6051 );
xor \U$5982 ( \6359 , \6358 , \6056 );
and \U$5983 ( \6360 , \6357 , \6359 );
xor \U$5984 ( \6361 , \6063 , \6067 );
xor \U$5985 ( \6362 , \6361 , \6072 );
and \U$5986 ( \6363 , \6359 , \6362 );
and \U$5987 ( \6364 , \6357 , \6362 );
or \U$5988 ( \6365 , \6360 , \6363 , \6364 );
and \U$5989 ( \6366 , \6355 , \6365 );
and \U$5990 ( \6367 , \6345 , \6365 );
or \U$5991 ( \6368 , \6356 , \6366 , \6367 );
and \U$5992 ( \6369 , \6335 , \6368 );
xor \U$5993 ( \6370 , \6081 , \6083 );
xor \U$5994 ( \6371 , \6370 , \6086 );
xor \U$5995 ( \6372 , \6091 , \6093 );
xor \U$5996 ( \6373 , \6372 , \6096 );
and \U$5997 ( \6374 , \6371 , \6373 );
xor \U$5998 ( \6375 , \6102 , \6104 );
and \U$5999 ( \6376 , \6373 , \6375 );
and \U$6000 ( \6377 , \6371 , \6375 );
or \U$6001 ( \6378 , \6374 , \6376 , \6377 );
and \U$6002 ( \6379 , \6368 , \6378 );
and \U$6003 ( \6380 , \6335 , \6378 );
or \U$6004 ( \6381 , \6369 , \6379 , \6380 );
xor \U$6005 ( \6382 , \5952 , \5970 );
xor \U$6006 ( \6383 , \6382 , \5987 );
xor \U$6007 ( \6384 , \6006 , \6022 );
xor \U$6008 ( \6385 , \6384 , \6039 );
and \U$6009 ( \6386 , \6383 , \6385 );
xnor \U$6010 ( \6387 , \6059 , \6075 );
and \U$6011 ( \6388 , \6385 , \6387 );
and \U$6012 ( \6389 , \6383 , \6387 );
or \U$6013 ( \6390 , \6386 , \6388 , \6389 );
xor \U$6014 ( \6391 , \6111 , \6113 );
xor \U$6015 ( \6392 , \6391 , \6116 );
and \U$6016 ( \6393 , \6390 , \6392 );
xor \U$6017 ( \6394 , \6124 , \6126 );
xor \U$6018 ( \6395 , \6394 , \6129 );
and \U$6019 ( \6396 , \6392 , \6395 );
and \U$6020 ( \6397 , \6390 , \6395 );
or \U$6021 ( \6398 , \6393 , \6396 , \6397 );
and \U$6022 ( \6399 , \6381 , \6398 );
xor \U$6023 ( \6400 , \5990 , \6042 );
xor \U$6024 ( \6401 , \6400 , \6076 );
xor \U$6025 ( \6402 , \6089 , \6099 );
xor \U$6026 ( \6403 , \6402 , \6105 );
and \U$6027 ( \6404 , \6401 , \6403 );
and \U$6028 ( \6405 , \6398 , \6404 );
and \U$6029 ( \6406 , \6381 , \6404 );
or \U$6030 ( \6407 , \6399 , \6405 , \6406 );
xor \U$6031 ( \6408 , \6079 , \6108 );
xor \U$6032 ( \6409 , \6408 , \6119 );
xor \U$6033 ( \6410 , \6132 , \6134 );
xor \U$6034 ( \6411 , \6410 , \6137 );
and \U$6035 ( \6412 , \6409 , \6411 );
xor \U$6036 ( \6413 , \6143 , \6145 );
xor \U$6037 ( \6414 , \6413 , \6148 );
and \U$6038 ( \6415 , \6411 , \6414 );
and \U$6039 ( \6416 , \6409 , \6414 );
or \U$6040 ( \6417 , \6412 , \6415 , \6416 );
and \U$6041 ( \6418 , \6407 , \6417 );
xor \U$6042 ( \6419 , \6156 , \6158 );
xor \U$6043 ( \6420 , \6419 , \6161 );
and \U$6044 ( \6421 , \6417 , \6420 );
and \U$6045 ( \6422 , \6407 , \6420 );
or \U$6046 ( \6423 , \6418 , \6421 , \6422 );
xor \U$6047 ( \6424 , \5891 , \5901 );
xor \U$6048 ( \6425 , \6424 , \5904 );
and \U$6049 ( \6426 , \6423 , \6425 );
xor \U$6050 ( \6427 , \6154 , \6164 );
xor \U$6051 ( \6428 , \6427 , \6167 );
and \U$6052 ( \6429 , \6425 , \6428 );
and \U$6053 ( \6430 , \6423 , \6428 );
or \U$6054 ( \6431 , \6426 , \6429 , \6430 );
xor \U$6055 ( \6432 , \6170 , \6172 );
xor \U$6056 ( \6433 , \6432 , \6175 );
and \U$6057 ( \6434 , \6431 , \6433 );
and \U$6058 ( \6435 , \6184 , \6434 );
xor \U$6059 ( \6436 , \6184 , \6434 );
xor \U$6060 ( \6437 , \6431 , \6433 );
xor \U$6061 ( \6438 , \6228 , \6232 );
xor \U$6062 ( \6439 , \6438 , \6237 );
xor \U$6063 ( \6440 , \6244 , \6248 );
xor \U$6064 ( \6441 , \6440 , \6253 );
and \U$6065 ( \6442 , \6439 , \6441 );
xor \U$6066 ( \6443 , \6261 , \6265 );
xor \U$6067 ( \6444 , \6443 , \6270 );
and \U$6068 ( \6445 , \6441 , \6444 );
and \U$6069 ( \6446 , \6439 , \6444 );
or \U$6070 ( \6447 , \6442 , \6445 , \6446 );
xor \U$6071 ( \6448 , \6281 , \6285 );
xor \U$6072 ( \6449 , \6448 , \6290 );
xor \U$6073 ( \6450 , \6300 , \6304 );
xor \U$6074 ( \6451 , \6450 , \6309 );
and \U$6075 ( \6452 , \6449 , \6451 );
xor \U$6076 ( \6453 , \6317 , \6321 );
xor \U$6077 ( \6454 , \6453 , \6326 );
and \U$6078 ( \6455 , \6451 , \6454 );
and \U$6079 ( \6456 , \6449 , \6454 );
or \U$6080 ( \6457 , \6452 , \6455 , \6456 );
and \U$6081 ( \6458 , \6447 , \6457 );
xor \U$6082 ( \6459 , \6188 , \6192 );
xor \U$6083 ( \6460 , \6459 , \6197 );
xor \U$6084 ( \6461 , \6204 , \6208 );
xor \U$6085 ( \6462 , \6461 , \6214 );
and \U$6086 ( \6463 , \6460 , \6462 );
not \U$6087 ( \6464 , \6220 );
and \U$6088 ( \6465 , \6462 , \6464 );
and \U$6089 ( \6466 , \6460 , \6464 );
or \U$6090 ( \6467 , \6463 , \6465 , \6466 );
and \U$6091 ( \6468 , \6457 , \6467 );
and \U$6092 ( \6469 , \6447 , \6467 );
or \U$6093 ( \6470 , \6458 , \6468 , \6469 );
and \U$6094 ( \6471 , \487 , \5242 );
and \U$6095 ( \6472 , \479 , \5240 );
nor \U$6096 ( \6473 , \6471 , \6472 );
xnor \U$6097 ( \6474 , \6473 , \5054 );
and \U$6098 ( \6475 , \561 , \4868 );
and \U$6099 ( \6476 , \556 , \4866 );
nor \U$6100 ( \6477 , \6475 , \6476 );
xnor \U$6101 ( \6478 , \6477 , \4636 );
and \U$6102 ( \6479 , \6474 , \6478 );
and \U$6103 ( \6480 , \666 , \4417 );
and \U$6104 ( \6481 , \615 , \4415 );
nor \U$6105 ( \6482 , \6480 , \6481 );
xnor \U$6106 ( \6483 , \6482 , \4274 );
and \U$6107 ( \6484 , \6478 , \6483 );
and \U$6108 ( \6485 , \6474 , \6483 );
or \U$6109 ( \6486 , \6479 , \6484 , \6485 );
buf \U$6110 ( \6487 , RIc225eb8_50);
buf \U$6111 ( \6488 , RIc225e40_51);
and \U$6112 ( \6489 , \6487 , \6488 );
not \U$6113 ( \6490 , \6489 );
and \U$6114 ( \6491 , \5954 , \6490 );
not \U$6115 ( \6492 , \6491 );
and \U$6116 ( \6493 , \392 , \6297 );
and \U$6117 ( \6494 , \378 , \6295 );
nor \U$6118 ( \6495 , \6493 , \6494 );
xnor \U$6119 ( \6496 , \6495 , \5957 );
and \U$6120 ( \6497 , \6492 , \6496 );
and \U$6121 ( \6498 , \431 , \5708 );
and \U$6122 ( \6499 , \410 , \5706 );
nor \U$6123 ( \6500 , \6498 , \6499 );
xnor \U$6124 ( \6501 , \6500 , \5467 );
and \U$6125 ( \6502 , \6496 , \6501 );
and \U$6126 ( \6503 , \6492 , \6501 );
or \U$6127 ( \6504 , \6497 , \6502 , \6503 );
and \U$6128 ( \6505 , \6486 , \6504 );
and \U$6129 ( \6506 , \771 , \4094 );
and \U$6130 ( \6507 , \743 , \4092 );
nor \U$6131 ( \6508 , \6506 , \6507 );
xnor \U$6132 ( \6509 , \6508 , \3848 );
and \U$6133 ( \6510 , \925 , \3699 );
and \U$6134 ( \6511 , \851 , \3697 );
nor \U$6135 ( \6512 , \6510 , \6511 );
xnor \U$6136 ( \6513 , \6512 , \3512 );
and \U$6137 ( \6514 , \6509 , \6513 );
and \U$6138 ( \6515 , \1050 , \3386 );
and \U$6139 ( \6516 , \987 , \3384 );
nor \U$6140 ( \6517 , \6515 , \6516 );
xnor \U$6141 ( \6518 , \6517 , \3181 );
and \U$6142 ( \6519 , \6513 , \6518 );
and \U$6143 ( \6520 , \6509 , \6518 );
or \U$6144 ( \6521 , \6514 , \6519 , \6520 );
and \U$6145 ( \6522 , \6504 , \6521 );
and \U$6146 ( \6523 , \6486 , \6521 );
or \U$6147 ( \6524 , \6505 , \6522 , \6523 );
and \U$6148 ( \6525 , \3951 , \888 );
and \U$6149 ( \6526 , \3743 , \886 );
nor \U$6150 ( \6527 , \6525 , \6526 );
xnor \U$6151 ( \6528 , \6527 , \816 );
and \U$6152 ( \6529 , \4078 , \754 );
and \U$6153 ( \6530 , \4073 , \752 );
nor \U$6154 ( \6531 , \6529 , \6530 );
xnor \U$6155 ( \6532 , \6531 , \711 );
and \U$6156 ( \6533 , \6528 , \6532 );
and \U$6157 ( \6534 , \4531 , \641 );
and \U$6158 ( \6535 , \4334 , \639 );
nor \U$6159 ( \6536 , \6534 , \6535 );
xnor \U$6160 ( \6537 , \6536 , \592 );
and \U$6161 ( \6538 , \6532 , \6537 );
and \U$6162 ( \6539 , \6528 , \6537 );
or \U$6163 ( \6540 , \6533 , \6538 , \6539 );
and \U$6164 ( \6541 , \4841 , \540 );
and \U$6165 ( \6542 , \4833 , \538 );
nor \U$6166 ( \6543 , \6541 , \6542 );
xnor \U$6167 ( \6544 , \6543 , \499 );
and \U$6168 ( \6545 , \5315 , \470 );
and \U$6169 ( \6546 , \5310 , \468 );
nor \U$6170 ( \6547 , \6545 , \6546 );
xnor \U$6171 ( \6548 , \6547 , \440 );
and \U$6172 ( \6549 , \6544 , \6548 );
and \U$6173 ( \6550 , \5838 , \422 );
and \U$6174 ( \6551 , \5579 , \420 );
nor \U$6175 ( \6552 , \6550 , \6551 );
xnor \U$6176 ( \6553 , \6552 , \403 );
and \U$6177 ( \6554 , \6548 , \6553 );
and \U$6178 ( \6555 , \6544 , \6553 );
or \U$6179 ( \6556 , \6549 , \6554 , \6555 );
and \U$6180 ( \6557 , \6540 , \6556 );
and \U$6181 ( \6558 , \6219 , \385 );
and \U$6182 ( \6559 , \6210 , \383 );
nor \U$6183 ( \6560 , \6558 , \6559 );
xnor \U$6184 ( \6561 , \6560 , \390 );
buf \U$6185 ( \6562 , RIc224130_113);
and \U$6186 ( \6563 , \6562 , \379 );
and \U$6187 ( \6564 , \6561 , \6563 );
and \U$6188 ( \6565 , \6556 , \6564 );
and \U$6189 ( \6566 , \6540 , \6564 );
or \U$6190 ( \6567 , \6557 , \6565 , \6566 );
and \U$6191 ( \6568 , \6524 , \6567 );
and \U$6192 ( \6569 , \1336 , \2980 );
and \U$6193 ( \6570 , \1248 , \2978 );
nor \U$6194 ( \6571 , \6569 , \6570 );
xnor \U$6195 ( \6572 , \6571 , \2831 );
and \U$6196 ( \6573 , \1446 , \2658 );
and \U$6197 ( \6574 , \1441 , \2656 );
nor \U$6198 ( \6575 , \6573 , \6574 );
xnor \U$6199 ( \6576 , \6575 , \2516 );
and \U$6200 ( \6577 , \6572 , \6576 );
and \U$6201 ( \6578 , \1677 , \2362 );
and \U$6202 ( \6579 , \1562 , \2360 );
nor \U$6203 ( \6580 , \6578 , \6579 );
xnor \U$6204 ( \6581 , \6580 , \2225 );
and \U$6205 ( \6582 , \6576 , \6581 );
and \U$6206 ( \6583 , \6572 , \6581 );
or \U$6207 ( \6584 , \6577 , \6582 , \6583 );
and \U$6208 ( \6585 , \1861 , \2156 );
and \U$6209 ( \6586 , \1853 , \2154 );
nor \U$6210 ( \6587 , \6585 , \6586 );
xnor \U$6211 ( \6588 , \6587 , \2004 );
and \U$6212 ( \6589 , \2109 , \1888 );
and \U$6213 ( \6590 , \2104 , \1886 );
nor \U$6214 ( \6591 , \6589 , \6590 );
xnor \U$6215 ( \6592 , \6591 , \1732 );
and \U$6216 ( \6593 , \6588 , \6592 );
and \U$6217 ( \6594 , \2439 , \1616 );
and \U$6218 ( \6595 , \2295 , \1614 );
nor \U$6219 ( \6596 , \6594 , \6595 );
xnor \U$6220 ( \6597 , \6596 , \1503 );
and \U$6221 ( \6598 , \6592 , \6597 );
and \U$6222 ( \6599 , \6588 , \6597 );
or \U$6223 ( \6600 , \6593 , \6598 , \6599 );
and \U$6224 ( \6601 , \6584 , \6600 );
and \U$6225 ( \6602 , \2728 , \1422 );
and \U$6226 ( \6603 , \2703 , \1420 );
nor \U$6227 ( \6604 , \6602 , \6603 );
xnor \U$6228 ( \6605 , \6604 , \1286 );
and \U$6229 ( \6606 , \3069 , \1222 );
and \U$6230 ( \6607 , \2902 , \1220 );
nor \U$6231 ( \6608 , \6606 , \6607 );
xnor \U$6232 ( \6609 , \6608 , \1144 );
and \U$6233 ( \6610 , \6605 , \6609 );
and \U$6234 ( \6611 , \3326 , \1058 );
and \U$6235 ( \6612 , \3207 , \1056 );
nor \U$6236 ( \6613 , \6611 , \6612 );
xnor \U$6237 ( \6614 , \6613 , \964 );
and \U$6238 ( \6615 , \6609 , \6614 );
and \U$6239 ( \6616 , \6605 , \6614 );
or \U$6240 ( \6617 , \6610 , \6615 , \6616 );
and \U$6241 ( \6618 , \6600 , \6617 );
and \U$6242 ( \6619 , \6584 , \6617 );
or \U$6243 ( \6620 , \6601 , \6618 , \6619 );
and \U$6244 ( \6621 , \6567 , \6620 );
and \U$6245 ( \6622 , \6524 , \6620 );
or \U$6246 ( \6623 , \6568 , \6621 , \6622 );
and \U$6247 ( \6624 , \6470 , \6623 );
xor \U$6248 ( \6625 , \6337 , \6339 );
xor \U$6249 ( \6626 , \6625 , \6342 );
xor \U$6250 ( \6627 , \6347 , \6349 );
xor \U$6251 ( \6628 , \6627 , \6352 );
and \U$6252 ( \6629 , \6626 , \6628 );
xor \U$6253 ( \6630 , \6357 , \6359 );
xor \U$6254 ( \6631 , \6630 , \6362 );
and \U$6255 ( \6632 , \6628 , \6631 );
and \U$6256 ( \6633 , \6626 , \6631 );
or \U$6257 ( \6634 , \6629 , \6632 , \6633 );
and \U$6258 ( \6635 , \6623 , \6634 );
and \U$6259 ( \6636 , \6470 , \6634 );
or \U$6260 ( \6637 , \6624 , \6635 , \6636 );
xor \U$6261 ( \6638 , \6200 , \6217 );
xor \U$6262 ( \6639 , \6638 , \6221 );
xor \U$6263 ( \6640 , \6240 , \6256 );
xor \U$6264 ( \6641 , \6640 , \6273 );
and \U$6265 ( \6642 , \6639 , \6641 );
xor \U$6266 ( \6643 , \6293 , \6312 );
xor \U$6267 ( \6644 , \6643 , \6329 );
and \U$6268 ( \6645 , \6641 , \6644 );
and \U$6269 ( \6646 , \6639 , \6644 );
or \U$6270 ( \6647 , \6642 , \6645 , \6646 );
xor \U$6271 ( \6648 , \6383 , \6385 );
xor \U$6272 ( \6649 , \6648 , \6387 );
and \U$6273 ( \6650 , \6647 , \6649 );
xor \U$6274 ( \6651 , \6371 , \6373 );
xor \U$6275 ( \6652 , \6651 , \6375 );
and \U$6276 ( \6653 , \6649 , \6652 );
and \U$6277 ( \6654 , \6647 , \6652 );
or \U$6278 ( \6655 , \6650 , \6653 , \6654 );
and \U$6279 ( \6656 , \6637 , \6655 );
xor \U$6280 ( \6657 , \6224 , \6276 );
xor \U$6281 ( \6658 , \6657 , \6332 );
xor \U$6282 ( \6659 , \6345 , \6355 );
xor \U$6283 ( \6660 , \6659 , \6365 );
and \U$6284 ( \6661 , \6658 , \6660 );
and \U$6285 ( \6662 , \6655 , \6661 );
and \U$6286 ( \6663 , \6637 , \6661 );
or \U$6287 ( \6664 , \6656 , \6662 , \6663 );
xor \U$6288 ( \6665 , \6335 , \6368 );
xor \U$6289 ( \6666 , \6665 , \6378 );
xor \U$6290 ( \6667 , \6390 , \6392 );
xor \U$6291 ( \6668 , \6667 , \6395 );
and \U$6292 ( \6669 , \6666 , \6668 );
xor \U$6293 ( \6670 , \6401 , \6403 );
and \U$6294 ( \6671 , \6668 , \6670 );
and \U$6295 ( \6672 , \6666 , \6670 );
or \U$6296 ( \6673 , \6669 , \6671 , \6672 );
and \U$6297 ( \6674 , \6664 , \6673 );
xor \U$6298 ( \6675 , \6409 , \6411 );
xor \U$6299 ( \6676 , \6675 , \6414 );
and \U$6300 ( \6677 , \6673 , \6676 );
and \U$6301 ( \6678 , \6664 , \6676 );
or \U$6302 ( \6679 , \6674 , \6677 , \6678 );
xor \U$6303 ( \6680 , \6122 , \6140 );
xor \U$6304 ( \6681 , \6680 , \6151 );
and \U$6305 ( \6682 , \6679 , \6681 );
xor \U$6306 ( \6683 , \6407 , \6417 );
xor \U$6307 ( \6684 , \6683 , \6420 );
and \U$6308 ( \6685 , \6681 , \6684 );
and \U$6309 ( \6686 , \6679 , \6684 );
or \U$6310 ( \6687 , \6682 , \6685 , \6686 );
xor \U$6311 ( \6688 , \6423 , \6425 );
xor \U$6312 ( \6689 , \6688 , \6428 );
and \U$6313 ( \6690 , \6687 , \6689 );
and \U$6314 ( \6691 , \6437 , \6690 );
xor \U$6315 ( \6692 , \6437 , \6690 );
xor \U$6316 ( \6693 , \6687 , \6689 );
xor \U$6317 ( \6694 , \6572 , \6576 );
xor \U$6318 ( \6695 , \6694 , \6581 );
xor \U$6319 ( \6696 , \6588 , \6592 );
xor \U$6320 ( \6697 , \6696 , \6597 );
and \U$6321 ( \6698 , \6695 , \6697 );
xor \U$6322 ( \6699 , \6605 , \6609 );
xor \U$6323 ( \6700 , \6699 , \6614 );
and \U$6324 ( \6701 , \6697 , \6700 );
and \U$6325 ( \6702 , \6695 , \6700 );
or \U$6326 ( \6703 , \6698 , \6701 , \6702 );
xor \U$6327 ( \6704 , \6474 , \6478 );
xor \U$6328 ( \6705 , \6704 , \6483 );
xor \U$6329 ( \6706 , \6492 , \6496 );
xor \U$6330 ( \6707 , \6706 , \6501 );
and \U$6331 ( \6708 , \6705 , \6707 );
xor \U$6332 ( \6709 , \6509 , \6513 );
xor \U$6333 ( \6710 , \6709 , \6518 );
and \U$6334 ( \6711 , \6707 , \6710 );
and \U$6335 ( \6712 , \6705 , \6710 );
or \U$6336 ( \6713 , \6708 , \6711 , \6712 );
and \U$6337 ( \6714 , \6703 , \6713 );
xor \U$6338 ( \6715 , \6528 , \6532 );
xor \U$6339 ( \6716 , \6715 , \6537 );
xor \U$6340 ( \6717 , \6544 , \6548 );
xor \U$6341 ( \6718 , \6717 , \6553 );
and \U$6342 ( \6719 , \6716 , \6718 );
xor \U$6343 ( \6720 , \6561 , \6563 );
and \U$6344 ( \6721 , \6718 , \6720 );
and \U$6345 ( \6722 , \6716 , \6720 );
or \U$6346 ( \6723 , \6719 , \6721 , \6722 );
and \U$6347 ( \6724 , \6713 , \6723 );
and \U$6348 ( \6725 , \6703 , \6723 );
or \U$6349 ( \6726 , \6714 , \6724 , \6725 );
and \U$6350 ( \6727 , \4073 , \888 );
and \U$6351 ( \6728 , \3951 , \886 );
nor \U$6352 ( \6729 , \6727 , \6728 );
xnor \U$6353 ( \6730 , \6729 , \816 );
and \U$6354 ( \6731 , \4334 , \754 );
and \U$6355 ( \6732 , \4078 , \752 );
nor \U$6356 ( \6733 , \6731 , \6732 );
xnor \U$6357 ( \6734 , \6733 , \711 );
and \U$6358 ( \6735 , \6730 , \6734 );
and \U$6359 ( \6736 , \4833 , \641 );
and \U$6360 ( \6737 , \4531 , \639 );
nor \U$6361 ( \6738 , \6736 , \6737 );
xnor \U$6362 ( \6739 , \6738 , \592 );
and \U$6363 ( \6740 , \6734 , \6739 );
and \U$6364 ( \6741 , \6730 , \6739 );
or \U$6365 ( \6742 , \6735 , \6740 , \6741 );
and \U$6366 ( \6743 , \5310 , \540 );
and \U$6367 ( \6744 , \4841 , \538 );
nor \U$6368 ( \6745 , \6743 , \6744 );
xnor \U$6369 ( \6746 , \6745 , \499 );
and \U$6370 ( \6747 , \5579 , \470 );
and \U$6371 ( \6748 , \5315 , \468 );
nor \U$6372 ( \6749 , \6747 , \6748 );
xnor \U$6373 ( \6750 , \6749 , \440 );
and \U$6374 ( \6751 , \6746 , \6750 );
and \U$6375 ( \6752 , \6210 , \422 );
and \U$6376 ( \6753 , \5838 , \420 );
nor \U$6377 ( \6754 , \6752 , \6753 );
xnor \U$6378 ( \6755 , \6754 , \403 );
and \U$6379 ( \6756 , \6750 , \6755 );
and \U$6380 ( \6757 , \6746 , \6755 );
or \U$6381 ( \6758 , \6751 , \6756 , \6757 );
and \U$6382 ( \6759 , \6742 , \6758 );
and \U$6383 ( \6760 , \6562 , \385 );
and \U$6384 ( \6761 , \6219 , \383 );
nor \U$6385 ( \6762 , \6760 , \6761 );
xnor \U$6386 ( \6763 , \6762 , \390 );
buf \U$6387 ( \6764 , RIc2240b8_114);
and \U$6388 ( \6765 , \6764 , \379 );
or \U$6389 ( \6766 , \6763 , \6765 );
and \U$6390 ( \6767 , \6758 , \6766 );
and \U$6391 ( \6768 , \6742 , \6766 );
or \U$6392 ( \6769 , \6759 , \6767 , \6768 );
and \U$6393 ( \6770 , \851 , \4094 );
and \U$6394 ( \6771 , \771 , \4092 );
nor \U$6395 ( \6772 , \6770 , \6771 );
xnor \U$6396 ( \6773 , \6772 , \3848 );
and \U$6397 ( \6774 , \987 , \3699 );
and \U$6398 ( \6775 , \925 , \3697 );
nor \U$6399 ( \6776 , \6774 , \6775 );
xnor \U$6400 ( \6777 , \6776 , \3512 );
and \U$6401 ( \6778 , \6773 , \6777 );
and \U$6402 ( \6779 , \1248 , \3386 );
and \U$6403 ( \6780 , \1050 , \3384 );
nor \U$6404 ( \6781 , \6779 , \6780 );
xnor \U$6405 ( \6782 , \6781 , \3181 );
and \U$6406 ( \6783 , \6777 , \6782 );
and \U$6407 ( \6784 , \6773 , \6782 );
or \U$6408 ( \6785 , \6778 , \6783 , \6784 );
and \U$6409 ( \6786 , \556 , \5242 );
and \U$6410 ( \6787 , \487 , \5240 );
nor \U$6411 ( \6788 , \6786 , \6787 );
xnor \U$6412 ( \6789 , \6788 , \5054 );
and \U$6413 ( \6790 , \615 , \4868 );
and \U$6414 ( \6791 , \561 , \4866 );
nor \U$6415 ( \6792 , \6790 , \6791 );
xnor \U$6416 ( \6793 , \6792 , \4636 );
and \U$6417 ( \6794 , \6789 , \6793 );
and \U$6418 ( \6795 , \743 , \4417 );
and \U$6419 ( \6796 , \666 , \4415 );
nor \U$6420 ( \6797 , \6795 , \6796 );
xnor \U$6421 ( \6798 , \6797 , \4274 );
and \U$6422 ( \6799 , \6793 , \6798 );
and \U$6423 ( \6800 , \6789 , \6798 );
or \U$6424 ( \6801 , \6794 , \6799 , \6800 );
and \U$6425 ( \6802 , \6785 , \6801 );
xor \U$6426 ( \6803 , \5954 , \6487 );
xor \U$6427 ( \6804 , \6487 , \6488 );
not \U$6428 ( \6805 , \6804 );
and \U$6429 ( \6806 , \6803 , \6805 );
and \U$6430 ( \6807 , \378 , \6806 );
not \U$6431 ( \6808 , \6807 );
xnor \U$6432 ( \6809 , \6808 , \6491 );
and \U$6433 ( \6810 , \410 , \6297 );
and \U$6434 ( \6811 , \392 , \6295 );
nor \U$6435 ( \6812 , \6810 , \6811 );
xnor \U$6436 ( \6813 , \6812 , \5957 );
and \U$6437 ( \6814 , \6809 , \6813 );
and \U$6438 ( \6815 , \479 , \5708 );
and \U$6439 ( \6816 , \431 , \5706 );
nor \U$6440 ( \6817 , \6815 , \6816 );
xnor \U$6441 ( \6818 , \6817 , \5467 );
and \U$6442 ( \6819 , \6813 , \6818 );
and \U$6443 ( \6820 , \6809 , \6818 );
or \U$6444 ( \6821 , \6814 , \6819 , \6820 );
and \U$6445 ( \6822 , \6801 , \6821 );
and \U$6446 ( \6823 , \6785 , \6821 );
or \U$6447 ( \6824 , \6802 , \6822 , \6823 );
and \U$6448 ( \6825 , \6769 , \6824 );
and \U$6449 ( \6826 , \2104 , \2156 );
and \U$6450 ( \6827 , \1861 , \2154 );
nor \U$6451 ( \6828 , \6826 , \6827 );
xnor \U$6452 ( \6829 , \6828 , \2004 );
and \U$6453 ( \6830 , \2295 , \1888 );
and \U$6454 ( \6831 , \2109 , \1886 );
nor \U$6455 ( \6832 , \6830 , \6831 );
xnor \U$6456 ( \6833 , \6832 , \1732 );
and \U$6457 ( \6834 , \6829 , \6833 );
and \U$6458 ( \6835 , \2703 , \1616 );
and \U$6459 ( \6836 , \2439 , \1614 );
nor \U$6460 ( \6837 , \6835 , \6836 );
xnor \U$6461 ( \6838 , \6837 , \1503 );
and \U$6462 ( \6839 , \6833 , \6838 );
and \U$6463 ( \6840 , \6829 , \6838 );
or \U$6464 ( \6841 , \6834 , \6839 , \6840 );
and \U$6465 ( \6842 , \2902 , \1422 );
and \U$6466 ( \6843 , \2728 , \1420 );
nor \U$6467 ( \6844 , \6842 , \6843 );
xnor \U$6468 ( \6845 , \6844 , \1286 );
and \U$6469 ( \6846 , \3207 , \1222 );
and \U$6470 ( \6847 , \3069 , \1220 );
nor \U$6471 ( \6848 , \6846 , \6847 );
xnor \U$6472 ( \6849 , \6848 , \1144 );
and \U$6473 ( \6850 , \6845 , \6849 );
and \U$6474 ( \6851 , \3743 , \1058 );
and \U$6475 ( \6852 , \3326 , \1056 );
nor \U$6476 ( \6853 , \6851 , \6852 );
xnor \U$6477 ( \6854 , \6853 , \964 );
and \U$6478 ( \6855 , \6849 , \6854 );
and \U$6479 ( \6856 , \6845 , \6854 );
or \U$6480 ( \6857 , \6850 , \6855 , \6856 );
and \U$6481 ( \6858 , \6841 , \6857 );
and \U$6482 ( \6859 , \1441 , \2980 );
and \U$6483 ( \6860 , \1336 , \2978 );
nor \U$6484 ( \6861 , \6859 , \6860 );
xnor \U$6485 ( \6862 , \6861 , \2831 );
and \U$6486 ( \6863 , \1562 , \2658 );
and \U$6487 ( \6864 , \1446 , \2656 );
nor \U$6488 ( \6865 , \6863 , \6864 );
xnor \U$6489 ( \6866 , \6865 , \2516 );
and \U$6490 ( \6867 , \6862 , \6866 );
and \U$6491 ( \6868 , \1853 , \2362 );
and \U$6492 ( \6869 , \1677 , \2360 );
nor \U$6493 ( \6870 , \6868 , \6869 );
xnor \U$6494 ( \6871 , \6870 , \2225 );
and \U$6495 ( \6872 , \6866 , \6871 );
and \U$6496 ( \6873 , \6862 , \6871 );
or \U$6497 ( \6874 , \6867 , \6872 , \6873 );
and \U$6498 ( \6875 , \6857 , \6874 );
and \U$6499 ( \6876 , \6841 , \6874 );
or \U$6500 ( \6877 , \6858 , \6875 , \6876 );
and \U$6501 ( \6878 , \6824 , \6877 );
and \U$6502 ( \6879 , \6769 , \6877 );
or \U$6503 ( \6880 , \6825 , \6878 , \6879 );
and \U$6504 ( \6881 , \6726 , \6880 );
xor \U$6505 ( \6882 , \6439 , \6441 );
xor \U$6506 ( \6883 , \6882 , \6444 );
xor \U$6507 ( \6884 , \6449 , \6451 );
xor \U$6508 ( \6885 , \6884 , \6454 );
and \U$6509 ( \6886 , \6883 , \6885 );
xor \U$6510 ( \6887 , \6460 , \6462 );
xor \U$6511 ( \6888 , \6887 , \6464 );
and \U$6512 ( \6889 , \6885 , \6888 );
and \U$6513 ( \6890 , \6883 , \6888 );
or \U$6514 ( \6891 , \6886 , \6889 , \6890 );
and \U$6515 ( \6892 , \6880 , \6891 );
and \U$6516 ( \6893 , \6726 , \6891 );
or \U$6517 ( \6894 , \6881 , \6892 , \6893 );
xor \U$6518 ( \6895 , \6486 , \6504 );
xor \U$6519 ( \6896 , \6895 , \6521 );
xor \U$6520 ( \6897 , \6540 , \6556 );
xor \U$6521 ( \6898 , \6897 , \6564 );
and \U$6522 ( \6899 , \6896 , \6898 );
xor \U$6523 ( \6900 , \6584 , \6600 );
xor \U$6524 ( \6901 , \6900 , \6617 );
and \U$6525 ( \6902 , \6898 , \6901 );
and \U$6526 ( \6903 , \6896 , \6901 );
or \U$6527 ( \6904 , \6899 , \6902 , \6903 );
xor \U$6528 ( \6905 , \6639 , \6641 );
xor \U$6529 ( \6906 , \6905 , \6644 );
and \U$6530 ( \6907 , \6904 , \6906 );
xor \U$6531 ( \6908 , \6626 , \6628 );
xor \U$6532 ( \6909 , \6908 , \6631 );
and \U$6533 ( \6910 , \6906 , \6909 );
and \U$6534 ( \6911 , \6904 , \6909 );
or \U$6535 ( \6912 , \6907 , \6910 , \6911 );
and \U$6536 ( \6913 , \6894 , \6912 );
xor \U$6537 ( \6914 , \6447 , \6457 );
xor \U$6538 ( \6915 , \6914 , \6467 );
xor \U$6539 ( \6916 , \6524 , \6567 );
xor \U$6540 ( \6917 , \6916 , \6620 );
and \U$6541 ( \6918 , \6915 , \6917 );
and \U$6542 ( \6919 , \6912 , \6918 );
and \U$6543 ( \6920 , \6894 , \6918 );
or \U$6544 ( \6921 , \6913 , \6919 , \6920 );
xor \U$6545 ( \6922 , \6470 , \6623 );
xor \U$6546 ( \6923 , \6922 , \6634 );
xor \U$6547 ( \6924 , \6647 , \6649 );
xor \U$6548 ( \6925 , \6924 , \6652 );
and \U$6549 ( \6926 , \6923 , \6925 );
xor \U$6550 ( \6927 , \6658 , \6660 );
and \U$6551 ( \6928 , \6925 , \6927 );
and \U$6552 ( \6929 , \6923 , \6927 );
or \U$6553 ( \6930 , \6926 , \6928 , \6929 );
and \U$6554 ( \6931 , \6921 , \6930 );
xor \U$6555 ( \6932 , \6666 , \6668 );
xor \U$6556 ( \6933 , \6932 , \6670 );
and \U$6557 ( \6934 , \6930 , \6933 );
and \U$6558 ( \6935 , \6921 , \6933 );
or \U$6559 ( \6936 , \6931 , \6934 , \6935 );
xor \U$6560 ( \6937 , \6381 , \6398 );
xor \U$6561 ( \6938 , \6937 , \6404 );
and \U$6562 ( \6939 , \6936 , \6938 );
xor \U$6563 ( \6940 , \6664 , \6673 );
xor \U$6564 ( \6941 , \6940 , \6676 );
and \U$6565 ( \6942 , \6938 , \6941 );
and \U$6566 ( \6943 , \6936 , \6941 );
or \U$6567 ( \6944 , \6939 , \6942 , \6943 );
xor \U$6568 ( \6945 , \6679 , \6681 );
xor \U$6569 ( \6946 , \6945 , \6684 );
and \U$6570 ( \6947 , \6944 , \6946 );
and \U$6571 ( \6948 , \6693 , \6947 );
xor \U$6572 ( \6949 , \6693 , \6947 );
xor \U$6573 ( \6950 , \6944 , \6946 );
and \U$6574 ( \6951 , \1336 , \3386 );
and \U$6575 ( \6952 , \1248 , \3384 );
nor \U$6576 ( \6953 , \6951 , \6952 );
xnor \U$6577 ( \6954 , \6953 , \3181 );
and \U$6578 ( \6955 , \1446 , \2980 );
and \U$6579 ( \6956 , \1441 , \2978 );
nor \U$6580 ( \6957 , \6955 , \6956 );
xnor \U$6581 ( \6958 , \6957 , \2831 );
and \U$6582 ( \6959 , \6954 , \6958 );
and \U$6583 ( \6960 , \1677 , \2658 );
and \U$6584 ( \6961 , \1562 , \2656 );
nor \U$6585 ( \6962 , \6960 , \6961 );
xnor \U$6586 ( \6963 , \6962 , \2516 );
and \U$6587 ( \6964 , \6958 , \6963 );
and \U$6588 ( \6965 , \6954 , \6963 );
or \U$6589 ( \6966 , \6959 , \6964 , \6965 );
and \U$6590 ( \6967 , \1861 , \2362 );
and \U$6591 ( \6968 , \1853 , \2360 );
nor \U$6592 ( \6969 , \6967 , \6968 );
xnor \U$6593 ( \6970 , \6969 , \2225 );
and \U$6594 ( \6971 , \2109 , \2156 );
and \U$6595 ( \6972 , \2104 , \2154 );
nor \U$6596 ( \6973 , \6971 , \6972 );
xnor \U$6597 ( \6974 , \6973 , \2004 );
and \U$6598 ( \6975 , \6970 , \6974 );
and \U$6599 ( \6976 , \2439 , \1888 );
and \U$6600 ( \6977 , \2295 , \1886 );
nor \U$6601 ( \6978 , \6976 , \6977 );
xnor \U$6602 ( \6979 , \6978 , \1732 );
and \U$6603 ( \6980 , \6974 , \6979 );
and \U$6604 ( \6981 , \6970 , \6979 );
or \U$6605 ( \6982 , \6975 , \6980 , \6981 );
and \U$6606 ( \6983 , \6966 , \6982 );
and \U$6607 ( \6984 , \2728 , \1616 );
and \U$6608 ( \6985 , \2703 , \1614 );
nor \U$6609 ( \6986 , \6984 , \6985 );
xnor \U$6610 ( \6987 , \6986 , \1503 );
and \U$6611 ( \6988 , \3069 , \1422 );
and \U$6612 ( \6989 , \2902 , \1420 );
nor \U$6613 ( \6990 , \6988 , \6989 );
xnor \U$6614 ( \6991 , \6990 , \1286 );
and \U$6615 ( \6992 , \6987 , \6991 );
and \U$6616 ( \6993 , \3326 , \1222 );
and \U$6617 ( \6994 , \3207 , \1220 );
nor \U$6618 ( \6995 , \6993 , \6994 );
xnor \U$6619 ( \6996 , \6995 , \1144 );
and \U$6620 ( \6997 , \6991 , \6996 );
and \U$6621 ( \6998 , \6987 , \6996 );
or \U$6622 ( \6999 , \6992 , \6997 , \6998 );
and \U$6623 ( \7000 , \6982 , \6999 );
and \U$6624 ( \7001 , \6966 , \6999 );
or \U$6625 ( \7002 , \6983 , \7000 , \7001 );
and \U$6626 ( \7003 , \487 , \5708 );
and \U$6627 ( \7004 , \479 , \5706 );
nor \U$6628 ( \7005 , \7003 , \7004 );
xnor \U$6629 ( \7006 , \7005 , \5467 );
and \U$6630 ( \7007 , \561 , \5242 );
and \U$6631 ( \7008 , \556 , \5240 );
nor \U$6632 ( \7009 , \7007 , \7008 );
xnor \U$6633 ( \7010 , \7009 , \5054 );
and \U$6634 ( \7011 , \7006 , \7010 );
and \U$6635 ( \7012 , \666 , \4868 );
and \U$6636 ( \7013 , \615 , \4866 );
nor \U$6637 ( \7014 , \7012 , \7013 );
xnor \U$6638 ( \7015 , \7014 , \4636 );
and \U$6639 ( \7016 , \7010 , \7015 );
and \U$6640 ( \7017 , \7006 , \7015 );
or \U$6641 ( \7018 , \7011 , \7016 , \7017 );
and \U$6642 ( \7019 , \771 , \4417 );
and \U$6643 ( \7020 , \743 , \4415 );
nor \U$6644 ( \7021 , \7019 , \7020 );
xnor \U$6645 ( \7022 , \7021 , \4274 );
and \U$6646 ( \7023 , \925 , \4094 );
and \U$6647 ( \7024 , \851 , \4092 );
nor \U$6648 ( \7025 , \7023 , \7024 );
xnor \U$6649 ( \7026 , \7025 , \3848 );
and \U$6650 ( \7027 , \7022 , \7026 );
and \U$6651 ( \7028 , \1050 , \3699 );
and \U$6652 ( \7029 , \987 , \3697 );
nor \U$6653 ( \7030 , \7028 , \7029 );
xnor \U$6654 ( \7031 , \7030 , \3512 );
and \U$6655 ( \7032 , \7026 , \7031 );
and \U$6656 ( \7033 , \7022 , \7031 );
or \U$6657 ( \7034 , \7027 , \7032 , \7033 );
and \U$6658 ( \7035 , \7018 , \7034 );
buf \U$6659 ( \7036 , RIc225dc8_52);
buf \U$6660 ( \7037 , RIc225d50_53);
and \U$6661 ( \7038 , \7036 , \7037 );
not \U$6662 ( \7039 , \7038 );
and \U$6663 ( \7040 , \6488 , \7039 );
not \U$6664 ( \7041 , \7040 );
and \U$6665 ( \7042 , \392 , \6806 );
and \U$6666 ( \7043 , \378 , \6804 );
nor \U$6667 ( \7044 , \7042 , \7043 );
xnor \U$6668 ( \7045 , \7044 , \6491 );
and \U$6669 ( \7046 , \7041 , \7045 );
and \U$6670 ( \7047 , \431 , \6297 );
and \U$6671 ( \7048 , \410 , \6295 );
nor \U$6672 ( \7049 , \7047 , \7048 );
xnor \U$6673 ( \7050 , \7049 , \5957 );
and \U$6674 ( \7051 , \7045 , \7050 );
and \U$6675 ( \7052 , \7041 , \7050 );
or \U$6676 ( \7053 , \7046 , \7051 , \7052 );
and \U$6677 ( \7054 , \7034 , \7053 );
and \U$6678 ( \7055 , \7018 , \7053 );
or \U$6679 ( \7056 , \7035 , \7054 , \7055 );
and \U$6680 ( \7057 , \7002 , \7056 );
and \U$6681 ( \7058 , \6219 , \422 );
and \U$6682 ( \7059 , \6210 , \420 );
nor \U$6683 ( \7060 , \7058 , \7059 );
xnor \U$6684 ( \7061 , \7060 , \403 );
and \U$6685 ( \7062 , \6764 , \385 );
and \U$6686 ( \7063 , \6562 , \383 );
nor \U$6687 ( \7064 , \7062 , \7063 );
xnor \U$6688 ( \7065 , \7064 , \390 );
and \U$6689 ( \7066 , \7061 , \7065 );
buf \U$6690 ( \7067 , RIc224040_115);
and \U$6691 ( \7068 , \7067 , \379 );
and \U$6692 ( \7069 , \7065 , \7068 );
and \U$6693 ( \7070 , \7061 , \7068 );
or \U$6694 ( \7071 , \7066 , \7069 , \7070 );
and \U$6695 ( \7072 , \3951 , \1058 );
and \U$6696 ( \7073 , \3743 , \1056 );
nor \U$6697 ( \7074 , \7072 , \7073 );
xnor \U$6698 ( \7075 , \7074 , \964 );
and \U$6699 ( \7076 , \4078 , \888 );
and \U$6700 ( \7077 , \4073 , \886 );
nor \U$6701 ( \7078 , \7076 , \7077 );
xnor \U$6702 ( \7079 , \7078 , \816 );
and \U$6703 ( \7080 , \7075 , \7079 );
and \U$6704 ( \7081 , \4531 , \754 );
and \U$6705 ( \7082 , \4334 , \752 );
nor \U$6706 ( \7083 , \7081 , \7082 );
xnor \U$6707 ( \7084 , \7083 , \711 );
and \U$6708 ( \7085 , \7079 , \7084 );
and \U$6709 ( \7086 , \7075 , \7084 );
or \U$6710 ( \7087 , \7080 , \7085 , \7086 );
and \U$6711 ( \7088 , \7071 , \7087 );
and \U$6712 ( \7089 , \4841 , \641 );
and \U$6713 ( \7090 , \4833 , \639 );
nor \U$6714 ( \7091 , \7089 , \7090 );
xnor \U$6715 ( \7092 , \7091 , \592 );
and \U$6716 ( \7093 , \5315 , \540 );
and \U$6717 ( \7094 , \5310 , \538 );
nor \U$6718 ( \7095 , \7093 , \7094 );
xnor \U$6719 ( \7096 , \7095 , \499 );
and \U$6720 ( \7097 , \7092 , \7096 );
and \U$6721 ( \7098 , \5838 , \470 );
and \U$6722 ( \7099 , \5579 , \468 );
nor \U$6723 ( \7100 , \7098 , \7099 );
xnor \U$6724 ( \7101 , \7100 , \440 );
and \U$6725 ( \7102 , \7096 , \7101 );
and \U$6726 ( \7103 , \7092 , \7101 );
or \U$6727 ( \7104 , \7097 , \7102 , \7103 );
and \U$6728 ( \7105 , \7087 , \7104 );
and \U$6729 ( \7106 , \7071 , \7104 );
or \U$6730 ( \7107 , \7088 , \7105 , \7106 );
and \U$6731 ( \7108 , \7056 , \7107 );
and \U$6732 ( \7109 , \7002 , \7107 );
or \U$6733 ( \7110 , \7057 , \7108 , \7109 );
xor \U$6734 ( \7111 , \6829 , \6833 );
xor \U$6735 ( \7112 , \7111 , \6838 );
xor \U$6736 ( \7113 , \6845 , \6849 );
xor \U$6737 ( \7114 , \7113 , \6854 );
and \U$6738 ( \7115 , \7112 , \7114 );
xor \U$6739 ( \7116 , \6862 , \6866 );
xor \U$6740 ( \7117 , \7116 , \6871 );
and \U$6741 ( \7118 , \7114 , \7117 );
and \U$6742 ( \7119 , \7112 , \7117 );
or \U$6743 ( \7120 , \7115 , \7118 , \7119 );
xor \U$6744 ( \7121 , \6773 , \6777 );
xor \U$6745 ( \7122 , \7121 , \6782 );
xor \U$6746 ( \7123 , \6789 , \6793 );
xor \U$6747 ( \7124 , \7123 , \6798 );
and \U$6748 ( \7125 , \7122 , \7124 );
xor \U$6749 ( \7126 , \6809 , \6813 );
xor \U$6750 ( \7127 , \7126 , \6818 );
and \U$6751 ( \7128 , \7124 , \7127 );
and \U$6752 ( \7129 , \7122 , \7127 );
or \U$6753 ( \7130 , \7125 , \7128 , \7129 );
and \U$6754 ( \7131 , \7120 , \7130 );
xor \U$6755 ( \7132 , \6730 , \6734 );
xor \U$6756 ( \7133 , \7132 , \6739 );
xor \U$6757 ( \7134 , \6746 , \6750 );
xor \U$6758 ( \7135 , \7134 , \6755 );
and \U$6759 ( \7136 , \7133 , \7135 );
xnor \U$6760 ( \7137 , \6763 , \6765 );
and \U$6761 ( \7138 , \7135 , \7137 );
and \U$6762 ( \7139 , \7133 , \7137 );
or \U$6763 ( \7140 , \7136 , \7138 , \7139 );
and \U$6764 ( \7141 , \7130 , \7140 );
and \U$6765 ( \7142 , \7120 , \7140 );
or \U$6766 ( \7143 , \7131 , \7141 , \7142 );
and \U$6767 ( \7144 , \7110 , \7143 );
xor \U$6768 ( \7145 , \6695 , \6697 );
xor \U$6769 ( \7146 , \7145 , \6700 );
xor \U$6770 ( \7147 , \6705 , \6707 );
xor \U$6771 ( \7148 , \7147 , \6710 );
and \U$6772 ( \7149 , \7146 , \7148 );
xor \U$6773 ( \7150 , \6716 , \6718 );
xor \U$6774 ( \7151 , \7150 , \6720 );
and \U$6775 ( \7152 , \7148 , \7151 );
and \U$6776 ( \7153 , \7146 , \7151 );
or \U$6777 ( \7154 , \7149 , \7152 , \7153 );
and \U$6778 ( \7155 , \7143 , \7154 );
and \U$6779 ( \7156 , \7110 , \7154 );
or \U$6780 ( \7157 , \7144 , \7155 , \7156 );
xor \U$6781 ( \7158 , \6742 , \6758 );
xor \U$6782 ( \7159 , \7158 , \6766 );
xor \U$6783 ( \7160 , \6785 , \6801 );
xor \U$6784 ( \7161 , \7160 , \6821 );
and \U$6785 ( \7162 , \7159 , \7161 );
xor \U$6786 ( \7163 , \6841 , \6857 );
xor \U$6787 ( \7164 , \7163 , \6874 );
and \U$6788 ( \7165 , \7161 , \7164 );
and \U$6789 ( \7166 , \7159 , \7164 );
or \U$6790 ( \7167 , \7162 , \7165 , \7166 );
xor \U$6791 ( \7168 , \6896 , \6898 );
xor \U$6792 ( \7169 , \7168 , \6901 );
and \U$6793 ( \7170 , \7167 , \7169 );
xor \U$6794 ( \7171 , \6883 , \6885 );
xor \U$6795 ( \7172 , \7171 , \6888 );
and \U$6796 ( \7173 , \7169 , \7172 );
and \U$6797 ( \7174 , \7167 , \7172 );
or \U$6798 ( \7175 , \7170 , \7173 , \7174 );
and \U$6799 ( \7176 , \7157 , \7175 );
xor \U$6800 ( \7177 , \6703 , \6713 );
xor \U$6801 ( \7178 , \7177 , \6723 );
xor \U$6802 ( \7179 , \6769 , \6824 );
xor \U$6803 ( \7180 , \7179 , \6877 );
and \U$6804 ( \7181 , \7178 , \7180 );
and \U$6805 ( \7182 , \7175 , \7181 );
and \U$6806 ( \7183 , \7157 , \7181 );
or \U$6807 ( \7184 , \7176 , \7182 , \7183 );
xor \U$6808 ( \7185 , \6726 , \6880 );
xor \U$6809 ( \7186 , \7185 , \6891 );
xor \U$6810 ( \7187 , \6904 , \6906 );
xor \U$6811 ( \7188 , \7187 , \6909 );
and \U$6812 ( \7189 , \7186 , \7188 );
xor \U$6813 ( \7190 , \6915 , \6917 );
and \U$6814 ( \7191 , \7188 , \7190 );
and \U$6815 ( \7192 , \7186 , \7190 );
or \U$6816 ( \7193 , \7189 , \7191 , \7192 );
and \U$6817 ( \7194 , \7184 , \7193 );
xor \U$6818 ( \7195 , \6923 , \6925 );
xor \U$6819 ( \7196 , \7195 , \6927 );
and \U$6820 ( \7197 , \7193 , \7196 );
and \U$6821 ( \7198 , \7184 , \7196 );
or \U$6822 ( \7199 , \7194 , \7197 , \7198 );
xor \U$6823 ( \7200 , \6637 , \6655 );
xor \U$6824 ( \7201 , \7200 , \6661 );
and \U$6825 ( \7202 , \7199 , \7201 );
xor \U$6826 ( \7203 , \6921 , \6930 );
xor \U$6827 ( \7204 , \7203 , \6933 );
and \U$6828 ( \7205 , \7201 , \7204 );
and \U$6829 ( \7206 , \7199 , \7204 );
or \U$6830 ( \7207 , \7202 , \7205 , \7206 );
xor \U$6831 ( \7208 , \6936 , \6938 );
xor \U$6832 ( \7209 , \7208 , \6941 );
and \U$6833 ( \7210 , \7207 , \7209 );
and \U$6834 ( \7211 , \6950 , \7210 );
xor \U$6835 ( \7212 , \6950 , \7210 );
xor \U$6836 ( \7213 , \7207 , \7209 );
and \U$6837 ( \7214 , \4073 , \1058 );
and \U$6838 ( \7215 , \3951 , \1056 );
nor \U$6839 ( \7216 , \7214 , \7215 );
xnor \U$6840 ( \7217 , \7216 , \964 );
and \U$6841 ( \7218 , \4334 , \888 );
and \U$6842 ( \7219 , \4078 , \886 );
nor \U$6843 ( \7220 , \7218 , \7219 );
xnor \U$6844 ( \7221 , \7220 , \816 );
and \U$6845 ( \7222 , \7217 , \7221 );
and \U$6846 ( \7223 , \4833 , \754 );
and \U$6847 ( \7224 , \4531 , \752 );
nor \U$6848 ( \7225 , \7223 , \7224 );
xnor \U$6849 ( \7226 , \7225 , \711 );
and \U$6850 ( \7227 , \7221 , \7226 );
and \U$6851 ( \7228 , \7217 , \7226 );
or \U$6852 ( \7229 , \7222 , \7227 , \7228 );
and \U$6853 ( \7230 , \6562 , \422 );
and \U$6854 ( \7231 , \6219 , \420 );
nor \U$6855 ( \7232 , \7230 , \7231 );
xnor \U$6856 ( \7233 , \7232 , \403 );
and \U$6857 ( \7234 , \7067 , \385 );
and \U$6858 ( \7235 , \6764 , \383 );
nor \U$6859 ( \7236 , \7234 , \7235 );
xnor \U$6860 ( \7237 , \7236 , \390 );
and \U$6861 ( \7238 , \7233 , \7237 );
buf \U$6862 ( \7239 , RIc223fc8_116);
and \U$6863 ( \7240 , \7239 , \379 );
and \U$6864 ( \7241 , \7237 , \7240 );
and \U$6865 ( \7242 , \7233 , \7240 );
or \U$6866 ( \7243 , \7238 , \7241 , \7242 );
and \U$6867 ( \7244 , \7229 , \7243 );
and \U$6868 ( \7245 , \5310 , \641 );
and \U$6869 ( \7246 , \4841 , \639 );
nor \U$6870 ( \7247 , \7245 , \7246 );
xnor \U$6871 ( \7248 , \7247 , \592 );
and \U$6872 ( \7249 , \5579 , \540 );
and \U$6873 ( \7250 , \5315 , \538 );
nor \U$6874 ( \7251 , \7249 , \7250 );
xnor \U$6875 ( \7252 , \7251 , \499 );
and \U$6876 ( \7253 , \7248 , \7252 );
and \U$6877 ( \7254 , \6210 , \470 );
and \U$6878 ( \7255 , \5838 , \468 );
nor \U$6879 ( \7256 , \7254 , \7255 );
xnor \U$6880 ( \7257 , \7256 , \440 );
and \U$6881 ( \7258 , \7252 , \7257 );
and \U$6882 ( \7259 , \7248 , \7257 );
or \U$6883 ( \7260 , \7253 , \7258 , \7259 );
and \U$6884 ( \7261 , \7243 , \7260 );
and \U$6885 ( \7262 , \7229 , \7260 );
or \U$6886 ( \7263 , \7244 , \7261 , \7262 );
and \U$6887 ( \7264 , \556 , \5708 );
and \U$6888 ( \7265 , \487 , \5706 );
nor \U$6889 ( \7266 , \7264 , \7265 );
xnor \U$6890 ( \7267 , \7266 , \5467 );
and \U$6891 ( \7268 , \615 , \5242 );
and \U$6892 ( \7269 , \561 , \5240 );
nor \U$6893 ( \7270 , \7268 , \7269 );
xnor \U$6894 ( \7271 , \7270 , \5054 );
and \U$6895 ( \7272 , \7267 , \7271 );
and \U$6896 ( \7273 , \743 , \4868 );
and \U$6897 ( \7274 , \666 , \4866 );
nor \U$6898 ( \7275 , \7273 , \7274 );
xnor \U$6899 ( \7276 , \7275 , \4636 );
and \U$6900 ( \7277 , \7271 , \7276 );
and \U$6901 ( \7278 , \7267 , \7276 );
or \U$6902 ( \7279 , \7272 , \7277 , \7278 );
and \U$6903 ( \7280 , \851 , \4417 );
and \U$6904 ( \7281 , \771 , \4415 );
nor \U$6905 ( \7282 , \7280 , \7281 );
xnor \U$6906 ( \7283 , \7282 , \4274 );
and \U$6907 ( \7284 , \987 , \4094 );
and \U$6908 ( \7285 , \925 , \4092 );
nor \U$6909 ( \7286 , \7284 , \7285 );
xnor \U$6910 ( \7287 , \7286 , \3848 );
and \U$6911 ( \7288 , \7283 , \7287 );
and \U$6912 ( \7289 , \1248 , \3699 );
and \U$6913 ( \7290 , \1050 , \3697 );
nor \U$6914 ( \7291 , \7289 , \7290 );
xnor \U$6915 ( \7292 , \7291 , \3512 );
and \U$6916 ( \7293 , \7287 , \7292 );
and \U$6917 ( \7294 , \7283 , \7292 );
or \U$6918 ( \7295 , \7288 , \7293 , \7294 );
and \U$6919 ( \7296 , \7279 , \7295 );
xor \U$6920 ( \7297 , \6488 , \7036 );
xor \U$6921 ( \7298 , \7036 , \7037 );
not \U$6922 ( \7299 , \7298 );
and \U$6923 ( \7300 , \7297 , \7299 );
and \U$6924 ( \7301 , \378 , \7300 );
not \U$6925 ( \7302 , \7301 );
xnor \U$6926 ( \7303 , \7302 , \7040 );
and \U$6927 ( \7304 , \410 , \6806 );
and \U$6928 ( \7305 , \392 , \6804 );
nor \U$6929 ( \7306 , \7304 , \7305 );
xnor \U$6930 ( \7307 , \7306 , \6491 );
and \U$6931 ( \7308 , \7303 , \7307 );
and \U$6932 ( \7309 , \479 , \6297 );
and \U$6933 ( \7310 , \431 , \6295 );
nor \U$6934 ( \7311 , \7309 , \7310 );
xnor \U$6935 ( \7312 , \7311 , \5957 );
and \U$6936 ( \7313 , \7307 , \7312 );
and \U$6937 ( \7314 , \7303 , \7312 );
or \U$6938 ( \7315 , \7308 , \7313 , \7314 );
and \U$6939 ( \7316 , \7295 , \7315 );
and \U$6940 ( \7317 , \7279 , \7315 );
or \U$6941 ( \7318 , \7296 , \7316 , \7317 );
and \U$6942 ( \7319 , \7263 , \7318 );
and \U$6943 ( \7320 , \1441 , \3386 );
and \U$6944 ( \7321 , \1336 , \3384 );
nor \U$6945 ( \7322 , \7320 , \7321 );
xnor \U$6946 ( \7323 , \7322 , \3181 );
and \U$6947 ( \7324 , \1562 , \2980 );
and \U$6948 ( \7325 , \1446 , \2978 );
nor \U$6949 ( \7326 , \7324 , \7325 );
xnor \U$6950 ( \7327 , \7326 , \2831 );
and \U$6951 ( \7328 , \7323 , \7327 );
and \U$6952 ( \7329 , \1853 , \2658 );
and \U$6953 ( \7330 , \1677 , \2656 );
nor \U$6954 ( \7331 , \7329 , \7330 );
xnor \U$6955 ( \7332 , \7331 , \2516 );
and \U$6956 ( \7333 , \7327 , \7332 );
and \U$6957 ( \7334 , \7323 , \7332 );
or \U$6958 ( \7335 , \7328 , \7333 , \7334 );
and \U$6959 ( \7336 , \2104 , \2362 );
and \U$6960 ( \7337 , \1861 , \2360 );
nor \U$6961 ( \7338 , \7336 , \7337 );
xnor \U$6962 ( \7339 , \7338 , \2225 );
and \U$6963 ( \7340 , \2295 , \2156 );
and \U$6964 ( \7341 , \2109 , \2154 );
nor \U$6965 ( \7342 , \7340 , \7341 );
xnor \U$6966 ( \7343 , \7342 , \2004 );
and \U$6967 ( \7344 , \7339 , \7343 );
and \U$6968 ( \7345 , \2703 , \1888 );
and \U$6969 ( \7346 , \2439 , \1886 );
nor \U$6970 ( \7347 , \7345 , \7346 );
xnor \U$6971 ( \7348 , \7347 , \1732 );
and \U$6972 ( \7349 , \7343 , \7348 );
and \U$6973 ( \7350 , \7339 , \7348 );
or \U$6974 ( \7351 , \7344 , \7349 , \7350 );
and \U$6975 ( \7352 , \7335 , \7351 );
and \U$6976 ( \7353 , \2902 , \1616 );
and \U$6977 ( \7354 , \2728 , \1614 );
nor \U$6978 ( \7355 , \7353 , \7354 );
xnor \U$6979 ( \7356 , \7355 , \1503 );
and \U$6980 ( \7357 , \3207 , \1422 );
and \U$6981 ( \7358 , \3069 , \1420 );
nor \U$6982 ( \7359 , \7357 , \7358 );
xnor \U$6983 ( \7360 , \7359 , \1286 );
and \U$6984 ( \7361 , \7356 , \7360 );
and \U$6985 ( \7362 , \3743 , \1222 );
and \U$6986 ( \7363 , \3326 , \1220 );
nor \U$6987 ( \7364 , \7362 , \7363 );
xnor \U$6988 ( \7365 , \7364 , \1144 );
and \U$6989 ( \7366 , \7360 , \7365 );
and \U$6990 ( \7367 , \7356 , \7365 );
or \U$6991 ( \7368 , \7361 , \7366 , \7367 );
and \U$6992 ( \7369 , \7351 , \7368 );
and \U$6993 ( \7370 , \7335 , \7368 );
or \U$6994 ( \7371 , \7352 , \7369 , \7370 );
and \U$6995 ( \7372 , \7318 , \7371 );
and \U$6996 ( \7373 , \7263 , \7371 );
or \U$6997 ( \7374 , \7319 , \7372 , \7373 );
xor \U$6998 ( \7375 , \7061 , \7065 );
xor \U$6999 ( \7376 , \7375 , \7068 );
xor \U$7000 ( \7377 , \7075 , \7079 );
xor \U$7001 ( \7378 , \7377 , \7084 );
and \U$7002 ( \7379 , \7376 , \7378 );
xor \U$7003 ( \7380 , \7092 , \7096 );
xor \U$7004 ( \7381 , \7380 , \7101 );
and \U$7005 ( \7382 , \7378 , \7381 );
and \U$7006 ( \7383 , \7376 , \7381 );
or \U$7007 ( \7384 , \7379 , \7382 , \7383 );
xor \U$7008 ( \7385 , \6954 , \6958 );
xor \U$7009 ( \7386 , \7385 , \6963 );
xor \U$7010 ( \7387 , \6970 , \6974 );
xor \U$7011 ( \7388 , \7387 , \6979 );
and \U$7012 ( \7389 , \7386 , \7388 );
xor \U$7013 ( \7390 , \6987 , \6991 );
xor \U$7014 ( \7391 , \7390 , \6996 );
and \U$7015 ( \7392 , \7388 , \7391 );
and \U$7016 ( \7393 , \7386 , \7391 );
or \U$7017 ( \7394 , \7389 , \7392 , \7393 );
and \U$7018 ( \7395 , \7384 , \7394 );
xor \U$7019 ( \7396 , \7006 , \7010 );
xor \U$7020 ( \7397 , \7396 , \7015 );
xor \U$7021 ( \7398 , \7022 , \7026 );
xor \U$7022 ( \7399 , \7398 , \7031 );
and \U$7023 ( \7400 , \7397 , \7399 );
xor \U$7024 ( \7401 , \7041 , \7045 );
xor \U$7025 ( \7402 , \7401 , \7050 );
and \U$7026 ( \7403 , \7399 , \7402 );
and \U$7027 ( \7404 , \7397 , \7402 );
or \U$7028 ( \7405 , \7400 , \7403 , \7404 );
and \U$7029 ( \7406 , \7394 , \7405 );
and \U$7030 ( \7407 , \7384 , \7405 );
or \U$7031 ( \7408 , \7395 , \7406 , \7407 );
and \U$7032 ( \7409 , \7374 , \7408 );
xor \U$7033 ( \7410 , \7112 , \7114 );
xor \U$7034 ( \7411 , \7410 , \7117 );
xor \U$7035 ( \7412 , \7122 , \7124 );
xor \U$7036 ( \7413 , \7412 , \7127 );
and \U$7037 ( \7414 , \7411 , \7413 );
xor \U$7038 ( \7415 , \7133 , \7135 );
xor \U$7039 ( \7416 , \7415 , \7137 );
and \U$7040 ( \7417 , \7413 , \7416 );
and \U$7041 ( \7418 , \7411 , \7416 );
or \U$7042 ( \7419 , \7414 , \7417 , \7418 );
and \U$7043 ( \7420 , \7408 , \7419 );
and \U$7044 ( \7421 , \7374 , \7419 );
or \U$7045 ( \7422 , \7409 , \7420 , \7421 );
xor \U$7046 ( \7423 , \6966 , \6982 );
xor \U$7047 ( \7424 , \7423 , \6999 );
xor \U$7048 ( \7425 , \7018 , \7034 );
xor \U$7049 ( \7426 , \7425 , \7053 );
and \U$7050 ( \7427 , \7424 , \7426 );
xor \U$7051 ( \7428 , \7071 , \7087 );
xor \U$7052 ( \7429 , \7428 , \7104 );
and \U$7053 ( \7430 , \7426 , \7429 );
and \U$7054 ( \7431 , \7424 , \7429 );
or \U$7055 ( \7432 , \7427 , \7430 , \7431 );
xor \U$7056 ( \7433 , \7159 , \7161 );
xor \U$7057 ( \7434 , \7433 , \7164 );
and \U$7058 ( \7435 , \7432 , \7434 );
xor \U$7059 ( \7436 , \7146 , \7148 );
xor \U$7060 ( \7437 , \7436 , \7151 );
and \U$7061 ( \7438 , \7434 , \7437 );
and \U$7062 ( \7439 , \7432 , \7437 );
or \U$7063 ( \7440 , \7435 , \7438 , \7439 );
and \U$7064 ( \7441 , \7422 , \7440 );
xor \U$7065 ( \7442 , \7002 , \7056 );
xor \U$7066 ( \7443 , \7442 , \7107 );
xor \U$7067 ( \7444 , \7120 , \7130 );
xor \U$7068 ( \7445 , \7444 , \7140 );
and \U$7069 ( \7446 , \7443 , \7445 );
and \U$7070 ( \7447 , \7440 , \7446 );
and \U$7071 ( \7448 , \7422 , \7446 );
or \U$7072 ( \7449 , \7441 , \7447 , \7448 );
xor \U$7073 ( \7450 , \7110 , \7143 );
xor \U$7074 ( \7451 , \7450 , \7154 );
xor \U$7075 ( \7452 , \7167 , \7169 );
xor \U$7076 ( \7453 , \7452 , \7172 );
and \U$7077 ( \7454 , \7451 , \7453 );
xor \U$7078 ( \7455 , \7178 , \7180 );
and \U$7079 ( \7456 , \7453 , \7455 );
and \U$7080 ( \7457 , \7451 , \7455 );
or \U$7081 ( \7458 , \7454 , \7456 , \7457 );
and \U$7082 ( \7459 , \7449 , \7458 );
xor \U$7083 ( \7460 , \7186 , \7188 );
xor \U$7084 ( \7461 , \7460 , \7190 );
and \U$7085 ( \7462 , \7458 , \7461 );
and \U$7086 ( \7463 , \7449 , \7461 );
or \U$7087 ( \7464 , \7459 , \7462 , \7463 );
xor \U$7088 ( \7465 , \6894 , \6912 );
xor \U$7089 ( \7466 , \7465 , \6918 );
and \U$7090 ( \7467 , \7464 , \7466 );
xor \U$7091 ( \7468 , \7184 , \7193 );
xor \U$7092 ( \7469 , \7468 , \7196 );
and \U$7093 ( \7470 , \7466 , \7469 );
and \U$7094 ( \7471 , \7464 , \7469 );
or \U$7095 ( \7472 , \7467 , \7470 , \7471 );
xor \U$7096 ( \7473 , \7199 , \7201 );
xor \U$7097 ( \7474 , \7473 , \7204 );
and \U$7098 ( \7475 , \7472 , \7474 );
and \U$7099 ( \7476 , \7213 , \7475 );
xor \U$7100 ( \7477 , \7213 , \7475 );
xor \U$7101 ( \7478 , \7472 , \7474 );
xor \U$7102 ( \7479 , \7267 , \7271 );
xor \U$7103 ( \7480 , \7479 , \7276 );
xor \U$7104 ( \7481 , \7323 , \7327 );
xor \U$7105 ( \7482 , \7481 , \7332 );
and \U$7106 ( \7483 , \7480 , \7482 );
xor \U$7107 ( \7484 , \7283 , \7287 );
xor \U$7108 ( \7485 , \7484 , \7292 );
and \U$7109 ( \7486 , \7482 , \7485 );
and \U$7110 ( \7487 , \7480 , \7485 );
or \U$7111 ( \7488 , \7483 , \7486 , \7487 );
xor \U$7112 ( \7489 , \7339 , \7343 );
xor \U$7113 ( \7490 , \7489 , \7348 );
xor \U$7114 ( \7491 , \7217 , \7221 );
xor \U$7115 ( \7492 , \7491 , \7226 );
and \U$7116 ( \7493 , \7490 , \7492 );
xor \U$7117 ( \7494 , \7356 , \7360 );
xor \U$7118 ( \7495 , \7494 , \7365 );
and \U$7119 ( \7496 , \7492 , \7495 );
and \U$7120 ( \7497 , \7490 , \7495 );
or \U$7121 ( \7498 , \7493 , \7496 , \7497 );
and \U$7122 ( \7499 , \7488 , \7498 );
xor \U$7123 ( \7500 , \7233 , \7237 );
xor \U$7124 ( \7501 , \7500 , \7240 );
xor \U$7125 ( \7502 , \7248 , \7252 );
xor \U$7126 ( \7503 , \7502 , \7257 );
or \U$7127 ( \7504 , \7501 , \7503 );
and \U$7128 ( \7505 , \7498 , \7504 );
and \U$7129 ( \7506 , \7488 , \7504 );
or \U$7130 ( \7507 , \7499 , \7505 , \7506 );
and \U$7131 ( \7508 , \1861 , \2658 );
and \U$7132 ( \7509 , \1853 , \2656 );
nor \U$7133 ( \7510 , \7508 , \7509 );
xnor \U$7134 ( \7511 , \7510 , \2516 );
and \U$7135 ( \7512 , \2109 , \2362 );
and \U$7136 ( \7513 , \2104 , \2360 );
nor \U$7137 ( \7514 , \7512 , \7513 );
xnor \U$7138 ( \7515 , \7514 , \2225 );
and \U$7139 ( \7516 , \7511 , \7515 );
and \U$7140 ( \7517 , \2439 , \2156 );
and \U$7141 ( \7518 , \2295 , \2154 );
nor \U$7142 ( \7519 , \7517 , \7518 );
xnor \U$7143 ( \7520 , \7519 , \2004 );
and \U$7144 ( \7521 , \7515 , \7520 );
and \U$7145 ( \7522 , \7511 , \7520 );
or \U$7146 ( \7523 , \7516 , \7521 , \7522 );
and \U$7147 ( \7524 , \1336 , \3699 );
and \U$7148 ( \7525 , \1248 , \3697 );
nor \U$7149 ( \7526 , \7524 , \7525 );
xnor \U$7150 ( \7527 , \7526 , \3512 );
and \U$7151 ( \7528 , \1446 , \3386 );
and \U$7152 ( \7529 , \1441 , \3384 );
nor \U$7153 ( \7530 , \7528 , \7529 );
xnor \U$7154 ( \7531 , \7530 , \3181 );
and \U$7155 ( \7532 , \7527 , \7531 );
and \U$7156 ( \7533 , \1677 , \2980 );
and \U$7157 ( \7534 , \1562 , \2978 );
nor \U$7158 ( \7535 , \7533 , \7534 );
xnor \U$7159 ( \7536 , \7535 , \2831 );
and \U$7160 ( \7537 , \7531 , \7536 );
and \U$7161 ( \7538 , \7527 , \7536 );
or \U$7162 ( \7539 , \7532 , \7537 , \7538 );
and \U$7163 ( \7540 , \7523 , \7539 );
and \U$7164 ( \7541 , \2728 , \1888 );
and \U$7165 ( \7542 , \2703 , \1886 );
nor \U$7166 ( \7543 , \7541 , \7542 );
xnor \U$7167 ( \7544 , \7543 , \1732 );
and \U$7168 ( \7545 , \3069 , \1616 );
and \U$7169 ( \7546 , \2902 , \1614 );
nor \U$7170 ( \7547 , \7545 , \7546 );
xnor \U$7171 ( \7548 , \7547 , \1503 );
and \U$7172 ( \7549 , \7544 , \7548 );
and \U$7173 ( \7550 , \3326 , \1422 );
and \U$7174 ( \7551 , \3207 , \1420 );
nor \U$7175 ( \7552 , \7550 , \7551 );
xnor \U$7176 ( \7553 , \7552 , \1286 );
and \U$7177 ( \7554 , \7548 , \7553 );
and \U$7178 ( \7555 , \7544 , \7553 );
or \U$7179 ( \7556 , \7549 , \7554 , \7555 );
and \U$7180 ( \7557 , \7539 , \7556 );
and \U$7181 ( \7558 , \7523 , \7556 );
or \U$7182 ( \7559 , \7540 , \7557 , \7558 );
and \U$7183 ( \7560 , \487 , \6297 );
and \U$7184 ( \7561 , \479 , \6295 );
nor \U$7185 ( \7562 , \7560 , \7561 );
xnor \U$7186 ( \7563 , \7562 , \5957 );
and \U$7187 ( \7564 , \561 , \5708 );
and \U$7188 ( \7565 , \556 , \5706 );
nor \U$7189 ( \7566 , \7564 , \7565 );
xnor \U$7190 ( \7567 , \7566 , \5467 );
and \U$7191 ( \7568 , \7563 , \7567 );
and \U$7192 ( \7569 , \666 , \5242 );
and \U$7193 ( \7570 , \615 , \5240 );
nor \U$7194 ( \7571 , \7569 , \7570 );
xnor \U$7195 ( \7572 , \7571 , \5054 );
and \U$7196 ( \7573 , \7567 , \7572 );
and \U$7197 ( \7574 , \7563 , \7572 );
or \U$7198 ( \7575 , \7568 , \7573 , \7574 );
buf \U$7199 ( \7576 , RIc225cd8_54);
buf \U$7200 ( \7577 , RIc225c60_55);
and \U$7201 ( \7578 , \7576 , \7577 );
not \U$7202 ( \7579 , \7578 );
and \U$7203 ( \7580 , \7037 , \7579 );
not \U$7204 ( \7581 , \7580 );
and \U$7205 ( \7582 , \392 , \7300 );
and \U$7206 ( \7583 , \378 , \7298 );
nor \U$7207 ( \7584 , \7582 , \7583 );
xnor \U$7208 ( \7585 , \7584 , \7040 );
and \U$7209 ( \7586 , \7581 , \7585 );
and \U$7210 ( \7587 , \431 , \6806 );
and \U$7211 ( \7588 , \410 , \6804 );
nor \U$7212 ( \7589 , \7587 , \7588 );
xnor \U$7213 ( \7590 , \7589 , \6491 );
and \U$7214 ( \7591 , \7585 , \7590 );
and \U$7215 ( \7592 , \7581 , \7590 );
or \U$7216 ( \7593 , \7586 , \7591 , \7592 );
and \U$7217 ( \7594 , \7575 , \7593 );
and \U$7218 ( \7595 , \771 , \4868 );
and \U$7219 ( \7596 , \743 , \4866 );
nor \U$7220 ( \7597 , \7595 , \7596 );
xnor \U$7221 ( \7598 , \7597 , \4636 );
and \U$7222 ( \7599 , \925 , \4417 );
and \U$7223 ( \7600 , \851 , \4415 );
nor \U$7224 ( \7601 , \7599 , \7600 );
xnor \U$7225 ( \7602 , \7601 , \4274 );
and \U$7226 ( \7603 , \7598 , \7602 );
and \U$7227 ( \7604 , \1050 , \4094 );
and \U$7228 ( \7605 , \987 , \4092 );
nor \U$7229 ( \7606 , \7604 , \7605 );
xnor \U$7230 ( \7607 , \7606 , \3848 );
and \U$7231 ( \7608 , \7602 , \7607 );
and \U$7232 ( \7609 , \7598 , \7607 );
or \U$7233 ( \7610 , \7603 , \7608 , \7609 );
and \U$7234 ( \7611 , \7593 , \7610 );
and \U$7235 ( \7612 , \7575 , \7610 );
or \U$7236 ( \7613 , \7594 , \7611 , \7612 );
and \U$7237 ( \7614 , \7559 , \7613 );
and \U$7238 ( \7615 , \3951 , \1222 );
and \U$7239 ( \7616 , \3743 , \1220 );
nor \U$7240 ( \7617 , \7615 , \7616 );
xnor \U$7241 ( \7618 , \7617 , \1144 );
and \U$7242 ( \7619 , \4078 , \1058 );
and \U$7243 ( \7620 , \4073 , \1056 );
nor \U$7244 ( \7621 , \7619 , \7620 );
xnor \U$7245 ( \7622 , \7621 , \964 );
and \U$7246 ( \7623 , \7618 , \7622 );
and \U$7247 ( \7624 , \4531 , \888 );
and \U$7248 ( \7625 , \4334 , \886 );
nor \U$7249 ( \7626 , \7624 , \7625 );
xnor \U$7250 ( \7627 , \7626 , \816 );
and \U$7251 ( \7628 , \7622 , \7627 );
and \U$7252 ( \7629 , \7618 , \7627 );
or \U$7253 ( \7630 , \7623 , \7628 , \7629 );
and \U$7254 ( \7631 , \4841 , \754 );
and \U$7255 ( \7632 , \4833 , \752 );
nor \U$7256 ( \7633 , \7631 , \7632 );
xnor \U$7257 ( \7634 , \7633 , \711 );
and \U$7258 ( \7635 , \5315 , \641 );
and \U$7259 ( \7636 , \5310 , \639 );
nor \U$7260 ( \7637 , \7635 , \7636 );
xnor \U$7261 ( \7638 , \7637 , \592 );
and \U$7262 ( \7639 , \7634 , \7638 );
and \U$7263 ( \7640 , \5838 , \540 );
and \U$7264 ( \7641 , \5579 , \538 );
nor \U$7265 ( \7642 , \7640 , \7641 );
xnor \U$7266 ( \7643 , \7642 , \499 );
and \U$7267 ( \7644 , \7638 , \7643 );
and \U$7268 ( \7645 , \7634 , \7643 );
or \U$7269 ( \7646 , \7639 , \7644 , \7645 );
and \U$7270 ( \7647 , \7630 , \7646 );
and \U$7271 ( \7648 , \6219 , \470 );
and \U$7272 ( \7649 , \6210 , \468 );
nor \U$7273 ( \7650 , \7648 , \7649 );
xnor \U$7274 ( \7651 , \7650 , \440 );
and \U$7275 ( \7652 , \6764 , \422 );
and \U$7276 ( \7653 , \6562 , \420 );
nor \U$7277 ( \7654 , \7652 , \7653 );
xnor \U$7278 ( \7655 , \7654 , \403 );
and \U$7279 ( \7656 , \7651 , \7655 );
and \U$7280 ( \7657 , \7239 , \385 );
and \U$7281 ( \7658 , \7067 , \383 );
nor \U$7282 ( \7659 , \7657 , \7658 );
xnor \U$7283 ( \7660 , \7659 , \390 );
and \U$7284 ( \7661 , \7655 , \7660 );
and \U$7285 ( \7662 , \7651 , \7660 );
or \U$7286 ( \7663 , \7656 , \7661 , \7662 );
and \U$7287 ( \7664 , \7646 , \7663 );
and \U$7288 ( \7665 , \7630 , \7663 );
or \U$7289 ( \7666 , \7647 , \7664 , \7665 );
and \U$7290 ( \7667 , \7613 , \7666 );
and \U$7291 ( \7668 , \7559 , \7666 );
or \U$7292 ( \7669 , \7614 , \7667 , \7668 );
and \U$7293 ( \7670 , \7507 , \7669 );
xor \U$7294 ( \7671 , \7376 , \7378 );
xor \U$7295 ( \7672 , \7671 , \7381 );
xor \U$7296 ( \7673 , \7386 , \7388 );
xor \U$7297 ( \7674 , \7673 , \7391 );
and \U$7298 ( \7675 , \7672 , \7674 );
xor \U$7299 ( \7676 , \7397 , \7399 );
xor \U$7300 ( \7677 , \7676 , \7402 );
and \U$7301 ( \7678 , \7674 , \7677 );
and \U$7302 ( \7679 , \7672 , \7677 );
or \U$7303 ( \7680 , \7675 , \7678 , \7679 );
and \U$7304 ( \7681 , \7669 , \7680 );
and \U$7305 ( \7682 , \7507 , \7680 );
or \U$7306 ( \7683 , \7670 , \7681 , \7682 );
xor \U$7307 ( \7684 , \7229 , \7243 );
xor \U$7308 ( \7685 , \7684 , \7260 );
xor \U$7309 ( \7686 , \7279 , \7295 );
xor \U$7310 ( \7687 , \7686 , \7315 );
and \U$7311 ( \7688 , \7685 , \7687 );
xor \U$7312 ( \7689 , \7335 , \7351 );
xor \U$7313 ( \7690 , \7689 , \7368 );
and \U$7314 ( \7691 , \7687 , \7690 );
and \U$7315 ( \7692 , \7685 , \7690 );
or \U$7316 ( \7693 , \7688 , \7691 , \7692 );
xor \U$7317 ( \7694 , \7424 , \7426 );
xor \U$7318 ( \7695 , \7694 , \7429 );
and \U$7319 ( \7696 , \7693 , \7695 );
xor \U$7320 ( \7697 , \7411 , \7413 );
xor \U$7321 ( \7698 , \7697 , \7416 );
and \U$7322 ( \7699 , \7695 , \7698 );
and \U$7323 ( \7700 , \7693 , \7698 );
or \U$7324 ( \7701 , \7696 , \7699 , \7700 );
and \U$7325 ( \7702 , \7683 , \7701 );
xor \U$7326 ( \7703 , \7263 , \7318 );
xor \U$7327 ( \7704 , \7703 , \7371 );
xor \U$7328 ( \7705 , \7384 , \7394 );
xor \U$7329 ( \7706 , \7705 , \7405 );
and \U$7330 ( \7707 , \7704 , \7706 );
and \U$7331 ( \7708 , \7701 , \7707 );
and \U$7332 ( \7709 , \7683 , \7707 );
or \U$7333 ( \7710 , \7702 , \7708 , \7709 );
xor \U$7334 ( \7711 , \7374 , \7408 );
xor \U$7335 ( \7712 , \7711 , \7419 );
xor \U$7336 ( \7713 , \7432 , \7434 );
xor \U$7337 ( \7714 , \7713 , \7437 );
and \U$7338 ( \7715 , \7712 , \7714 );
xor \U$7339 ( \7716 , \7443 , \7445 );
and \U$7340 ( \7717 , \7714 , \7716 );
and \U$7341 ( \7718 , \7712 , \7716 );
or \U$7342 ( \7719 , \7715 , \7717 , \7718 );
and \U$7343 ( \7720 , \7710 , \7719 );
xor \U$7344 ( \7721 , \7451 , \7453 );
xor \U$7345 ( \7722 , \7721 , \7455 );
and \U$7346 ( \7723 , \7719 , \7722 );
and \U$7347 ( \7724 , \7710 , \7722 );
or \U$7348 ( \7725 , \7720 , \7723 , \7724 );
xor \U$7349 ( \7726 , \7157 , \7175 );
xor \U$7350 ( \7727 , \7726 , \7181 );
and \U$7351 ( \7728 , \7725 , \7727 );
xor \U$7352 ( \7729 , \7449 , \7458 );
xor \U$7353 ( \7730 , \7729 , \7461 );
and \U$7354 ( \7731 , \7727 , \7730 );
and \U$7355 ( \7732 , \7725 , \7730 );
or \U$7356 ( \7733 , \7728 , \7731 , \7732 );
xor \U$7357 ( \7734 , \7464 , \7466 );
xor \U$7358 ( \7735 , \7734 , \7469 );
and \U$7359 ( \7736 , \7733 , \7735 );
and \U$7360 ( \7737 , \7478 , \7736 );
xor \U$7361 ( \7738 , \7478 , \7736 );
xor \U$7362 ( \7739 , \7733 , \7735 );
and \U$7363 ( \7740 , \4073 , \1222 );
and \U$7364 ( \7741 , \3951 , \1220 );
nor \U$7365 ( \7742 , \7740 , \7741 );
xnor \U$7366 ( \7743 , \7742 , \1144 );
and \U$7367 ( \7744 , \4334 , \1058 );
and \U$7368 ( \7745 , \4078 , \1056 );
nor \U$7369 ( \7746 , \7744 , \7745 );
xnor \U$7370 ( \7747 , \7746 , \964 );
and \U$7371 ( \7748 , \7743 , \7747 );
and \U$7372 ( \7749 , \4833 , \888 );
and \U$7373 ( \7750 , \4531 , \886 );
nor \U$7374 ( \7751 , \7749 , \7750 );
xnor \U$7375 ( \7752 , \7751 , \816 );
and \U$7376 ( \7753 , \7747 , \7752 );
and \U$7377 ( \7754 , \7743 , \7752 );
or \U$7378 ( \7755 , \7748 , \7753 , \7754 );
and \U$7379 ( \7756 , \6562 , \470 );
and \U$7380 ( \7757 , \6219 , \468 );
nor \U$7381 ( \7758 , \7756 , \7757 );
xnor \U$7382 ( \7759 , \7758 , \440 );
and \U$7383 ( \7760 , \7067 , \422 );
and \U$7384 ( \7761 , \6764 , \420 );
nor \U$7385 ( \7762 , \7760 , \7761 );
xnor \U$7386 ( \7763 , \7762 , \403 );
and \U$7387 ( \7764 , \7759 , \7763 );
buf \U$7388 ( \7765 , RIc223f50_117);
and \U$7389 ( \7766 , \7765 , \385 );
and \U$7390 ( \7767 , \7239 , \383 );
nor \U$7391 ( \7768 , \7766 , \7767 );
xnor \U$7392 ( \7769 , \7768 , \390 );
and \U$7393 ( \7770 , \7763 , \7769 );
and \U$7394 ( \7771 , \7759 , \7769 );
or \U$7395 ( \7772 , \7764 , \7770 , \7771 );
and \U$7396 ( \7773 , \7755 , \7772 );
and \U$7397 ( \7774 , \5310 , \754 );
and \U$7398 ( \7775 , \4841 , \752 );
nor \U$7399 ( \7776 , \7774 , \7775 );
xnor \U$7400 ( \7777 , \7776 , \711 );
and \U$7401 ( \7778 , \5579 , \641 );
and \U$7402 ( \7779 , \5315 , \639 );
nor \U$7403 ( \7780 , \7778 , \7779 );
xnor \U$7404 ( \7781 , \7780 , \592 );
and \U$7405 ( \7782 , \7777 , \7781 );
and \U$7406 ( \7783 , \6210 , \540 );
and \U$7407 ( \7784 , \5838 , \538 );
nor \U$7408 ( \7785 , \7783 , \7784 );
xnor \U$7409 ( \7786 , \7785 , \499 );
and \U$7410 ( \7787 , \7781 , \7786 );
and \U$7411 ( \7788 , \7777 , \7786 );
or \U$7412 ( \7789 , \7782 , \7787 , \7788 );
and \U$7413 ( \7790 , \7772 , \7789 );
and \U$7414 ( \7791 , \7755 , \7789 );
or \U$7415 ( \7792 , \7773 , \7790 , \7791 );
and \U$7416 ( \7793 , \556 , \6297 );
and \U$7417 ( \7794 , \487 , \6295 );
nor \U$7418 ( \7795 , \7793 , \7794 );
xnor \U$7419 ( \7796 , \7795 , \5957 );
and \U$7420 ( \7797 , \615 , \5708 );
and \U$7421 ( \7798 , \561 , \5706 );
nor \U$7422 ( \7799 , \7797 , \7798 );
xnor \U$7423 ( \7800 , \7799 , \5467 );
and \U$7424 ( \7801 , \7796 , \7800 );
and \U$7425 ( \7802 , \743 , \5242 );
and \U$7426 ( \7803 , \666 , \5240 );
nor \U$7427 ( \7804 , \7802 , \7803 );
xnor \U$7428 ( \7805 , \7804 , \5054 );
and \U$7429 ( \7806 , \7800 , \7805 );
and \U$7430 ( \7807 , \7796 , \7805 );
or \U$7431 ( \7808 , \7801 , \7806 , \7807 );
and \U$7432 ( \7809 , \851 , \4868 );
and \U$7433 ( \7810 , \771 , \4866 );
nor \U$7434 ( \7811 , \7809 , \7810 );
xnor \U$7435 ( \7812 , \7811 , \4636 );
and \U$7436 ( \7813 , \987 , \4417 );
and \U$7437 ( \7814 , \925 , \4415 );
nor \U$7438 ( \7815 , \7813 , \7814 );
xnor \U$7439 ( \7816 , \7815 , \4274 );
and \U$7440 ( \7817 , \7812 , \7816 );
and \U$7441 ( \7818 , \1248 , \4094 );
and \U$7442 ( \7819 , \1050 , \4092 );
nor \U$7443 ( \7820 , \7818 , \7819 );
xnor \U$7444 ( \7821 , \7820 , \3848 );
and \U$7445 ( \7822 , \7816 , \7821 );
and \U$7446 ( \7823 , \7812 , \7821 );
or \U$7447 ( \7824 , \7817 , \7822 , \7823 );
and \U$7448 ( \7825 , \7808 , \7824 );
xor \U$7449 ( \7826 , \7037 , \7576 );
xor \U$7450 ( \7827 , \7576 , \7577 );
not \U$7451 ( \7828 , \7827 );
and \U$7452 ( \7829 , \7826 , \7828 );
and \U$7453 ( \7830 , \378 , \7829 );
not \U$7454 ( \7831 , \7830 );
xnor \U$7455 ( \7832 , \7831 , \7580 );
and \U$7456 ( \7833 , \410 , \7300 );
and \U$7457 ( \7834 , \392 , \7298 );
nor \U$7458 ( \7835 , \7833 , \7834 );
xnor \U$7459 ( \7836 , \7835 , \7040 );
and \U$7460 ( \7837 , \7832 , \7836 );
and \U$7461 ( \7838 , \479 , \6806 );
and \U$7462 ( \7839 , \431 , \6804 );
nor \U$7463 ( \7840 , \7838 , \7839 );
xnor \U$7464 ( \7841 , \7840 , \6491 );
and \U$7465 ( \7842 , \7836 , \7841 );
and \U$7466 ( \7843 , \7832 , \7841 );
or \U$7467 ( \7844 , \7837 , \7842 , \7843 );
and \U$7468 ( \7845 , \7824 , \7844 );
and \U$7469 ( \7846 , \7808 , \7844 );
or \U$7470 ( \7847 , \7825 , \7845 , \7846 );
and \U$7471 ( \7848 , \7792 , \7847 );
and \U$7472 ( \7849 , \2902 , \1888 );
and \U$7473 ( \7850 , \2728 , \1886 );
nor \U$7474 ( \7851 , \7849 , \7850 );
xnor \U$7475 ( \7852 , \7851 , \1732 );
and \U$7476 ( \7853 , \3207 , \1616 );
and \U$7477 ( \7854 , \3069 , \1614 );
nor \U$7478 ( \7855 , \7853 , \7854 );
xnor \U$7479 ( \7856 , \7855 , \1503 );
and \U$7480 ( \7857 , \7852 , \7856 );
and \U$7481 ( \7858 , \3743 , \1422 );
and \U$7482 ( \7859 , \3326 , \1420 );
nor \U$7483 ( \7860 , \7858 , \7859 );
xnor \U$7484 ( \7861 , \7860 , \1286 );
and \U$7485 ( \7862 , \7856 , \7861 );
and \U$7486 ( \7863 , \7852 , \7861 );
or \U$7487 ( \7864 , \7857 , \7862 , \7863 );
and \U$7488 ( \7865 , \1441 , \3699 );
and \U$7489 ( \7866 , \1336 , \3697 );
nor \U$7490 ( \7867 , \7865 , \7866 );
xnor \U$7491 ( \7868 , \7867 , \3512 );
and \U$7492 ( \7869 , \1562 , \3386 );
and \U$7493 ( \7870 , \1446 , \3384 );
nor \U$7494 ( \7871 , \7869 , \7870 );
xnor \U$7495 ( \7872 , \7871 , \3181 );
and \U$7496 ( \7873 , \7868 , \7872 );
and \U$7497 ( \7874 , \1853 , \2980 );
and \U$7498 ( \7875 , \1677 , \2978 );
nor \U$7499 ( \7876 , \7874 , \7875 );
xnor \U$7500 ( \7877 , \7876 , \2831 );
and \U$7501 ( \7878 , \7872 , \7877 );
and \U$7502 ( \7879 , \7868 , \7877 );
or \U$7503 ( \7880 , \7873 , \7878 , \7879 );
and \U$7504 ( \7881 , \7864 , \7880 );
and \U$7505 ( \7882 , \2104 , \2658 );
and \U$7506 ( \7883 , \1861 , \2656 );
nor \U$7507 ( \7884 , \7882 , \7883 );
xnor \U$7508 ( \7885 , \7884 , \2516 );
and \U$7509 ( \7886 , \2295 , \2362 );
and \U$7510 ( \7887 , \2109 , \2360 );
nor \U$7511 ( \7888 , \7886 , \7887 );
xnor \U$7512 ( \7889 , \7888 , \2225 );
and \U$7513 ( \7890 , \7885 , \7889 );
and \U$7514 ( \7891 , \2703 , \2156 );
and \U$7515 ( \7892 , \2439 , \2154 );
nor \U$7516 ( \7893 , \7891 , \7892 );
xnor \U$7517 ( \7894 , \7893 , \2004 );
and \U$7518 ( \7895 , \7889 , \7894 );
and \U$7519 ( \7896 , \7885 , \7894 );
or \U$7520 ( \7897 , \7890 , \7895 , \7896 );
and \U$7521 ( \7898 , \7880 , \7897 );
and \U$7522 ( \7899 , \7864 , \7897 );
or \U$7523 ( \7900 , \7881 , \7898 , \7899 );
and \U$7524 ( \7901 , \7847 , \7900 );
and \U$7525 ( \7902 , \7792 , \7900 );
or \U$7526 ( \7903 , \7848 , \7901 , \7902 );
xor \U$7527 ( \7904 , \7563 , \7567 );
xor \U$7528 ( \7905 , \7904 , \7572 );
xor \U$7529 ( \7906 , \7527 , \7531 );
xor \U$7530 ( \7907 , \7906 , \7536 );
and \U$7531 ( \7908 , \7905 , \7907 );
xor \U$7532 ( \7909 , \7598 , \7602 );
xor \U$7533 ( \7910 , \7909 , \7607 );
and \U$7534 ( \7911 , \7907 , \7910 );
and \U$7535 ( \7912 , \7905 , \7910 );
or \U$7536 ( \7913 , \7908 , \7911 , \7912 );
and \U$7537 ( \7914 , \7765 , \379 );
xor \U$7538 ( \7915 , \7634 , \7638 );
xor \U$7539 ( \7916 , \7915 , \7643 );
and \U$7540 ( \7917 , \7914 , \7916 );
xor \U$7541 ( \7918 , \7651 , \7655 );
xor \U$7542 ( \7919 , \7918 , \7660 );
and \U$7543 ( \7920 , \7916 , \7919 );
and \U$7544 ( \7921 , \7914 , \7919 );
or \U$7545 ( \7922 , \7917 , \7920 , \7921 );
and \U$7546 ( \7923 , \7913 , \7922 );
xor \U$7547 ( \7924 , \7618 , \7622 );
xor \U$7548 ( \7925 , \7924 , \7627 );
xor \U$7549 ( \7926 , \7511 , \7515 );
xor \U$7550 ( \7927 , \7926 , \7520 );
and \U$7551 ( \7928 , \7925 , \7927 );
xor \U$7552 ( \7929 , \7544 , \7548 );
xor \U$7553 ( \7930 , \7929 , \7553 );
and \U$7554 ( \7931 , \7927 , \7930 );
and \U$7555 ( \7932 , \7925 , \7930 );
or \U$7556 ( \7933 , \7928 , \7931 , \7932 );
and \U$7557 ( \7934 , \7922 , \7933 );
and \U$7558 ( \7935 , \7913 , \7933 );
or \U$7559 ( \7936 , \7923 , \7934 , \7935 );
and \U$7560 ( \7937 , \7903 , \7936 );
xor \U$7561 ( \7938 , \7303 , \7307 );
xor \U$7562 ( \7939 , \7938 , \7312 );
xor \U$7563 ( \7940 , \7480 , \7482 );
xor \U$7564 ( \7941 , \7940 , \7485 );
and \U$7565 ( \7942 , \7939 , \7941 );
xor \U$7566 ( \7943 , \7490 , \7492 );
xor \U$7567 ( \7944 , \7943 , \7495 );
and \U$7568 ( \7945 , \7941 , \7944 );
and \U$7569 ( \7946 , \7939 , \7944 );
or \U$7570 ( \7947 , \7942 , \7945 , \7946 );
and \U$7571 ( \7948 , \7936 , \7947 );
and \U$7572 ( \7949 , \7903 , \7947 );
or \U$7573 ( \7950 , \7937 , \7948 , \7949 );
xor \U$7574 ( \7951 , \7523 , \7539 );
xor \U$7575 ( \7952 , \7951 , \7556 );
xor \U$7576 ( \7953 , \7630 , \7646 );
xor \U$7577 ( \7954 , \7953 , \7663 );
and \U$7578 ( \7955 , \7952 , \7954 );
xnor \U$7579 ( \7956 , \7501 , \7503 );
and \U$7580 ( \7957 , \7954 , \7956 );
and \U$7581 ( \7958 , \7952 , \7956 );
or \U$7582 ( \7959 , \7955 , \7957 , \7958 );
xor \U$7583 ( \7960 , \7685 , \7687 );
xor \U$7584 ( \7961 , \7960 , \7690 );
and \U$7585 ( \7962 , \7959 , \7961 );
xor \U$7586 ( \7963 , \7672 , \7674 );
xor \U$7587 ( \7964 , \7963 , \7677 );
and \U$7588 ( \7965 , \7961 , \7964 );
and \U$7589 ( \7966 , \7959 , \7964 );
or \U$7590 ( \7967 , \7962 , \7965 , \7966 );
and \U$7591 ( \7968 , \7950 , \7967 );
xor \U$7592 ( \7969 , \7488 , \7498 );
xor \U$7593 ( \7970 , \7969 , \7504 );
xor \U$7594 ( \7971 , \7559 , \7613 );
xor \U$7595 ( \7972 , \7971 , \7666 );
and \U$7596 ( \7973 , \7970 , \7972 );
and \U$7597 ( \7974 , \7967 , \7973 );
and \U$7598 ( \7975 , \7950 , \7973 );
or \U$7599 ( \7976 , \7968 , \7974 , \7975 );
xor \U$7600 ( \7977 , \7507 , \7669 );
xor \U$7601 ( \7978 , \7977 , \7680 );
xor \U$7602 ( \7979 , \7693 , \7695 );
xor \U$7603 ( \7980 , \7979 , \7698 );
and \U$7604 ( \7981 , \7978 , \7980 );
xor \U$7605 ( \7982 , \7704 , \7706 );
and \U$7606 ( \7983 , \7980 , \7982 );
and \U$7607 ( \7984 , \7978 , \7982 );
or \U$7608 ( \7985 , \7981 , \7983 , \7984 );
and \U$7609 ( \7986 , \7976 , \7985 );
xor \U$7610 ( \7987 , \7712 , \7714 );
xor \U$7611 ( \7988 , \7987 , \7716 );
and \U$7612 ( \7989 , \7985 , \7988 );
and \U$7613 ( \7990 , \7976 , \7988 );
or \U$7614 ( \7991 , \7986 , \7989 , \7990 );
xor \U$7615 ( \7992 , \7422 , \7440 );
xor \U$7616 ( \7993 , \7992 , \7446 );
and \U$7617 ( \7994 , \7991 , \7993 );
xor \U$7618 ( \7995 , \7710 , \7719 );
xor \U$7619 ( \7996 , \7995 , \7722 );
and \U$7620 ( \7997 , \7993 , \7996 );
and \U$7621 ( \7998 , \7991 , \7996 );
or \U$7622 ( \7999 , \7994 , \7997 , \7998 );
xor \U$7623 ( \8000 , \7725 , \7727 );
xor \U$7624 ( \8001 , \8000 , \7730 );
and \U$7625 ( \8002 , \7999 , \8001 );
and \U$7626 ( \8003 , \7739 , \8002 );
xor \U$7627 ( \8004 , \7739 , \8002 );
xor \U$7628 ( \8005 , \7999 , \8001 );
and \U$7629 ( \8006 , \2728 , \2156 );
and \U$7630 ( \8007 , \2703 , \2154 );
nor \U$7631 ( \8008 , \8006 , \8007 );
xnor \U$7632 ( \8009 , \8008 , \2004 );
and \U$7633 ( \8010 , \3069 , \1888 );
and \U$7634 ( \8011 , \2902 , \1886 );
nor \U$7635 ( \8012 , \8010 , \8011 );
xnor \U$7636 ( \8013 , \8012 , \1732 );
and \U$7637 ( \8014 , \8009 , \8013 );
and \U$7638 ( \8015 , \3326 , \1616 );
and \U$7639 ( \8016 , \3207 , \1614 );
nor \U$7640 ( \8017 , \8015 , \8016 );
xnor \U$7641 ( \8018 , \8017 , \1503 );
and \U$7642 ( \8019 , \8013 , \8018 );
and \U$7643 ( \8020 , \8009 , \8018 );
or \U$7644 ( \8021 , \8014 , \8019 , \8020 );
and \U$7645 ( \8022 , \1336 , \4094 );
and \U$7646 ( \8023 , \1248 , \4092 );
nor \U$7647 ( \8024 , \8022 , \8023 );
xnor \U$7648 ( \8025 , \8024 , \3848 );
and \U$7649 ( \8026 , \1446 , \3699 );
and \U$7650 ( \8027 , \1441 , \3697 );
nor \U$7651 ( \8028 , \8026 , \8027 );
xnor \U$7652 ( \8029 , \8028 , \3512 );
and \U$7653 ( \8030 , \8025 , \8029 );
and \U$7654 ( \8031 , \1677 , \3386 );
and \U$7655 ( \8032 , \1562 , \3384 );
nor \U$7656 ( \8033 , \8031 , \8032 );
xnor \U$7657 ( \8034 , \8033 , \3181 );
and \U$7658 ( \8035 , \8029 , \8034 );
and \U$7659 ( \8036 , \8025 , \8034 );
or \U$7660 ( \8037 , \8030 , \8035 , \8036 );
and \U$7661 ( \8038 , \8021 , \8037 );
and \U$7662 ( \8039 , \1861 , \2980 );
and \U$7663 ( \8040 , \1853 , \2978 );
nor \U$7664 ( \8041 , \8039 , \8040 );
xnor \U$7665 ( \8042 , \8041 , \2831 );
and \U$7666 ( \8043 , \2109 , \2658 );
and \U$7667 ( \8044 , \2104 , \2656 );
nor \U$7668 ( \8045 , \8043 , \8044 );
xnor \U$7669 ( \8046 , \8045 , \2516 );
and \U$7670 ( \8047 , \8042 , \8046 );
and \U$7671 ( \8048 , \2439 , \2362 );
and \U$7672 ( \8049 , \2295 , \2360 );
nor \U$7673 ( \8050 , \8048 , \8049 );
xnor \U$7674 ( \8051 , \8050 , \2225 );
and \U$7675 ( \8052 , \8046 , \8051 );
and \U$7676 ( \8053 , \8042 , \8051 );
or \U$7677 ( \8054 , \8047 , \8052 , \8053 );
and \U$7678 ( \8055 , \8037 , \8054 );
and \U$7679 ( \8056 , \8021 , \8054 );
or \U$7680 ( \8057 , \8038 , \8055 , \8056 );
and \U$7681 ( \8058 , \771 , \5242 );
and \U$7682 ( \8059 , \743 , \5240 );
nor \U$7683 ( \8060 , \8058 , \8059 );
xnor \U$7684 ( \8061 , \8060 , \5054 );
and \U$7685 ( \8062 , \925 , \4868 );
and \U$7686 ( \8063 , \851 , \4866 );
nor \U$7687 ( \8064 , \8062 , \8063 );
xnor \U$7688 ( \8065 , \8064 , \4636 );
and \U$7689 ( \8066 , \8061 , \8065 );
and \U$7690 ( \8067 , \1050 , \4417 );
and \U$7691 ( \8068 , \987 , \4415 );
nor \U$7692 ( \8069 , \8067 , \8068 );
xnor \U$7693 ( \8070 , \8069 , \4274 );
and \U$7694 ( \8071 , \8065 , \8070 );
and \U$7695 ( \8072 , \8061 , \8070 );
or \U$7696 ( \8073 , \8066 , \8071 , \8072 );
buf \U$7697 ( \8074 , RIc225be8_56);
buf \U$7698 ( \8075 , RIc225b70_57);
and \U$7699 ( \8076 , \8074 , \8075 );
not \U$7700 ( \8077 , \8076 );
and \U$7701 ( \8078 , \7577 , \8077 );
not \U$7702 ( \8079 , \8078 );
and \U$7703 ( \8080 , \392 , \7829 );
and \U$7704 ( \8081 , \378 , \7827 );
nor \U$7705 ( \8082 , \8080 , \8081 );
xnor \U$7706 ( \8083 , \8082 , \7580 );
and \U$7707 ( \8084 , \8079 , \8083 );
and \U$7708 ( \8085 , \431 , \7300 );
and \U$7709 ( \8086 , \410 , \7298 );
nor \U$7710 ( \8087 , \8085 , \8086 );
xnor \U$7711 ( \8088 , \8087 , \7040 );
and \U$7712 ( \8089 , \8083 , \8088 );
and \U$7713 ( \8090 , \8079 , \8088 );
or \U$7714 ( \8091 , \8084 , \8089 , \8090 );
and \U$7715 ( \8092 , \8073 , \8091 );
and \U$7716 ( \8093 , \487 , \6806 );
and \U$7717 ( \8094 , \479 , \6804 );
nor \U$7718 ( \8095 , \8093 , \8094 );
xnor \U$7719 ( \8096 , \8095 , \6491 );
and \U$7720 ( \8097 , \561 , \6297 );
and \U$7721 ( \8098 , \556 , \6295 );
nor \U$7722 ( \8099 , \8097 , \8098 );
xnor \U$7723 ( \8100 , \8099 , \5957 );
and \U$7724 ( \8101 , \8096 , \8100 );
and \U$7725 ( \8102 , \666 , \5708 );
and \U$7726 ( \8103 , \615 , \5706 );
nor \U$7727 ( \8104 , \8102 , \8103 );
xnor \U$7728 ( \8105 , \8104 , \5467 );
and \U$7729 ( \8106 , \8100 , \8105 );
and \U$7730 ( \8107 , \8096 , \8105 );
or \U$7731 ( \8108 , \8101 , \8106 , \8107 );
and \U$7732 ( \8109 , \8091 , \8108 );
and \U$7733 ( \8110 , \8073 , \8108 );
or \U$7734 ( \8111 , \8092 , \8109 , \8110 );
and \U$7735 ( \8112 , \8057 , \8111 );
and \U$7736 ( \8113 , \4841 , \888 );
and \U$7737 ( \8114 , \4833 , \886 );
nor \U$7738 ( \8115 , \8113 , \8114 );
xnor \U$7739 ( \8116 , \8115 , \816 );
and \U$7740 ( \8117 , \5315 , \754 );
and \U$7741 ( \8118 , \5310 , \752 );
nor \U$7742 ( \8119 , \8117 , \8118 );
xnor \U$7743 ( \8120 , \8119 , \711 );
and \U$7744 ( \8121 , \8116 , \8120 );
and \U$7745 ( \8122 , \5838 , \641 );
and \U$7746 ( \8123 , \5579 , \639 );
nor \U$7747 ( \8124 , \8122 , \8123 );
xnor \U$7748 ( \8125 , \8124 , \592 );
and \U$7749 ( \8126 , \8120 , \8125 );
and \U$7750 ( \8127 , \8116 , \8125 );
or \U$7751 ( \8128 , \8121 , \8126 , \8127 );
and \U$7752 ( \8129 , \6219 , \540 );
and \U$7753 ( \8130 , \6210 , \538 );
nor \U$7754 ( \8131 , \8129 , \8130 );
xnor \U$7755 ( \8132 , \8131 , \499 );
and \U$7756 ( \8133 , \6764 , \470 );
and \U$7757 ( \8134 , \6562 , \468 );
nor \U$7758 ( \8135 , \8133 , \8134 );
xnor \U$7759 ( \8136 , \8135 , \440 );
and \U$7760 ( \8137 , \8132 , \8136 );
and \U$7761 ( \8138 , \7239 , \422 );
and \U$7762 ( \8139 , \7067 , \420 );
nor \U$7763 ( \8140 , \8138 , \8139 );
xnor \U$7764 ( \8141 , \8140 , \403 );
and \U$7765 ( \8142 , \8136 , \8141 );
and \U$7766 ( \8143 , \8132 , \8141 );
or \U$7767 ( \8144 , \8137 , \8142 , \8143 );
and \U$7768 ( \8145 , \8128 , \8144 );
and \U$7769 ( \8146 , \3951 , \1422 );
and \U$7770 ( \8147 , \3743 , \1420 );
nor \U$7771 ( \8148 , \8146 , \8147 );
xnor \U$7772 ( \8149 , \8148 , \1286 );
and \U$7773 ( \8150 , \4078 , \1222 );
and \U$7774 ( \8151 , \4073 , \1220 );
nor \U$7775 ( \8152 , \8150 , \8151 );
xnor \U$7776 ( \8153 , \8152 , \1144 );
and \U$7777 ( \8154 , \8149 , \8153 );
and \U$7778 ( \8155 , \4531 , \1058 );
and \U$7779 ( \8156 , \4334 , \1056 );
nor \U$7780 ( \8157 , \8155 , \8156 );
xnor \U$7781 ( \8158 , \8157 , \964 );
and \U$7782 ( \8159 , \8153 , \8158 );
and \U$7783 ( \8160 , \8149 , \8158 );
or \U$7784 ( \8161 , \8154 , \8159 , \8160 );
and \U$7785 ( \8162 , \8144 , \8161 );
and \U$7786 ( \8163 , \8128 , \8161 );
or \U$7787 ( \8164 , \8145 , \8162 , \8163 );
and \U$7788 ( \8165 , \8111 , \8164 );
and \U$7789 ( \8166 , \8057 , \8164 );
or \U$7790 ( \8167 , \8112 , \8165 , \8166 );
xor \U$7791 ( \8168 , \7743 , \7747 );
xor \U$7792 ( \8169 , \8168 , \7752 );
xor \U$7793 ( \8170 , \7852 , \7856 );
xor \U$7794 ( \8171 , \8170 , \7861 );
and \U$7795 ( \8172 , \8169 , \8171 );
xor \U$7796 ( \8173 , \7777 , \7781 );
xor \U$7797 ( \8174 , \8173 , \7786 );
and \U$7798 ( \8175 , \8171 , \8174 );
and \U$7799 ( \8176 , \8169 , \8174 );
or \U$7800 ( \8177 , \8172 , \8175 , \8176 );
xor \U$7801 ( \8178 , \7812 , \7816 );
xor \U$7802 ( \8179 , \8178 , \7821 );
xor \U$7803 ( \8180 , \7868 , \7872 );
xor \U$7804 ( \8181 , \8180 , \7877 );
and \U$7805 ( \8182 , \8179 , \8181 );
xor \U$7806 ( \8183 , \7885 , \7889 );
xor \U$7807 ( \8184 , \8183 , \7894 );
and \U$7808 ( \8185 , \8181 , \8184 );
and \U$7809 ( \8186 , \8179 , \8184 );
or \U$7810 ( \8187 , \8182 , \8185 , \8186 );
and \U$7811 ( \8188 , \8177 , \8187 );
buf \U$7812 ( \8189 , RIc223ed8_118);
and \U$7813 ( \8190 , \8189 , \379 );
xor \U$7814 ( \8191 , \7759 , \7763 );
xor \U$7815 ( \8192 , \8191 , \7769 );
or \U$7816 ( \8193 , \8190 , \8192 );
and \U$7817 ( \8194 , \8187 , \8193 );
and \U$7818 ( \8195 , \8177 , \8193 );
or \U$7819 ( \8196 , \8188 , \8194 , \8195 );
and \U$7820 ( \8197 , \8167 , \8196 );
xor \U$7821 ( \8198 , \7581 , \7585 );
xor \U$7822 ( \8199 , \8198 , \7590 );
xor \U$7823 ( \8200 , \7905 , \7907 );
xor \U$7824 ( \8201 , \8200 , \7910 );
and \U$7825 ( \8202 , \8199 , \8201 );
xor \U$7826 ( \8203 , \7925 , \7927 );
xor \U$7827 ( \8204 , \8203 , \7930 );
and \U$7828 ( \8205 , \8201 , \8204 );
and \U$7829 ( \8206 , \8199 , \8204 );
or \U$7830 ( \8207 , \8202 , \8205 , \8206 );
and \U$7831 ( \8208 , \8196 , \8207 );
and \U$7832 ( \8209 , \8167 , \8207 );
or \U$7833 ( \8210 , \8197 , \8208 , \8209 );
xor \U$7834 ( \8211 , \7792 , \7847 );
xor \U$7835 ( \8212 , \8211 , \7900 );
xor \U$7836 ( \8213 , \7913 , \7922 );
xor \U$7837 ( \8214 , \8213 , \7933 );
and \U$7838 ( \8215 , \8212 , \8214 );
xor \U$7839 ( \8216 , \7939 , \7941 );
xor \U$7840 ( \8217 , \8216 , \7944 );
and \U$7841 ( \8218 , \8214 , \8217 );
and \U$7842 ( \8219 , \8212 , \8217 );
or \U$7843 ( \8220 , \8215 , \8218 , \8219 );
and \U$7844 ( \8221 , \8210 , \8220 );
xor \U$7845 ( \8222 , \7755 , \7772 );
xor \U$7846 ( \8223 , \8222 , \7789 );
xor \U$7847 ( \8224 , \7864 , \7880 );
xor \U$7848 ( \8225 , \8224 , \7897 );
and \U$7849 ( \8226 , \8223 , \8225 );
xor \U$7850 ( \8227 , \7914 , \7916 );
xor \U$7851 ( \8228 , \8227 , \7919 );
and \U$7852 ( \8229 , \8225 , \8228 );
and \U$7853 ( \8230 , \8223 , \8228 );
or \U$7854 ( \8231 , \8226 , \8229 , \8230 );
xor \U$7855 ( \8232 , \7575 , \7593 );
xor \U$7856 ( \8233 , \8232 , \7610 );
and \U$7857 ( \8234 , \8231 , \8233 );
xor \U$7858 ( \8235 , \7952 , \7954 );
xor \U$7859 ( \8236 , \8235 , \7956 );
and \U$7860 ( \8237 , \8233 , \8236 );
and \U$7861 ( \8238 , \8231 , \8236 );
or \U$7862 ( \8239 , \8234 , \8237 , \8238 );
and \U$7863 ( \8240 , \8220 , \8239 );
and \U$7864 ( \8241 , \8210 , \8239 );
or \U$7865 ( \8242 , \8221 , \8240 , \8241 );
xor \U$7866 ( \8243 , \7903 , \7936 );
xor \U$7867 ( \8244 , \8243 , \7947 );
xor \U$7868 ( \8245 , \7959 , \7961 );
xor \U$7869 ( \8246 , \8245 , \7964 );
and \U$7870 ( \8247 , \8244 , \8246 );
xor \U$7871 ( \8248 , \7970 , \7972 );
and \U$7872 ( \8249 , \8246 , \8248 );
and \U$7873 ( \8250 , \8244 , \8248 );
or \U$7874 ( \8251 , \8247 , \8249 , \8250 );
and \U$7875 ( \8252 , \8242 , \8251 );
xor \U$7876 ( \8253 , \7978 , \7980 );
xor \U$7877 ( \8254 , \8253 , \7982 );
and \U$7878 ( \8255 , \8251 , \8254 );
and \U$7879 ( \8256 , \8242 , \8254 );
or \U$7880 ( \8257 , \8252 , \8255 , \8256 );
xor \U$7881 ( \8258 , \7683 , \7701 );
xor \U$7882 ( \8259 , \8258 , \7707 );
and \U$7883 ( \8260 , \8257 , \8259 );
xor \U$7884 ( \8261 , \7976 , \7985 );
xor \U$7885 ( \8262 , \8261 , \7988 );
and \U$7886 ( \8263 , \8259 , \8262 );
and \U$7887 ( \8264 , \8257 , \8262 );
or \U$7888 ( \8265 , \8260 , \8263 , \8264 );
xor \U$7889 ( \8266 , \7991 , \7993 );
xor \U$7890 ( \8267 , \8266 , \7996 );
and \U$7891 ( \8268 , \8265 , \8267 );
and \U$7892 ( \8269 , \8005 , \8268 );
xor \U$7893 ( \8270 , \8005 , \8268 );
xor \U$7894 ( \8271 , \8265 , \8267 );
and \U$7895 ( \8272 , \2104 , \2980 );
and \U$7896 ( \8273 , \1861 , \2978 );
nor \U$7897 ( \8274 , \8272 , \8273 );
xnor \U$7898 ( \8275 , \8274 , \2831 );
and \U$7899 ( \8276 , \2295 , \2658 );
and \U$7900 ( \8277 , \2109 , \2656 );
nor \U$7901 ( \8278 , \8276 , \8277 );
xnor \U$7902 ( \8279 , \8278 , \2516 );
and \U$7903 ( \8280 , \8275 , \8279 );
and \U$7904 ( \8281 , \2703 , \2362 );
and \U$7905 ( \8282 , \2439 , \2360 );
nor \U$7906 ( \8283 , \8281 , \8282 );
xnor \U$7907 ( \8284 , \8283 , \2225 );
and \U$7908 ( \8285 , \8279 , \8284 );
and \U$7909 ( \8286 , \8275 , \8284 );
or \U$7910 ( \8287 , \8280 , \8285 , \8286 );
and \U$7911 ( \8288 , \2902 , \2156 );
and \U$7912 ( \8289 , \2728 , \2154 );
nor \U$7913 ( \8290 , \8288 , \8289 );
xnor \U$7914 ( \8291 , \8290 , \2004 );
and \U$7915 ( \8292 , \3207 , \1888 );
and \U$7916 ( \8293 , \3069 , \1886 );
nor \U$7917 ( \8294 , \8292 , \8293 );
xnor \U$7918 ( \8295 , \8294 , \1732 );
and \U$7919 ( \8296 , \8291 , \8295 );
and \U$7920 ( \8297 , \3743 , \1616 );
and \U$7921 ( \8298 , \3326 , \1614 );
nor \U$7922 ( \8299 , \8297 , \8298 );
xnor \U$7923 ( \8300 , \8299 , \1503 );
and \U$7924 ( \8301 , \8295 , \8300 );
and \U$7925 ( \8302 , \8291 , \8300 );
or \U$7926 ( \8303 , \8296 , \8301 , \8302 );
and \U$7927 ( \8304 , \8287 , \8303 );
and \U$7928 ( \8305 , \1441 , \4094 );
and \U$7929 ( \8306 , \1336 , \4092 );
nor \U$7930 ( \8307 , \8305 , \8306 );
xnor \U$7931 ( \8308 , \8307 , \3848 );
and \U$7932 ( \8309 , \1562 , \3699 );
and \U$7933 ( \8310 , \1446 , \3697 );
nor \U$7934 ( \8311 , \8309 , \8310 );
xnor \U$7935 ( \8312 , \8311 , \3512 );
and \U$7936 ( \8313 , \8308 , \8312 );
and \U$7937 ( \8314 , \1853 , \3386 );
and \U$7938 ( \8315 , \1677 , \3384 );
nor \U$7939 ( \8316 , \8314 , \8315 );
xnor \U$7940 ( \8317 , \8316 , \3181 );
and \U$7941 ( \8318 , \8312 , \8317 );
and \U$7942 ( \8319 , \8308 , \8317 );
or \U$7943 ( \8320 , \8313 , \8318 , \8319 );
and \U$7944 ( \8321 , \8303 , \8320 );
and \U$7945 ( \8322 , \8287 , \8320 );
or \U$7946 ( \8323 , \8304 , \8321 , \8322 );
and \U$7947 ( \8324 , \5310 , \888 );
and \U$7948 ( \8325 , \4841 , \886 );
nor \U$7949 ( \8326 , \8324 , \8325 );
xnor \U$7950 ( \8327 , \8326 , \816 );
and \U$7951 ( \8328 , \5579 , \754 );
and \U$7952 ( \8329 , \5315 , \752 );
nor \U$7953 ( \8330 , \8328 , \8329 );
xnor \U$7954 ( \8331 , \8330 , \711 );
and \U$7955 ( \8332 , \8327 , \8331 );
and \U$7956 ( \8333 , \6210 , \641 );
and \U$7957 ( \8334 , \5838 , \639 );
nor \U$7958 ( \8335 , \8333 , \8334 );
xnor \U$7959 ( \8336 , \8335 , \592 );
and \U$7960 ( \8337 , \8331 , \8336 );
and \U$7961 ( \8338 , \8327 , \8336 );
or \U$7962 ( \8339 , \8332 , \8337 , \8338 );
and \U$7963 ( \8340 , \4073 , \1422 );
and \U$7964 ( \8341 , \3951 , \1420 );
nor \U$7965 ( \8342 , \8340 , \8341 );
xnor \U$7966 ( \8343 , \8342 , \1286 );
and \U$7967 ( \8344 , \4334 , \1222 );
and \U$7968 ( \8345 , \4078 , \1220 );
nor \U$7969 ( \8346 , \8344 , \8345 );
xnor \U$7970 ( \8347 , \8346 , \1144 );
and \U$7971 ( \8348 , \8343 , \8347 );
and \U$7972 ( \8349 , \4833 , \1058 );
and \U$7973 ( \8350 , \4531 , \1056 );
nor \U$7974 ( \8351 , \8349 , \8350 );
xnor \U$7975 ( \8352 , \8351 , \964 );
and \U$7976 ( \8353 , \8347 , \8352 );
and \U$7977 ( \8354 , \8343 , \8352 );
or \U$7978 ( \8355 , \8348 , \8353 , \8354 );
and \U$7979 ( \8356 , \8339 , \8355 );
and \U$7980 ( \8357 , \6562 , \540 );
and \U$7981 ( \8358 , \6219 , \538 );
nor \U$7982 ( \8359 , \8357 , \8358 );
xnor \U$7983 ( \8360 , \8359 , \499 );
and \U$7984 ( \8361 , \7067 , \470 );
and \U$7985 ( \8362 , \6764 , \468 );
nor \U$7986 ( \8363 , \8361 , \8362 );
xnor \U$7987 ( \8364 , \8363 , \440 );
and \U$7988 ( \8365 , \8360 , \8364 );
and \U$7989 ( \8366 , \7765 , \422 );
and \U$7990 ( \8367 , \7239 , \420 );
nor \U$7991 ( \8368 , \8366 , \8367 );
xnor \U$7992 ( \8369 , \8368 , \403 );
and \U$7993 ( \8370 , \8364 , \8369 );
and \U$7994 ( \8371 , \8360 , \8369 );
or \U$7995 ( \8372 , \8365 , \8370 , \8371 );
and \U$7996 ( \8373 , \8355 , \8372 );
and \U$7997 ( \8374 , \8339 , \8372 );
or \U$7998 ( \8375 , \8356 , \8373 , \8374 );
and \U$7999 ( \8376 , \8323 , \8375 );
and \U$8000 ( \8377 , \851 , \5242 );
and \U$8001 ( \8378 , \771 , \5240 );
nor \U$8002 ( \8379 , \8377 , \8378 );
xnor \U$8003 ( \8380 , \8379 , \5054 );
and \U$8004 ( \8381 , \987 , \4868 );
and \U$8005 ( \8382 , \925 , \4866 );
nor \U$8006 ( \8383 , \8381 , \8382 );
xnor \U$8007 ( \8384 , \8383 , \4636 );
and \U$8008 ( \8385 , \8380 , \8384 );
and \U$8009 ( \8386 , \1248 , \4417 );
and \U$8010 ( \8387 , \1050 , \4415 );
nor \U$8011 ( \8388 , \8386 , \8387 );
xnor \U$8012 ( \8389 , \8388 , \4274 );
and \U$8013 ( \8390 , \8384 , \8389 );
and \U$8014 ( \8391 , \8380 , \8389 );
or \U$8015 ( \8392 , \8385 , \8390 , \8391 );
xor \U$8016 ( \8393 , \7577 , \8074 );
xor \U$8017 ( \8394 , \8074 , \8075 );
not \U$8018 ( \8395 , \8394 );
and \U$8019 ( \8396 , \8393 , \8395 );
and \U$8020 ( \8397 , \378 , \8396 );
not \U$8021 ( \8398 , \8397 );
xnor \U$8022 ( \8399 , \8398 , \8078 );
and \U$8023 ( \8400 , \410 , \7829 );
and \U$8024 ( \8401 , \392 , \7827 );
nor \U$8025 ( \8402 , \8400 , \8401 );
xnor \U$8026 ( \8403 , \8402 , \7580 );
and \U$8027 ( \8404 , \8399 , \8403 );
and \U$8028 ( \8405 , \479 , \7300 );
and \U$8029 ( \8406 , \431 , \7298 );
nor \U$8030 ( \8407 , \8405 , \8406 );
xnor \U$8031 ( \8408 , \8407 , \7040 );
and \U$8032 ( \8409 , \8403 , \8408 );
and \U$8033 ( \8410 , \8399 , \8408 );
or \U$8034 ( \8411 , \8404 , \8409 , \8410 );
and \U$8035 ( \8412 , \8392 , \8411 );
and \U$8036 ( \8413 , \556 , \6806 );
and \U$8037 ( \8414 , \487 , \6804 );
nor \U$8038 ( \8415 , \8413 , \8414 );
xnor \U$8039 ( \8416 , \8415 , \6491 );
and \U$8040 ( \8417 , \615 , \6297 );
and \U$8041 ( \8418 , \561 , \6295 );
nor \U$8042 ( \8419 , \8417 , \8418 );
xnor \U$8043 ( \8420 , \8419 , \5957 );
and \U$8044 ( \8421 , \8416 , \8420 );
and \U$8045 ( \8422 , \743 , \5708 );
and \U$8046 ( \8423 , \666 , \5706 );
nor \U$8047 ( \8424 , \8422 , \8423 );
xnor \U$8048 ( \8425 , \8424 , \5467 );
and \U$8049 ( \8426 , \8420 , \8425 );
and \U$8050 ( \8427 , \8416 , \8425 );
or \U$8051 ( \8428 , \8421 , \8426 , \8427 );
and \U$8052 ( \8429 , \8411 , \8428 );
and \U$8053 ( \8430 , \8392 , \8428 );
or \U$8054 ( \8431 , \8412 , \8429 , \8430 );
and \U$8055 ( \8432 , \8375 , \8431 );
and \U$8056 ( \8433 , \8323 , \8431 );
or \U$8057 ( \8434 , \8376 , \8432 , \8433 );
buf \U$8058 ( \8435 , RIc223e60_119);
and \U$8059 ( \8436 , \8435 , \385 );
and \U$8060 ( \8437 , \8189 , \383 );
nor \U$8061 ( \8438 , \8436 , \8437 );
xnor \U$8062 ( \8439 , \8438 , \390 );
buf \U$8063 ( \8440 , RIc223de8_120);
and \U$8064 ( \8441 , \8440 , \379 );
or \U$8065 ( \8442 , \8439 , \8441 );
and \U$8066 ( \8443 , \8189 , \385 );
and \U$8067 ( \8444 , \7765 , \383 );
nor \U$8068 ( \8445 , \8443 , \8444 );
xnor \U$8069 ( \8446 , \8445 , \390 );
and \U$8070 ( \8447 , \8442 , \8446 );
and \U$8071 ( \8448 , \8435 , \379 );
and \U$8072 ( \8449 , \8446 , \8448 );
and \U$8073 ( \8450 , \8442 , \8448 );
or \U$8074 ( \8451 , \8447 , \8449 , \8450 );
xor \U$8075 ( \8452 , \8116 , \8120 );
xor \U$8076 ( \8453 , \8452 , \8125 );
xor \U$8077 ( \8454 , \8132 , \8136 );
xor \U$8078 ( \8455 , \8454 , \8141 );
and \U$8079 ( \8456 , \8453 , \8455 );
xor \U$8080 ( \8457 , \8149 , \8153 );
xor \U$8081 ( \8458 , \8457 , \8158 );
and \U$8082 ( \8459 , \8455 , \8458 );
and \U$8083 ( \8460 , \8453 , \8458 );
or \U$8084 ( \8461 , \8456 , \8459 , \8460 );
and \U$8085 ( \8462 , \8451 , \8461 );
xor \U$8086 ( \8463 , \8009 , \8013 );
xor \U$8087 ( \8464 , \8463 , \8018 );
xor \U$8088 ( \8465 , \8025 , \8029 );
xor \U$8089 ( \8466 , \8465 , \8034 );
and \U$8090 ( \8467 , \8464 , \8466 );
xor \U$8091 ( \8468 , \8042 , \8046 );
xor \U$8092 ( \8469 , \8468 , \8051 );
and \U$8093 ( \8470 , \8466 , \8469 );
and \U$8094 ( \8471 , \8464 , \8469 );
or \U$8095 ( \8472 , \8467 , \8470 , \8471 );
and \U$8096 ( \8473 , \8461 , \8472 );
and \U$8097 ( \8474 , \8451 , \8472 );
or \U$8098 ( \8475 , \8462 , \8473 , \8474 );
and \U$8099 ( \8476 , \8434 , \8475 );
xor \U$8100 ( \8477 , \8061 , \8065 );
xor \U$8101 ( \8478 , \8477 , \8070 );
xor \U$8102 ( \8479 , \8079 , \8083 );
xor \U$8103 ( \8480 , \8479 , \8088 );
and \U$8104 ( \8481 , \8478 , \8480 );
xor \U$8105 ( \8482 , \8096 , \8100 );
xor \U$8106 ( \8483 , \8482 , \8105 );
and \U$8107 ( \8484 , \8480 , \8483 );
and \U$8108 ( \8485 , \8478 , \8483 );
or \U$8109 ( \8486 , \8481 , \8484 , \8485 );
xor \U$8110 ( \8487 , \7796 , \7800 );
xor \U$8111 ( \8488 , \8487 , \7805 );
and \U$8112 ( \8489 , \8486 , \8488 );
xor \U$8113 ( \8490 , \7832 , \7836 );
xor \U$8114 ( \8491 , \8490 , \7841 );
and \U$8115 ( \8492 , \8488 , \8491 );
and \U$8116 ( \8493 , \8486 , \8491 );
or \U$8117 ( \8494 , \8489 , \8492 , \8493 );
and \U$8118 ( \8495 , \8475 , \8494 );
and \U$8119 ( \8496 , \8434 , \8494 );
or \U$8120 ( \8497 , \8476 , \8495 , \8496 );
xor \U$8121 ( \8498 , \8021 , \8037 );
xor \U$8122 ( \8499 , \8498 , \8054 );
xor \U$8123 ( \8500 , \8073 , \8091 );
xor \U$8124 ( \8501 , \8500 , \8108 );
and \U$8125 ( \8502 , \8499 , \8501 );
xor \U$8126 ( \8503 , \8128 , \8144 );
xor \U$8127 ( \8504 , \8503 , \8161 );
and \U$8128 ( \8505 , \8501 , \8504 );
and \U$8129 ( \8506 , \8499 , \8504 );
or \U$8130 ( \8507 , \8502 , \8505 , \8506 );
xor \U$8131 ( \8508 , \8169 , \8171 );
xor \U$8132 ( \8509 , \8508 , \8174 );
xor \U$8133 ( \8510 , \8179 , \8181 );
xor \U$8134 ( \8511 , \8510 , \8184 );
and \U$8135 ( \8512 , \8509 , \8511 );
xnor \U$8136 ( \8513 , \8190 , \8192 );
and \U$8137 ( \8514 , \8511 , \8513 );
and \U$8138 ( \8515 , \8509 , \8513 );
or \U$8139 ( \8516 , \8512 , \8514 , \8515 );
and \U$8140 ( \8517 , \8507 , \8516 );
xor \U$8141 ( \8518 , \7808 , \7824 );
xor \U$8142 ( \8519 , \8518 , \7844 );
and \U$8143 ( \8520 , \8516 , \8519 );
and \U$8144 ( \8521 , \8507 , \8519 );
or \U$8145 ( \8522 , \8517 , \8520 , \8521 );
and \U$8146 ( \8523 , \8497 , \8522 );
xor \U$8147 ( \8524 , \8177 , \8187 );
xor \U$8148 ( \8525 , \8524 , \8193 );
xor \U$8149 ( \8526 , \8223 , \8225 );
xor \U$8150 ( \8527 , \8526 , \8228 );
and \U$8151 ( \8528 , \8525 , \8527 );
xor \U$8152 ( \8529 , \8199 , \8201 );
xor \U$8153 ( \8530 , \8529 , \8204 );
and \U$8154 ( \8531 , \8527 , \8530 );
and \U$8155 ( \8532 , \8525 , \8530 );
or \U$8156 ( \8533 , \8528 , \8531 , \8532 );
and \U$8157 ( \8534 , \8522 , \8533 );
and \U$8158 ( \8535 , \8497 , \8533 );
or \U$8159 ( \8536 , \8523 , \8534 , \8535 );
xor \U$8160 ( \8537 , \8167 , \8196 );
xor \U$8161 ( \8538 , \8537 , \8207 );
xor \U$8162 ( \8539 , \8212 , \8214 );
xor \U$8163 ( \8540 , \8539 , \8217 );
and \U$8164 ( \8541 , \8538 , \8540 );
xor \U$8165 ( \8542 , \8231 , \8233 );
xor \U$8166 ( \8543 , \8542 , \8236 );
and \U$8167 ( \8544 , \8540 , \8543 );
and \U$8168 ( \8545 , \8538 , \8543 );
or \U$8169 ( \8546 , \8541 , \8544 , \8545 );
and \U$8170 ( \8547 , \8536 , \8546 );
xor \U$8171 ( \8548 , \8244 , \8246 );
xor \U$8172 ( \8549 , \8548 , \8248 );
and \U$8173 ( \8550 , \8546 , \8549 );
and \U$8174 ( \8551 , \8536 , \8549 );
or \U$8175 ( \8552 , \8547 , \8550 , \8551 );
xor \U$8176 ( \8553 , \7950 , \7967 );
xor \U$8177 ( \8554 , \8553 , \7973 );
and \U$8178 ( \8555 , \8552 , \8554 );
xor \U$8179 ( \8556 , \8242 , \8251 );
xor \U$8180 ( \8557 , \8556 , \8254 );
and \U$8181 ( \8558 , \8554 , \8557 );
and \U$8182 ( \8559 , \8552 , \8557 );
or \U$8183 ( \8560 , \8555 , \8558 , \8559 );
xor \U$8184 ( \8561 , \8257 , \8259 );
xor \U$8185 ( \8562 , \8561 , \8262 );
and \U$8186 ( \8563 , \8560 , \8562 );
and \U$8187 ( \8564 , \8271 , \8563 );
xor \U$8188 ( \8565 , \8271 , \8563 );
xor \U$8189 ( \8566 , \8560 , \8562 );
and \U$8190 ( \8567 , \487 , \7300 );
and \U$8191 ( \8568 , \479 , \7298 );
nor \U$8192 ( \8569 , \8567 , \8568 );
xnor \U$8193 ( \8570 , \8569 , \7040 );
and \U$8194 ( \8571 , \561 , \6806 );
and \U$8195 ( \8572 , \556 , \6804 );
nor \U$8196 ( \8573 , \8571 , \8572 );
xnor \U$8197 ( \8574 , \8573 , \6491 );
and \U$8198 ( \8575 , \8570 , \8574 );
and \U$8199 ( \8576 , \666 , \6297 );
and \U$8200 ( \8577 , \615 , \6295 );
nor \U$8201 ( \8578 , \8576 , \8577 );
xnor \U$8202 ( \8579 , \8578 , \5957 );
and \U$8203 ( \8580 , \8574 , \8579 );
and \U$8204 ( \8581 , \8570 , \8579 );
or \U$8205 ( \8582 , \8575 , \8580 , \8581 );
buf \U$8206 ( \8583 , RIc225af8_58);
buf \U$8207 ( \8584 , RIc225a80_59);
and \U$8208 ( \8585 , \8583 , \8584 );
not \U$8209 ( \8586 , \8585 );
and \U$8210 ( \8587 , \8075 , \8586 );
not \U$8211 ( \8588 , \8587 );
and \U$8212 ( \8589 , \392 , \8396 );
and \U$8213 ( \8590 , \378 , \8394 );
nor \U$8214 ( \8591 , \8589 , \8590 );
xnor \U$8215 ( \8592 , \8591 , \8078 );
and \U$8216 ( \8593 , \8588 , \8592 );
and \U$8217 ( \8594 , \431 , \7829 );
and \U$8218 ( \8595 , \410 , \7827 );
nor \U$8219 ( \8596 , \8594 , \8595 );
xnor \U$8220 ( \8597 , \8596 , \7580 );
and \U$8221 ( \8598 , \8592 , \8597 );
and \U$8222 ( \8599 , \8588 , \8597 );
or \U$8223 ( \8600 , \8593 , \8598 , \8599 );
and \U$8224 ( \8601 , \8582 , \8600 );
and \U$8225 ( \8602 , \771 , \5708 );
and \U$8226 ( \8603 , \743 , \5706 );
nor \U$8227 ( \8604 , \8602 , \8603 );
xnor \U$8228 ( \8605 , \8604 , \5467 );
and \U$8229 ( \8606 , \925 , \5242 );
and \U$8230 ( \8607 , \851 , \5240 );
nor \U$8231 ( \8608 , \8606 , \8607 );
xnor \U$8232 ( \8609 , \8608 , \5054 );
and \U$8233 ( \8610 , \8605 , \8609 );
and \U$8234 ( \8611 , \1050 , \4868 );
and \U$8235 ( \8612 , \987 , \4866 );
nor \U$8236 ( \8613 , \8611 , \8612 );
xnor \U$8237 ( \8614 , \8613 , \4636 );
and \U$8238 ( \8615 , \8609 , \8614 );
and \U$8239 ( \8616 , \8605 , \8614 );
or \U$8240 ( \8617 , \8610 , \8615 , \8616 );
and \U$8241 ( \8618 , \8600 , \8617 );
and \U$8242 ( \8619 , \8582 , \8617 );
or \U$8243 ( \8620 , \8601 , \8618 , \8619 );
and \U$8244 ( \8621 , \2728 , \2362 );
and \U$8245 ( \8622 , \2703 , \2360 );
nor \U$8246 ( \8623 , \8621 , \8622 );
xnor \U$8247 ( \8624 , \8623 , \2225 );
and \U$8248 ( \8625 , \3069 , \2156 );
and \U$8249 ( \8626 , \2902 , \2154 );
nor \U$8250 ( \8627 , \8625 , \8626 );
xnor \U$8251 ( \8628 , \8627 , \2004 );
and \U$8252 ( \8629 , \8624 , \8628 );
and \U$8253 ( \8630 , \3326 , \1888 );
and \U$8254 ( \8631 , \3207 , \1886 );
nor \U$8255 ( \8632 , \8630 , \8631 );
xnor \U$8256 ( \8633 , \8632 , \1732 );
and \U$8257 ( \8634 , \8628 , \8633 );
and \U$8258 ( \8635 , \8624 , \8633 );
or \U$8259 ( \8636 , \8629 , \8634 , \8635 );
and \U$8260 ( \8637 , \1861 , \3386 );
and \U$8261 ( \8638 , \1853 , \3384 );
nor \U$8262 ( \8639 , \8637 , \8638 );
xnor \U$8263 ( \8640 , \8639 , \3181 );
and \U$8264 ( \8641 , \2109 , \2980 );
and \U$8265 ( \8642 , \2104 , \2978 );
nor \U$8266 ( \8643 , \8641 , \8642 );
xnor \U$8267 ( \8644 , \8643 , \2831 );
and \U$8268 ( \8645 , \8640 , \8644 );
and \U$8269 ( \8646 , \2439 , \2658 );
and \U$8270 ( \8647 , \2295 , \2656 );
nor \U$8271 ( \8648 , \8646 , \8647 );
xnor \U$8272 ( \8649 , \8648 , \2516 );
and \U$8273 ( \8650 , \8644 , \8649 );
and \U$8274 ( \8651 , \8640 , \8649 );
or \U$8275 ( \8652 , \8645 , \8650 , \8651 );
and \U$8276 ( \8653 , \8636 , \8652 );
and \U$8277 ( \8654 , \1336 , \4417 );
and \U$8278 ( \8655 , \1248 , \4415 );
nor \U$8279 ( \8656 , \8654 , \8655 );
xnor \U$8280 ( \8657 , \8656 , \4274 );
and \U$8281 ( \8658 , \1446 , \4094 );
and \U$8282 ( \8659 , \1441 , \4092 );
nor \U$8283 ( \8660 , \8658 , \8659 );
xnor \U$8284 ( \8661 , \8660 , \3848 );
and \U$8285 ( \8662 , \8657 , \8661 );
and \U$8286 ( \8663 , \1677 , \3699 );
and \U$8287 ( \8664 , \1562 , \3697 );
nor \U$8288 ( \8665 , \8663 , \8664 );
xnor \U$8289 ( \8666 , \8665 , \3512 );
and \U$8290 ( \8667 , \8661 , \8666 );
and \U$8291 ( \8668 , \8657 , \8666 );
or \U$8292 ( \8669 , \8662 , \8667 , \8668 );
and \U$8293 ( \8670 , \8652 , \8669 );
and \U$8294 ( \8671 , \8636 , \8669 );
or \U$8295 ( \8672 , \8653 , \8670 , \8671 );
and \U$8296 ( \8673 , \8620 , \8672 );
and \U$8297 ( \8674 , \4841 , \1058 );
and \U$8298 ( \8675 , \4833 , \1056 );
nor \U$8299 ( \8676 , \8674 , \8675 );
xnor \U$8300 ( \8677 , \8676 , \964 );
and \U$8301 ( \8678 , \5315 , \888 );
and \U$8302 ( \8679 , \5310 , \886 );
nor \U$8303 ( \8680 , \8678 , \8679 );
xnor \U$8304 ( \8681 , \8680 , \816 );
and \U$8305 ( \8682 , \8677 , \8681 );
and \U$8306 ( \8683 , \5838 , \754 );
and \U$8307 ( \8684 , \5579 , \752 );
nor \U$8308 ( \8685 , \8683 , \8684 );
xnor \U$8309 ( \8686 , \8685 , \711 );
and \U$8310 ( \8687 , \8681 , \8686 );
and \U$8311 ( \8688 , \8677 , \8686 );
or \U$8312 ( \8689 , \8682 , \8687 , \8688 );
and \U$8313 ( \8690 , \3951 , \1616 );
and \U$8314 ( \8691 , \3743 , \1614 );
nor \U$8315 ( \8692 , \8690 , \8691 );
xnor \U$8316 ( \8693 , \8692 , \1503 );
and \U$8317 ( \8694 , \4078 , \1422 );
and \U$8318 ( \8695 , \4073 , \1420 );
nor \U$8319 ( \8696 , \8694 , \8695 );
xnor \U$8320 ( \8697 , \8696 , \1286 );
and \U$8321 ( \8698 , \8693 , \8697 );
and \U$8322 ( \8699 , \4531 , \1222 );
and \U$8323 ( \8700 , \4334 , \1220 );
nor \U$8324 ( \8701 , \8699 , \8700 );
xnor \U$8325 ( \8702 , \8701 , \1144 );
and \U$8326 ( \8703 , \8697 , \8702 );
and \U$8327 ( \8704 , \8693 , \8702 );
or \U$8328 ( \8705 , \8698 , \8703 , \8704 );
and \U$8329 ( \8706 , \8689 , \8705 );
and \U$8330 ( \8707 , \6219 , \641 );
and \U$8331 ( \8708 , \6210 , \639 );
nor \U$8332 ( \8709 , \8707 , \8708 );
xnor \U$8333 ( \8710 , \8709 , \592 );
and \U$8334 ( \8711 , \6764 , \540 );
and \U$8335 ( \8712 , \6562 , \538 );
nor \U$8336 ( \8713 , \8711 , \8712 );
xnor \U$8337 ( \8714 , \8713 , \499 );
and \U$8338 ( \8715 , \8710 , \8714 );
and \U$8339 ( \8716 , \7239 , \470 );
and \U$8340 ( \8717 , \7067 , \468 );
nor \U$8341 ( \8718 , \8716 , \8717 );
xnor \U$8342 ( \8719 , \8718 , \440 );
and \U$8343 ( \8720 , \8714 , \8719 );
and \U$8344 ( \8721 , \8710 , \8719 );
or \U$8345 ( \8722 , \8715 , \8720 , \8721 );
and \U$8346 ( \8723 , \8705 , \8722 );
and \U$8347 ( \8724 , \8689 , \8722 );
or \U$8348 ( \8725 , \8706 , \8723 , \8724 );
and \U$8349 ( \8726 , \8672 , \8725 );
and \U$8350 ( \8727 , \8620 , \8725 );
or \U$8351 ( \8728 , \8673 , \8726 , \8727 );
xor \U$8352 ( \8729 , \8275 , \8279 );
xor \U$8353 ( \8730 , \8729 , \8284 );
xor \U$8354 ( \8731 , \8380 , \8384 );
xor \U$8355 ( \8732 , \8731 , \8389 );
and \U$8356 ( \8733 , \8730 , \8732 );
xor \U$8357 ( \8734 , \8308 , \8312 );
xor \U$8358 ( \8735 , \8734 , \8317 );
and \U$8359 ( \8736 , \8732 , \8735 );
and \U$8360 ( \8737 , \8730 , \8735 );
or \U$8361 ( \8738 , \8733 , \8736 , \8737 );
xor \U$8362 ( \8739 , \8291 , \8295 );
xor \U$8363 ( \8740 , \8739 , \8300 );
xor \U$8364 ( \8741 , \8327 , \8331 );
xor \U$8365 ( \8742 , \8741 , \8336 );
and \U$8366 ( \8743 , \8740 , \8742 );
xor \U$8367 ( \8744 , \8343 , \8347 );
xor \U$8368 ( \8745 , \8744 , \8352 );
and \U$8369 ( \8746 , \8742 , \8745 );
and \U$8370 ( \8747 , \8740 , \8745 );
or \U$8371 ( \8748 , \8743 , \8746 , \8747 );
and \U$8372 ( \8749 , \8738 , \8748 );
and \U$8373 ( \8750 , \8189 , \422 );
and \U$8374 ( \8751 , \7765 , \420 );
nor \U$8375 ( \8752 , \8750 , \8751 );
xnor \U$8376 ( \8753 , \8752 , \403 );
and \U$8377 ( \8754 , \8440 , \385 );
and \U$8378 ( \8755 , \8435 , \383 );
nor \U$8379 ( \8756 , \8754 , \8755 );
xnor \U$8380 ( \8757 , \8756 , \390 );
and \U$8381 ( \8758 , \8753 , \8757 );
buf \U$8382 ( \8759 , RIc223d70_121);
and \U$8383 ( \8760 , \8759 , \379 );
and \U$8384 ( \8761 , \8757 , \8760 );
and \U$8385 ( \8762 , \8753 , \8760 );
or \U$8386 ( \8763 , \8758 , \8761 , \8762 );
xor \U$8387 ( \8764 , \8360 , \8364 );
xor \U$8388 ( \8765 , \8764 , \8369 );
and \U$8389 ( \8766 , \8763 , \8765 );
xnor \U$8390 ( \8767 , \8439 , \8441 );
and \U$8391 ( \8768 , \8765 , \8767 );
and \U$8392 ( \8769 , \8763 , \8767 );
or \U$8393 ( \8770 , \8766 , \8768 , \8769 );
and \U$8394 ( \8771 , \8748 , \8770 );
and \U$8395 ( \8772 , \8738 , \8770 );
or \U$8396 ( \8773 , \8749 , \8771 , \8772 );
and \U$8397 ( \8774 , \8728 , \8773 );
xor \U$8398 ( \8775 , \8453 , \8455 );
xor \U$8399 ( \8776 , \8775 , \8458 );
xor \U$8400 ( \8777 , \8464 , \8466 );
xor \U$8401 ( \8778 , \8777 , \8469 );
and \U$8402 ( \8779 , \8776 , \8778 );
xor \U$8403 ( \8780 , \8478 , \8480 );
xor \U$8404 ( \8781 , \8780 , \8483 );
and \U$8405 ( \8782 , \8778 , \8781 );
and \U$8406 ( \8783 , \8776 , \8781 );
or \U$8407 ( \8784 , \8779 , \8782 , \8783 );
and \U$8408 ( \8785 , \8773 , \8784 );
and \U$8409 ( \8786 , \8728 , \8784 );
or \U$8410 ( \8787 , \8774 , \8785 , \8786 );
xor \U$8411 ( \8788 , \8323 , \8375 );
xor \U$8412 ( \8789 , \8788 , \8431 );
xor \U$8413 ( \8790 , \8451 , \8461 );
xor \U$8414 ( \8791 , \8790 , \8472 );
and \U$8415 ( \8792 , \8789 , \8791 );
xor \U$8416 ( \8793 , \8486 , \8488 );
xor \U$8417 ( \8794 , \8793 , \8491 );
and \U$8418 ( \8795 , \8791 , \8794 );
and \U$8419 ( \8796 , \8789 , \8794 );
or \U$8420 ( \8797 , \8792 , \8795 , \8796 );
and \U$8421 ( \8798 , \8787 , \8797 );
xor \U$8422 ( \8799 , \8287 , \8303 );
xor \U$8423 ( \8800 , \8799 , \8320 );
xor \U$8424 ( \8801 , \8339 , \8355 );
xor \U$8425 ( \8802 , \8801 , \8372 );
and \U$8426 ( \8803 , \8800 , \8802 );
xor \U$8427 ( \8804 , \8442 , \8446 );
xor \U$8428 ( \8805 , \8804 , \8448 );
and \U$8429 ( \8806 , \8802 , \8805 );
and \U$8430 ( \8807 , \8800 , \8805 );
or \U$8431 ( \8808 , \8803 , \8806 , \8807 );
xor \U$8432 ( \8809 , \8499 , \8501 );
xor \U$8433 ( \8810 , \8809 , \8504 );
and \U$8434 ( \8811 , \8808 , \8810 );
xor \U$8435 ( \8812 , \8509 , \8511 );
xor \U$8436 ( \8813 , \8812 , \8513 );
and \U$8437 ( \8814 , \8810 , \8813 );
and \U$8438 ( \8815 , \8808 , \8813 );
or \U$8439 ( \8816 , \8811 , \8814 , \8815 );
and \U$8440 ( \8817 , \8797 , \8816 );
and \U$8441 ( \8818 , \8787 , \8816 );
or \U$8442 ( \8819 , \8798 , \8817 , \8818 );
xor \U$8443 ( \8820 , \8057 , \8111 );
xor \U$8444 ( \8821 , \8820 , \8164 );
xor \U$8445 ( \8822 , \8507 , \8516 );
xor \U$8446 ( \8823 , \8822 , \8519 );
and \U$8447 ( \8824 , \8821 , \8823 );
xor \U$8448 ( \8825 , \8525 , \8527 );
xor \U$8449 ( \8826 , \8825 , \8530 );
and \U$8450 ( \8827 , \8823 , \8826 );
and \U$8451 ( \8828 , \8821 , \8826 );
or \U$8452 ( \8829 , \8824 , \8827 , \8828 );
and \U$8453 ( \8830 , \8819 , \8829 );
xor \U$8454 ( \8831 , \8538 , \8540 );
xor \U$8455 ( \8832 , \8831 , \8543 );
and \U$8456 ( \8833 , \8829 , \8832 );
and \U$8457 ( \8834 , \8819 , \8832 );
or \U$8458 ( \8835 , \8830 , \8833 , \8834 );
xor \U$8459 ( \8836 , \8210 , \8220 );
xor \U$8460 ( \8837 , \8836 , \8239 );
and \U$8461 ( \8838 , \8835 , \8837 );
xor \U$8462 ( \8839 , \8536 , \8546 );
xor \U$8463 ( \8840 , \8839 , \8549 );
and \U$8464 ( \8841 , \8837 , \8840 );
and \U$8465 ( \8842 , \8835 , \8840 );
or \U$8466 ( \8843 , \8838 , \8841 , \8842 );
xor \U$8467 ( \8844 , \8552 , \8554 );
xor \U$8468 ( \8845 , \8844 , \8557 );
and \U$8469 ( \8846 , \8843 , \8845 );
and \U$8470 ( \8847 , \8566 , \8846 );
xor \U$8471 ( \8848 , \8566 , \8846 );
xor \U$8472 ( \8849 , \8843 , \8845 );
and \U$8473 ( \8850 , \2902 , \2362 );
and \U$8474 ( \8851 , \2728 , \2360 );
nor \U$8475 ( \8852 , \8850 , \8851 );
xnor \U$8476 ( \8853 , \8852 , \2225 );
and \U$8477 ( \8854 , \3207 , \2156 );
and \U$8478 ( \8855 , \3069 , \2154 );
nor \U$8479 ( \8856 , \8854 , \8855 );
xnor \U$8480 ( \8857 , \8856 , \2004 );
and \U$8481 ( \8858 , \8853 , \8857 );
and \U$8482 ( \8859 , \3743 , \1888 );
and \U$8483 ( \8860 , \3326 , \1886 );
nor \U$8484 ( \8861 , \8859 , \8860 );
xnor \U$8485 ( \8862 , \8861 , \1732 );
and \U$8486 ( \8863 , \8857 , \8862 );
and \U$8487 ( \8864 , \8853 , \8862 );
or \U$8488 ( \8865 , \8858 , \8863 , \8864 );
and \U$8489 ( \8866 , \1441 , \4417 );
and \U$8490 ( \8867 , \1336 , \4415 );
nor \U$8491 ( \8868 , \8866 , \8867 );
xnor \U$8492 ( \8869 , \8868 , \4274 );
and \U$8493 ( \8870 , \1562 , \4094 );
and \U$8494 ( \8871 , \1446 , \4092 );
nor \U$8495 ( \8872 , \8870 , \8871 );
xnor \U$8496 ( \8873 , \8872 , \3848 );
and \U$8497 ( \8874 , \8869 , \8873 );
and \U$8498 ( \8875 , \1853 , \3699 );
and \U$8499 ( \8876 , \1677 , \3697 );
nor \U$8500 ( \8877 , \8875 , \8876 );
xnor \U$8501 ( \8878 , \8877 , \3512 );
and \U$8502 ( \8879 , \8873 , \8878 );
and \U$8503 ( \8880 , \8869 , \8878 );
or \U$8504 ( \8881 , \8874 , \8879 , \8880 );
and \U$8505 ( \8882 , \8865 , \8881 );
and \U$8506 ( \8883 , \2104 , \3386 );
and \U$8507 ( \8884 , \1861 , \3384 );
nor \U$8508 ( \8885 , \8883 , \8884 );
xnor \U$8509 ( \8886 , \8885 , \3181 );
and \U$8510 ( \8887 , \2295 , \2980 );
and \U$8511 ( \8888 , \2109 , \2978 );
nor \U$8512 ( \8889 , \8887 , \8888 );
xnor \U$8513 ( \8890 , \8889 , \2831 );
and \U$8514 ( \8891 , \8886 , \8890 );
and \U$8515 ( \8892 , \2703 , \2658 );
and \U$8516 ( \8893 , \2439 , \2656 );
nor \U$8517 ( \8894 , \8892 , \8893 );
xnor \U$8518 ( \8895 , \8894 , \2516 );
and \U$8519 ( \8896 , \8890 , \8895 );
and \U$8520 ( \8897 , \8886 , \8895 );
or \U$8521 ( \8898 , \8891 , \8896 , \8897 );
and \U$8522 ( \8899 , \8881 , \8898 );
and \U$8523 ( \8900 , \8865 , \8898 );
or \U$8524 ( \8901 , \8882 , \8899 , \8900 );
and \U$8525 ( \8902 , \6562 , \641 );
and \U$8526 ( \8903 , \6219 , \639 );
nor \U$8527 ( \8904 , \8902 , \8903 );
xnor \U$8528 ( \8905 , \8904 , \592 );
and \U$8529 ( \8906 , \7067 , \540 );
and \U$8530 ( \8907 , \6764 , \538 );
nor \U$8531 ( \8908 , \8906 , \8907 );
xnor \U$8532 ( \8909 , \8908 , \499 );
and \U$8533 ( \8910 , \8905 , \8909 );
and \U$8534 ( \8911 , \7765 , \470 );
and \U$8535 ( \8912 , \7239 , \468 );
nor \U$8536 ( \8913 , \8911 , \8912 );
xnor \U$8537 ( \8914 , \8913 , \440 );
and \U$8538 ( \8915 , \8909 , \8914 );
and \U$8539 ( \8916 , \8905 , \8914 );
or \U$8540 ( \8917 , \8910 , \8915 , \8916 );
and \U$8541 ( \8918 , \5310 , \1058 );
and \U$8542 ( \8919 , \4841 , \1056 );
nor \U$8543 ( \8920 , \8918 , \8919 );
xnor \U$8544 ( \8921 , \8920 , \964 );
and \U$8545 ( \8922 , \5579 , \888 );
and \U$8546 ( \8923 , \5315 , \886 );
nor \U$8547 ( \8924 , \8922 , \8923 );
xnor \U$8548 ( \8925 , \8924 , \816 );
and \U$8549 ( \8926 , \8921 , \8925 );
and \U$8550 ( \8927 , \6210 , \754 );
and \U$8551 ( \8928 , \5838 , \752 );
nor \U$8552 ( \8929 , \8927 , \8928 );
xnor \U$8553 ( \8930 , \8929 , \711 );
and \U$8554 ( \8931 , \8925 , \8930 );
and \U$8555 ( \8932 , \8921 , \8930 );
or \U$8556 ( \8933 , \8926 , \8931 , \8932 );
and \U$8557 ( \8934 , \8917 , \8933 );
and \U$8558 ( \8935 , \4073 , \1616 );
and \U$8559 ( \8936 , \3951 , \1614 );
nor \U$8560 ( \8937 , \8935 , \8936 );
xnor \U$8561 ( \8938 , \8937 , \1503 );
and \U$8562 ( \8939 , \4334 , \1422 );
and \U$8563 ( \8940 , \4078 , \1420 );
nor \U$8564 ( \8941 , \8939 , \8940 );
xnor \U$8565 ( \8942 , \8941 , \1286 );
and \U$8566 ( \8943 , \8938 , \8942 );
and \U$8567 ( \8944 , \4833 , \1222 );
and \U$8568 ( \8945 , \4531 , \1220 );
nor \U$8569 ( \8946 , \8944 , \8945 );
xnor \U$8570 ( \8947 , \8946 , \1144 );
and \U$8571 ( \8948 , \8942 , \8947 );
and \U$8572 ( \8949 , \8938 , \8947 );
or \U$8573 ( \8950 , \8943 , \8948 , \8949 );
and \U$8574 ( \8951 , \8933 , \8950 );
and \U$8575 ( \8952 , \8917 , \8950 );
or \U$8576 ( \8953 , \8934 , \8951 , \8952 );
and \U$8577 ( \8954 , \8901 , \8953 );
xor \U$8578 ( \8955 , \8075 , \8583 );
xor \U$8579 ( \8956 , \8583 , \8584 );
not \U$8580 ( \8957 , \8956 );
and \U$8581 ( \8958 , \8955 , \8957 );
and \U$8582 ( \8959 , \378 , \8958 );
not \U$8583 ( \8960 , \8959 );
xnor \U$8584 ( \8961 , \8960 , \8587 );
and \U$8585 ( \8962 , \410 , \8396 );
and \U$8586 ( \8963 , \392 , \8394 );
nor \U$8587 ( \8964 , \8962 , \8963 );
xnor \U$8588 ( \8965 , \8964 , \8078 );
and \U$8589 ( \8966 , \8961 , \8965 );
and \U$8590 ( \8967 , \479 , \7829 );
and \U$8591 ( \8968 , \431 , \7827 );
nor \U$8592 ( \8969 , \8967 , \8968 );
xnor \U$8593 ( \8970 , \8969 , \7580 );
and \U$8594 ( \8971 , \8965 , \8970 );
and \U$8595 ( \8972 , \8961 , \8970 );
or \U$8596 ( \8973 , \8966 , \8971 , \8972 );
and \U$8597 ( \8974 , \851 , \5708 );
and \U$8598 ( \8975 , \771 , \5706 );
nor \U$8599 ( \8976 , \8974 , \8975 );
xnor \U$8600 ( \8977 , \8976 , \5467 );
and \U$8601 ( \8978 , \987 , \5242 );
and \U$8602 ( \8979 , \925 , \5240 );
nor \U$8603 ( \8980 , \8978 , \8979 );
xnor \U$8604 ( \8981 , \8980 , \5054 );
and \U$8605 ( \8982 , \8977 , \8981 );
and \U$8606 ( \8983 , \1248 , \4868 );
and \U$8607 ( \8984 , \1050 , \4866 );
nor \U$8608 ( \8985 , \8983 , \8984 );
xnor \U$8609 ( \8986 , \8985 , \4636 );
and \U$8610 ( \8987 , \8981 , \8986 );
and \U$8611 ( \8988 , \8977 , \8986 );
or \U$8612 ( \8989 , \8982 , \8987 , \8988 );
and \U$8613 ( \8990 , \8973 , \8989 );
and \U$8614 ( \8991 , \556 , \7300 );
and \U$8615 ( \8992 , \487 , \7298 );
nor \U$8616 ( \8993 , \8991 , \8992 );
xnor \U$8617 ( \8994 , \8993 , \7040 );
and \U$8618 ( \8995 , \615 , \6806 );
and \U$8619 ( \8996 , \561 , \6804 );
nor \U$8620 ( \8997 , \8995 , \8996 );
xnor \U$8621 ( \8998 , \8997 , \6491 );
and \U$8622 ( \8999 , \8994 , \8998 );
and \U$8623 ( \9000 , \743 , \6297 );
and \U$8624 ( \9001 , \666 , \6295 );
nor \U$8625 ( \9002 , \9000 , \9001 );
xnor \U$8626 ( \9003 , \9002 , \5957 );
and \U$8627 ( \9004 , \8998 , \9003 );
and \U$8628 ( \9005 , \8994 , \9003 );
or \U$8629 ( \9006 , \8999 , \9004 , \9005 );
and \U$8630 ( \9007 , \8989 , \9006 );
and \U$8631 ( \9008 , \8973 , \9006 );
or \U$8632 ( \9009 , \8990 , \9007 , \9008 );
and \U$8633 ( \9010 , \8953 , \9009 );
and \U$8634 ( \9011 , \8901 , \9009 );
or \U$8635 ( \9012 , \8954 , \9010 , \9011 );
xor \U$8636 ( \9013 , \8605 , \8609 );
xor \U$8637 ( \9014 , \9013 , \8614 );
xor \U$8638 ( \9015 , \8640 , \8644 );
xor \U$8639 ( \9016 , \9015 , \8649 );
and \U$8640 ( \9017 , \9014 , \9016 );
xor \U$8641 ( \9018 , \8657 , \8661 );
xor \U$8642 ( \9019 , \9018 , \8666 );
and \U$8643 ( \9020 , \9016 , \9019 );
and \U$8644 ( \9021 , \9014 , \9019 );
or \U$8645 ( \9022 , \9017 , \9020 , \9021 );
xor \U$8646 ( \9023 , \8624 , \8628 );
xor \U$8647 ( \9024 , \9023 , \8633 );
xor \U$8648 ( \9025 , \8677 , \8681 );
xor \U$8649 ( \9026 , \9025 , \8686 );
and \U$8650 ( \9027 , \9024 , \9026 );
xor \U$8651 ( \9028 , \8693 , \8697 );
xor \U$8652 ( \9029 , \9028 , \8702 );
and \U$8653 ( \9030 , \9026 , \9029 );
and \U$8654 ( \9031 , \9024 , \9029 );
or \U$8655 ( \9032 , \9027 , \9030 , \9031 );
and \U$8656 ( \9033 , \9022 , \9032 );
and \U$8657 ( \9034 , \8435 , \422 );
and \U$8658 ( \9035 , \8189 , \420 );
nor \U$8659 ( \9036 , \9034 , \9035 );
xnor \U$8660 ( \9037 , \9036 , \403 );
and \U$8661 ( \9038 , \8759 , \385 );
and \U$8662 ( \9039 , \8440 , \383 );
nor \U$8663 ( \9040 , \9038 , \9039 );
xnor \U$8664 ( \9041 , \9040 , \390 );
and \U$8665 ( \9042 , \9037 , \9041 );
buf \U$8666 ( \9043 , RIc223cf8_122);
and \U$8667 ( \9044 , \9043 , \379 );
and \U$8668 ( \9045 , \9041 , \9044 );
and \U$8669 ( \9046 , \9037 , \9044 );
or \U$8670 ( \9047 , \9042 , \9045 , \9046 );
xor \U$8671 ( \9048 , \8753 , \8757 );
xor \U$8672 ( \9049 , \9048 , \8760 );
and \U$8673 ( \9050 , \9047 , \9049 );
xor \U$8674 ( \9051 , \8710 , \8714 );
xor \U$8675 ( \9052 , \9051 , \8719 );
and \U$8676 ( \9053 , \9049 , \9052 );
and \U$8677 ( \9054 , \9047 , \9052 );
or \U$8678 ( \9055 , \9050 , \9053 , \9054 );
and \U$8679 ( \9056 , \9032 , \9055 );
and \U$8680 ( \9057 , \9022 , \9055 );
or \U$8681 ( \9058 , \9033 , \9056 , \9057 );
and \U$8682 ( \9059 , \9012 , \9058 );
xor \U$8683 ( \9060 , \8399 , \8403 );
xor \U$8684 ( \9061 , \9060 , \8408 );
xor \U$8685 ( \9062 , \8416 , \8420 );
xor \U$8686 ( \9063 , \9062 , \8425 );
and \U$8687 ( \9064 , \9061 , \9063 );
xor \U$8688 ( \9065 , \8730 , \8732 );
xor \U$8689 ( \9066 , \9065 , \8735 );
and \U$8690 ( \9067 , \9063 , \9066 );
and \U$8691 ( \9068 , \9061 , \9066 );
or \U$8692 ( \9069 , \9064 , \9067 , \9068 );
and \U$8693 ( \9070 , \9058 , \9069 );
and \U$8694 ( \9071 , \9012 , \9069 );
or \U$8695 ( \9072 , \9059 , \9070 , \9071 );
xor \U$8696 ( \9073 , \8689 , \8705 );
xor \U$8697 ( \9074 , \9073 , \8722 );
xor \U$8698 ( \9075 , \8740 , \8742 );
xor \U$8699 ( \9076 , \9075 , \8745 );
and \U$8700 ( \9077 , \9074 , \9076 );
xor \U$8701 ( \9078 , \8763 , \8765 );
xor \U$8702 ( \9079 , \9078 , \8767 );
and \U$8703 ( \9080 , \9076 , \9079 );
and \U$8704 ( \9081 , \9074 , \9079 );
or \U$8705 ( \9082 , \9077 , \9080 , \9081 );
xor \U$8706 ( \9083 , \8392 , \8411 );
xor \U$8707 ( \9084 , \9083 , \8428 );
and \U$8708 ( \9085 , \9082 , \9084 );
xor \U$8709 ( \9086 , \8800 , \8802 );
xor \U$8710 ( \9087 , \9086 , \8805 );
and \U$8711 ( \9088 , \9084 , \9087 );
and \U$8712 ( \9089 , \9082 , \9087 );
or \U$8713 ( \9090 , \9085 , \9088 , \9089 );
and \U$8714 ( \9091 , \9072 , \9090 );
xor \U$8715 ( \9092 , \8620 , \8672 );
xor \U$8716 ( \9093 , \9092 , \8725 );
xor \U$8717 ( \9094 , \8738 , \8748 );
xor \U$8718 ( \9095 , \9094 , \8770 );
and \U$8719 ( \9096 , \9093 , \9095 );
xor \U$8720 ( \9097 , \8776 , \8778 );
xor \U$8721 ( \9098 , \9097 , \8781 );
and \U$8722 ( \9099 , \9095 , \9098 );
and \U$8723 ( \9100 , \9093 , \9098 );
or \U$8724 ( \9101 , \9096 , \9099 , \9100 );
and \U$8725 ( \9102 , \9090 , \9101 );
and \U$8726 ( \9103 , \9072 , \9101 );
or \U$8727 ( \9104 , \9091 , \9102 , \9103 );
xor \U$8728 ( \9105 , \8728 , \8773 );
xor \U$8729 ( \9106 , \9105 , \8784 );
xor \U$8730 ( \9107 , \8789 , \8791 );
xor \U$8731 ( \9108 , \9107 , \8794 );
and \U$8732 ( \9109 , \9106 , \9108 );
xor \U$8733 ( \9110 , \8808 , \8810 );
xor \U$8734 ( \9111 , \9110 , \8813 );
and \U$8735 ( \9112 , \9108 , \9111 );
and \U$8736 ( \9113 , \9106 , \9111 );
or \U$8737 ( \9114 , \9109 , \9112 , \9113 );
and \U$8738 ( \9115 , \9104 , \9114 );
xor \U$8739 ( \9116 , \8434 , \8475 );
xor \U$8740 ( \9117 , \9116 , \8494 );
and \U$8741 ( \9118 , \9114 , \9117 );
and \U$8742 ( \9119 , \9104 , \9117 );
or \U$8743 ( \9120 , \9115 , \9118 , \9119 );
xor \U$8744 ( \9121 , \8787 , \8797 );
xor \U$8745 ( \9122 , \9121 , \8816 );
xor \U$8746 ( \9123 , \8821 , \8823 );
xor \U$8747 ( \9124 , \9123 , \8826 );
and \U$8748 ( \9125 , \9122 , \9124 );
and \U$8749 ( \9126 , \9120 , \9125 );
xor \U$8750 ( \9127 , \8497 , \8522 );
xor \U$8751 ( \9128 , \9127 , \8533 );
and \U$8752 ( \9129 , \9125 , \9128 );
and \U$8753 ( \9130 , \9120 , \9128 );
or \U$8754 ( \9131 , \9126 , \9129 , \9130 );
xor \U$8755 ( \9132 , \8835 , \8837 );
xor \U$8756 ( \9133 , \9132 , \8840 );
and \U$8757 ( \9134 , \9131 , \9133 );
and \U$8758 ( \9135 , \8849 , \9134 );
xor \U$8759 ( \9136 , \8849 , \9134 );
xor \U$8760 ( \9137 , \9131 , \9133 );
xor \U$8761 ( \9138 , \8905 , \8909 );
xor \U$8762 ( \9139 , \9138 , \8914 );
xor \U$8763 ( \9140 , \8921 , \8925 );
xor \U$8764 ( \9141 , \9140 , \8930 );
and \U$8765 ( \9142 , \9139 , \9141 );
xor \U$8766 ( \9143 , \8938 , \8942 );
xor \U$8767 ( \9144 , \9143 , \8947 );
and \U$8768 ( \9145 , \9141 , \9144 );
and \U$8769 ( \9146 , \9139 , \9144 );
or \U$8770 ( \9147 , \9142 , \9145 , \9146 );
xor \U$8771 ( \9148 , \8853 , \8857 );
xor \U$8772 ( \9149 , \9148 , \8862 );
xor \U$8773 ( \9150 , \8869 , \8873 );
xor \U$8774 ( \9151 , \9150 , \8878 );
and \U$8775 ( \9152 , \9149 , \9151 );
xor \U$8776 ( \9153 , \8886 , \8890 );
xor \U$8777 ( \9154 , \9153 , \8895 );
and \U$8778 ( \9155 , \9151 , \9154 );
and \U$8779 ( \9156 , \9149 , \9154 );
or \U$8780 ( \9157 , \9152 , \9155 , \9156 );
and \U$8781 ( \9158 , \9147 , \9157 );
and \U$8782 ( \9159 , \8189 , \470 );
and \U$8783 ( \9160 , \7765 , \468 );
nor \U$8784 ( \9161 , \9159 , \9160 );
xnor \U$8785 ( \9162 , \9161 , \440 );
and \U$8786 ( \9163 , \8440 , \422 );
and \U$8787 ( \9164 , \8435 , \420 );
nor \U$8788 ( \9165 , \9163 , \9164 );
xnor \U$8789 ( \9166 , \9165 , \403 );
and \U$8790 ( \9167 , \9162 , \9166 );
and \U$8791 ( \9168 , \9043 , \385 );
and \U$8792 ( \9169 , \8759 , \383 );
nor \U$8793 ( \9170 , \9168 , \9169 );
xnor \U$8794 ( \9171 , \9170 , \390 );
and \U$8795 ( \9172 , \9166 , \9171 );
and \U$8796 ( \9173 , \9162 , \9171 );
or \U$8797 ( \9174 , \9167 , \9172 , \9173 );
xor \U$8798 ( \9175 , \9037 , \9041 );
xor \U$8799 ( \9176 , \9175 , \9044 );
or \U$8800 ( \9177 , \9174 , \9176 );
and \U$8801 ( \9178 , \9157 , \9177 );
and \U$8802 ( \9179 , \9147 , \9177 );
or \U$8803 ( \9180 , \9158 , \9178 , \9179 );
buf \U$8804 ( \9181 , RIc225a08_60);
buf \U$8805 ( \9182 , RIc225990_61);
and \U$8806 ( \9183 , \9181 , \9182 );
not \U$8807 ( \9184 , \9183 );
and \U$8808 ( \9185 , \8584 , \9184 );
not \U$8809 ( \9186 , \9185 );
and \U$8810 ( \9187 , \392 , \8958 );
and \U$8811 ( \9188 , \378 , \8956 );
nor \U$8812 ( \9189 , \9187 , \9188 );
xnor \U$8813 ( \9190 , \9189 , \8587 );
and \U$8814 ( \9191 , \9186 , \9190 );
and \U$8815 ( \9192 , \431 , \8396 );
and \U$8816 ( \9193 , \410 , \8394 );
nor \U$8817 ( \9194 , \9192 , \9193 );
xnor \U$8818 ( \9195 , \9194 , \8078 );
and \U$8819 ( \9196 , \9190 , \9195 );
and \U$8820 ( \9197 , \9186 , \9195 );
or \U$8821 ( \9198 , \9191 , \9196 , \9197 );
and \U$8822 ( \9199 , \771 , \6297 );
and \U$8823 ( \9200 , \743 , \6295 );
nor \U$8824 ( \9201 , \9199 , \9200 );
xnor \U$8825 ( \9202 , \9201 , \5957 );
and \U$8826 ( \9203 , \925 , \5708 );
and \U$8827 ( \9204 , \851 , \5706 );
nor \U$8828 ( \9205 , \9203 , \9204 );
xnor \U$8829 ( \9206 , \9205 , \5467 );
and \U$8830 ( \9207 , \9202 , \9206 );
and \U$8831 ( \9208 , \1050 , \5242 );
and \U$8832 ( \9209 , \987 , \5240 );
nor \U$8833 ( \9210 , \9208 , \9209 );
xnor \U$8834 ( \9211 , \9210 , \5054 );
and \U$8835 ( \9212 , \9206 , \9211 );
and \U$8836 ( \9213 , \9202 , \9211 );
or \U$8837 ( \9214 , \9207 , \9212 , \9213 );
and \U$8838 ( \9215 , \9198 , \9214 );
and \U$8839 ( \9216 , \487 , \7829 );
and \U$8840 ( \9217 , \479 , \7827 );
nor \U$8841 ( \9218 , \9216 , \9217 );
xnor \U$8842 ( \9219 , \9218 , \7580 );
and \U$8843 ( \9220 , \561 , \7300 );
and \U$8844 ( \9221 , \556 , \7298 );
nor \U$8845 ( \9222 , \9220 , \9221 );
xnor \U$8846 ( \9223 , \9222 , \7040 );
and \U$8847 ( \9224 , \9219 , \9223 );
and \U$8848 ( \9225 , \666 , \6806 );
and \U$8849 ( \9226 , \615 , \6804 );
nor \U$8850 ( \9227 , \9225 , \9226 );
xnor \U$8851 ( \9228 , \9227 , \6491 );
and \U$8852 ( \9229 , \9223 , \9228 );
and \U$8853 ( \9230 , \9219 , \9228 );
or \U$8854 ( \9231 , \9224 , \9229 , \9230 );
and \U$8855 ( \9232 , \9214 , \9231 );
and \U$8856 ( \9233 , \9198 , \9231 );
or \U$8857 ( \9234 , \9215 , \9232 , \9233 );
and \U$8858 ( \9235 , \1861 , \3699 );
and \U$8859 ( \9236 , \1853 , \3697 );
nor \U$8860 ( \9237 , \9235 , \9236 );
xnor \U$8861 ( \9238 , \9237 , \3512 );
and \U$8862 ( \9239 , \2109 , \3386 );
and \U$8863 ( \9240 , \2104 , \3384 );
nor \U$8864 ( \9241 , \9239 , \9240 );
xnor \U$8865 ( \9242 , \9241 , \3181 );
and \U$8866 ( \9243 , \9238 , \9242 );
and \U$8867 ( \9244 , \2439 , \2980 );
and \U$8868 ( \9245 , \2295 , \2978 );
nor \U$8869 ( \9246 , \9244 , \9245 );
xnor \U$8870 ( \9247 , \9246 , \2831 );
and \U$8871 ( \9248 , \9242 , \9247 );
and \U$8872 ( \9249 , \9238 , \9247 );
or \U$8873 ( \9250 , \9243 , \9248 , \9249 );
and \U$8874 ( \9251 , \2728 , \2658 );
and \U$8875 ( \9252 , \2703 , \2656 );
nor \U$8876 ( \9253 , \9251 , \9252 );
xnor \U$8877 ( \9254 , \9253 , \2516 );
and \U$8878 ( \9255 , \3069 , \2362 );
and \U$8879 ( \9256 , \2902 , \2360 );
nor \U$8880 ( \9257 , \9255 , \9256 );
xnor \U$8881 ( \9258 , \9257 , \2225 );
and \U$8882 ( \9259 , \9254 , \9258 );
and \U$8883 ( \9260 , \3326 , \2156 );
and \U$8884 ( \9261 , \3207 , \2154 );
nor \U$8885 ( \9262 , \9260 , \9261 );
xnor \U$8886 ( \9263 , \9262 , \2004 );
and \U$8887 ( \9264 , \9258 , \9263 );
and \U$8888 ( \9265 , \9254 , \9263 );
or \U$8889 ( \9266 , \9259 , \9264 , \9265 );
and \U$8890 ( \9267 , \9250 , \9266 );
and \U$8891 ( \9268 , \1336 , \4868 );
and \U$8892 ( \9269 , \1248 , \4866 );
nor \U$8893 ( \9270 , \9268 , \9269 );
xnor \U$8894 ( \9271 , \9270 , \4636 );
and \U$8895 ( \9272 , \1446 , \4417 );
and \U$8896 ( \9273 , \1441 , \4415 );
nor \U$8897 ( \9274 , \9272 , \9273 );
xnor \U$8898 ( \9275 , \9274 , \4274 );
and \U$8899 ( \9276 , \9271 , \9275 );
and \U$8900 ( \9277 , \1677 , \4094 );
and \U$8901 ( \9278 , \1562 , \4092 );
nor \U$8902 ( \9279 , \9277 , \9278 );
xnor \U$8903 ( \9280 , \9279 , \3848 );
and \U$8904 ( \9281 , \9275 , \9280 );
and \U$8905 ( \9282 , \9271 , \9280 );
or \U$8906 ( \9283 , \9276 , \9281 , \9282 );
and \U$8907 ( \9284 , \9266 , \9283 );
and \U$8908 ( \9285 , \9250 , \9283 );
or \U$8909 ( \9286 , \9267 , \9284 , \9285 );
and \U$8910 ( \9287 , \9234 , \9286 );
and \U$8911 ( \9288 , \6219 , \754 );
and \U$8912 ( \9289 , \6210 , \752 );
nor \U$8913 ( \9290 , \9288 , \9289 );
xnor \U$8914 ( \9291 , \9290 , \711 );
and \U$8915 ( \9292 , \6764 , \641 );
and \U$8916 ( \9293 , \6562 , \639 );
nor \U$8917 ( \9294 , \9292 , \9293 );
xnor \U$8918 ( \9295 , \9294 , \592 );
and \U$8919 ( \9296 , \9291 , \9295 );
and \U$8920 ( \9297 , \7239 , \540 );
and \U$8921 ( \9298 , \7067 , \538 );
nor \U$8922 ( \9299 , \9297 , \9298 );
xnor \U$8923 ( \9300 , \9299 , \499 );
and \U$8924 ( \9301 , \9295 , \9300 );
and \U$8925 ( \9302 , \9291 , \9300 );
or \U$8926 ( \9303 , \9296 , \9301 , \9302 );
and \U$8927 ( \9304 , \4841 , \1222 );
and \U$8928 ( \9305 , \4833 , \1220 );
nor \U$8929 ( \9306 , \9304 , \9305 );
xnor \U$8930 ( \9307 , \9306 , \1144 );
and \U$8931 ( \9308 , \5315 , \1058 );
and \U$8932 ( \9309 , \5310 , \1056 );
nor \U$8933 ( \9310 , \9308 , \9309 );
xnor \U$8934 ( \9311 , \9310 , \964 );
and \U$8935 ( \9312 , \9307 , \9311 );
and \U$8936 ( \9313 , \5838 , \888 );
and \U$8937 ( \9314 , \5579 , \886 );
nor \U$8938 ( \9315 , \9313 , \9314 );
xnor \U$8939 ( \9316 , \9315 , \816 );
and \U$8940 ( \9317 , \9311 , \9316 );
and \U$8941 ( \9318 , \9307 , \9316 );
or \U$8942 ( \9319 , \9312 , \9317 , \9318 );
and \U$8943 ( \9320 , \9303 , \9319 );
and \U$8944 ( \9321 , \3951 , \1888 );
and \U$8945 ( \9322 , \3743 , \1886 );
nor \U$8946 ( \9323 , \9321 , \9322 );
xnor \U$8947 ( \9324 , \9323 , \1732 );
and \U$8948 ( \9325 , \4078 , \1616 );
and \U$8949 ( \9326 , \4073 , \1614 );
nor \U$8950 ( \9327 , \9325 , \9326 );
xnor \U$8951 ( \9328 , \9327 , \1503 );
and \U$8952 ( \9329 , \9324 , \9328 );
and \U$8953 ( \9330 , \4531 , \1422 );
and \U$8954 ( \9331 , \4334 , \1420 );
nor \U$8955 ( \9332 , \9330 , \9331 );
xnor \U$8956 ( \9333 , \9332 , \1286 );
and \U$8957 ( \9334 , \9328 , \9333 );
and \U$8958 ( \9335 , \9324 , \9333 );
or \U$8959 ( \9336 , \9329 , \9334 , \9335 );
and \U$8960 ( \9337 , \9319 , \9336 );
and \U$8961 ( \9338 , \9303 , \9336 );
or \U$8962 ( \9339 , \9320 , \9337 , \9338 );
and \U$8963 ( \9340 , \9286 , \9339 );
and \U$8964 ( \9341 , \9234 , \9339 );
or \U$8965 ( \9342 , \9287 , \9340 , \9341 );
and \U$8966 ( \9343 , \9180 , \9342 );
xor \U$8967 ( \9344 , \8961 , \8965 );
xor \U$8968 ( \9345 , \9344 , \8970 );
xor \U$8969 ( \9346 , \8977 , \8981 );
xor \U$8970 ( \9347 , \9346 , \8986 );
and \U$8971 ( \9348 , \9345 , \9347 );
xor \U$8972 ( \9349 , \8994 , \8998 );
xor \U$8973 ( \9350 , \9349 , \9003 );
and \U$8974 ( \9351 , \9347 , \9350 );
and \U$8975 ( \9352 , \9345 , \9350 );
or \U$8976 ( \9353 , \9348 , \9351 , \9352 );
xor \U$8977 ( \9354 , \8570 , \8574 );
xor \U$8978 ( \9355 , \9354 , \8579 );
and \U$8979 ( \9356 , \9353 , \9355 );
xor \U$8980 ( \9357 , \8588 , \8592 );
xor \U$8981 ( \9358 , \9357 , \8597 );
and \U$8982 ( \9359 , \9355 , \9358 );
and \U$8983 ( \9360 , \9353 , \9358 );
or \U$8984 ( \9361 , \9356 , \9359 , \9360 );
and \U$8985 ( \9362 , \9342 , \9361 );
and \U$8986 ( \9363 , \9180 , \9361 );
or \U$8987 ( \9364 , \9343 , \9362 , \9363 );
xor \U$8988 ( \9365 , \8865 , \8881 );
xor \U$8989 ( \9366 , \9365 , \8898 );
xor \U$8990 ( \9367 , \8917 , \8933 );
xor \U$8991 ( \9368 , \9367 , \8950 );
and \U$8992 ( \9369 , \9366 , \9368 );
xor \U$8993 ( \9370 , \8973 , \8989 );
xor \U$8994 ( \9371 , \9370 , \9006 );
and \U$8995 ( \9372 , \9368 , \9371 );
and \U$8996 ( \9373 , \9366 , \9371 );
or \U$8997 ( \9374 , \9369 , \9372 , \9373 );
xor \U$8998 ( \9375 , \9014 , \9016 );
xor \U$8999 ( \9376 , \9375 , \9019 );
xor \U$9000 ( \9377 , \9024 , \9026 );
xor \U$9001 ( \9378 , \9377 , \9029 );
and \U$9002 ( \9379 , \9376 , \9378 );
xor \U$9003 ( \9380 , \9047 , \9049 );
xor \U$9004 ( \9381 , \9380 , \9052 );
and \U$9005 ( \9382 , \9378 , \9381 );
and \U$9006 ( \9383 , \9376 , \9381 );
or \U$9007 ( \9384 , \9379 , \9382 , \9383 );
and \U$9008 ( \9385 , \9374 , \9384 );
xor \U$9009 ( \9386 , \8636 , \8652 );
xor \U$9010 ( \9387 , \9386 , \8669 );
and \U$9011 ( \9388 , \9384 , \9387 );
and \U$9012 ( \9389 , \9374 , \9387 );
or \U$9013 ( \9390 , \9385 , \9388 , \9389 );
and \U$9014 ( \9391 , \9364 , \9390 );
xor \U$9015 ( \9392 , \8582 , \8600 );
xor \U$9016 ( \9393 , \9392 , \8617 );
xor \U$9017 ( \9394 , \9061 , \9063 );
xor \U$9018 ( \9395 , \9394 , \9066 );
and \U$9019 ( \9396 , \9393 , \9395 );
xor \U$9020 ( \9397 , \9074 , \9076 );
xor \U$9021 ( \9398 , \9397 , \9079 );
and \U$9022 ( \9399 , \9395 , \9398 );
and \U$9023 ( \9400 , \9393 , \9398 );
or \U$9024 ( \9401 , \9396 , \9399 , \9400 );
and \U$9025 ( \9402 , \9390 , \9401 );
and \U$9026 ( \9403 , \9364 , \9401 );
or \U$9027 ( \9404 , \9391 , \9402 , \9403 );
xor \U$9028 ( \9405 , \9012 , \9058 );
xor \U$9029 ( \9406 , \9405 , \9069 );
xor \U$9030 ( \9407 , \9082 , \9084 );
xor \U$9031 ( \9408 , \9407 , \9087 );
and \U$9032 ( \9409 , \9406 , \9408 );
xor \U$9033 ( \9410 , \9093 , \9095 );
xor \U$9034 ( \9411 , \9410 , \9098 );
and \U$9035 ( \9412 , \9408 , \9411 );
and \U$9036 ( \9413 , \9406 , \9411 );
or \U$9037 ( \9414 , \9409 , \9412 , \9413 );
and \U$9038 ( \9415 , \9404 , \9414 );
xor \U$9039 ( \9416 , \9106 , \9108 );
xor \U$9040 ( \9417 , \9416 , \9111 );
and \U$9041 ( \9418 , \9414 , \9417 );
and \U$9042 ( \9419 , \9404 , \9417 );
or \U$9043 ( \9420 , \9415 , \9418 , \9419 );
xor \U$9044 ( \9421 , \9104 , \9114 );
xor \U$9045 ( \9422 , \9421 , \9117 );
and \U$9046 ( \9423 , \9420 , \9422 );
xor \U$9047 ( \9424 , \9122 , \9124 );
and \U$9048 ( \9425 , \9422 , \9424 );
and \U$9049 ( \9426 , \9420 , \9424 );
or \U$9050 ( \9427 , \9423 , \9425 , \9426 );
xor \U$9051 ( \9428 , \9120 , \9125 );
xor \U$9052 ( \9429 , \9428 , \9128 );
and \U$9053 ( \9430 , \9427 , \9429 );
xor \U$9054 ( \9431 , \8819 , \8829 );
xor \U$9055 ( \9432 , \9431 , \8832 );
and \U$9056 ( \9433 , \9429 , \9432 );
and \U$9057 ( \9434 , \9427 , \9432 );
or \U$9058 ( \9435 , \9430 , \9433 , \9434 );
and \U$9059 ( \9436 , \9137 , \9435 );
xor \U$9060 ( \9437 , \9137 , \9435 );
xor \U$9061 ( \9438 , \9427 , \9429 );
xor \U$9062 ( \9439 , \9438 , \9432 );
and \U$9063 ( \9440 , \5310 , \1222 );
and \U$9064 ( \9441 , \4841 , \1220 );
nor \U$9065 ( \9442 , \9440 , \9441 );
xnor \U$9066 ( \9443 , \9442 , \1144 );
and \U$9067 ( \9444 , \5579 , \1058 );
and \U$9068 ( \9445 , \5315 , \1056 );
nor \U$9069 ( \9446 , \9444 , \9445 );
xnor \U$9070 ( \9447 , \9446 , \964 );
and \U$9071 ( \9448 , \9443 , \9447 );
and \U$9072 ( \9449 , \6210 , \888 );
and \U$9073 ( \9450 , \5838 , \886 );
nor \U$9074 ( \9451 , \9449 , \9450 );
xnor \U$9075 ( \9452 , \9451 , \816 );
and \U$9076 ( \9453 , \9447 , \9452 );
and \U$9077 ( \9454 , \9443 , \9452 );
or \U$9078 ( \9455 , \9448 , \9453 , \9454 );
and \U$9079 ( \9456 , \4073 , \1888 );
and \U$9080 ( \9457 , \3951 , \1886 );
nor \U$9081 ( \9458 , \9456 , \9457 );
xnor \U$9082 ( \9459 , \9458 , \1732 );
and \U$9083 ( \9460 , \4334 , \1616 );
and \U$9084 ( \9461 , \4078 , \1614 );
nor \U$9085 ( \9462 , \9460 , \9461 );
xnor \U$9086 ( \9463 , \9462 , \1503 );
and \U$9087 ( \9464 , \9459 , \9463 );
and \U$9088 ( \9465 , \4833 , \1422 );
and \U$9089 ( \9466 , \4531 , \1420 );
nor \U$9090 ( \9467 , \9465 , \9466 );
xnor \U$9091 ( \9468 , \9467 , \1286 );
and \U$9092 ( \9469 , \9463 , \9468 );
and \U$9093 ( \9470 , \9459 , \9468 );
or \U$9094 ( \9471 , \9464 , \9469 , \9470 );
and \U$9095 ( \9472 , \9455 , \9471 );
and \U$9096 ( \9473 , \6562 , \754 );
and \U$9097 ( \9474 , \6219 , \752 );
nor \U$9098 ( \9475 , \9473 , \9474 );
xnor \U$9099 ( \9476 , \9475 , \711 );
and \U$9100 ( \9477 , \7067 , \641 );
and \U$9101 ( \9478 , \6764 , \639 );
nor \U$9102 ( \9479 , \9477 , \9478 );
xnor \U$9103 ( \9480 , \9479 , \592 );
and \U$9104 ( \9481 , \9476 , \9480 );
and \U$9105 ( \9482 , \7765 , \540 );
and \U$9106 ( \9483 , \7239 , \538 );
nor \U$9107 ( \9484 , \9482 , \9483 );
xnor \U$9108 ( \9485 , \9484 , \499 );
and \U$9109 ( \9486 , \9480 , \9485 );
and \U$9110 ( \9487 , \9476 , \9485 );
or \U$9111 ( \9488 , \9481 , \9486 , \9487 );
and \U$9112 ( \9489 , \9471 , \9488 );
and \U$9113 ( \9490 , \9455 , \9488 );
or \U$9114 ( \9491 , \9472 , \9489 , \9490 );
xor \U$9115 ( \9492 , \8584 , \9181 );
xor \U$9116 ( \9493 , \9181 , \9182 );
not \U$9117 ( \9494 , \9493 );
and \U$9118 ( \9495 , \9492 , \9494 );
and \U$9119 ( \9496 , \378 , \9495 );
not \U$9120 ( \9497 , \9496 );
xnor \U$9121 ( \9498 , \9497 , \9185 );
and \U$9122 ( \9499 , \410 , \8958 );
and \U$9123 ( \9500 , \392 , \8956 );
nor \U$9124 ( \9501 , \9499 , \9500 );
xnor \U$9125 ( \9502 , \9501 , \8587 );
and \U$9126 ( \9503 , \9498 , \9502 );
and \U$9127 ( \9504 , \479 , \8396 );
and \U$9128 ( \9505 , \431 , \8394 );
nor \U$9129 ( \9506 , \9504 , \9505 );
xnor \U$9130 ( \9507 , \9506 , \8078 );
and \U$9131 ( \9508 , \9502 , \9507 );
and \U$9132 ( \9509 , \9498 , \9507 );
or \U$9133 ( \9510 , \9503 , \9508 , \9509 );
and \U$9134 ( \9511 , \851 , \6297 );
and \U$9135 ( \9512 , \771 , \6295 );
nor \U$9136 ( \9513 , \9511 , \9512 );
xnor \U$9137 ( \9514 , \9513 , \5957 );
and \U$9138 ( \9515 , \987 , \5708 );
and \U$9139 ( \9516 , \925 , \5706 );
nor \U$9140 ( \9517 , \9515 , \9516 );
xnor \U$9141 ( \9518 , \9517 , \5467 );
and \U$9142 ( \9519 , \9514 , \9518 );
and \U$9143 ( \9520 , \1248 , \5242 );
and \U$9144 ( \9521 , \1050 , \5240 );
nor \U$9145 ( \9522 , \9520 , \9521 );
xnor \U$9146 ( \9523 , \9522 , \5054 );
and \U$9147 ( \9524 , \9518 , \9523 );
and \U$9148 ( \9525 , \9514 , \9523 );
or \U$9149 ( \9526 , \9519 , \9524 , \9525 );
and \U$9150 ( \9527 , \9510 , \9526 );
and \U$9151 ( \9528 , \556 , \7829 );
and \U$9152 ( \9529 , \487 , \7827 );
nor \U$9153 ( \9530 , \9528 , \9529 );
xnor \U$9154 ( \9531 , \9530 , \7580 );
and \U$9155 ( \9532 , \615 , \7300 );
and \U$9156 ( \9533 , \561 , \7298 );
nor \U$9157 ( \9534 , \9532 , \9533 );
xnor \U$9158 ( \9535 , \9534 , \7040 );
and \U$9159 ( \9536 , \9531 , \9535 );
and \U$9160 ( \9537 , \743 , \6806 );
and \U$9161 ( \9538 , \666 , \6804 );
nor \U$9162 ( \9539 , \9537 , \9538 );
xnor \U$9163 ( \9540 , \9539 , \6491 );
and \U$9164 ( \9541 , \9535 , \9540 );
and \U$9165 ( \9542 , \9531 , \9540 );
or \U$9166 ( \9543 , \9536 , \9541 , \9542 );
and \U$9167 ( \9544 , \9526 , \9543 );
and \U$9168 ( \9545 , \9510 , \9543 );
or \U$9169 ( \9546 , \9527 , \9544 , \9545 );
and \U$9170 ( \9547 , \9491 , \9546 );
and \U$9171 ( \9548 , \1441 , \4868 );
and \U$9172 ( \9549 , \1336 , \4866 );
nor \U$9173 ( \9550 , \9548 , \9549 );
xnor \U$9174 ( \9551 , \9550 , \4636 );
and \U$9175 ( \9552 , \1562 , \4417 );
and \U$9176 ( \9553 , \1446 , \4415 );
nor \U$9177 ( \9554 , \9552 , \9553 );
xnor \U$9178 ( \9555 , \9554 , \4274 );
and \U$9179 ( \9556 , \9551 , \9555 );
and \U$9180 ( \9557 , \1853 , \4094 );
and \U$9181 ( \9558 , \1677 , \4092 );
nor \U$9182 ( \9559 , \9557 , \9558 );
xnor \U$9183 ( \9560 , \9559 , \3848 );
and \U$9184 ( \9561 , \9555 , \9560 );
and \U$9185 ( \9562 , \9551 , \9560 );
or \U$9186 ( \9563 , \9556 , \9561 , \9562 );
and \U$9187 ( \9564 , \2902 , \2658 );
and \U$9188 ( \9565 , \2728 , \2656 );
nor \U$9189 ( \9566 , \9564 , \9565 );
xnor \U$9190 ( \9567 , \9566 , \2516 );
and \U$9191 ( \9568 , \3207 , \2362 );
and \U$9192 ( \9569 , \3069 , \2360 );
nor \U$9193 ( \9570 , \9568 , \9569 );
xnor \U$9194 ( \9571 , \9570 , \2225 );
and \U$9195 ( \9572 , \9567 , \9571 );
and \U$9196 ( \9573 , \3743 , \2156 );
and \U$9197 ( \9574 , \3326 , \2154 );
nor \U$9198 ( \9575 , \9573 , \9574 );
xnor \U$9199 ( \9576 , \9575 , \2004 );
and \U$9200 ( \9577 , \9571 , \9576 );
and \U$9201 ( \9578 , \9567 , \9576 );
or \U$9202 ( \9579 , \9572 , \9577 , \9578 );
and \U$9203 ( \9580 , \9563 , \9579 );
and \U$9204 ( \9581 , \2104 , \3699 );
and \U$9205 ( \9582 , \1861 , \3697 );
nor \U$9206 ( \9583 , \9581 , \9582 );
xnor \U$9207 ( \9584 , \9583 , \3512 );
and \U$9208 ( \9585 , \2295 , \3386 );
and \U$9209 ( \9586 , \2109 , \3384 );
nor \U$9210 ( \9587 , \9585 , \9586 );
xnor \U$9211 ( \9588 , \9587 , \3181 );
and \U$9212 ( \9589 , \9584 , \9588 );
and \U$9213 ( \9590 , \2703 , \2980 );
and \U$9214 ( \9591 , \2439 , \2978 );
nor \U$9215 ( \9592 , \9590 , \9591 );
xnor \U$9216 ( \9593 , \9592 , \2831 );
and \U$9217 ( \9594 , \9588 , \9593 );
and \U$9218 ( \9595 , \9584 , \9593 );
or \U$9219 ( \9596 , \9589 , \9594 , \9595 );
and \U$9220 ( \9597 , \9579 , \9596 );
and \U$9221 ( \9598 , \9563 , \9596 );
or \U$9222 ( \9599 , \9580 , \9597 , \9598 );
and \U$9223 ( \9600 , \9546 , \9599 );
and \U$9224 ( \9601 , \9491 , \9599 );
or \U$9225 ( \9602 , \9547 , \9600 , \9601 );
and \U$9226 ( \9603 , \8435 , \470 );
and \U$9227 ( \9604 , \8189 , \468 );
nor \U$9228 ( \9605 , \9603 , \9604 );
xnor \U$9229 ( \9606 , \9605 , \440 );
and \U$9230 ( \9607 , \8759 , \422 );
and \U$9231 ( \9608 , \8440 , \420 );
nor \U$9232 ( \9609 , \9607 , \9608 );
xnor \U$9233 ( \9610 , \9609 , \403 );
and \U$9234 ( \9611 , \9606 , \9610 );
buf \U$9235 ( \9612 , RIc223c80_123);
and \U$9236 ( \9613 , \9612 , \385 );
and \U$9237 ( \9614 , \9043 , \383 );
nor \U$9238 ( \9615 , \9613 , \9614 );
xnor \U$9239 ( \9616 , \9615 , \390 );
and \U$9240 ( \9617 , \9610 , \9616 );
and \U$9241 ( \9618 , \9606 , \9616 );
or \U$9242 ( \9619 , \9611 , \9617 , \9618 );
buf \U$9243 ( \9620 , RIc223c08_124);
and \U$9244 ( \9621 , \9620 , \379 );
buf \U$9245 ( \9622 , \9621 );
and \U$9246 ( \9623 , \9619 , \9622 );
and \U$9247 ( \9624 , \9612 , \379 );
and \U$9248 ( \9625 , \9622 , \9624 );
and \U$9249 ( \9626 , \9619 , \9624 );
or \U$9250 ( \9627 , \9623 , \9625 , \9626 );
xor \U$9251 ( \9628 , \9162 , \9166 );
xor \U$9252 ( \9629 , \9628 , \9171 );
xor \U$9253 ( \9630 , \9291 , \9295 );
xor \U$9254 ( \9631 , \9630 , \9300 );
and \U$9255 ( \9632 , \9629 , \9631 );
xor \U$9256 ( \9633 , \9307 , \9311 );
xor \U$9257 ( \9634 , \9633 , \9316 );
and \U$9258 ( \9635 , \9631 , \9634 );
and \U$9259 ( \9636 , \9629 , \9634 );
or \U$9260 ( \9637 , \9632 , \9635 , \9636 );
and \U$9261 ( \9638 , \9627 , \9637 );
xor \U$9262 ( \9639 , \9324 , \9328 );
xor \U$9263 ( \9640 , \9639 , \9333 );
xor \U$9264 ( \9641 , \9238 , \9242 );
xor \U$9265 ( \9642 , \9641 , \9247 );
and \U$9266 ( \9643 , \9640 , \9642 );
xor \U$9267 ( \9644 , \9254 , \9258 );
xor \U$9268 ( \9645 , \9644 , \9263 );
and \U$9269 ( \9646 , \9642 , \9645 );
and \U$9270 ( \9647 , \9640 , \9645 );
or \U$9271 ( \9648 , \9643 , \9646 , \9647 );
and \U$9272 ( \9649 , \9637 , \9648 );
and \U$9273 ( \9650 , \9627 , \9648 );
or \U$9274 ( \9651 , \9638 , \9649 , \9650 );
and \U$9275 ( \9652 , \9602 , \9651 );
xor \U$9276 ( \9653 , \9202 , \9206 );
xor \U$9277 ( \9654 , \9653 , \9211 );
xor \U$9278 ( \9655 , \9219 , \9223 );
xor \U$9279 ( \9656 , \9655 , \9228 );
and \U$9280 ( \9657 , \9654 , \9656 );
xor \U$9281 ( \9658 , \9271 , \9275 );
xor \U$9282 ( \9659 , \9658 , \9280 );
and \U$9283 ( \9660 , \9656 , \9659 );
and \U$9284 ( \9661 , \9654 , \9659 );
or \U$9285 ( \9662 , \9657 , \9660 , \9661 );
xor \U$9286 ( \9663 , \9345 , \9347 );
xor \U$9287 ( \9664 , \9663 , \9350 );
and \U$9288 ( \9665 , \9662 , \9664 );
xor \U$9289 ( \9666 , \9149 , \9151 );
xor \U$9290 ( \9667 , \9666 , \9154 );
and \U$9291 ( \9668 , \9664 , \9667 );
and \U$9292 ( \9669 , \9662 , \9667 );
or \U$9293 ( \9670 , \9665 , \9668 , \9669 );
and \U$9294 ( \9671 , \9651 , \9670 );
and \U$9295 ( \9672 , \9602 , \9670 );
or \U$9296 ( \9673 , \9652 , \9671 , \9672 );
xor \U$9297 ( \9674 , \9147 , \9157 );
xor \U$9298 ( \9675 , \9674 , \9177 );
xor \U$9299 ( \9676 , \9234 , \9286 );
xor \U$9300 ( \9677 , \9676 , \9339 );
and \U$9301 ( \9678 , \9675 , \9677 );
xor \U$9302 ( \9679 , \9353 , \9355 );
xor \U$9303 ( \9680 , \9679 , \9358 );
and \U$9304 ( \9681 , \9677 , \9680 );
and \U$9305 ( \9682 , \9675 , \9680 );
or \U$9306 ( \9683 , \9678 , \9681 , \9682 );
and \U$9307 ( \9684 , \9673 , \9683 );
xor \U$9308 ( \9685 , \9303 , \9319 );
xor \U$9309 ( \9686 , \9685 , \9336 );
xor \U$9310 ( \9687 , \9139 , \9141 );
xor \U$9311 ( \9688 , \9687 , \9144 );
and \U$9312 ( \9689 , \9686 , \9688 );
xnor \U$9313 ( \9690 , \9174 , \9176 );
and \U$9314 ( \9691 , \9688 , \9690 );
and \U$9315 ( \9692 , \9686 , \9690 );
or \U$9316 ( \9693 , \9689 , \9691 , \9692 );
xor \U$9317 ( \9694 , \9366 , \9368 );
xor \U$9318 ( \9695 , \9694 , \9371 );
and \U$9319 ( \9696 , \9693 , \9695 );
xor \U$9320 ( \9697 , \9376 , \9378 );
xor \U$9321 ( \9698 , \9697 , \9381 );
and \U$9322 ( \9699 , \9695 , \9698 );
and \U$9323 ( \9700 , \9693 , \9698 );
or \U$9324 ( \9701 , \9696 , \9699 , \9700 );
and \U$9325 ( \9702 , \9683 , \9701 );
and \U$9326 ( \9703 , \9673 , \9701 );
or \U$9327 ( \9704 , \9684 , \9702 , \9703 );
xor \U$9328 ( \9705 , \8901 , \8953 );
xor \U$9329 ( \9706 , \9705 , \9009 );
xor \U$9330 ( \9707 , \9022 , \9032 );
xor \U$9331 ( \9708 , \9707 , \9055 );
and \U$9332 ( \9709 , \9706 , \9708 );
xor \U$9333 ( \9710 , \9393 , \9395 );
xor \U$9334 ( \9711 , \9710 , \9398 );
and \U$9335 ( \9712 , \9708 , \9711 );
and \U$9336 ( \9713 , \9706 , \9711 );
or \U$9337 ( \9714 , \9709 , \9712 , \9713 );
and \U$9338 ( \9715 , \9704 , \9714 );
xor \U$9339 ( \9716 , \9406 , \9408 );
xor \U$9340 ( \9717 , \9716 , \9411 );
and \U$9341 ( \9718 , \9714 , \9717 );
and \U$9342 ( \9719 , \9704 , \9717 );
or \U$9343 ( \9720 , \9715 , \9718 , \9719 );
xor \U$9344 ( \9721 , \9072 , \9090 );
xor \U$9345 ( \9722 , \9721 , \9101 );
and \U$9346 ( \9723 , \9720 , \9722 );
xor \U$9347 ( \9724 , \9404 , \9414 );
xor \U$9348 ( \9725 , \9724 , \9417 );
and \U$9349 ( \9726 , \9722 , \9725 );
and \U$9350 ( \9727 , \9720 , \9725 );
or \U$9351 ( \9728 , \9723 , \9726 , \9727 );
xor \U$9352 ( \9729 , \9420 , \9422 );
xor \U$9353 ( \9730 , \9729 , \9424 );
and \U$9354 ( \9731 , \9728 , \9730 );
and \U$9355 ( \9732 , \9439 , \9731 );
xor \U$9356 ( \9733 , \9439 , \9731 );
xor \U$9357 ( \9734 , \9728 , \9730 );
and \U$9358 ( \9735 , \2728 , \2980 );
and \U$9359 ( \9736 , \2703 , \2978 );
nor \U$9360 ( \9737 , \9735 , \9736 );
xnor \U$9361 ( \9738 , \9737 , \2831 );
and \U$9362 ( \9739 , \3069 , \2658 );
and \U$9363 ( \9740 , \2902 , \2656 );
nor \U$9364 ( \9741 , \9739 , \9740 );
xnor \U$9365 ( \9742 , \9741 , \2516 );
and \U$9366 ( \9743 , \9738 , \9742 );
and \U$9367 ( \9744 , \3326 , \2362 );
and \U$9368 ( \9745 , \3207 , \2360 );
nor \U$9369 ( \9746 , \9744 , \9745 );
xnor \U$9370 ( \9747 , \9746 , \2225 );
and \U$9371 ( \9748 , \9742 , \9747 );
and \U$9372 ( \9749 , \9738 , \9747 );
or \U$9373 ( \9750 , \9743 , \9748 , \9749 );
and \U$9374 ( \9751 , \1861 , \4094 );
and \U$9375 ( \9752 , \1853 , \4092 );
nor \U$9376 ( \9753 , \9751 , \9752 );
xnor \U$9377 ( \9754 , \9753 , \3848 );
and \U$9378 ( \9755 , \2109 , \3699 );
and \U$9379 ( \9756 , \2104 , \3697 );
nor \U$9380 ( \9757 , \9755 , \9756 );
xnor \U$9381 ( \9758 , \9757 , \3512 );
and \U$9382 ( \9759 , \9754 , \9758 );
and \U$9383 ( \9760 , \2439 , \3386 );
and \U$9384 ( \9761 , \2295 , \3384 );
nor \U$9385 ( \9762 , \9760 , \9761 );
xnor \U$9386 ( \9763 , \9762 , \3181 );
and \U$9387 ( \9764 , \9758 , \9763 );
and \U$9388 ( \9765 , \9754 , \9763 );
or \U$9389 ( \9766 , \9759 , \9764 , \9765 );
and \U$9390 ( \9767 , \9750 , \9766 );
and \U$9391 ( \9768 , \1336 , \5242 );
and \U$9392 ( \9769 , \1248 , \5240 );
nor \U$9393 ( \9770 , \9768 , \9769 );
xnor \U$9394 ( \9771 , \9770 , \5054 );
and \U$9395 ( \9772 , \1446 , \4868 );
and \U$9396 ( \9773 , \1441 , \4866 );
nor \U$9397 ( \9774 , \9772 , \9773 );
xnor \U$9398 ( \9775 , \9774 , \4636 );
and \U$9399 ( \9776 , \9771 , \9775 );
and \U$9400 ( \9777 , \1677 , \4417 );
and \U$9401 ( \9778 , \1562 , \4415 );
nor \U$9402 ( \9779 , \9777 , \9778 );
xnor \U$9403 ( \9780 , \9779 , \4274 );
and \U$9404 ( \9781 , \9775 , \9780 );
and \U$9405 ( \9782 , \9771 , \9780 );
or \U$9406 ( \9783 , \9776 , \9781 , \9782 );
and \U$9407 ( \9784 , \9766 , \9783 );
and \U$9408 ( \9785 , \9750 , \9783 );
or \U$9409 ( \9786 , \9767 , \9784 , \9785 );
and \U$9410 ( \9787 , \771 , \6806 );
and \U$9411 ( \9788 , \743 , \6804 );
nor \U$9412 ( \9789 , \9787 , \9788 );
xnor \U$9413 ( \9790 , \9789 , \6491 );
and \U$9414 ( \9791 , \925 , \6297 );
and \U$9415 ( \9792 , \851 , \6295 );
nor \U$9416 ( \9793 , \9791 , \9792 );
xnor \U$9417 ( \9794 , \9793 , \5957 );
and \U$9418 ( \9795 , \9790 , \9794 );
and \U$9419 ( \9796 , \1050 , \5708 );
and \U$9420 ( \9797 , \987 , \5706 );
nor \U$9421 ( \9798 , \9796 , \9797 );
xnor \U$9422 ( \9799 , \9798 , \5467 );
and \U$9423 ( \9800 , \9794 , \9799 );
and \U$9424 ( \9801 , \9790 , \9799 );
or \U$9425 ( \9802 , \9795 , \9800 , \9801 );
and \U$9426 ( \9803 , \487 , \8396 );
and \U$9427 ( \9804 , \479 , \8394 );
nor \U$9428 ( \9805 , \9803 , \9804 );
xnor \U$9429 ( \9806 , \9805 , \8078 );
and \U$9430 ( \9807 , \561 , \7829 );
and \U$9431 ( \9808 , \556 , \7827 );
nor \U$9432 ( \9809 , \9807 , \9808 );
xnor \U$9433 ( \9810 , \9809 , \7580 );
and \U$9434 ( \9811 , \9806 , \9810 );
and \U$9435 ( \9812 , \666 , \7300 );
and \U$9436 ( \9813 , \615 , \7298 );
nor \U$9437 ( \9814 , \9812 , \9813 );
xnor \U$9438 ( \9815 , \9814 , \7040 );
and \U$9439 ( \9816 , \9810 , \9815 );
and \U$9440 ( \9817 , \9806 , \9815 );
or \U$9441 ( \9818 , \9811 , \9816 , \9817 );
and \U$9442 ( \9819 , \9802 , \9818 );
buf \U$9443 ( \9820 , RIc225918_62);
buf \U$9444 ( \9821 , RIc2258a0_63);
and \U$9445 ( \9822 , \9820 , \9821 );
not \U$9446 ( \9823 , \9822 );
and \U$9447 ( \9824 , \9182 , \9823 );
not \U$9448 ( \9825 , \9824 );
and \U$9449 ( \9826 , \392 , \9495 );
and \U$9450 ( \9827 , \378 , \9493 );
nor \U$9451 ( \9828 , \9826 , \9827 );
xnor \U$9452 ( \9829 , \9828 , \9185 );
and \U$9453 ( \9830 , \9825 , \9829 );
and \U$9454 ( \9831 , \431 , \8958 );
and \U$9455 ( \9832 , \410 , \8956 );
nor \U$9456 ( \9833 , \9831 , \9832 );
xnor \U$9457 ( \9834 , \9833 , \8587 );
and \U$9458 ( \9835 , \9829 , \9834 );
and \U$9459 ( \9836 , \9825 , \9834 );
or \U$9460 ( \9837 , \9830 , \9835 , \9836 );
and \U$9461 ( \9838 , \9818 , \9837 );
and \U$9462 ( \9839 , \9802 , \9837 );
or \U$9463 ( \9840 , \9819 , \9838 , \9839 );
and \U$9464 ( \9841 , \9786 , \9840 );
and \U$9465 ( \9842 , \6219 , \888 );
and \U$9466 ( \9843 , \6210 , \886 );
nor \U$9467 ( \9844 , \9842 , \9843 );
xnor \U$9468 ( \9845 , \9844 , \816 );
and \U$9469 ( \9846 , \6764 , \754 );
and \U$9470 ( \9847 , \6562 , \752 );
nor \U$9471 ( \9848 , \9846 , \9847 );
xnor \U$9472 ( \9849 , \9848 , \711 );
and \U$9473 ( \9850 , \9845 , \9849 );
and \U$9474 ( \9851 , \7239 , \641 );
and \U$9475 ( \9852 , \7067 , \639 );
nor \U$9476 ( \9853 , \9851 , \9852 );
xnor \U$9477 ( \9854 , \9853 , \592 );
and \U$9478 ( \9855 , \9849 , \9854 );
and \U$9479 ( \9856 , \9845 , \9854 );
or \U$9480 ( \9857 , \9850 , \9855 , \9856 );
and \U$9481 ( \9858 , \4841 , \1422 );
and \U$9482 ( \9859 , \4833 , \1420 );
nor \U$9483 ( \9860 , \9858 , \9859 );
xnor \U$9484 ( \9861 , \9860 , \1286 );
and \U$9485 ( \9862 , \5315 , \1222 );
and \U$9486 ( \9863 , \5310 , \1220 );
nor \U$9487 ( \9864 , \9862 , \9863 );
xnor \U$9488 ( \9865 , \9864 , \1144 );
and \U$9489 ( \9866 , \9861 , \9865 );
and \U$9490 ( \9867 , \5838 , \1058 );
and \U$9491 ( \9868 , \5579 , \1056 );
nor \U$9492 ( \9869 , \9867 , \9868 );
xnor \U$9493 ( \9870 , \9869 , \964 );
and \U$9494 ( \9871 , \9865 , \9870 );
and \U$9495 ( \9872 , \9861 , \9870 );
or \U$9496 ( \9873 , \9866 , \9871 , \9872 );
and \U$9497 ( \9874 , \9857 , \9873 );
and \U$9498 ( \9875 , \3951 , \2156 );
and \U$9499 ( \9876 , \3743 , \2154 );
nor \U$9500 ( \9877 , \9875 , \9876 );
xnor \U$9501 ( \9878 , \9877 , \2004 );
and \U$9502 ( \9879 , \4078 , \1888 );
and \U$9503 ( \9880 , \4073 , \1886 );
nor \U$9504 ( \9881 , \9879 , \9880 );
xnor \U$9505 ( \9882 , \9881 , \1732 );
and \U$9506 ( \9883 , \9878 , \9882 );
and \U$9507 ( \9884 , \4531 , \1616 );
and \U$9508 ( \9885 , \4334 , \1614 );
nor \U$9509 ( \9886 , \9884 , \9885 );
xnor \U$9510 ( \9887 , \9886 , \1503 );
and \U$9511 ( \9888 , \9882 , \9887 );
and \U$9512 ( \9889 , \9878 , \9887 );
or \U$9513 ( \9890 , \9883 , \9888 , \9889 );
and \U$9514 ( \9891 , \9873 , \9890 );
and \U$9515 ( \9892 , \9857 , \9890 );
or \U$9516 ( \9893 , \9874 , \9891 , \9892 );
and \U$9517 ( \9894 , \9840 , \9893 );
and \U$9518 ( \9895 , \9786 , \9893 );
or \U$9519 ( \9896 , \9841 , \9894 , \9895 );
xor \U$9520 ( \9897 , \9551 , \9555 );
xor \U$9521 ( \9898 , \9897 , \9560 );
xor \U$9522 ( \9899 , \9567 , \9571 );
xor \U$9523 ( \9900 , \9899 , \9576 );
and \U$9524 ( \9901 , \9898 , \9900 );
xor \U$9525 ( \9902 , \9584 , \9588 );
xor \U$9526 ( \9903 , \9902 , \9593 );
and \U$9527 ( \9904 , \9900 , \9903 );
and \U$9528 ( \9905 , \9898 , \9903 );
or \U$9529 ( \9906 , \9901 , \9904 , \9905 );
xor \U$9530 ( \9907 , \9443 , \9447 );
xor \U$9531 ( \9908 , \9907 , \9452 );
xor \U$9532 ( \9909 , \9459 , \9463 );
xor \U$9533 ( \9910 , \9909 , \9468 );
and \U$9534 ( \9911 , \9908 , \9910 );
xor \U$9535 ( \9912 , \9476 , \9480 );
xor \U$9536 ( \9913 , \9912 , \9485 );
and \U$9537 ( \9914 , \9910 , \9913 );
and \U$9538 ( \9915 , \9908 , \9913 );
or \U$9539 ( \9916 , \9911 , \9914 , \9915 );
and \U$9540 ( \9917 , \9906 , \9916 );
and \U$9541 ( \9918 , \8189 , \540 );
and \U$9542 ( \9919 , \7765 , \538 );
nor \U$9543 ( \9920 , \9918 , \9919 );
xnor \U$9544 ( \9921 , \9920 , \499 );
and \U$9545 ( \9922 , \8440 , \470 );
and \U$9546 ( \9923 , \8435 , \468 );
nor \U$9547 ( \9924 , \9922 , \9923 );
xnor \U$9548 ( \9925 , \9924 , \440 );
and \U$9549 ( \9926 , \9921 , \9925 );
and \U$9550 ( \9927 , \9043 , \422 );
and \U$9551 ( \9928 , \8759 , \420 );
nor \U$9552 ( \9929 , \9927 , \9928 );
xnor \U$9553 ( \9930 , \9929 , \403 );
and \U$9554 ( \9931 , \9925 , \9930 );
and \U$9555 ( \9932 , \9921 , \9930 );
or \U$9556 ( \9933 , \9926 , \9931 , \9932 );
xor \U$9557 ( \9934 , \9606 , \9610 );
xor \U$9558 ( \9935 , \9934 , \9616 );
and \U$9559 ( \9936 , \9933 , \9935 );
not \U$9560 ( \9937 , \9621 );
and \U$9561 ( \9938 , \9935 , \9937 );
and \U$9562 ( \9939 , \9933 , \9937 );
or \U$9563 ( \9940 , \9936 , \9938 , \9939 );
and \U$9564 ( \9941 , \9916 , \9940 );
and \U$9565 ( \9942 , \9906 , \9940 );
or \U$9566 ( \9943 , \9917 , \9941 , \9942 );
and \U$9567 ( \9944 , \9896 , \9943 );
xor \U$9568 ( \9945 , \9498 , \9502 );
xor \U$9569 ( \9946 , \9945 , \9507 );
xor \U$9570 ( \9947 , \9514 , \9518 );
xor \U$9571 ( \9948 , \9947 , \9523 );
and \U$9572 ( \9949 , \9946 , \9948 );
xor \U$9573 ( \9950 , \9531 , \9535 );
xor \U$9574 ( \9951 , \9950 , \9540 );
and \U$9575 ( \9952 , \9948 , \9951 );
and \U$9576 ( \9953 , \9946 , \9951 );
or \U$9577 ( \9954 , \9949 , \9952 , \9953 );
xor \U$9578 ( \9955 , \9186 , \9190 );
xor \U$9579 ( \9956 , \9955 , \9195 );
and \U$9580 ( \9957 , \9954 , \9956 );
xor \U$9581 ( \9958 , \9654 , \9656 );
xor \U$9582 ( \9959 , \9958 , \9659 );
and \U$9583 ( \9960 , \9956 , \9959 );
and \U$9584 ( \9961 , \9954 , \9959 );
or \U$9585 ( \9962 , \9957 , \9960 , \9961 );
and \U$9586 ( \9963 , \9943 , \9962 );
and \U$9587 ( \9964 , \9896 , \9962 );
or \U$9588 ( \9965 , \9944 , \9963 , \9964 );
xor \U$9589 ( \9966 , \9455 , \9471 );
xor \U$9590 ( \9967 , \9966 , \9488 );
xor \U$9591 ( \9968 , \9510 , \9526 );
xor \U$9592 ( \9969 , \9968 , \9543 );
and \U$9593 ( \9970 , \9967 , \9969 );
xor \U$9594 ( \9971 , \9563 , \9579 );
xor \U$9595 ( \9972 , \9971 , \9596 );
and \U$9596 ( \9973 , \9969 , \9972 );
and \U$9597 ( \9974 , \9967 , \9972 );
or \U$9598 ( \9975 , \9970 , \9973 , \9974 );
xor \U$9599 ( \9976 , \9619 , \9622 );
xor \U$9600 ( \9977 , \9976 , \9624 );
xor \U$9601 ( \9978 , \9629 , \9631 );
xor \U$9602 ( \9979 , \9978 , \9634 );
and \U$9603 ( \9980 , \9977 , \9979 );
xor \U$9604 ( \9981 , \9640 , \9642 );
xor \U$9605 ( \9982 , \9981 , \9645 );
and \U$9606 ( \9983 , \9979 , \9982 );
and \U$9607 ( \9984 , \9977 , \9982 );
or \U$9608 ( \9985 , \9980 , \9983 , \9984 );
and \U$9609 ( \9986 , \9975 , \9985 );
xor \U$9610 ( \9987 , \9250 , \9266 );
xor \U$9611 ( \9988 , \9987 , \9283 );
and \U$9612 ( \9989 , \9985 , \9988 );
and \U$9613 ( \9990 , \9975 , \9988 );
or \U$9614 ( \9991 , \9986 , \9989 , \9990 );
and \U$9615 ( \9992 , \9965 , \9991 );
xor \U$9616 ( \9993 , \9198 , \9214 );
xor \U$9617 ( \9994 , \9993 , \9231 );
xor \U$9618 ( \9995 , \9662 , \9664 );
xor \U$9619 ( \9996 , \9995 , \9667 );
and \U$9620 ( \9997 , \9994 , \9996 );
xor \U$9621 ( \9998 , \9686 , \9688 );
xor \U$9622 ( \9999 , \9998 , \9690 );
and \U$9623 ( \10000 , \9996 , \9999 );
and \U$9624 ( \10001 , \9994 , \9999 );
or \U$9625 ( \10002 , \9997 , \10000 , \10001 );
and \U$9626 ( \10003 , \9991 , \10002 );
and \U$9627 ( \10004 , \9965 , \10002 );
or \U$9628 ( \10005 , \9992 , \10003 , \10004 );
xor \U$9629 ( \10006 , \9602 , \9651 );
xor \U$9630 ( \10007 , \10006 , \9670 );
xor \U$9631 ( \10008 , \9675 , \9677 );
xor \U$9632 ( \10009 , \10008 , \9680 );
and \U$9633 ( \10010 , \10007 , \10009 );
xor \U$9634 ( \10011 , \9693 , \9695 );
xor \U$9635 ( \10012 , \10011 , \9698 );
and \U$9636 ( \10013 , \10009 , \10012 );
and \U$9637 ( \10014 , \10007 , \10012 );
or \U$9638 ( \10015 , \10010 , \10013 , \10014 );
and \U$9639 ( \10016 , \10005 , \10015 );
xor \U$9640 ( \10017 , \9374 , \9384 );
xor \U$9641 ( \10018 , \10017 , \9387 );
and \U$9642 ( \10019 , \10015 , \10018 );
and \U$9643 ( \10020 , \10005 , \10018 );
or \U$9644 ( \10021 , \10016 , \10019 , \10020 );
xor \U$9645 ( \10022 , \9180 , \9342 );
xor \U$9646 ( \10023 , \10022 , \9361 );
xor \U$9647 ( \10024 , \9673 , \9683 );
xor \U$9648 ( \10025 , \10024 , \9701 );
and \U$9649 ( \10026 , \10023 , \10025 );
xor \U$9650 ( \10027 , \9706 , \9708 );
xor \U$9651 ( \10028 , \10027 , \9711 );
and \U$9652 ( \10029 , \10025 , \10028 );
and \U$9653 ( \10030 , \10023 , \10028 );
or \U$9654 ( \10031 , \10026 , \10029 , \10030 );
and \U$9655 ( \10032 , \10021 , \10031 );
xor \U$9656 ( \10033 , \9364 , \9390 );
xor \U$9657 ( \10034 , \10033 , \9401 );
and \U$9658 ( \10035 , \10031 , \10034 );
and \U$9659 ( \10036 , \10021 , \10034 );
or \U$9660 ( \10037 , \10032 , \10035 , \10036 );
xor \U$9661 ( \10038 , \9720 , \9722 );
xor \U$9662 ( \10039 , \10038 , \9725 );
and \U$9663 ( \10040 , \10037 , \10039 );
and \U$9664 ( \10041 , \9734 , \10040 );
xor \U$9665 ( \10042 , \9734 , \10040 );
xor \U$9666 ( \10043 , \10037 , \10039 );
and \U$9667 ( \10044 , \851 , \6806 );
and \U$9668 ( \10045 , \771 , \6804 );
nor \U$9669 ( \10046 , \10044 , \10045 );
xnor \U$9670 ( \10047 , \10046 , \6491 );
and \U$9671 ( \10048 , \987 , \6297 );
and \U$9672 ( \10049 , \925 , \6295 );
nor \U$9673 ( \10050 , \10048 , \10049 );
xnor \U$9674 ( \10051 , \10050 , \5957 );
and \U$9675 ( \10052 , \10047 , \10051 );
and \U$9676 ( \10053 , \1248 , \5708 );
and \U$9677 ( \10054 , \1050 , \5706 );
nor \U$9678 ( \10055 , \10053 , \10054 );
xnor \U$9679 ( \10056 , \10055 , \5467 );
and \U$9680 ( \10057 , \10051 , \10056 );
and \U$9681 ( \10058 , \10047 , \10056 );
or \U$9682 ( \10059 , \10052 , \10057 , \10058 );
xor \U$9683 ( \10060 , \9182 , \9820 );
xor \U$9684 ( \10061 , \9820 , \9821 );
not \U$9685 ( \10062 , \10061 );
and \U$9686 ( \10063 , \10060 , \10062 );
and \U$9687 ( \10064 , \378 , \10063 );
not \U$9688 ( \10065 , \10064 );
xnor \U$9689 ( \10066 , \10065 , \9824 );
and \U$9690 ( \10067 , \410 , \9495 );
and \U$9691 ( \10068 , \392 , \9493 );
nor \U$9692 ( \10069 , \10067 , \10068 );
xnor \U$9693 ( \10070 , \10069 , \9185 );
and \U$9694 ( \10071 , \10066 , \10070 );
and \U$9695 ( \10072 , \479 , \8958 );
and \U$9696 ( \10073 , \431 , \8956 );
nor \U$9697 ( \10074 , \10072 , \10073 );
xnor \U$9698 ( \10075 , \10074 , \8587 );
and \U$9699 ( \10076 , \10070 , \10075 );
and \U$9700 ( \10077 , \10066 , \10075 );
or \U$9701 ( \10078 , \10071 , \10076 , \10077 );
and \U$9702 ( \10079 , \10059 , \10078 );
and \U$9703 ( \10080 , \556 , \8396 );
and \U$9704 ( \10081 , \487 , \8394 );
nor \U$9705 ( \10082 , \10080 , \10081 );
xnor \U$9706 ( \10083 , \10082 , \8078 );
and \U$9707 ( \10084 , \615 , \7829 );
and \U$9708 ( \10085 , \561 , \7827 );
nor \U$9709 ( \10086 , \10084 , \10085 );
xnor \U$9710 ( \10087 , \10086 , \7580 );
and \U$9711 ( \10088 , \10083 , \10087 );
and \U$9712 ( \10089 , \743 , \7300 );
and \U$9713 ( \10090 , \666 , \7298 );
nor \U$9714 ( \10091 , \10089 , \10090 );
xnor \U$9715 ( \10092 , \10091 , \7040 );
and \U$9716 ( \10093 , \10087 , \10092 );
and \U$9717 ( \10094 , \10083 , \10092 );
or \U$9718 ( \10095 , \10088 , \10093 , \10094 );
and \U$9719 ( \10096 , \10078 , \10095 );
and \U$9720 ( \10097 , \10059 , \10095 );
or \U$9721 ( \10098 , \10079 , \10096 , \10097 );
and \U$9722 ( \10099 , \6562 , \888 );
and \U$9723 ( \10100 , \6219 , \886 );
nor \U$9724 ( \10101 , \10099 , \10100 );
xnor \U$9725 ( \10102 , \10101 , \816 );
and \U$9726 ( \10103 , \7067 , \754 );
and \U$9727 ( \10104 , \6764 , \752 );
nor \U$9728 ( \10105 , \10103 , \10104 );
xnor \U$9729 ( \10106 , \10105 , \711 );
and \U$9730 ( \10107 , \10102 , \10106 );
and \U$9731 ( \10108 , \7765 , \641 );
and \U$9732 ( \10109 , \7239 , \639 );
nor \U$9733 ( \10110 , \10108 , \10109 );
xnor \U$9734 ( \10111 , \10110 , \592 );
and \U$9735 ( \10112 , \10106 , \10111 );
and \U$9736 ( \10113 , \10102 , \10111 );
or \U$9737 ( \10114 , \10107 , \10112 , \10113 );
and \U$9738 ( \10115 , \4073 , \2156 );
and \U$9739 ( \10116 , \3951 , \2154 );
nor \U$9740 ( \10117 , \10115 , \10116 );
xnor \U$9741 ( \10118 , \10117 , \2004 );
and \U$9742 ( \10119 , \4334 , \1888 );
and \U$9743 ( \10120 , \4078 , \1886 );
nor \U$9744 ( \10121 , \10119 , \10120 );
xnor \U$9745 ( \10122 , \10121 , \1732 );
and \U$9746 ( \10123 , \10118 , \10122 );
and \U$9747 ( \10124 , \4833 , \1616 );
and \U$9748 ( \10125 , \4531 , \1614 );
nor \U$9749 ( \10126 , \10124 , \10125 );
xnor \U$9750 ( \10127 , \10126 , \1503 );
and \U$9751 ( \10128 , \10122 , \10127 );
and \U$9752 ( \10129 , \10118 , \10127 );
or \U$9753 ( \10130 , \10123 , \10128 , \10129 );
and \U$9754 ( \10131 , \10114 , \10130 );
and \U$9755 ( \10132 , \5310 , \1422 );
and \U$9756 ( \10133 , \4841 , \1420 );
nor \U$9757 ( \10134 , \10132 , \10133 );
xnor \U$9758 ( \10135 , \10134 , \1286 );
and \U$9759 ( \10136 , \5579 , \1222 );
and \U$9760 ( \10137 , \5315 , \1220 );
nor \U$9761 ( \10138 , \10136 , \10137 );
xnor \U$9762 ( \10139 , \10138 , \1144 );
and \U$9763 ( \10140 , \10135 , \10139 );
and \U$9764 ( \10141 , \6210 , \1058 );
and \U$9765 ( \10142 , \5838 , \1056 );
nor \U$9766 ( \10143 , \10141 , \10142 );
xnor \U$9767 ( \10144 , \10143 , \964 );
and \U$9768 ( \10145 , \10139 , \10144 );
and \U$9769 ( \10146 , \10135 , \10144 );
or \U$9770 ( \10147 , \10140 , \10145 , \10146 );
and \U$9771 ( \10148 , \10130 , \10147 );
and \U$9772 ( \10149 , \10114 , \10147 );
or \U$9773 ( \10150 , \10131 , \10148 , \10149 );
and \U$9774 ( \10151 , \10098 , \10150 );
and \U$9775 ( \10152 , \1441 , \5242 );
and \U$9776 ( \10153 , \1336 , \5240 );
nor \U$9777 ( \10154 , \10152 , \10153 );
xnor \U$9778 ( \10155 , \10154 , \5054 );
and \U$9779 ( \10156 , \1562 , \4868 );
and \U$9780 ( \10157 , \1446 , \4866 );
nor \U$9781 ( \10158 , \10156 , \10157 );
xnor \U$9782 ( \10159 , \10158 , \4636 );
and \U$9783 ( \10160 , \10155 , \10159 );
and \U$9784 ( \10161 , \1853 , \4417 );
and \U$9785 ( \10162 , \1677 , \4415 );
nor \U$9786 ( \10163 , \10161 , \10162 );
xnor \U$9787 ( \10164 , \10163 , \4274 );
and \U$9788 ( \10165 , \10159 , \10164 );
and \U$9789 ( \10166 , \10155 , \10164 );
or \U$9790 ( \10167 , \10160 , \10165 , \10166 );
and \U$9791 ( \10168 , \2902 , \2980 );
and \U$9792 ( \10169 , \2728 , \2978 );
nor \U$9793 ( \10170 , \10168 , \10169 );
xnor \U$9794 ( \10171 , \10170 , \2831 );
and \U$9795 ( \10172 , \3207 , \2658 );
and \U$9796 ( \10173 , \3069 , \2656 );
nor \U$9797 ( \10174 , \10172 , \10173 );
xnor \U$9798 ( \10175 , \10174 , \2516 );
and \U$9799 ( \10176 , \10171 , \10175 );
and \U$9800 ( \10177 , \3743 , \2362 );
and \U$9801 ( \10178 , \3326 , \2360 );
nor \U$9802 ( \10179 , \10177 , \10178 );
xnor \U$9803 ( \10180 , \10179 , \2225 );
and \U$9804 ( \10181 , \10175 , \10180 );
and \U$9805 ( \10182 , \10171 , \10180 );
or \U$9806 ( \10183 , \10176 , \10181 , \10182 );
and \U$9807 ( \10184 , \10167 , \10183 );
and \U$9808 ( \10185 , \2104 , \4094 );
and \U$9809 ( \10186 , \1861 , \4092 );
nor \U$9810 ( \10187 , \10185 , \10186 );
xnor \U$9811 ( \10188 , \10187 , \3848 );
and \U$9812 ( \10189 , \2295 , \3699 );
and \U$9813 ( \10190 , \2109 , \3697 );
nor \U$9814 ( \10191 , \10189 , \10190 );
xnor \U$9815 ( \10192 , \10191 , \3512 );
and \U$9816 ( \10193 , \10188 , \10192 );
and \U$9817 ( \10194 , \2703 , \3386 );
and \U$9818 ( \10195 , \2439 , \3384 );
nor \U$9819 ( \10196 , \10194 , \10195 );
xnor \U$9820 ( \10197 , \10196 , \3181 );
and \U$9821 ( \10198 , \10192 , \10197 );
and \U$9822 ( \10199 , \10188 , \10197 );
or \U$9823 ( \10200 , \10193 , \10198 , \10199 );
and \U$9824 ( \10201 , \10183 , \10200 );
and \U$9825 ( \10202 , \10167 , \10200 );
or \U$9826 ( \10203 , \10184 , \10201 , \10202 );
and \U$9827 ( \10204 , \10150 , \10203 );
and \U$9828 ( \10205 , \10098 , \10203 );
or \U$9829 ( \10206 , \10151 , \10204 , \10205 );
and \U$9830 ( \10207 , \8435 , \540 );
and \U$9831 ( \10208 , \8189 , \538 );
nor \U$9832 ( \10209 , \10207 , \10208 );
xnor \U$9833 ( \10210 , \10209 , \499 );
and \U$9834 ( \10211 , \8759 , \470 );
and \U$9835 ( \10212 , \8440 , \468 );
nor \U$9836 ( \10213 , \10211 , \10212 );
xnor \U$9837 ( \10214 , \10213 , \440 );
and \U$9838 ( \10215 , \10210 , \10214 );
and \U$9839 ( \10216 , \9612 , \422 );
and \U$9840 ( \10217 , \9043 , \420 );
nor \U$9841 ( \10218 , \10216 , \10217 );
xnor \U$9842 ( \10219 , \10218 , \403 );
and \U$9843 ( \10220 , \10214 , \10219 );
and \U$9844 ( \10221 , \10210 , \10219 );
or \U$9845 ( \10222 , \10215 , \10220 , \10221 );
buf \U$9846 ( \10223 , RIc223b90_125);
and \U$9847 ( \10224 , \10223 , \385 );
and \U$9848 ( \10225 , \9620 , \383 );
nor \U$9849 ( \10226 , \10224 , \10225 );
xnor \U$9850 ( \10227 , \10226 , \390 );
buf \U$9851 ( \10228 , RIc223b18_126);
and \U$9852 ( \10229 , \10228 , \379 );
or \U$9853 ( \10230 , \10227 , \10229 );
and \U$9854 ( \10231 , \10222 , \10230 );
and \U$9855 ( \10232 , \9620 , \385 );
and \U$9856 ( \10233 , \9612 , \383 );
nor \U$9857 ( \10234 , \10232 , \10233 );
xnor \U$9858 ( \10235 , \10234 , \390 );
and \U$9859 ( \10236 , \10230 , \10235 );
and \U$9860 ( \10237 , \10222 , \10235 );
or \U$9861 ( \10238 , \10231 , \10236 , \10237 );
and \U$9862 ( \10239 , \10223 , \379 );
xor \U$9863 ( \10240 , \9845 , \9849 );
xor \U$9864 ( \10241 , \10240 , \9854 );
and \U$9865 ( \10242 , \10239 , \10241 );
xor \U$9866 ( \10243 , \9921 , \9925 );
xor \U$9867 ( \10244 , \10243 , \9930 );
and \U$9868 ( \10245 , \10241 , \10244 );
and \U$9869 ( \10246 , \10239 , \10244 );
or \U$9870 ( \10247 , \10242 , \10245 , \10246 );
and \U$9871 ( \10248 , \10238 , \10247 );
xor \U$9872 ( \10249 , \9738 , \9742 );
xor \U$9873 ( \10250 , \10249 , \9747 );
xor \U$9874 ( \10251 , \9861 , \9865 );
xor \U$9875 ( \10252 , \10251 , \9870 );
and \U$9876 ( \10253 , \10250 , \10252 );
xor \U$9877 ( \10254 , \9878 , \9882 );
xor \U$9878 ( \10255 , \10254 , \9887 );
and \U$9879 ( \10256 , \10252 , \10255 );
and \U$9880 ( \10257 , \10250 , \10255 );
or \U$9881 ( \10258 , \10253 , \10256 , \10257 );
and \U$9882 ( \10259 , \10247 , \10258 );
and \U$9883 ( \10260 , \10238 , \10258 );
or \U$9884 ( \10261 , \10248 , \10259 , \10260 );
and \U$9885 ( \10262 , \10206 , \10261 );
xor \U$9886 ( \10263 , \9790 , \9794 );
xor \U$9887 ( \10264 , \10263 , \9799 );
xor \U$9888 ( \10265 , \9754 , \9758 );
xor \U$9889 ( \10266 , \10265 , \9763 );
and \U$9890 ( \10267 , \10264 , \10266 );
xor \U$9891 ( \10268 , \9771 , \9775 );
xor \U$9892 ( \10269 , \10268 , \9780 );
and \U$9893 ( \10270 , \10266 , \10269 );
and \U$9894 ( \10271 , \10264 , \10269 );
or \U$9895 ( \10272 , \10267 , \10270 , \10271 );
xor \U$9896 ( \10273 , \9806 , \9810 );
xor \U$9897 ( \10274 , \10273 , \9815 );
xor \U$9898 ( \10275 , \9825 , \9829 );
xor \U$9899 ( \10276 , \10275 , \9834 );
and \U$9900 ( \10277 , \10274 , \10276 );
and \U$9901 ( \10278 , \10272 , \10277 );
xor \U$9902 ( \10279 , \9946 , \9948 );
xor \U$9903 ( \10280 , \10279 , \9951 );
and \U$9904 ( \10281 , \10277 , \10280 );
and \U$9905 ( \10282 , \10272 , \10280 );
or \U$9906 ( \10283 , \10278 , \10281 , \10282 );
and \U$9907 ( \10284 , \10261 , \10283 );
and \U$9908 ( \10285 , \10206 , \10283 );
or \U$9909 ( \10286 , \10262 , \10284 , \10285 );
xor \U$9910 ( \10287 , \9750 , \9766 );
xor \U$9911 ( \10288 , \10287 , \9783 );
xor \U$9912 ( \10289 , \9802 , \9818 );
xor \U$9913 ( \10290 , \10289 , \9837 );
and \U$9914 ( \10291 , \10288 , \10290 );
xor \U$9915 ( \10292 , \9857 , \9873 );
xor \U$9916 ( \10293 , \10292 , \9890 );
and \U$9917 ( \10294 , \10290 , \10293 );
and \U$9918 ( \10295 , \10288 , \10293 );
or \U$9919 ( \10296 , \10291 , \10294 , \10295 );
xor \U$9920 ( \10297 , \9898 , \9900 );
xor \U$9921 ( \10298 , \10297 , \9903 );
xor \U$9922 ( \10299 , \9908 , \9910 );
xor \U$9923 ( \10300 , \10299 , \9913 );
and \U$9924 ( \10301 , \10298 , \10300 );
xor \U$9925 ( \10302 , \9933 , \9935 );
xor \U$9926 ( \10303 , \10302 , \9937 );
and \U$9927 ( \10304 , \10300 , \10303 );
and \U$9928 ( \10305 , \10298 , \10303 );
or \U$9929 ( \10306 , \10301 , \10304 , \10305 );
and \U$9930 ( \10307 , \10296 , \10306 );
xor \U$9931 ( \10308 , \9967 , \9969 );
xor \U$9932 ( \10309 , \10308 , \9972 );
and \U$9933 ( \10310 , \10306 , \10309 );
and \U$9934 ( \10311 , \10296 , \10309 );
or \U$9935 ( \10312 , \10307 , \10310 , \10311 );
and \U$9936 ( \10313 , \10286 , \10312 );
xor \U$9937 ( \10314 , \9906 , \9916 );
xor \U$9938 ( \10315 , \10314 , \9940 );
xor \U$9939 ( \10316 , \9977 , \9979 );
xor \U$9940 ( \10317 , \10316 , \9982 );
and \U$9941 ( \10318 , \10315 , \10317 );
xor \U$9942 ( \10319 , \9954 , \9956 );
xor \U$9943 ( \10320 , \10319 , \9959 );
and \U$9944 ( \10321 , \10317 , \10320 );
and \U$9945 ( \10322 , \10315 , \10320 );
or \U$9946 ( \10323 , \10318 , \10321 , \10322 );
and \U$9947 ( \10324 , \10312 , \10323 );
and \U$9948 ( \10325 , \10286 , \10323 );
or \U$9949 ( \10326 , \10313 , \10324 , \10325 );
xor \U$9950 ( \10327 , \9491 , \9546 );
xor \U$9951 ( \10328 , \10327 , \9599 );
xor \U$9952 ( \10329 , \9627 , \9637 );
xor \U$9953 ( \10330 , \10329 , \9648 );
and \U$9954 ( \10331 , \10328 , \10330 );
xor \U$9955 ( \10332 , \9994 , \9996 );
xor \U$9956 ( \10333 , \10332 , \9999 );
and \U$9957 ( \10334 , \10330 , \10333 );
and \U$9958 ( \10335 , \10328 , \10333 );
or \U$9959 ( \10336 , \10331 , \10334 , \10335 );
and \U$9960 ( \10337 , \10326 , \10336 );
xor \U$9961 ( \10338 , \10007 , \10009 );
xor \U$9962 ( \10339 , \10338 , \10012 );
and \U$9963 ( \10340 , \10336 , \10339 );
and \U$9964 ( \10341 , \10326 , \10339 );
or \U$9965 ( \10342 , \10337 , \10340 , \10341 );
xor \U$9966 ( \10343 , \10005 , \10015 );
xor \U$9967 ( \10344 , \10343 , \10018 );
and \U$9968 ( \10345 , \10342 , \10344 );
xor \U$9969 ( \10346 , \10023 , \10025 );
xor \U$9970 ( \10347 , \10346 , \10028 );
and \U$9971 ( \10348 , \10344 , \10347 );
and \U$9972 ( \10349 , \10342 , \10347 );
or \U$9973 ( \10350 , \10345 , \10348 , \10349 );
xor \U$9974 ( \10351 , \10021 , \10031 );
xor \U$9975 ( \10352 , \10351 , \10034 );
and \U$9976 ( \10353 , \10350 , \10352 );
xor \U$9977 ( \10354 , \9704 , \9714 );
xor \U$9978 ( \10355 , \10354 , \9717 );
and \U$9979 ( \10356 , \10352 , \10355 );
and \U$9980 ( \10357 , \10350 , \10355 );
or \U$9981 ( \10358 , \10353 , \10356 , \10357 );
and \U$9982 ( \10359 , \10043 , \10358 );
xor \U$9983 ( \10360 , \10043 , \10358 );
xor \U$9984 ( \10361 , \10350 , \10352 );
xor \U$9985 ( \10362 , \10361 , \10355 );
xor \U$9986 ( \10363 , \10171 , \10175 );
xor \U$9987 ( \10364 , \10363 , \10180 );
xor \U$9988 ( \10365 , \10188 , \10192 );
xor \U$9989 ( \10366 , \10365 , \10197 );
and \U$9990 ( \10367 , \10364 , \10366 );
xor \U$9991 ( \10368 , \10118 , \10122 );
xor \U$9992 ( \10369 , \10368 , \10127 );
and \U$9993 ( \10370 , \10366 , \10369 );
and \U$9994 ( \10371 , \10364 , \10369 );
or \U$9995 ( \10372 , \10367 , \10370 , \10371 );
xor \U$9996 ( \10373 , \10102 , \10106 );
xor \U$9997 ( \10374 , \10373 , \10111 );
xor \U$9998 ( \10375 , \10210 , \10214 );
xor \U$9999 ( \10376 , \10375 , \10219 );
and \U$10000 ( \10377 , \10374 , \10376 );
xor \U$10001 ( \10378 , \10135 , \10139 );
xor \U$10002 ( \10379 , \10378 , \10144 );
and \U$10003 ( \10380 , \10376 , \10379 );
and \U$10004 ( \10381 , \10374 , \10379 );
or \U$10005 ( \10382 , \10377 , \10380 , \10381 );
and \U$10006 ( \10383 , \10372 , \10382 );
and \U$10007 ( \10384 , \8189 , \641 );
and \U$10008 ( \10385 , \7765 , \639 );
nor \U$10009 ( \10386 , \10384 , \10385 );
xnor \U$10010 ( \10387 , \10386 , \592 );
and \U$10011 ( \10388 , \8440 , \540 );
and \U$10012 ( \10389 , \8435 , \538 );
nor \U$10013 ( \10390 , \10388 , \10389 );
xnor \U$10014 ( \10391 , \10390 , \499 );
and \U$10015 ( \10392 , \10387 , \10391 );
and \U$10016 ( \10393 , \9043 , \470 );
and \U$10017 ( \10394 , \8759 , \468 );
nor \U$10018 ( \10395 , \10393 , \10394 );
xnor \U$10019 ( \10396 , \10395 , \440 );
and \U$10020 ( \10397 , \10391 , \10396 );
and \U$10021 ( \10398 , \10387 , \10396 );
or \U$10022 ( \10399 , \10392 , \10397 , \10398 );
and \U$10023 ( \10400 , \9620 , \422 );
and \U$10024 ( \10401 , \9612 , \420 );
nor \U$10025 ( \10402 , \10400 , \10401 );
xnor \U$10026 ( \10403 , \10402 , \403 );
and \U$10027 ( \10404 , \10228 , \385 );
and \U$10028 ( \10405 , \10223 , \383 );
nor \U$10029 ( \10406 , \10404 , \10405 );
xnor \U$10030 ( \10407 , \10406 , \390 );
and \U$10031 ( \10408 , \10403 , \10407 );
buf \U$10032 ( \10409 , RIc2294a0_127);
and \U$10033 ( \10410 , \10409 , \379 );
and \U$10034 ( \10411 , \10407 , \10410 );
and \U$10035 ( \10412 , \10403 , \10410 );
or \U$10036 ( \10413 , \10408 , \10411 , \10412 );
and \U$10037 ( \10414 , \10399 , \10413 );
xnor \U$10038 ( \10415 , \10227 , \10229 );
and \U$10039 ( \10416 , \10413 , \10415 );
and \U$10040 ( \10417 , \10399 , \10415 );
or \U$10041 ( \10418 , \10414 , \10416 , \10417 );
and \U$10042 ( \10419 , \10382 , \10418 );
and \U$10043 ( \10420 , \10372 , \10418 );
or \U$10044 ( \10421 , \10383 , \10419 , \10420 );
not \U$10045 ( \10422 , \9821 );
and \U$10046 ( \10423 , \392 , \10063 );
and \U$10047 ( \10424 , \378 , \10061 );
nor \U$10048 ( \10425 , \10423 , \10424 );
xnor \U$10049 ( \10426 , \10425 , \9824 );
and \U$10050 ( \10427 , \10422 , \10426 );
and \U$10051 ( \10428 , \431 , \9495 );
and \U$10052 ( \10429 , \410 , \9493 );
nor \U$10053 ( \10430 , \10428 , \10429 );
xnor \U$10054 ( \10431 , \10430 , \9185 );
and \U$10055 ( \10432 , \10426 , \10431 );
and \U$10056 ( \10433 , \10422 , \10431 );
or \U$10057 ( \10434 , \10427 , \10432 , \10433 );
and \U$10058 ( \10435 , \487 , \8958 );
and \U$10059 ( \10436 , \479 , \8956 );
nor \U$10060 ( \10437 , \10435 , \10436 );
xnor \U$10061 ( \10438 , \10437 , \8587 );
and \U$10062 ( \10439 , \561 , \8396 );
and \U$10063 ( \10440 , \556 , \8394 );
nor \U$10064 ( \10441 , \10439 , \10440 );
xnor \U$10065 ( \10442 , \10441 , \8078 );
and \U$10066 ( \10443 , \10438 , \10442 );
and \U$10067 ( \10444 , \666 , \7829 );
and \U$10068 ( \10445 , \615 , \7827 );
nor \U$10069 ( \10446 , \10444 , \10445 );
xnor \U$10070 ( \10447 , \10446 , \7580 );
and \U$10071 ( \10448 , \10442 , \10447 );
and \U$10072 ( \10449 , \10438 , \10447 );
or \U$10073 ( \10450 , \10443 , \10448 , \10449 );
and \U$10074 ( \10451 , \10434 , \10450 );
and \U$10075 ( \10452 , \771 , \7300 );
and \U$10076 ( \10453 , \743 , \7298 );
nor \U$10077 ( \10454 , \10452 , \10453 );
xnor \U$10078 ( \10455 , \10454 , \7040 );
and \U$10079 ( \10456 , \925 , \6806 );
and \U$10080 ( \10457 , \851 , \6804 );
nor \U$10081 ( \10458 , \10456 , \10457 );
xnor \U$10082 ( \10459 , \10458 , \6491 );
and \U$10083 ( \10460 , \10455 , \10459 );
and \U$10084 ( \10461 , \1050 , \6297 );
and \U$10085 ( \10462 , \987 , \6295 );
nor \U$10086 ( \10463 , \10461 , \10462 );
xnor \U$10087 ( \10464 , \10463 , \5957 );
and \U$10088 ( \10465 , \10459 , \10464 );
and \U$10089 ( \10466 , \10455 , \10464 );
or \U$10090 ( \10467 , \10460 , \10465 , \10466 );
and \U$10091 ( \10468 , \10450 , \10467 );
and \U$10092 ( \10469 , \10434 , \10467 );
or \U$10093 ( \10470 , \10451 , \10468 , \10469 );
and \U$10094 ( \10471 , \4841 , \1616 );
and \U$10095 ( \10472 , \4833 , \1614 );
nor \U$10096 ( \10473 , \10471 , \10472 );
xnor \U$10097 ( \10474 , \10473 , \1503 );
and \U$10098 ( \10475 , \5315 , \1422 );
and \U$10099 ( \10476 , \5310 , \1420 );
nor \U$10100 ( \10477 , \10475 , \10476 );
xnor \U$10101 ( \10478 , \10477 , \1286 );
and \U$10102 ( \10479 , \10474 , \10478 );
and \U$10103 ( \10480 , \5838 , \1222 );
and \U$10104 ( \10481 , \5579 , \1220 );
nor \U$10105 ( \10482 , \10480 , \10481 );
xnor \U$10106 ( \10483 , \10482 , \1144 );
and \U$10107 ( \10484 , \10478 , \10483 );
and \U$10108 ( \10485 , \10474 , \10483 );
or \U$10109 ( \10486 , \10479 , \10484 , \10485 );
and \U$10110 ( \10487 , \3951 , \2362 );
and \U$10111 ( \10488 , \3743 , \2360 );
nor \U$10112 ( \10489 , \10487 , \10488 );
xnor \U$10113 ( \10490 , \10489 , \2225 );
and \U$10114 ( \10491 , \4078 , \2156 );
and \U$10115 ( \10492 , \4073 , \2154 );
nor \U$10116 ( \10493 , \10491 , \10492 );
xnor \U$10117 ( \10494 , \10493 , \2004 );
and \U$10118 ( \10495 , \10490 , \10494 );
and \U$10119 ( \10496 , \4531 , \1888 );
and \U$10120 ( \10497 , \4334 , \1886 );
nor \U$10121 ( \10498 , \10496 , \10497 );
xnor \U$10122 ( \10499 , \10498 , \1732 );
and \U$10123 ( \10500 , \10494 , \10499 );
and \U$10124 ( \10501 , \10490 , \10499 );
or \U$10125 ( \10502 , \10495 , \10500 , \10501 );
and \U$10126 ( \10503 , \10486 , \10502 );
and \U$10127 ( \10504 , \6219 , \1058 );
and \U$10128 ( \10505 , \6210 , \1056 );
nor \U$10129 ( \10506 , \10504 , \10505 );
xnor \U$10130 ( \10507 , \10506 , \964 );
and \U$10131 ( \10508 , \6764 , \888 );
and \U$10132 ( \10509 , \6562 , \886 );
nor \U$10133 ( \10510 , \10508 , \10509 );
xnor \U$10134 ( \10511 , \10510 , \816 );
and \U$10135 ( \10512 , \10507 , \10511 );
and \U$10136 ( \10513 , \7239 , \754 );
and \U$10137 ( \10514 , \7067 , \752 );
nor \U$10138 ( \10515 , \10513 , \10514 );
xnor \U$10139 ( \10516 , \10515 , \711 );
and \U$10140 ( \10517 , \10511 , \10516 );
and \U$10141 ( \10518 , \10507 , \10516 );
or \U$10142 ( \10519 , \10512 , \10517 , \10518 );
and \U$10143 ( \10520 , \10502 , \10519 );
and \U$10144 ( \10521 , \10486 , \10519 );
or \U$10145 ( \10522 , \10503 , \10520 , \10521 );
and \U$10146 ( \10523 , \10470 , \10522 );
and \U$10147 ( \10524 , \1861 , \4417 );
and \U$10148 ( \10525 , \1853 , \4415 );
nor \U$10149 ( \10526 , \10524 , \10525 );
xnor \U$10150 ( \10527 , \10526 , \4274 );
and \U$10151 ( \10528 , \2109 , \4094 );
and \U$10152 ( \10529 , \2104 , \4092 );
nor \U$10153 ( \10530 , \10528 , \10529 );
xnor \U$10154 ( \10531 , \10530 , \3848 );
and \U$10155 ( \10532 , \10527 , \10531 );
and \U$10156 ( \10533 , \2439 , \3699 );
and \U$10157 ( \10534 , \2295 , \3697 );
nor \U$10158 ( \10535 , \10533 , \10534 );
xnor \U$10159 ( \10536 , \10535 , \3512 );
and \U$10160 ( \10537 , \10531 , \10536 );
and \U$10161 ( \10538 , \10527 , \10536 );
or \U$10162 ( \10539 , \10532 , \10537 , \10538 );
and \U$10163 ( \10540 , \2728 , \3386 );
and \U$10164 ( \10541 , \2703 , \3384 );
nor \U$10165 ( \10542 , \10540 , \10541 );
xnor \U$10166 ( \10543 , \10542 , \3181 );
and \U$10167 ( \10544 , \3069 , \2980 );
and \U$10168 ( \10545 , \2902 , \2978 );
nor \U$10169 ( \10546 , \10544 , \10545 );
xnor \U$10170 ( \10547 , \10546 , \2831 );
and \U$10171 ( \10548 , \10543 , \10547 );
and \U$10172 ( \10549 , \3326 , \2658 );
and \U$10173 ( \10550 , \3207 , \2656 );
nor \U$10174 ( \10551 , \10549 , \10550 );
xnor \U$10175 ( \10552 , \10551 , \2516 );
and \U$10176 ( \10553 , \10547 , \10552 );
and \U$10177 ( \10554 , \10543 , \10552 );
or \U$10178 ( \10555 , \10548 , \10553 , \10554 );
and \U$10179 ( \10556 , \10539 , \10555 );
and \U$10180 ( \10557 , \1336 , \5708 );
and \U$10181 ( \10558 , \1248 , \5706 );
nor \U$10182 ( \10559 , \10557 , \10558 );
xnor \U$10183 ( \10560 , \10559 , \5467 );
and \U$10184 ( \10561 , \1446 , \5242 );
and \U$10185 ( \10562 , \1441 , \5240 );
nor \U$10186 ( \10563 , \10561 , \10562 );
xnor \U$10187 ( \10564 , \10563 , \5054 );
and \U$10188 ( \10565 , \10560 , \10564 );
and \U$10189 ( \10566 , \1677 , \4868 );
and \U$10190 ( \10567 , \1562 , \4866 );
nor \U$10191 ( \10568 , \10566 , \10567 );
xnor \U$10192 ( \10569 , \10568 , \4636 );
and \U$10193 ( \10570 , \10564 , \10569 );
and \U$10194 ( \10571 , \10560 , \10569 );
or \U$10195 ( \10572 , \10565 , \10570 , \10571 );
and \U$10196 ( \10573 , \10555 , \10572 );
and \U$10197 ( \10574 , \10539 , \10572 );
or \U$10198 ( \10575 , \10556 , \10573 , \10574 );
and \U$10199 ( \10576 , \10522 , \10575 );
and \U$10200 ( \10577 , \10470 , \10575 );
or \U$10201 ( \10578 , \10523 , \10576 , \10577 );
and \U$10202 ( \10579 , \10421 , \10578 );
xor \U$10203 ( \10580 , \10155 , \10159 );
xor \U$10204 ( \10581 , \10580 , \10164 );
xor \U$10205 ( \10582 , \10047 , \10051 );
xor \U$10206 ( \10583 , \10582 , \10056 );
and \U$10207 ( \10584 , \10581 , \10583 );
xor \U$10208 ( \10585 , \10083 , \10087 );
xor \U$10209 ( \10586 , \10585 , \10092 );
and \U$10210 ( \10587 , \10583 , \10586 );
and \U$10211 ( \10588 , \10581 , \10586 );
or \U$10212 ( \10589 , \10584 , \10587 , \10588 );
xor \U$10213 ( \10590 , \10264 , \10266 );
xor \U$10214 ( \10591 , \10590 , \10269 );
and \U$10215 ( \10592 , \10589 , \10591 );
xor \U$10216 ( \10593 , \10274 , \10276 );
and \U$10217 ( \10594 , \10591 , \10593 );
and \U$10218 ( \10595 , \10589 , \10593 );
or \U$10219 ( \10596 , \10592 , \10594 , \10595 );
and \U$10220 ( \10597 , \10578 , \10596 );
and \U$10221 ( \10598 , \10421 , \10596 );
or \U$10222 ( \10599 , \10579 , \10597 , \10598 );
xor \U$10223 ( \10600 , \10059 , \10078 );
xor \U$10224 ( \10601 , \10600 , \10095 );
xor \U$10225 ( \10602 , \10114 , \10130 );
xor \U$10226 ( \10603 , \10602 , \10147 );
and \U$10227 ( \10604 , \10601 , \10603 );
xor \U$10228 ( \10605 , \10167 , \10183 );
xor \U$10229 ( \10606 , \10605 , \10200 );
and \U$10230 ( \10607 , \10603 , \10606 );
and \U$10231 ( \10608 , \10601 , \10606 );
or \U$10232 ( \10609 , \10604 , \10607 , \10608 );
xor \U$10233 ( \10610 , \10222 , \10230 );
xor \U$10234 ( \10611 , \10610 , \10235 );
xor \U$10235 ( \10612 , \10239 , \10241 );
xor \U$10236 ( \10613 , \10612 , \10244 );
and \U$10237 ( \10614 , \10611 , \10613 );
xor \U$10238 ( \10615 , \10250 , \10252 );
xor \U$10239 ( \10616 , \10615 , \10255 );
and \U$10240 ( \10617 , \10613 , \10616 );
and \U$10241 ( \10618 , \10611 , \10616 );
or \U$10242 ( \10619 , \10614 , \10617 , \10618 );
and \U$10243 ( \10620 , \10609 , \10619 );
xor \U$10244 ( \10621 , \10288 , \10290 );
xor \U$10245 ( \10622 , \10621 , \10293 );
and \U$10246 ( \10623 , \10619 , \10622 );
and \U$10247 ( \10624 , \10609 , \10622 );
or \U$10248 ( \10625 , \10620 , \10623 , \10624 );
and \U$10249 ( \10626 , \10599 , \10625 );
xor \U$10250 ( \10627 , \10238 , \10247 );
xor \U$10251 ( \10628 , \10627 , \10258 );
xor \U$10252 ( \10629 , \10272 , \10277 );
xor \U$10253 ( \10630 , \10629 , \10280 );
and \U$10254 ( \10631 , \10628 , \10630 );
xor \U$10255 ( \10632 , \10298 , \10300 );
xor \U$10256 ( \10633 , \10632 , \10303 );
and \U$10257 ( \10634 , \10630 , \10633 );
and \U$10258 ( \10635 , \10628 , \10633 );
or \U$10259 ( \10636 , \10631 , \10634 , \10635 );
and \U$10260 ( \10637 , \10625 , \10636 );
and \U$10261 ( \10638 , \10599 , \10636 );
or \U$10262 ( \10639 , \10626 , \10637 , \10638 );
xor \U$10263 ( \10640 , \9786 , \9840 );
xor \U$10264 ( \10641 , \10640 , \9893 );
xor \U$10265 ( \10642 , \10296 , \10306 );
xor \U$10266 ( \10643 , \10642 , \10309 );
and \U$10267 ( \10644 , \10641 , \10643 );
xor \U$10268 ( \10645 , \10315 , \10317 );
xor \U$10269 ( \10646 , \10645 , \10320 );
and \U$10270 ( \10647 , \10643 , \10646 );
and \U$10271 ( \10648 , \10641 , \10646 );
or \U$10272 ( \10649 , \10644 , \10647 , \10648 );
and \U$10273 ( \10650 , \10639 , \10649 );
xor \U$10274 ( \10651 , \9975 , \9985 );
xor \U$10275 ( \10652 , \10651 , \9988 );
and \U$10276 ( \10653 , \10649 , \10652 );
and \U$10277 ( \10654 , \10639 , \10652 );
or \U$10278 ( \10655 , \10650 , \10653 , \10654 );
xor \U$10279 ( \10656 , \9896 , \9943 );
xor \U$10280 ( \10657 , \10656 , \9962 );
xor \U$10281 ( \10658 , \10286 , \10312 );
xor \U$10282 ( \10659 , \10658 , \10323 );
and \U$10283 ( \10660 , \10657 , \10659 );
xor \U$10284 ( \10661 , \10328 , \10330 );
xor \U$10285 ( \10662 , \10661 , \10333 );
and \U$10286 ( \10663 , \10659 , \10662 );
and \U$10287 ( \10664 , \10657 , \10662 );
or \U$10288 ( \10665 , \10660 , \10663 , \10664 );
and \U$10289 ( \10666 , \10655 , \10665 );
xor \U$10290 ( \10667 , \9965 , \9991 );
xor \U$10291 ( \10668 , \10667 , \10002 );
and \U$10292 ( \10669 , \10665 , \10668 );
and \U$10293 ( \10670 , \10655 , \10668 );
or \U$10294 ( \10671 , \10666 , \10669 , \10670 );
xor \U$10295 ( \10672 , \10342 , \10344 );
xor \U$10296 ( \10673 , \10672 , \10347 );
and \U$10297 ( \10674 , \10671 , \10673 );
and \U$10298 ( \10675 , \10362 , \10674 );
xor \U$10299 ( \10676 , \10362 , \10674 );
xor \U$10300 ( \10677 , \10671 , \10673 );
xor \U$10301 ( \10678 , \10474 , \10478 );
xor \U$10302 ( \10679 , \10678 , \10483 );
xor \U$10303 ( \10680 , \10490 , \10494 );
xor \U$10304 ( \10681 , \10680 , \10499 );
and \U$10305 ( \10682 , \10679 , \10681 );
xor \U$10306 ( \10683 , \10543 , \10547 );
xor \U$10307 ( \10684 , \10683 , \10552 );
and \U$10308 ( \10685 , \10681 , \10684 );
and \U$10309 ( \10686 , \10679 , \10684 );
or \U$10310 ( \10687 , \10682 , \10685 , \10686 );
xor \U$10311 ( \10688 , \10387 , \10391 );
xor \U$10312 ( \10689 , \10688 , \10396 );
xor \U$10313 ( \10690 , \10403 , \10407 );
xor \U$10314 ( \10691 , \10690 , \10410 );
and \U$10315 ( \10692 , \10689 , \10691 );
xor \U$10316 ( \10693 , \10507 , \10511 );
xor \U$10317 ( \10694 , \10693 , \10516 );
and \U$10318 ( \10695 , \10691 , \10694 );
and \U$10319 ( \10696 , \10689 , \10694 );
or \U$10320 ( \10697 , \10692 , \10695 , \10696 );
and \U$10321 ( \10698 , \10687 , \10697 );
and \U$10322 ( \10699 , \7765 , \754 );
and \U$10323 ( \10700 , \7239 , \752 );
nor \U$10324 ( \10701 , \10699 , \10700 );
xnor \U$10325 ( \10702 , \10701 , \711 );
and \U$10326 ( \10703 , \8435 , \641 );
and \U$10327 ( \10704 , \8189 , \639 );
nor \U$10328 ( \10705 , \10703 , \10704 );
xnor \U$10329 ( \10706 , \10705 , \592 );
and \U$10330 ( \10707 , \10702 , \10706 );
and \U$10331 ( \10708 , \8759 , \540 );
and \U$10332 ( \10709 , \8440 , \538 );
nor \U$10333 ( \10710 , \10708 , \10709 );
xnor \U$10334 ( \10711 , \10710 , \499 );
and \U$10335 ( \10712 , \10706 , \10711 );
and \U$10336 ( \10713 , \10702 , \10711 );
or \U$10337 ( \10714 , \10707 , \10712 , \10713 );
and \U$10338 ( \10715 , \9612 , \470 );
and \U$10339 ( \10716 , \9043 , \468 );
nor \U$10340 ( \10717 , \10715 , \10716 );
xnor \U$10341 ( \10718 , \10717 , \440 );
and \U$10342 ( \10719 , \10223 , \422 );
and \U$10343 ( \10720 , \9620 , \420 );
nor \U$10344 ( \10721 , \10719 , \10720 );
xnor \U$10345 ( \10722 , \10721 , \403 );
and \U$10346 ( \10723 , \10718 , \10722 );
and \U$10347 ( \10724 , \10409 , \385 );
and \U$10348 ( \10725 , \10228 , \383 );
nor \U$10349 ( \10726 , \10724 , \10725 );
xnor \U$10350 ( \10727 , \10726 , \390 );
and \U$10351 ( \10728 , \10722 , \10727 );
and \U$10352 ( \10729 , \10718 , \10727 );
or \U$10353 ( \10730 , \10723 , \10728 , \10729 );
or \U$10354 ( \10731 , \10714 , \10730 );
and \U$10355 ( \10732 , \10697 , \10731 );
and \U$10356 ( \10733 , \10687 , \10731 );
or \U$10357 ( \10734 , \10698 , \10732 , \10733 );
and \U$10358 ( \10735 , \4833 , \1888 );
and \U$10359 ( \10736 , \4531 , \1886 );
nor \U$10360 ( \10737 , \10735 , \10736 );
xnor \U$10361 ( \10738 , \10737 , \1732 );
and \U$10362 ( \10739 , \5310 , \1616 );
and \U$10363 ( \10740 , \4841 , \1614 );
nor \U$10364 ( \10741 , \10739 , \10740 );
xnor \U$10365 ( \10742 , \10741 , \1503 );
and \U$10366 ( \10743 , \10738 , \10742 );
and \U$10367 ( \10744 , \5579 , \1422 );
and \U$10368 ( \10745 , \5315 , \1420 );
nor \U$10369 ( \10746 , \10744 , \10745 );
xnor \U$10370 ( \10747 , \10746 , \1286 );
and \U$10371 ( \10748 , \10742 , \10747 );
and \U$10372 ( \10749 , \10738 , \10747 );
or \U$10373 ( \10750 , \10743 , \10748 , \10749 );
and \U$10374 ( \10751 , \6210 , \1222 );
and \U$10375 ( \10752 , \5838 , \1220 );
nor \U$10376 ( \10753 , \10751 , \10752 );
xnor \U$10377 ( \10754 , \10753 , \1144 );
and \U$10378 ( \10755 , \6562 , \1058 );
and \U$10379 ( \10756 , \6219 , \1056 );
nor \U$10380 ( \10757 , \10755 , \10756 );
xnor \U$10381 ( \10758 , \10757 , \964 );
and \U$10382 ( \10759 , \10754 , \10758 );
and \U$10383 ( \10760 , \7067 , \888 );
and \U$10384 ( \10761 , \6764 , \886 );
nor \U$10385 ( \10762 , \10760 , \10761 );
xnor \U$10386 ( \10763 , \10762 , \816 );
and \U$10387 ( \10764 , \10758 , \10763 );
and \U$10388 ( \10765 , \10754 , \10763 );
or \U$10389 ( \10766 , \10759 , \10764 , \10765 );
and \U$10390 ( \10767 , \10750 , \10766 );
and \U$10391 ( \10768 , \3743 , \2658 );
and \U$10392 ( \10769 , \3326 , \2656 );
nor \U$10393 ( \10770 , \10768 , \10769 );
xnor \U$10394 ( \10771 , \10770 , \2516 );
and \U$10395 ( \10772 , \4073 , \2362 );
and \U$10396 ( \10773 , \3951 , \2360 );
nor \U$10397 ( \10774 , \10772 , \10773 );
xnor \U$10398 ( \10775 , \10774 , \2225 );
and \U$10399 ( \10776 , \10771 , \10775 );
and \U$10400 ( \10777 , \4334 , \2156 );
and \U$10401 ( \10778 , \4078 , \2154 );
nor \U$10402 ( \10779 , \10777 , \10778 );
xnor \U$10403 ( \10780 , \10779 , \2004 );
and \U$10404 ( \10781 , \10775 , \10780 );
and \U$10405 ( \10782 , \10771 , \10780 );
or \U$10406 ( \10783 , \10776 , \10781 , \10782 );
and \U$10407 ( \10784 , \10766 , \10783 );
and \U$10408 ( \10785 , \10750 , \10783 );
or \U$10409 ( \10786 , \10767 , \10784 , \10785 );
and \U$10410 ( \10787 , \1853 , \4868 );
and \U$10411 ( \10788 , \1677 , \4866 );
nor \U$10412 ( \10789 , \10787 , \10788 );
xnor \U$10413 ( \10790 , \10789 , \4636 );
and \U$10414 ( \10791 , \2104 , \4417 );
and \U$10415 ( \10792 , \1861 , \4415 );
nor \U$10416 ( \10793 , \10791 , \10792 );
xnor \U$10417 ( \10794 , \10793 , \4274 );
and \U$10418 ( \10795 , \10790 , \10794 );
and \U$10419 ( \10796 , \2295 , \4094 );
and \U$10420 ( \10797 , \2109 , \4092 );
nor \U$10421 ( \10798 , \10796 , \10797 );
xnor \U$10422 ( \10799 , \10798 , \3848 );
and \U$10423 ( \10800 , \10794 , \10799 );
and \U$10424 ( \10801 , \10790 , \10799 );
or \U$10425 ( \10802 , \10795 , \10800 , \10801 );
and \U$10426 ( \10803 , \2703 , \3699 );
and \U$10427 ( \10804 , \2439 , \3697 );
nor \U$10428 ( \10805 , \10803 , \10804 );
xnor \U$10429 ( \10806 , \10805 , \3512 );
and \U$10430 ( \10807 , \2902 , \3386 );
and \U$10431 ( \10808 , \2728 , \3384 );
nor \U$10432 ( \10809 , \10807 , \10808 );
xnor \U$10433 ( \10810 , \10809 , \3181 );
and \U$10434 ( \10811 , \10806 , \10810 );
and \U$10435 ( \10812 , \3207 , \2980 );
and \U$10436 ( \10813 , \3069 , \2978 );
nor \U$10437 ( \10814 , \10812 , \10813 );
xnor \U$10438 ( \10815 , \10814 , \2831 );
and \U$10439 ( \10816 , \10810 , \10815 );
and \U$10440 ( \10817 , \10806 , \10815 );
or \U$10441 ( \10818 , \10811 , \10816 , \10817 );
and \U$10442 ( \10819 , \10802 , \10818 );
and \U$10443 ( \10820 , \1248 , \6297 );
and \U$10444 ( \10821 , \1050 , \6295 );
nor \U$10445 ( \10822 , \10820 , \10821 );
xnor \U$10446 ( \10823 , \10822 , \5957 );
and \U$10447 ( \10824 , \1441 , \5708 );
and \U$10448 ( \10825 , \1336 , \5706 );
nor \U$10449 ( \10826 , \10824 , \10825 );
xnor \U$10450 ( \10827 , \10826 , \5467 );
and \U$10451 ( \10828 , \10823 , \10827 );
and \U$10452 ( \10829 , \1562 , \5242 );
and \U$10453 ( \10830 , \1446 , \5240 );
nor \U$10454 ( \10831 , \10829 , \10830 );
xnor \U$10455 ( \10832 , \10831 , \5054 );
and \U$10456 ( \10833 , \10827 , \10832 );
and \U$10457 ( \10834 , \10823 , \10832 );
or \U$10458 ( \10835 , \10828 , \10833 , \10834 );
and \U$10459 ( \10836 , \10818 , \10835 );
and \U$10460 ( \10837 , \10802 , \10835 );
or \U$10461 ( \10838 , \10819 , \10836 , \10837 );
and \U$10462 ( \10839 , \10786 , \10838 );
and \U$10463 ( \10840 , \479 , \9495 );
and \U$10464 ( \10841 , \431 , \9493 );
nor \U$10465 ( \10842 , \10840 , \10841 );
xnor \U$10466 ( \10843 , \10842 , \9185 );
and \U$10467 ( \10844 , \556 , \8958 );
and \U$10468 ( \10845 , \487 , \8956 );
nor \U$10469 ( \10846 , \10844 , \10845 );
xnor \U$10470 ( \10847 , \10846 , \8587 );
and \U$10471 ( \10848 , \10843 , \10847 );
and \U$10472 ( \10849 , \615 , \8396 );
and \U$10473 ( \10850 , \561 , \8394 );
nor \U$10474 ( \10851 , \10849 , \10850 );
xnor \U$10475 ( \10852 , \10851 , \8078 );
and \U$10476 ( \10853 , \10847 , \10852 );
and \U$10477 ( \10854 , \10843 , \10852 );
or \U$10478 ( \10855 , \10848 , \10853 , \10854 );
and \U$10479 ( \10856 , \743 , \7829 );
and \U$10480 ( \10857 , \666 , \7827 );
nor \U$10481 ( \10858 , \10856 , \10857 );
xnor \U$10482 ( \10859 , \10858 , \7580 );
and \U$10483 ( \10860 , \851 , \7300 );
and \U$10484 ( \10861 , \771 , \7298 );
nor \U$10485 ( \10862 , \10860 , \10861 );
xnor \U$10486 ( \10863 , \10862 , \7040 );
and \U$10487 ( \10864 , \10859 , \10863 );
and \U$10488 ( \10865 , \987 , \6806 );
and \U$10489 ( \10866 , \925 , \6804 );
nor \U$10490 ( \10867 , \10865 , \10866 );
xnor \U$10491 ( \10868 , \10867 , \6491 );
and \U$10492 ( \10869 , \10863 , \10868 );
and \U$10493 ( \10870 , \10859 , \10868 );
or \U$10494 ( \10871 , \10864 , \10869 , \10870 );
and \U$10495 ( \10872 , \10855 , \10871 );
buf \U$10496 ( \10873 , RIc225828_64);
xor \U$10497 ( \10874 , \9821 , \10873 );
not \U$10498 ( \10875 , \10873 );
and \U$10499 ( \10876 , \10874 , \10875 );
and \U$10500 ( \10877 , \378 , \10876 );
not \U$10501 ( \10878 , \10877 );
xnor \U$10502 ( \10879 , \10878 , \9821 );
and \U$10503 ( \10880 , \410 , \10063 );
and \U$10504 ( \10881 , \392 , \10061 );
nor \U$10505 ( \10882 , \10880 , \10881 );
xnor \U$10506 ( \10883 , \10882 , \9824 );
and \U$10507 ( \10884 , \10879 , \10883 );
and \U$10508 ( \10885 , \10871 , \10884 );
and \U$10509 ( \10886 , \10855 , \10884 );
or \U$10510 ( \10887 , \10872 , \10885 , \10886 );
and \U$10511 ( \10888 , \10838 , \10887 );
and \U$10512 ( \10889 , \10786 , \10887 );
or \U$10513 ( \10890 , \10839 , \10888 , \10889 );
and \U$10514 ( \10891 , \10734 , \10890 );
xor \U$10515 ( \10892 , \10527 , \10531 );
xor \U$10516 ( \10893 , \10892 , \10536 );
xor \U$10517 ( \10894 , \10455 , \10459 );
xor \U$10518 ( \10895 , \10894 , \10464 );
and \U$10519 ( \10896 , \10893 , \10895 );
xor \U$10520 ( \10897 , \10560 , \10564 );
xor \U$10521 ( \10898 , \10897 , \10569 );
and \U$10522 ( \10899 , \10895 , \10898 );
and \U$10523 ( \10900 , \10893 , \10898 );
or \U$10524 ( \10901 , \10896 , \10899 , \10900 );
xor \U$10525 ( \10902 , \10422 , \10426 );
xor \U$10526 ( \10903 , \10902 , \10431 );
xor \U$10527 ( \10904 , \10438 , \10442 );
xor \U$10528 ( \10905 , \10904 , \10447 );
and \U$10529 ( \10906 , \10903 , \10905 );
and \U$10530 ( \10907 , \10901 , \10906 );
xor \U$10531 ( \10908 , \10066 , \10070 );
xor \U$10532 ( \10909 , \10908 , \10075 );
and \U$10533 ( \10910 , \10906 , \10909 );
and \U$10534 ( \10911 , \10901 , \10909 );
or \U$10535 ( \10912 , \10907 , \10910 , \10911 );
and \U$10536 ( \10913 , \10890 , \10912 );
and \U$10537 ( \10914 , \10734 , \10912 );
or \U$10538 ( \10915 , \10891 , \10913 , \10914 );
xor \U$10539 ( \10916 , \10581 , \10583 );
xor \U$10540 ( \10917 , \10916 , \10586 );
xor \U$10541 ( \10918 , \10364 , \10366 );
xor \U$10542 ( \10919 , \10918 , \10369 );
and \U$10543 ( \10920 , \10917 , \10919 );
xor \U$10544 ( \10921 , \10374 , \10376 );
xor \U$10545 ( \10922 , \10921 , \10379 );
and \U$10546 ( \10923 , \10919 , \10922 );
and \U$10547 ( \10924 , \10917 , \10922 );
or \U$10548 ( \10925 , \10920 , \10923 , \10924 );
xor \U$10549 ( \10926 , \10486 , \10502 );
xor \U$10550 ( \10927 , \10926 , \10519 );
xor \U$10551 ( \10928 , \10539 , \10555 );
xor \U$10552 ( \10929 , \10928 , \10572 );
and \U$10553 ( \10930 , \10927 , \10929 );
xor \U$10554 ( \10931 , \10399 , \10413 );
xor \U$10555 ( \10932 , \10931 , \10415 );
and \U$10556 ( \10933 , \10929 , \10932 );
and \U$10557 ( \10934 , \10927 , \10932 );
or \U$10558 ( \10935 , \10930 , \10933 , \10934 );
and \U$10559 ( \10936 , \10925 , \10935 );
xor \U$10560 ( \10937 , \10601 , \10603 );
xor \U$10561 ( \10938 , \10937 , \10606 );
and \U$10562 ( \10939 , \10935 , \10938 );
and \U$10563 ( \10940 , \10925 , \10938 );
or \U$10564 ( \10941 , \10936 , \10939 , \10940 );
and \U$10565 ( \10942 , \10915 , \10941 );
xor \U$10566 ( \10943 , \10372 , \10382 );
xor \U$10567 ( \10944 , \10943 , \10418 );
xor \U$10568 ( \10945 , \10611 , \10613 );
xor \U$10569 ( \10946 , \10945 , \10616 );
and \U$10570 ( \10947 , \10944 , \10946 );
xor \U$10571 ( \10948 , \10589 , \10591 );
xor \U$10572 ( \10949 , \10948 , \10593 );
and \U$10573 ( \10950 , \10946 , \10949 );
and \U$10574 ( \10951 , \10944 , \10949 );
or \U$10575 ( \10952 , \10947 , \10950 , \10951 );
and \U$10576 ( \10953 , \10941 , \10952 );
and \U$10577 ( \10954 , \10915 , \10952 );
or \U$10578 ( \10955 , \10942 , \10953 , \10954 );
xor \U$10579 ( \10956 , \10098 , \10150 );
xor \U$10580 ( \10957 , \10956 , \10203 );
xor \U$10581 ( \10958 , \10609 , \10619 );
xor \U$10582 ( \10959 , \10958 , \10622 );
and \U$10583 ( \10960 , \10957 , \10959 );
xor \U$10584 ( \10961 , \10628 , \10630 );
xor \U$10585 ( \10962 , \10961 , \10633 );
and \U$10586 ( \10963 , \10959 , \10962 );
and \U$10587 ( \10964 , \10957 , \10962 );
or \U$10588 ( \10965 , \10960 , \10963 , \10964 );
and \U$10589 ( \10966 , \10955 , \10965 );
xor \U$10590 ( \10967 , \10206 , \10261 );
xor \U$10591 ( \10968 , \10967 , \10283 );
and \U$10592 ( \10969 , \10965 , \10968 );
and \U$10593 ( \10970 , \10955 , \10968 );
or \U$10594 ( \10971 , \10966 , \10969 , \10970 );
xor \U$10595 ( \10972 , \10639 , \10649 );
xor \U$10596 ( \10973 , \10972 , \10652 );
and \U$10597 ( \10974 , \10971 , \10973 );
xor \U$10598 ( \10975 , \10657 , \10659 );
xor \U$10599 ( \10976 , \10975 , \10662 );
and \U$10600 ( \10977 , \10973 , \10976 );
and \U$10601 ( \10978 , \10971 , \10976 );
or \U$10602 ( \10979 , \10974 , \10977 , \10978 );
xor \U$10603 ( \10980 , \10655 , \10665 );
xor \U$10604 ( \10981 , \10980 , \10668 );
and \U$10605 ( \10982 , \10979 , \10981 );
xor \U$10606 ( \10983 , \10326 , \10336 );
xor \U$10607 ( \10984 , \10983 , \10339 );
and \U$10608 ( \10985 , \10981 , \10984 );
and \U$10609 ( \10986 , \10979 , \10984 );
or \U$10610 ( \10987 , \10982 , \10985 , \10986 );
and \U$10611 ( \10988 , \10677 , \10987 );
xor \U$10612 ( \10989 , \10677 , \10987 );
xor \U$10613 ( \10990 , \10979 , \10981 );
xor \U$10614 ( \10991 , \10990 , \10984 );
xor \U$10615 ( \10992 , \10738 , \10742 );
xor \U$10616 ( \10993 , \10992 , \10747 );
xor \U$10617 ( \10994 , \10702 , \10706 );
xor \U$10618 ( \10995 , \10994 , \10711 );
and \U$10619 ( \10996 , \10993 , \10995 );
xor \U$10620 ( \10997 , \10754 , \10758 );
xor \U$10621 ( \10998 , \10997 , \10763 );
and \U$10622 ( \10999 , \10995 , \10998 );
and \U$10623 ( \11000 , \10993 , \10998 );
or \U$10624 ( \11001 , \10996 , \10999 , \11000 );
xor \U$10625 ( \11002 , \10790 , \10794 );
xor \U$10626 ( \11003 , \11002 , \10799 );
xor \U$10627 ( \11004 , \10806 , \10810 );
xor \U$10628 ( \11005 , \11004 , \10815 );
and \U$10629 ( \11006 , \11003 , \11005 );
xor \U$10630 ( \11007 , \10771 , \10775 );
xor \U$10631 ( \11008 , \11007 , \10780 );
and \U$10632 ( \11009 , \11005 , \11008 );
and \U$10633 ( \11010 , \11003 , \11008 );
or \U$10634 ( \11011 , \11006 , \11009 , \11010 );
and \U$10635 ( \11012 , \11001 , \11011 );
and \U$10636 ( \11013 , \8440 , \641 );
and \U$10637 ( \11014 , \8435 , \639 );
nor \U$10638 ( \11015 , \11013 , \11014 );
xnor \U$10639 ( \11016 , \11015 , \592 );
and \U$10640 ( \11017 , \9043 , \540 );
and \U$10641 ( \11018 , \8759 , \538 );
nor \U$10642 ( \11019 , \11017 , \11018 );
xnor \U$10643 ( \11020 , \11019 , \499 );
and \U$10644 ( \11021 , \11016 , \11020 );
and \U$10645 ( \11022 , \9620 , \470 );
and \U$10646 ( \11023 , \9612 , \468 );
nor \U$10647 ( \11024 , \11022 , \11023 );
xnor \U$10648 ( \11025 , \11024 , \440 );
and \U$10649 ( \11026 , \11020 , \11025 );
and \U$10650 ( \11027 , \11016 , \11025 );
or \U$10651 ( \11028 , \11021 , \11026 , \11027 );
buf \U$10652 ( \11029 , RIc229518_128);
nand \U$10653 ( \11030 , \11029 , \379 );
not \U$10654 ( \11031 , \11030 );
and \U$10655 ( \11032 , \11028 , \11031 );
xor \U$10656 ( \11033 , \10718 , \10722 );
xor \U$10657 ( \11034 , \11033 , \10727 );
and \U$10658 ( \11035 , \11031 , \11034 );
and \U$10659 ( \11036 , \11028 , \11034 );
or \U$10660 ( \11037 , \11032 , \11035 , \11036 );
and \U$10661 ( \11038 , \11011 , \11037 );
and \U$10662 ( \11039 , \11001 , \11037 );
or \U$10663 ( \11040 , \11012 , \11038 , \11039 );
and \U$10664 ( \11041 , \2109 , \4417 );
and \U$10665 ( \11042 , \2104 , \4415 );
nor \U$10666 ( \11043 , \11041 , \11042 );
xnor \U$10667 ( \11044 , \11043 , \4274 );
and \U$10668 ( \11045 , \2439 , \4094 );
and \U$10669 ( \11046 , \2295 , \4092 );
nor \U$10670 ( \11047 , \11045 , \11046 );
xnor \U$10671 ( \11048 , \11047 , \3848 );
and \U$10672 ( \11049 , \11044 , \11048 );
and \U$10673 ( \11050 , \2728 , \3699 );
and \U$10674 ( \11051 , \2703 , \3697 );
nor \U$10675 ( \11052 , \11050 , \11051 );
xnor \U$10676 ( \11053 , \11052 , \3512 );
and \U$10677 ( \11054 , \11048 , \11053 );
and \U$10678 ( \11055 , \11044 , \11053 );
or \U$10679 ( \11056 , \11049 , \11054 , \11055 );
and \U$10680 ( \11057 , \1446 , \5708 );
and \U$10681 ( \11058 , \1441 , \5706 );
nor \U$10682 ( \11059 , \11057 , \11058 );
xnor \U$10683 ( \11060 , \11059 , \5467 );
and \U$10684 ( \11061 , \1677 , \5242 );
and \U$10685 ( \11062 , \1562 , \5240 );
nor \U$10686 ( \11063 , \11061 , \11062 );
xnor \U$10687 ( \11064 , \11063 , \5054 );
and \U$10688 ( \11065 , \11060 , \11064 );
and \U$10689 ( \11066 , \1861 , \4868 );
and \U$10690 ( \11067 , \1853 , \4866 );
nor \U$10691 ( \11068 , \11066 , \11067 );
xnor \U$10692 ( \11069 , \11068 , \4636 );
and \U$10693 ( \11070 , \11064 , \11069 );
and \U$10694 ( \11071 , \11060 , \11069 );
or \U$10695 ( \11072 , \11065 , \11070 , \11071 );
and \U$10696 ( \11073 , \11056 , \11072 );
and \U$10697 ( \11074 , \3069 , \3386 );
and \U$10698 ( \11075 , \2902 , \3384 );
nor \U$10699 ( \11076 , \11074 , \11075 );
xnor \U$10700 ( \11077 , \11076 , \3181 );
and \U$10701 ( \11078 , \3326 , \2980 );
and \U$10702 ( \11079 , \3207 , \2978 );
nor \U$10703 ( \11080 , \11078 , \11079 );
xnor \U$10704 ( \11081 , \11080 , \2831 );
and \U$10705 ( \11082 , \11077 , \11081 );
and \U$10706 ( \11083 , \3951 , \2658 );
and \U$10707 ( \11084 , \3743 , \2656 );
nor \U$10708 ( \11085 , \11083 , \11084 );
xnor \U$10709 ( \11086 , \11085 , \2516 );
and \U$10710 ( \11087 , \11081 , \11086 );
and \U$10711 ( \11088 , \11077 , \11086 );
or \U$10712 ( \11089 , \11082 , \11087 , \11088 );
and \U$10713 ( \11090 , \11072 , \11089 );
and \U$10714 ( \11091 , \11056 , \11089 );
or \U$10715 ( \11092 , \11073 , \11090 , \11091 );
and \U$10716 ( \11093 , \925 , \7300 );
and \U$10717 ( \11094 , \851 , \7298 );
nor \U$10718 ( \11095 , \11093 , \11094 );
xnor \U$10719 ( \11096 , \11095 , \7040 );
and \U$10720 ( \11097 , \1050 , \6806 );
and \U$10721 ( \11098 , \987 , \6804 );
nor \U$10722 ( \11099 , \11097 , \11098 );
xnor \U$10723 ( \11100 , \11099 , \6491 );
and \U$10724 ( \11101 , \11096 , \11100 );
and \U$10725 ( \11102 , \1336 , \6297 );
and \U$10726 ( \11103 , \1248 , \6295 );
nor \U$10727 ( \11104 , \11102 , \11103 );
xnor \U$10728 ( \11105 , \11104 , \5957 );
and \U$10729 ( \11106 , \11100 , \11105 );
and \U$10730 ( \11107 , \11096 , \11105 );
or \U$10731 ( \11108 , \11101 , \11106 , \11107 );
and \U$10732 ( \11109 , \561 , \8958 );
and \U$10733 ( \11110 , \556 , \8956 );
nor \U$10734 ( \11111 , \11109 , \11110 );
xnor \U$10735 ( \11112 , \11111 , \8587 );
and \U$10736 ( \11113 , \666 , \8396 );
and \U$10737 ( \11114 , \615 , \8394 );
nor \U$10738 ( \11115 , \11113 , \11114 );
xnor \U$10739 ( \11116 , \11115 , \8078 );
and \U$10740 ( \11117 , \11112 , \11116 );
and \U$10741 ( \11118 , \771 , \7829 );
and \U$10742 ( \11119 , \743 , \7827 );
nor \U$10743 ( \11120 , \11118 , \11119 );
xnor \U$10744 ( \11121 , \11120 , \7580 );
and \U$10745 ( \11122 , \11116 , \11121 );
and \U$10746 ( \11123 , \11112 , \11121 );
or \U$10747 ( \11124 , \11117 , \11122 , \11123 );
and \U$10748 ( \11125 , \11108 , \11124 );
and \U$10749 ( \11126 , \392 , \10876 );
and \U$10750 ( \11127 , \378 , \10873 );
nor \U$10751 ( \11128 , \11126 , \11127 );
xnor \U$10752 ( \11129 , \11128 , \9821 );
and \U$10753 ( \11130 , \431 , \10063 );
and \U$10754 ( \11131 , \410 , \10061 );
nor \U$10755 ( \11132 , \11130 , \11131 );
xnor \U$10756 ( \11133 , \11132 , \9824 );
and \U$10757 ( \11134 , \11129 , \11133 );
and \U$10758 ( \11135 , \487 , \9495 );
and \U$10759 ( \11136 , \479 , \9493 );
nor \U$10760 ( \11137 , \11135 , \11136 );
xnor \U$10761 ( \11138 , \11137 , \9185 );
and \U$10762 ( \11139 , \11133 , \11138 );
and \U$10763 ( \11140 , \11129 , \11138 );
or \U$10764 ( \11141 , \11134 , \11139 , \11140 );
and \U$10765 ( \11142 , \11124 , \11141 );
and \U$10766 ( \11143 , \11108 , \11141 );
or \U$10767 ( \11144 , \11125 , \11142 , \11143 );
and \U$10768 ( \11145 , \11092 , \11144 );
and \U$10769 ( \11146 , \5315 , \1616 );
and \U$10770 ( \11147 , \5310 , \1614 );
nor \U$10771 ( \11148 , \11146 , \11147 );
xnor \U$10772 ( \11149 , \11148 , \1503 );
and \U$10773 ( \11150 , \5838 , \1422 );
and \U$10774 ( \11151 , \5579 , \1420 );
nor \U$10775 ( \11152 , \11150 , \11151 );
xnor \U$10776 ( \11153 , \11152 , \1286 );
and \U$10777 ( \11154 , \11149 , \11153 );
and \U$10778 ( \11155 , \6219 , \1222 );
and \U$10779 ( \11156 , \6210 , \1220 );
nor \U$10780 ( \11157 , \11155 , \11156 );
xnor \U$10781 ( \11158 , \11157 , \1144 );
and \U$10782 ( \11159 , \11153 , \11158 );
and \U$10783 ( \11160 , \11149 , \11158 );
or \U$10784 ( \11161 , \11154 , \11159 , \11160 );
and \U$10785 ( \11162 , \4078 , \2362 );
and \U$10786 ( \11163 , \4073 , \2360 );
nor \U$10787 ( \11164 , \11162 , \11163 );
xnor \U$10788 ( \11165 , \11164 , \2225 );
and \U$10789 ( \11166 , \4531 , \2156 );
and \U$10790 ( \11167 , \4334 , \2154 );
nor \U$10791 ( \11168 , \11166 , \11167 );
xnor \U$10792 ( \11169 , \11168 , \2004 );
and \U$10793 ( \11170 , \11165 , \11169 );
and \U$10794 ( \11171 , \4841 , \1888 );
and \U$10795 ( \11172 , \4833 , \1886 );
nor \U$10796 ( \11173 , \11171 , \11172 );
xnor \U$10797 ( \11174 , \11173 , \1732 );
and \U$10798 ( \11175 , \11169 , \11174 );
and \U$10799 ( \11176 , \11165 , \11174 );
or \U$10800 ( \11177 , \11170 , \11175 , \11176 );
and \U$10801 ( \11178 , \11161 , \11177 );
and \U$10802 ( \11179 , \6764 , \1058 );
and \U$10803 ( \11180 , \6562 , \1056 );
nor \U$10804 ( \11181 , \11179 , \11180 );
xnor \U$10805 ( \11182 , \11181 , \964 );
and \U$10806 ( \11183 , \7239 , \888 );
and \U$10807 ( \11184 , \7067 , \886 );
nor \U$10808 ( \11185 , \11183 , \11184 );
xnor \U$10809 ( \11186 , \11185 , \816 );
and \U$10810 ( \11187 , \11182 , \11186 );
and \U$10811 ( \11188 , \8189 , \754 );
and \U$10812 ( \11189 , \7765 , \752 );
nor \U$10813 ( \11190 , \11188 , \11189 );
xnor \U$10814 ( \11191 , \11190 , \711 );
and \U$10815 ( \11192 , \11186 , \11191 );
and \U$10816 ( \11193 , \11182 , \11191 );
or \U$10817 ( \11194 , \11187 , \11192 , \11193 );
and \U$10818 ( \11195 , \11177 , \11194 );
and \U$10819 ( \11196 , \11161 , \11194 );
or \U$10820 ( \11197 , \11178 , \11195 , \11196 );
and \U$10821 ( \11198 , \11144 , \11197 );
and \U$10822 ( \11199 , \11092 , \11197 );
or \U$10823 ( \11200 , \11145 , \11198 , \11199 );
and \U$10824 ( \11201 , \11040 , \11200 );
xor \U$10825 ( \11202 , \10843 , \10847 );
xor \U$10826 ( \11203 , \11202 , \10852 );
xor \U$10827 ( \11204 , \10859 , \10863 );
xor \U$10828 ( \11205 , \11204 , \10868 );
and \U$10829 ( \11206 , \11203 , \11205 );
xor \U$10830 ( \11207 , \10823 , \10827 );
xor \U$10831 ( \11208 , \11207 , \10832 );
and \U$10832 ( \11209 , \11205 , \11208 );
and \U$10833 ( \11210 , \11203 , \11208 );
or \U$10834 ( \11211 , \11206 , \11209 , \11210 );
xor \U$10835 ( \11212 , \10893 , \10895 );
xor \U$10836 ( \11213 , \11212 , \10898 );
and \U$10837 ( \11214 , \11211 , \11213 );
xor \U$10838 ( \11215 , \10903 , \10905 );
and \U$10839 ( \11216 , \11213 , \11215 );
and \U$10840 ( \11217 , \11211 , \11215 );
or \U$10841 ( \11218 , \11214 , \11216 , \11217 );
and \U$10842 ( \11219 , \11200 , \11218 );
and \U$10843 ( \11220 , \11040 , \11218 );
or \U$10844 ( \11221 , \11201 , \11219 , \11220 );
xor \U$10845 ( \11222 , \10750 , \10766 );
xor \U$10846 ( \11223 , \11222 , \10783 );
xor \U$10847 ( \11224 , \10802 , \10818 );
xor \U$10848 ( \11225 , \11224 , \10835 );
and \U$10849 ( \11226 , \11223 , \11225 );
xor \U$10850 ( \11227 , \10855 , \10871 );
xor \U$10851 ( \11228 , \11227 , \10884 );
and \U$10852 ( \11229 , \11225 , \11228 );
and \U$10853 ( \11230 , \11223 , \11228 );
or \U$10854 ( \11231 , \11226 , \11229 , \11230 );
xor \U$10855 ( \11232 , \10679 , \10681 );
xor \U$10856 ( \11233 , \11232 , \10684 );
xor \U$10857 ( \11234 , \10689 , \10691 );
xor \U$10858 ( \11235 , \11234 , \10694 );
and \U$10859 ( \11236 , \11233 , \11235 );
xnor \U$10860 ( \11237 , \10714 , \10730 );
and \U$10861 ( \11238 , \11235 , \11237 );
and \U$10862 ( \11239 , \11233 , \11237 );
or \U$10863 ( \11240 , \11236 , \11238 , \11239 );
and \U$10864 ( \11241 , \11231 , \11240 );
xor \U$10865 ( \11242 , \10434 , \10450 );
xor \U$10866 ( \11243 , \11242 , \10467 );
and \U$10867 ( \11244 , \11240 , \11243 );
and \U$10868 ( \11245 , \11231 , \11243 );
or \U$10869 ( \11246 , \11241 , \11244 , \11245 );
and \U$10870 ( \11247 , \11221 , \11246 );
xor \U$10871 ( \11248 , \10901 , \10906 );
xor \U$10872 ( \11249 , \11248 , \10909 );
xor \U$10873 ( \11250 , \10917 , \10919 );
xor \U$10874 ( \11251 , \11250 , \10922 );
and \U$10875 ( \11252 , \11249 , \11251 );
xor \U$10876 ( \11253 , \10927 , \10929 );
xor \U$10877 ( \11254 , \11253 , \10932 );
and \U$10878 ( \11255 , \11251 , \11254 );
and \U$10879 ( \11256 , \11249 , \11254 );
or \U$10880 ( \11257 , \11252 , \11255 , \11256 );
and \U$10881 ( \11258 , \11246 , \11257 );
and \U$10882 ( \11259 , \11221 , \11257 );
or \U$10883 ( \11260 , \11247 , \11258 , \11259 );
xor \U$10884 ( \11261 , \10470 , \10522 );
xor \U$10885 ( \11262 , \11261 , \10575 );
xor \U$10886 ( \11263 , \10925 , \10935 );
xor \U$10887 ( \11264 , \11263 , \10938 );
and \U$10888 ( \11265 , \11262 , \11264 );
xor \U$10889 ( \11266 , \10944 , \10946 );
xor \U$10890 ( \11267 , \11266 , \10949 );
and \U$10891 ( \11268 , \11264 , \11267 );
and \U$10892 ( \11269 , \11262 , \11267 );
or \U$10893 ( \11270 , \11265 , \11268 , \11269 );
and \U$10894 ( \11271 , \11260 , \11270 );
xor \U$10895 ( \11272 , \10421 , \10578 );
xor \U$10896 ( \11273 , \11272 , \10596 );
and \U$10897 ( \11274 , \11270 , \11273 );
and \U$10898 ( \11275 , \11260 , \11273 );
or \U$10899 ( \11276 , \11271 , \11274 , \11275 );
xor \U$10900 ( \11277 , \10915 , \10941 );
xor \U$10901 ( \11278 , \11277 , \10952 );
xor \U$10902 ( \11279 , \10957 , \10959 );
xor \U$10903 ( \11280 , \11279 , \10962 );
and \U$10904 ( \11281 , \11278 , \11280 );
and \U$10905 ( \11282 , \11276 , \11281 );
xor \U$10906 ( \11283 , \10641 , \10643 );
xor \U$10907 ( \11284 , \11283 , \10646 );
and \U$10908 ( \11285 , \11281 , \11284 );
and \U$10909 ( \11286 , \11276 , \11284 );
or \U$10910 ( \11287 , \11282 , \11285 , \11286 );
xor \U$10911 ( \11288 , \10599 , \10625 );
xor \U$10912 ( \11289 , \11288 , \10636 );
xor \U$10913 ( \11290 , \10955 , \10965 );
xor \U$10914 ( \11291 , \11290 , \10968 );
and \U$10915 ( \11292 , \11289 , \11291 );
and \U$10916 ( \11293 , \11287 , \11292 );
xor \U$10917 ( \11294 , \10971 , \10973 );
xor \U$10918 ( \11295 , \11294 , \10976 );
and \U$10919 ( \11296 , \11292 , \11295 );
and \U$10920 ( \11297 , \11287 , \11295 );
or \U$10921 ( \11298 , \11293 , \11296 , \11297 );
and \U$10922 ( \11299 , \10991 , \11298 );
xor \U$10923 ( \11300 , \10991 , \11298 );
xor \U$10924 ( \11301 , \11287 , \11292 );
xor \U$10925 ( \11302 , \11301 , \11295 );
and \U$10926 ( \11303 , \10223 , \470 );
and \U$10927 ( \11304 , \9620 , \468 );
nor \U$10928 ( \11305 , \11303 , \11304 );
xnor \U$10929 ( \11306 , \11305 , \440 );
and \U$10930 ( \11307 , \10409 , \422 );
and \U$10931 ( \11308 , \10228 , \420 );
nor \U$10932 ( \11309 , \11307 , \11308 );
xnor \U$10933 ( \11310 , \11309 , \403 );
and \U$10934 ( \11311 , \11306 , \11310 );
nand \U$10935 ( \11312 , \11029 , \383 );
xnor \U$10936 ( \11313 , \11312 , \390 );
and \U$10937 ( \11314 , \11310 , \11313 );
and \U$10938 ( \11315 , \11306 , \11313 );
or \U$10939 ( \11316 , \11311 , \11314 , \11315 );
and \U$10940 ( \11317 , \8435 , \754 );
and \U$10941 ( \11318 , \8189 , \752 );
nor \U$10942 ( \11319 , \11317 , \11318 );
xnor \U$10943 ( \11320 , \11319 , \711 );
and \U$10944 ( \11321 , \8759 , \641 );
and \U$10945 ( \11322 , \8440 , \639 );
nor \U$10946 ( \11323 , \11321 , \11322 );
xnor \U$10947 ( \11324 , \11323 , \592 );
and \U$10948 ( \11325 , \11320 , \11324 );
and \U$10949 ( \11326 , \9612 , \540 );
and \U$10950 ( \11327 , \9043 , \538 );
nor \U$10951 ( \11328 , \11326 , \11327 );
xnor \U$10952 ( \11329 , \11328 , \499 );
and \U$10953 ( \11330 , \11324 , \11329 );
and \U$10954 ( \11331 , \11320 , \11329 );
or \U$10955 ( \11332 , \11325 , \11330 , \11331 );
and \U$10956 ( \11333 , \11316 , \11332 );
and \U$10957 ( \11334 , \10228 , \422 );
and \U$10958 ( \11335 , \10223 , \420 );
nor \U$10959 ( \11336 , \11334 , \11335 );
xnor \U$10960 ( \11337 , \11336 , \403 );
and \U$10961 ( \11338 , \11332 , \11337 );
and \U$10962 ( \11339 , \11316 , \11337 );
or \U$10963 ( \11340 , \11333 , \11338 , \11339 );
and \U$10964 ( \11341 , \11029 , \385 );
and \U$10965 ( \11342 , \10409 , \383 );
nor \U$10966 ( \11343 , \11341 , \11342 );
xnor \U$10967 ( \11344 , \11343 , \390 );
xor \U$10968 ( \11345 , \11182 , \11186 );
xor \U$10969 ( \11346 , \11345 , \11191 );
and \U$10970 ( \11347 , \11344 , \11346 );
xor \U$10971 ( \11348 , \11016 , \11020 );
xor \U$10972 ( \11349 , \11348 , \11025 );
and \U$10973 ( \11350 , \11346 , \11349 );
and \U$10974 ( \11351 , \11344 , \11349 );
or \U$10975 ( \11352 , \11347 , \11350 , \11351 );
and \U$10976 ( \11353 , \11340 , \11352 );
xor \U$10977 ( \11354 , \11149 , \11153 );
xor \U$10978 ( \11355 , \11354 , \11158 );
xor \U$10979 ( \11356 , \11165 , \11169 );
xor \U$10980 ( \11357 , \11356 , \11174 );
and \U$10981 ( \11358 , \11355 , \11357 );
xor \U$10982 ( \11359 , \11077 , \11081 );
xor \U$10983 ( \11360 , \11359 , \11086 );
and \U$10984 ( \11361 , \11357 , \11360 );
and \U$10985 ( \11362 , \11355 , \11360 );
or \U$10986 ( \11363 , \11358 , \11361 , \11362 );
and \U$10987 ( \11364 , \11352 , \11363 );
and \U$10988 ( \11365 , \11340 , \11363 );
or \U$10989 ( \11366 , \11353 , \11364 , \11365 );
and \U$10990 ( \11367 , \5310 , \1888 );
and \U$10991 ( \11368 , \4841 , \1886 );
nor \U$10992 ( \11369 , \11367 , \11368 );
xnor \U$10993 ( \11370 , \11369 , \1732 );
and \U$10994 ( \11371 , \5579 , \1616 );
and \U$10995 ( \11372 , \5315 , \1614 );
nor \U$10996 ( \11373 , \11371 , \11372 );
xnor \U$10997 ( \11374 , \11373 , \1503 );
and \U$10998 ( \11375 , \11370 , \11374 );
and \U$10999 ( \11376 , \6210 , \1422 );
and \U$11000 ( \11377 , \5838 , \1420 );
nor \U$11001 ( \11378 , \11376 , \11377 );
xnor \U$11002 ( \11379 , \11378 , \1286 );
and \U$11003 ( \11380 , \11374 , \11379 );
and \U$11004 ( \11381 , \11370 , \11379 );
or \U$11005 ( \11382 , \11375 , \11380 , \11381 );
and \U$11006 ( \11383 , \4073 , \2658 );
and \U$11007 ( \11384 , \3951 , \2656 );
nor \U$11008 ( \11385 , \11383 , \11384 );
xnor \U$11009 ( \11386 , \11385 , \2516 );
and \U$11010 ( \11387 , \4334 , \2362 );
and \U$11011 ( \11388 , \4078 , \2360 );
nor \U$11012 ( \11389 , \11387 , \11388 );
xnor \U$11013 ( \11390 , \11389 , \2225 );
and \U$11014 ( \11391 , \11386 , \11390 );
and \U$11015 ( \11392 , \4833 , \2156 );
and \U$11016 ( \11393 , \4531 , \2154 );
nor \U$11017 ( \11394 , \11392 , \11393 );
xnor \U$11018 ( \11395 , \11394 , \2004 );
and \U$11019 ( \11396 , \11390 , \11395 );
and \U$11020 ( \11397 , \11386 , \11395 );
or \U$11021 ( \11398 , \11391 , \11396 , \11397 );
and \U$11022 ( \11399 , \11382 , \11398 );
and \U$11023 ( \11400 , \6562 , \1222 );
and \U$11024 ( \11401 , \6219 , \1220 );
nor \U$11025 ( \11402 , \11400 , \11401 );
xnor \U$11026 ( \11403 , \11402 , \1144 );
and \U$11027 ( \11404 , \7067 , \1058 );
and \U$11028 ( \11405 , \6764 , \1056 );
nor \U$11029 ( \11406 , \11404 , \11405 );
xnor \U$11030 ( \11407 , \11406 , \964 );
and \U$11031 ( \11408 , \11403 , \11407 );
and \U$11032 ( \11409 , \7765 , \888 );
and \U$11033 ( \11410 , \7239 , \886 );
nor \U$11034 ( \11411 , \11409 , \11410 );
xnor \U$11035 ( \11412 , \11411 , \816 );
and \U$11036 ( \11413 , \11407 , \11412 );
and \U$11037 ( \11414 , \11403 , \11412 );
or \U$11038 ( \11415 , \11408 , \11413 , \11414 );
and \U$11039 ( \11416 , \11398 , \11415 );
and \U$11040 ( \11417 , \11382 , \11415 );
or \U$11041 ( \11418 , \11399 , \11416 , \11417 );
and \U$11042 ( \11419 , \851 , \7829 );
and \U$11043 ( \11420 , \771 , \7827 );
nor \U$11044 ( \11421 , \11419 , \11420 );
xnor \U$11045 ( \11422 , \11421 , \7580 );
and \U$11046 ( \11423 , \987 , \7300 );
and \U$11047 ( \11424 , \925 , \7298 );
nor \U$11048 ( \11425 , \11423 , \11424 );
xnor \U$11049 ( \11426 , \11425 , \7040 );
and \U$11050 ( \11427 , \11422 , \11426 );
and \U$11051 ( \11428 , \1248 , \6806 );
and \U$11052 ( \11429 , \1050 , \6804 );
nor \U$11053 ( \11430 , \11428 , \11429 );
xnor \U$11054 ( \11431 , \11430 , \6491 );
and \U$11055 ( \11432 , \11426 , \11431 );
and \U$11056 ( \11433 , \11422 , \11431 );
or \U$11057 ( \11434 , \11427 , \11432 , \11433 );
and \U$11058 ( \11435 , \410 , \10876 );
and \U$11059 ( \11436 , \392 , \10873 );
nor \U$11060 ( \11437 , \11435 , \11436 );
xnor \U$11061 ( \11438 , \11437 , \9821 );
and \U$11062 ( \11439 , \479 , \10063 );
and \U$11063 ( \11440 , \431 , \10061 );
nor \U$11064 ( \11441 , \11439 , \11440 );
xnor \U$11065 ( \11442 , \11441 , \9824 );
and \U$11066 ( \11443 , \11438 , \11442 );
and \U$11067 ( \11444 , \11442 , \390 );
and \U$11068 ( \11445 , \11438 , \390 );
or \U$11069 ( \11446 , \11443 , \11444 , \11445 );
and \U$11070 ( \11447 , \11434 , \11446 );
and \U$11071 ( \11448 , \556 , \9495 );
and \U$11072 ( \11449 , \487 , \9493 );
nor \U$11073 ( \11450 , \11448 , \11449 );
xnor \U$11074 ( \11451 , \11450 , \9185 );
and \U$11075 ( \11452 , \615 , \8958 );
and \U$11076 ( \11453 , \561 , \8956 );
nor \U$11077 ( \11454 , \11452 , \11453 );
xnor \U$11078 ( \11455 , \11454 , \8587 );
and \U$11079 ( \11456 , \11451 , \11455 );
and \U$11080 ( \11457 , \743 , \8396 );
and \U$11081 ( \11458 , \666 , \8394 );
nor \U$11082 ( \11459 , \11457 , \11458 );
xnor \U$11083 ( \11460 , \11459 , \8078 );
and \U$11084 ( \11461 , \11455 , \11460 );
and \U$11085 ( \11462 , \11451 , \11460 );
or \U$11086 ( \11463 , \11456 , \11461 , \11462 );
and \U$11087 ( \11464 , \11446 , \11463 );
and \U$11088 ( \11465 , \11434 , \11463 );
or \U$11089 ( \11466 , \11447 , \11464 , \11465 );
and \U$11090 ( \11467 , \11418 , \11466 );
and \U$11091 ( \11468 , \2104 , \4868 );
and \U$11092 ( \11469 , \1861 , \4866 );
nor \U$11093 ( \11470 , \11468 , \11469 );
xnor \U$11094 ( \11471 , \11470 , \4636 );
and \U$11095 ( \11472 , \2295 , \4417 );
and \U$11096 ( \11473 , \2109 , \4415 );
nor \U$11097 ( \11474 , \11472 , \11473 );
xnor \U$11098 ( \11475 , \11474 , \4274 );
and \U$11099 ( \11476 , \11471 , \11475 );
and \U$11100 ( \11477 , \2703 , \4094 );
and \U$11101 ( \11478 , \2439 , \4092 );
nor \U$11102 ( \11479 , \11477 , \11478 );
xnor \U$11103 ( \11480 , \11479 , \3848 );
and \U$11104 ( \11481 , \11475 , \11480 );
and \U$11105 ( \11482 , \11471 , \11480 );
or \U$11106 ( \11483 , \11476 , \11481 , \11482 );
and \U$11107 ( \11484 , \1441 , \6297 );
and \U$11108 ( \11485 , \1336 , \6295 );
nor \U$11109 ( \11486 , \11484 , \11485 );
xnor \U$11110 ( \11487 , \11486 , \5957 );
and \U$11111 ( \11488 , \1562 , \5708 );
and \U$11112 ( \11489 , \1446 , \5706 );
nor \U$11113 ( \11490 , \11488 , \11489 );
xnor \U$11114 ( \11491 , \11490 , \5467 );
and \U$11115 ( \11492 , \11487 , \11491 );
and \U$11116 ( \11493 , \1853 , \5242 );
and \U$11117 ( \11494 , \1677 , \5240 );
nor \U$11118 ( \11495 , \11493 , \11494 );
xnor \U$11119 ( \11496 , \11495 , \5054 );
and \U$11120 ( \11497 , \11491 , \11496 );
and \U$11121 ( \11498 , \11487 , \11496 );
or \U$11122 ( \11499 , \11492 , \11497 , \11498 );
and \U$11123 ( \11500 , \11483 , \11499 );
and \U$11124 ( \11501 , \2902 , \3699 );
and \U$11125 ( \11502 , \2728 , \3697 );
nor \U$11126 ( \11503 , \11501 , \11502 );
xnor \U$11127 ( \11504 , \11503 , \3512 );
and \U$11128 ( \11505 , \3207 , \3386 );
and \U$11129 ( \11506 , \3069 , \3384 );
nor \U$11130 ( \11507 , \11505 , \11506 );
xnor \U$11131 ( \11508 , \11507 , \3181 );
and \U$11132 ( \11509 , \11504 , \11508 );
and \U$11133 ( \11510 , \3743 , \2980 );
and \U$11134 ( \11511 , \3326 , \2978 );
nor \U$11135 ( \11512 , \11510 , \11511 );
xnor \U$11136 ( \11513 , \11512 , \2831 );
and \U$11137 ( \11514 , \11508 , \11513 );
and \U$11138 ( \11515 , \11504 , \11513 );
or \U$11139 ( \11516 , \11509 , \11514 , \11515 );
and \U$11140 ( \11517 , \11499 , \11516 );
and \U$11141 ( \11518 , \11483 , \11516 );
or \U$11142 ( \11519 , \11500 , \11517 , \11518 );
and \U$11143 ( \11520 , \11466 , \11519 );
and \U$11144 ( \11521 , \11418 , \11519 );
or \U$11145 ( \11522 , \11467 , \11520 , \11521 );
and \U$11146 ( \11523 , \11366 , \11522 );
xor \U$11147 ( \11524 , \11044 , \11048 );
xor \U$11148 ( \11525 , \11524 , \11053 );
xor \U$11149 ( \11526 , \11060 , \11064 );
xor \U$11150 ( \11527 , \11526 , \11069 );
and \U$11151 ( \11528 , \11525 , \11527 );
xor \U$11152 ( \11529 , \11096 , \11100 );
xor \U$11153 ( \11530 , \11529 , \11105 );
and \U$11154 ( \11531 , \11527 , \11530 );
and \U$11155 ( \11532 , \11525 , \11530 );
or \U$11156 ( \11533 , \11528 , \11531 , \11532 );
xor \U$11157 ( \11534 , \11112 , \11116 );
xor \U$11158 ( \11535 , \11534 , \11121 );
xor \U$11159 ( \11536 , \11129 , \11133 );
xor \U$11160 ( \11537 , \11536 , \11138 );
and \U$11161 ( \11538 , \11535 , \11537 );
and \U$11162 ( \11539 , \11533 , \11538 );
xor \U$11163 ( \11540 , \10879 , \10883 );
and \U$11164 ( \11541 , \11538 , \11540 );
and \U$11165 ( \11542 , \11533 , \11540 );
or \U$11166 ( \11543 , \11539 , \11541 , \11542 );
and \U$11167 ( \11544 , \11522 , \11543 );
and \U$11168 ( \11545 , \11366 , \11543 );
or \U$11169 ( \11546 , \11523 , \11544 , \11545 );
xor \U$11170 ( \11547 , \11056 , \11072 );
xor \U$11171 ( \11548 , \11547 , \11089 );
xor \U$11172 ( \11549 , \11161 , \11177 );
xor \U$11173 ( \11550 , \11549 , \11194 );
and \U$11174 ( \11551 , \11548 , \11550 );
xor \U$11175 ( \11552 , \11028 , \11031 );
xor \U$11176 ( \11553 , \11552 , \11034 );
and \U$11177 ( \11554 , \11550 , \11553 );
and \U$11178 ( \11555 , \11548 , \11553 );
or \U$11179 ( \11556 , \11551 , \11554 , \11555 );
xor \U$11180 ( \11557 , \11203 , \11205 );
xor \U$11181 ( \11558 , \11557 , \11208 );
xor \U$11182 ( \11559 , \10993 , \10995 );
xor \U$11183 ( \11560 , \11559 , \10998 );
and \U$11184 ( \11561 , \11558 , \11560 );
xor \U$11185 ( \11562 , \11003 , \11005 );
xor \U$11186 ( \11563 , \11562 , \11008 );
and \U$11187 ( \11564 , \11560 , \11563 );
and \U$11188 ( \11565 , \11558 , \11563 );
or \U$11189 ( \11566 , \11561 , \11564 , \11565 );
and \U$11190 ( \11567 , \11556 , \11566 );
xor \U$11191 ( \11568 , \11223 , \11225 );
xor \U$11192 ( \11569 , \11568 , \11228 );
and \U$11193 ( \11570 , \11566 , \11569 );
and \U$11194 ( \11571 , \11556 , \11569 );
or \U$11195 ( \11572 , \11567 , \11570 , \11571 );
and \U$11196 ( \11573 , \11546 , \11572 );
xor \U$11197 ( \11574 , \11001 , \11011 );
xor \U$11198 ( \11575 , \11574 , \11037 );
xor \U$11199 ( \11576 , \11233 , \11235 );
xor \U$11200 ( \11577 , \11576 , \11237 );
and \U$11201 ( \11578 , \11575 , \11577 );
xor \U$11202 ( \11579 , \11211 , \11213 );
xor \U$11203 ( \11580 , \11579 , \11215 );
and \U$11204 ( \11581 , \11577 , \11580 );
and \U$11205 ( \11582 , \11575 , \11580 );
or \U$11206 ( \11583 , \11578 , \11581 , \11582 );
and \U$11207 ( \11584 , \11572 , \11583 );
and \U$11208 ( \11585 , \11546 , \11583 );
or \U$11209 ( \11586 , \11573 , \11584 , \11585 );
xor \U$11210 ( \11587 , \10687 , \10697 );
xor \U$11211 ( \11588 , \11587 , \10731 );
xor \U$11212 ( \11589 , \10786 , \10838 );
xor \U$11213 ( \11590 , \11589 , \10887 );
and \U$11214 ( \11591 , \11588 , \11590 );
xor \U$11215 ( \11592 , \11249 , \11251 );
xor \U$11216 ( \11593 , \11592 , \11254 );
and \U$11217 ( \11594 , \11590 , \11593 );
and \U$11218 ( \11595 , \11588 , \11593 );
or \U$11219 ( \11596 , \11591 , \11594 , \11595 );
and \U$11220 ( \11597 , \11586 , \11596 );
xor \U$11221 ( \11598 , \10734 , \10890 );
xor \U$11222 ( \11599 , \11598 , \10912 );
and \U$11223 ( \11600 , \11596 , \11599 );
and \U$11224 ( \11601 , \11586 , \11599 );
or \U$11225 ( \11602 , \11597 , \11600 , \11601 );
xor \U$11226 ( \11603 , \11260 , \11270 );
xor \U$11227 ( \11604 , \11603 , \11273 );
and \U$11228 ( \11605 , \11602 , \11604 );
xor \U$11229 ( \11606 , \11278 , \11280 );
and \U$11230 ( \11607 , \11604 , \11606 );
and \U$11231 ( \11608 , \11602 , \11606 );
or \U$11232 ( \11609 , \11605 , \11607 , \11608 );
xor \U$11233 ( \11610 , \11276 , \11281 );
xor \U$11234 ( \11611 , \11610 , \11284 );
and \U$11235 ( \11612 , \11609 , \11611 );
xor \U$11236 ( \11613 , \11289 , \11291 );
and \U$11237 ( \11614 , \11611 , \11613 );
and \U$11238 ( \11615 , \11609 , \11613 );
or \U$11239 ( \11616 , \11612 , \11614 , \11615 );
and \U$11240 ( \11617 , \11302 , \11616 );
xor \U$11241 ( \11618 , \11302 , \11616 );
xor \U$11242 ( \11619 , \11609 , \11611 );
xor \U$11243 ( \11620 , \11619 , \11613 );
and \U$11244 ( \11621 , \666 , \8958 );
and \U$11245 ( \11622 , \615 , \8956 );
nor \U$11246 ( \11623 , \11621 , \11622 );
xnor \U$11247 ( \11624 , \11623 , \8587 );
and \U$11248 ( \11625 , \771 , \8396 );
and \U$11249 ( \11626 , \743 , \8394 );
nor \U$11250 ( \11627 , \11625 , \11626 );
xnor \U$11251 ( \11628 , \11627 , \8078 );
and \U$11252 ( \11629 , \11624 , \11628 );
and \U$11253 ( \11630 , \925 , \7829 );
and \U$11254 ( \11631 , \851 , \7827 );
nor \U$11255 ( \11632 , \11630 , \11631 );
xnor \U$11256 ( \11633 , \11632 , \7580 );
and \U$11257 ( \11634 , \11628 , \11633 );
and \U$11258 ( \11635 , \11624 , \11633 );
or \U$11259 ( \11636 , \11629 , \11634 , \11635 );
and \U$11260 ( \11637 , \431 , \10876 );
and \U$11261 ( \11638 , \410 , \10873 );
nor \U$11262 ( \11639 , \11637 , \11638 );
xnor \U$11263 ( \11640 , \11639 , \9821 );
and \U$11264 ( \11641 , \487 , \10063 );
and \U$11265 ( \11642 , \479 , \10061 );
nor \U$11266 ( \11643 , \11641 , \11642 );
xnor \U$11267 ( \11644 , \11643 , \9824 );
and \U$11268 ( \11645 , \11640 , \11644 );
and \U$11269 ( \11646 , \561 , \9495 );
and \U$11270 ( \11647 , \556 , \9493 );
nor \U$11271 ( \11648 , \11646 , \11647 );
xnor \U$11272 ( \11649 , \11648 , \9185 );
and \U$11273 ( \11650 , \11644 , \11649 );
and \U$11274 ( \11651 , \11640 , \11649 );
or \U$11275 ( \11652 , \11645 , \11650 , \11651 );
and \U$11276 ( \11653 , \11636 , \11652 );
and \U$11277 ( \11654 , \1050 , \7300 );
and \U$11278 ( \11655 , \987 , \7298 );
nor \U$11279 ( \11656 , \11654 , \11655 );
xnor \U$11280 ( \11657 , \11656 , \7040 );
and \U$11281 ( \11658 , \1336 , \6806 );
and \U$11282 ( \11659 , \1248 , \6804 );
nor \U$11283 ( \11660 , \11658 , \11659 );
xnor \U$11284 ( \11661 , \11660 , \6491 );
and \U$11285 ( \11662 , \11657 , \11661 );
and \U$11286 ( \11663 , \1446 , \6297 );
and \U$11287 ( \11664 , \1441 , \6295 );
nor \U$11288 ( \11665 , \11663 , \11664 );
xnor \U$11289 ( \11666 , \11665 , \5957 );
and \U$11290 ( \11667 , \11661 , \11666 );
and \U$11291 ( \11668 , \11657 , \11666 );
or \U$11292 ( \11669 , \11662 , \11667 , \11668 );
and \U$11293 ( \11670 , \11652 , \11669 );
and \U$11294 ( \11671 , \11636 , \11669 );
or \U$11295 ( \11672 , \11653 , \11670 , \11671 );
and \U$11296 ( \11673 , \5838 , \1616 );
and \U$11297 ( \11674 , \5579 , \1614 );
nor \U$11298 ( \11675 , \11673 , \11674 );
xnor \U$11299 ( \11676 , \11675 , \1503 );
and \U$11300 ( \11677 , \6219 , \1422 );
and \U$11301 ( \11678 , \6210 , \1420 );
nor \U$11302 ( \11679 , \11677 , \11678 );
xnor \U$11303 ( \11680 , \11679 , \1286 );
and \U$11304 ( \11681 , \11676 , \11680 );
and \U$11305 ( \11682 , \6764 , \1222 );
and \U$11306 ( \11683 , \6562 , \1220 );
nor \U$11307 ( \11684 , \11682 , \11683 );
xnor \U$11308 ( \11685 , \11684 , \1144 );
and \U$11309 ( \11686 , \11680 , \11685 );
and \U$11310 ( \11687 , \11676 , \11685 );
or \U$11311 ( \11688 , \11681 , \11686 , \11687 );
and \U$11312 ( \11689 , \7239 , \1058 );
and \U$11313 ( \11690 , \7067 , \1056 );
nor \U$11314 ( \11691 , \11689 , \11690 );
xnor \U$11315 ( \11692 , \11691 , \964 );
and \U$11316 ( \11693 , \8189 , \888 );
and \U$11317 ( \11694 , \7765 , \886 );
nor \U$11318 ( \11695 , \11693 , \11694 );
xnor \U$11319 ( \11696 , \11695 , \816 );
and \U$11320 ( \11697 , \11692 , \11696 );
and \U$11321 ( \11698 , \8440 , \754 );
and \U$11322 ( \11699 , \8435 , \752 );
nor \U$11323 ( \11700 , \11698 , \11699 );
xnor \U$11324 ( \11701 , \11700 , \711 );
and \U$11325 ( \11702 , \11696 , \11701 );
and \U$11326 ( \11703 , \11692 , \11701 );
or \U$11327 ( \11704 , \11697 , \11702 , \11703 );
and \U$11328 ( \11705 , \11688 , \11704 );
and \U$11329 ( \11706 , \4531 , \2362 );
and \U$11330 ( \11707 , \4334 , \2360 );
nor \U$11331 ( \11708 , \11706 , \11707 );
xnor \U$11332 ( \11709 , \11708 , \2225 );
and \U$11333 ( \11710 , \4841 , \2156 );
and \U$11334 ( \11711 , \4833 , \2154 );
nor \U$11335 ( \11712 , \11710 , \11711 );
xnor \U$11336 ( \11713 , \11712 , \2004 );
and \U$11337 ( \11714 , \11709 , \11713 );
and \U$11338 ( \11715 , \5315 , \1888 );
and \U$11339 ( \11716 , \5310 , \1886 );
nor \U$11340 ( \11717 , \11715 , \11716 );
xnor \U$11341 ( \11718 , \11717 , \1732 );
and \U$11342 ( \11719 , \11713 , \11718 );
and \U$11343 ( \11720 , \11709 , \11718 );
or \U$11344 ( \11721 , \11714 , \11719 , \11720 );
and \U$11345 ( \11722 , \11704 , \11721 );
and \U$11346 ( \11723 , \11688 , \11721 );
or \U$11347 ( \11724 , \11705 , \11722 , \11723 );
and \U$11348 ( \11725 , \11672 , \11724 );
and \U$11349 ( \11726 , \1677 , \5708 );
and \U$11350 ( \11727 , \1562 , \5706 );
nor \U$11351 ( \11728 , \11726 , \11727 );
xnor \U$11352 ( \11729 , \11728 , \5467 );
and \U$11353 ( \11730 , \1861 , \5242 );
and \U$11354 ( \11731 , \1853 , \5240 );
nor \U$11355 ( \11732 , \11730 , \11731 );
xnor \U$11356 ( \11733 , \11732 , \5054 );
and \U$11357 ( \11734 , \11729 , \11733 );
and \U$11358 ( \11735 , \2109 , \4868 );
and \U$11359 ( \11736 , \2104 , \4866 );
nor \U$11360 ( \11737 , \11735 , \11736 );
xnor \U$11361 ( \11738 , \11737 , \4636 );
and \U$11362 ( \11739 , \11733 , \11738 );
and \U$11363 ( \11740 , \11729 , \11738 );
or \U$11364 ( \11741 , \11734 , \11739 , \11740 );
and \U$11365 ( \11742 , \3326 , \3386 );
and \U$11366 ( \11743 , \3207 , \3384 );
nor \U$11367 ( \11744 , \11742 , \11743 );
xnor \U$11368 ( \11745 , \11744 , \3181 );
and \U$11369 ( \11746 , \3951 , \2980 );
and \U$11370 ( \11747 , \3743 , \2978 );
nor \U$11371 ( \11748 , \11746 , \11747 );
xnor \U$11372 ( \11749 , \11748 , \2831 );
and \U$11373 ( \11750 , \11745 , \11749 );
and \U$11374 ( \11751 , \4078 , \2658 );
and \U$11375 ( \11752 , \4073 , \2656 );
nor \U$11376 ( \11753 , \11751 , \11752 );
xnor \U$11377 ( \11754 , \11753 , \2516 );
and \U$11378 ( \11755 , \11749 , \11754 );
and \U$11379 ( \11756 , \11745 , \11754 );
or \U$11380 ( \11757 , \11750 , \11755 , \11756 );
and \U$11381 ( \11758 , \11741 , \11757 );
and \U$11382 ( \11759 , \2439 , \4417 );
and \U$11383 ( \11760 , \2295 , \4415 );
nor \U$11384 ( \11761 , \11759 , \11760 );
xnor \U$11385 ( \11762 , \11761 , \4274 );
and \U$11386 ( \11763 , \2728 , \4094 );
and \U$11387 ( \11764 , \2703 , \4092 );
nor \U$11388 ( \11765 , \11763 , \11764 );
xnor \U$11389 ( \11766 , \11765 , \3848 );
and \U$11390 ( \11767 , \11762 , \11766 );
and \U$11391 ( \11768 , \3069 , \3699 );
and \U$11392 ( \11769 , \2902 , \3697 );
nor \U$11393 ( \11770 , \11768 , \11769 );
xnor \U$11394 ( \11771 , \11770 , \3512 );
and \U$11395 ( \11772 , \11766 , \11771 );
and \U$11396 ( \11773 , \11762 , \11771 );
or \U$11397 ( \11774 , \11767 , \11772 , \11773 );
and \U$11398 ( \11775 , \11757 , \11774 );
and \U$11399 ( \11776 , \11741 , \11774 );
or \U$11400 ( \11777 , \11758 , \11775 , \11776 );
and \U$11401 ( \11778 , \11724 , \11777 );
and \U$11402 ( \11779 , \11672 , \11777 );
or \U$11403 ( \11780 , \11725 , \11778 , \11779 );
xor \U$11404 ( \11781 , \11471 , \11475 );
xor \U$11405 ( \11782 , \11781 , \11480 );
xor \U$11406 ( \11783 , \11487 , \11491 );
xor \U$11407 ( \11784 , \11783 , \11496 );
and \U$11408 ( \11785 , \11782 , \11784 );
xor \U$11409 ( \11786 , \11504 , \11508 );
xor \U$11410 ( \11787 , \11786 , \11513 );
and \U$11411 ( \11788 , \11784 , \11787 );
and \U$11412 ( \11789 , \11782 , \11787 );
or \U$11413 ( \11790 , \11785 , \11788 , \11789 );
and \U$11414 ( \11791 , \9043 , \641 );
and \U$11415 ( \11792 , \8759 , \639 );
nor \U$11416 ( \11793 , \11791 , \11792 );
xnor \U$11417 ( \11794 , \11793 , \592 );
and \U$11418 ( \11795 , \9620 , \540 );
and \U$11419 ( \11796 , \9612 , \538 );
nor \U$11420 ( \11797 , \11795 , \11796 );
xnor \U$11421 ( \11798 , \11797 , \499 );
and \U$11422 ( \11799 , \11794 , \11798 );
and \U$11423 ( \11800 , \10228 , \470 );
and \U$11424 ( \11801 , \10223 , \468 );
nor \U$11425 ( \11802 , \11800 , \11801 );
xnor \U$11426 ( \11803 , \11802 , \440 );
and \U$11427 ( \11804 , \11798 , \11803 );
and \U$11428 ( \11805 , \11794 , \11803 );
or \U$11429 ( \11806 , \11799 , \11804 , \11805 );
xor \U$11430 ( \11807 , \11306 , \11310 );
xor \U$11431 ( \11808 , \11807 , \11313 );
and \U$11432 ( \11809 , \11806 , \11808 );
xor \U$11433 ( \11810 , \11320 , \11324 );
xor \U$11434 ( \11811 , \11810 , \11329 );
and \U$11435 ( \11812 , \11808 , \11811 );
and \U$11436 ( \11813 , \11806 , \11811 );
or \U$11437 ( \11814 , \11809 , \11812 , \11813 );
and \U$11438 ( \11815 , \11790 , \11814 );
xor \U$11439 ( \11816 , \11370 , \11374 );
xor \U$11440 ( \11817 , \11816 , \11379 );
xor \U$11441 ( \11818 , \11386 , \11390 );
xor \U$11442 ( \11819 , \11818 , \11395 );
and \U$11443 ( \11820 , \11817 , \11819 );
xor \U$11444 ( \11821 , \11403 , \11407 );
xor \U$11445 ( \11822 , \11821 , \11412 );
and \U$11446 ( \11823 , \11819 , \11822 );
and \U$11447 ( \11824 , \11817 , \11822 );
or \U$11448 ( \11825 , \11820 , \11823 , \11824 );
and \U$11449 ( \11826 , \11814 , \11825 );
and \U$11450 ( \11827 , \11790 , \11825 );
or \U$11451 ( \11828 , \11815 , \11826 , \11827 );
and \U$11452 ( \11829 , \11780 , \11828 );
xor \U$11453 ( \11830 , \11422 , \11426 );
xor \U$11454 ( \11831 , \11830 , \11431 );
xor \U$11455 ( \11832 , \11438 , \11442 );
xor \U$11456 ( \11833 , \11832 , \390 );
and \U$11457 ( \11834 , \11831 , \11833 );
xor \U$11458 ( \11835 , \11451 , \11455 );
xor \U$11459 ( \11836 , \11835 , \11460 );
and \U$11460 ( \11837 , \11833 , \11836 );
and \U$11461 ( \11838 , \11831 , \11836 );
or \U$11462 ( \11839 , \11834 , \11837 , \11838 );
xor \U$11463 ( \11840 , \11525 , \11527 );
xor \U$11464 ( \11841 , \11840 , \11530 );
and \U$11465 ( \11842 , \11839 , \11841 );
xor \U$11466 ( \11843 , \11535 , \11537 );
and \U$11467 ( \11844 , \11841 , \11843 );
and \U$11468 ( \11845 , \11839 , \11843 );
or \U$11469 ( \11846 , \11842 , \11844 , \11845 );
and \U$11470 ( \11847 , \11828 , \11846 );
and \U$11471 ( \11848 , \11780 , \11846 );
or \U$11472 ( \11849 , \11829 , \11847 , \11848 );
xor \U$11473 ( \11850 , \11382 , \11398 );
xor \U$11474 ( \11851 , \11850 , \11415 );
xor \U$11475 ( \11852 , \11434 , \11446 );
xor \U$11476 ( \11853 , \11852 , \11463 );
and \U$11477 ( \11854 , \11851 , \11853 );
xor \U$11478 ( \11855 , \11483 , \11499 );
xor \U$11479 ( \11856 , \11855 , \11516 );
and \U$11480 ( \11857 , \11853 , \11856 );
and \U$11481 ( \11858 , \11851 , \11856 );
or \U$11482 ( \11859 , \11854 , \11857 , \11858 );
xor \U$11483 ( \11860 , \11316 , \11332 );
xor \U$11484 ( \11861 , \11860 , \11337 );
xor \U$11485 ( \11862 , \11344 , \11346 );
xor \U$11486 ( \11863 , \11862 , \11349 );
and \U$11487 ( \11864 , \11861 , \11863 );
xor \U$11488 ( \11865 , \11355 , \11357 );
xor \U$11489 ( \11866 , \11865 , \11360 );
and \U$11490 ( \11867 , \11863 , \11866 );
and \U$11491 ( \11868 , \11861 , \11866 );
or \U$11492 ( \11869 , \11864 , \11867 , \11868 );
and \U$11493 ( \11870 , \11859 , \11869 );
xor \U$11494 ( \11871 , \11108 , \11124 );
xor \U$11495 ( \11872 , \11871 , \11141 );
and \U$11496 ( \11873 , \11869 , \11872 );
and \U$11497 ( \11874 , \11859 , \11872 );
or \U$11498 ( \11875 , \11870 , \11873 , \11874 );
and \U$11499 ( \11876 , \11849 , \11875 );
xor \U$11500 ( \11877 , \11548 , \11550 );
xor \U$11501 ( \11878 , \11877 , \11553 );
xor \U$11502 ( \11879 , \11558 , \11560 );
xor \U$11503 ( \11880 , \11879 , \11563 );
and \U$11504 ( \11881 , \11878 , \11880 );
xor \U$11505 ( \11882 , \11533 , \11538 );
xor \U$11506 ( \11883 , \11882 , \11540 );
and \U$11507 ( \11884 , \11880 , \11883 );
and \U$11508 ( \11885 , \11878 , \11883 );
or \U$11509 ( \11886 , \11881 , \11884 , \11885 );
and \U$11510 ( \11887 , \11875 , \11886 );
and \U$11511 ( \11888 , \11849 , \11886 );
or \U$11512 ( \11889 , \11876 , \11887 , \11888 );
xor \U$11513 ( \11890 , \11092 , \11144 );
xor \U$11514 ( \11891 , \11890 , \11197 );
xor \U$11515 ( \11892 , \11556 , \11566 );
xor \U$11516 ( \11893 , \11892 , \11569 );
and \U$11517 ( \11894 , \11891 , \11893 );
xor \U$11518 ( \11895 , \11575 , \11577 );
xor \U$11519 ( \11896 , \11895 , \11580 );
and \U$11520 ( \11897 , \11893 , \11896 );
and \U$11521 ( \11898 , \11891 , \11896 );
or \U$11522 ( \11899 , \11894 , \11897 , \11898 );
and \U$11523 ( \11900 , \11889 , \11899 );
xor \U$11524 ( \11901 , \11231 , \11240 );
xor \U$11525 ( \11902 , \11901 , \11243 );
and \U$11526 ( \11903 , \11899 , \11902 );
and \U$11527 ( \11904 , \11889 , \11902 );
or \U$11528 ( \11905 , \11900 , \11903 , \11904 );
xor \U$11529 ( \11906 , \11040 , \11200 );
xor \U$11530 ( \11907 , \11906 , \11218 );
xor \U$11531 ( \11908 , \11546 , \11572 );
xor \U$11532 ( \11909 , \11908 , \11583 );
and \U$11533 ( \11910 , \11907 , \11909 );
xor \U$11534 ( \11911 , \11588 , \11590 );
xor \U$11535 ( \11912 , \11911 , \11593 );
and \U$11536 ( \11913 , \11909 , \11912 );
and \U$11537 ( \11914 , \11907 , \11912 );
or \U$11538 ( \11915 , \11910 , \11913 , \11914 );
and \U$11539 ( \11916 , \11905 , \11915 );
xor \U$11540 ( \11917 , \11262 , \11264 );
xor \U$11541 ( \11918 , \11917 , \11267 );
and \U$11542 ( \11919 , \11915 , \11918 );
and \U$11543 ( \11920 , \11905 , \11918 );
or \U$11544 ( \11921 , \11916 , \11919 , \11920 );
xor \U$11545 ( \11922 , \11221 , \11246 );
xor \U$11546 ( \11923 , \11922 , \11257 );
xor \U$11547 ( \11924 , \11586 , \11596 );
xor \U$11548 ( \11925 , \11924 , \11599 );
and \U$11549 ( \11926 , \11923 , \11925 );
and \U$11550 ( \11927 , \11921 , \11926 );
xor \U$11551 ( \11928 , \11602 , \11604 );
xor \U$11552 ( \11929 , \11928 , \11606 );
and \U$11553 ( \11930 , \11926 , \11929 );
and \U$11554 ( \11931 , \11921 , \11929 );
or \U$11555 ( \11932 , \11927 , \11930 , \11931 );
and \U$11556 ( \11933 , \11620 , \11932 );
xor \U$11557 ( \11934 , \11620 , \11932 );
xor \U$11558 ( \11935 , \11921 , \11926 );
xor \U$11559 ( \11936 , \11935 , \11929 );
and \U$11560 ( \11937 , \7067 , \1222 );
and \U$11561 ( \11938 , \6764 , \1220 );
nor \U$11562 ( \11939 , \11937 , \11938 );
xnor \U$11563 ( \11940 , \11939 , \1144 );
and \U$11564 ( \11941 , \7765 , \1058 );
and \U$11565 ( \11942 , \7239 , \1056 );
nor \U$11566 ( \11943 , \11941 , \11942 );
xnor \U$11567 ( \11944 , \11943 , \964 );
and \U$11568 ( \11945 , \11940 , \11944 );
and \U$11569 ( \11946 , \8435 , \888 );
and \U$11570 ( \11947 , \8189 , \886 );
nor \U$11571 ( \11948 , \11946 , \11947 );
xnor \U$11572 ( \11949 , \11948 , \816 );
and \U$11573 ( \11950 , \11944 , \11949 );
and \U$11574 ( \11951 , \11940 , \11949 );
or \U$11575 ( \11952 , \11945 , \11950 , \11951 );
and \U$11576 ( \11953 , \4334 , \2658 );
and \U$11577 ( \11954 , \4078 , \2656 );
nor \U$11578 ( \11955 , \11953 , \11954 );
xnor \U$11579 ( \11956 , \11955 , \2516 );
and \U$11580 ( \11957 , \4833 , \2362 );
and \U$11581 ( \11958 , \4531 , \2360 );
nor \U$11582 ( \11959 , \11957 , \11958 );
xnor \U$11583 ( \11960 , \11959 , \2225 );
and \U$11584 ( \11961 , \11956 , \11960 );
and \U$11585 ( \11962 , \5310 , \2156 );
and \U$11586 ( \11963 , \4841 , \2154 );
nor \U$11587 ( \11964 , \11962 , \11963 );
xnor \U$11588 ( \11965 , \11964 , \2004 );
and \U$11589 ( \11966 , \11960 , \11965 );
and \U$11590 ( \11967 , \11956 , \11965 );
or \U$11591 ( \11968 , \11961 , \11966 , \11967 );
and \U$11592 ( \11969 , \11952 , \11968 );
and \U$11593 ( \11970 , \5579 , \1888 );
and \U$11594 ( \11971 , \5315 , \1886 );
nor \U$11595 ( \11972 , \11970 , \11971 );
xnor \U$11596 ( \11973 , \11972 , \1732 );
and \U$11597 ( \11974 , \6210 , \1616 );
and \U$11598 ( \11975 , \5838 , \1614 );
nor \U$11599 ( \11976 , \11974 , \11975 );
xnor \U$11600 ( \11977 , \11976 , \1503 );
and \U$11601 ( \11978 , \11973 , \11977 );
and \U$11602 ( \11979 , \6562 , \1422 );
and \U$11603 ( \11980 , \6219 , \1420 );
nor \U$11604 ( \11981 , \11979 , \11980 );
xnor \U$11605 ( \11982 , \11981 , \1286 );
and \U$11606 ( \11983 , \11977 , \11982 );
and \U$11607 ( \11984 , \11973 , \11982 );
or \U$11608 ( \11985 , \11978 , \11983 , \11984 );
and \U$11609 ( \11986 , \11968 , \11985 );
and \U$11610 ( \11987 , \11952 , \11985 );
or \U$11611 ( \11988 , \11969 , \11986 , \11987 );
and \U$11612 ( \11989 , \987 , \7829 );
and \U$11613 ( \11990 , \925 , \7827 );
nor \U$11614 ( \11991 , \11989 , \11990 );
xnor \U$11615 ( \11992 , \11991 , \7580 );
and \U$11616 ( \11993 , \1248 , \7300 );
and \U$11617 ( \11994 , \1050 , \7298 );
nor \U$11618 ( \11995 , \11993 , \11994 );
xnor \U$11619 ( \11996 , \11995 , \7040 );
and \U$11620 ( \11997 , \11992 , \11996 );
and \U$11621 ( \11998 , \1441 , \6806 );
and \U$11622 ( \11999 , \1336 , \6804 );
nor \U$11623 ( \12000 , \11998 , \11999 );
xnor \U$11624 ( \12001 , \12000 , \6491 );
and \U$11625 ( \12002 , \11996 , \12001 );
and \U$11626 ( \12003 , \11992 , \12001 );
or \U$11627 ( \12004 , \11997 , \12002 , \12003 );
and \U$11628 ( \12005 , \615 , \9495 );
and \U$11629 ( \12006 , \561 , \9493 );
nor \U$11630 ( \12007 , \12005 , \12006 );
xnor \U$11631 ( \12008 , \12007 , \9185 );
and \U$11632 ( \12009 , \743 , \8958 );
and \U$11633 ( \12010 , \666 , \8956 );
nor \U$11634 ( \12011 , \12009 , \12010 );
xnor \U$11635 ( \12012 , \12011 , \8587 );
and \U$11636 ( \12013 , \12008 , \12012 );
and \U$11637 ( \12014 , \851 , \8396 );
and \U$11638 ( \12015 , \771 , \8394 );
nor \U$11639 ( \12016 , \12014 , \12015 );
xnor \U$11640 ( \12017 , \12016 , \8078 );
and \U$11641 ( \12018 , \12012 , \12017 );
and \U$11642 ( \12019 , \12008 , \12017 );
or \U$11643 ( \12020 , \12013 , \12018 , \12019 );
and \U$11644 ( \12021 , \12004 , \12020 );
and \U$11645 ( \12022 , \479 , \10876 );
and \U$11646 ( \12023 , \431 , \10873 );
nor \U$11647 ( \12024 , \12022 , \12023 );
xnor \U$11648 ( \12025 , \12024 , \9821 );
and \U$11649 ( \12026 , \556 , \10063 );
and \U$11650 ( \12027 , \487 , \10061 );
nor \U$11651 ( \12028 , \12026 , \12027 );
xnor \U$11652 ( \12029 , \12028 , \9824 );
and \U$11653 ( \12030 , \12025 , \12029 );
and \U$11654 ( \12031 , \12029 , \403 );
and \U$11655 ( \12032 , \12025 , \403 );
or \U$11656 ( \12033 , \12030 , \12031 , \12032 );
and \U$11657 ( \12034 , \12020 , \12033 );
and \U$11658 ( \12035 , \12004 , \12033 );
or \U$11659 ( \12036 , \12021 , \12034 , \12035 );
and \U$11660 ( \12037 , \11988 , \12036 );
and \U$11661 ( \12038 , \1562 , \6297 );
and \U$11662 ( \12039 , \1446 , \6295 );
nor \U$11663 ( \12040 , \12038 , \12039 );
xnor \U$11664 ( \12041 , \12040 , \5957 );
and \U$11665 ( \12042 , \1853 , \5708 );
and \U$11666 ( \12043 , \1677 , \5706 );
nor \U$11667 ( \12044 , \12042 , \12043 );
xnor \U$11668 ( \12045 , \12044 , \5467 );
and \U$11669 ( \12046 , \12041 , \12045 );
and \U$11670 ( \12047 , \2104 , \5242 );
and \U$11671 ( \12048 , \1861 , \5240 );
nor \U$11672 ( \12049 , \12047 , \12048 );
xnor \U$11673 ( \12050 , \12049 , \5054 );
and \U$11674 ( \12051 , \12045 , \12050 );
and \U$11675 ( \12052 , \12041 , \12050 );
or \U$11676 ( \12053 , \12046 , \12051 , \12052 );
and \U$11677 ( \12054 , \2295 , \4868 );
and \U$11678 ( \12055 , \2109 , \4866 );
nor \U$11679 ( \12056 , \12054 , \12055 );
xnor \U$11680 ( \12057 , \12056 , \4636 );
and \U$11681 ( \12058 , \2703 , \4417 );
and \U$11682 ( \12059 , \2439 , \4415 );
nor \U$11683 ( \12060 , \12058 , \12059 );
xnor \U$11684 ( \12061 , \12060 , \4274 );
and \U$11685 ( \12062 , \12057 , \12061 );
and \U$11686 ( \12063 , \2902 , \4094 );
and \U$11687 ( \12064 , \2728 , \4092 );
nor \U$11688 ( \12065 , \12063 , \12064 );
xnor \U$11689 ( \12066 , \12065 , \3848 );
and \U$11690 ( \12067 , \12061 , \12066 );
and \U$11691 ( \12068 , \12057 , \12066 );
or \U$11692 ( \12069 , \12062 , \12067 , \12068 );
and \U$11693 ( \12070 , \12053 , \12069 );
and \U$11694 ( \12071 , \3207 , \3699 );
and \U$11695 ( \12072 , \3069 , \3697 );
nor \U$11696 ( \12073 , \12071 , \12072 );
xnor \U$11697 ( \12074 , \12073 , \3512 );
and \U$11698 ( \12075 , \3743 , \3386 );
and \U$11699 ( \12076 , \3326 , \3384 );
nor \U$11700 ( \12077 , \12075 , \12076 );
xnor \U$11701 ( \12078 , \12077 , \3181 );
and \U$11702 ( \12079 , \12074 , \12078 );
and \U$11703 ( \12080 , \4073 , \2980 );
and \U$11704 ( \12081 , \3951 , \2978 );
nor \U$11705 ( \12082 , \12080 , \12081 );
xnor \U$11706 ( \12083 , \12082 , \2831 );
and \U$11707 ( \12084 , \12078 , \12083 );
and \U$11708 ( \12085 , \12074 , \12083 );
or \U$11709 ( \12086 , \12079 , \12084 , \12085 );
and \U$11710 ( \12087 , \12069 , \12086 );
and \U$11711 ( \12088 , \12053 , \12086 );
or \U$11712 ( \12089 , \12070 , \12087 , \12088 );
and \U$11713 ( \12090 , \12036 , \12089 );
and \U$11714 ( \12091 , \11988 , \12089 );
or \U$11715 ( \12092 , \12037 , \12090 , \12091 );
and \U$11716 ( \12093 , \8759 , \754 );
and \U$11717 ( \12094 , \8440 , \752 );
nor \U$11718 ( \12095 , \12093 , \12094 );
xnor \U$11719 ( \12096 , \12095 , \711 );
and \U$11720 ( \12097 , \9612 , \641 );
and \U$11721 ( \12098 , \9043 , \639 );
nor \U$11722 ( \12099 , \12097 , \12098 );
xnor \U$11723 ( \12100 , \12099 , \592 );
and \U$11724 ( \12101 , \12096 , \12100 );
and \U$11725 ( \12102 , \10223 , \540 );
and \U$11726 ( \12103 , \9620 , \538 );
nor \U$11727 ( \12104 , \12102 , \12103 );
xnor \U$11728 ( \12105 , \12104 , \499 );
and \U$11729 ( \12106 , \12100 , \12105 );
and \U$11730 ( \12107 , \12096 , \12105 );
or \U$11731 ( \12108 , \12101 , \12106 , \12107 );
and \U$11732 ( \12109 , \10409 , \470 );
and \U$11733 ( \12110 , \10228 , \468 );
nor \U$11734 ( \12111 , \12109 , \12110 );
xnor \U$11735 ( \12112 , \12111 , \440 );
nand \U$11736 ( \12113 , \11029 , \420 );
xnor \U$11737 ( \12114 , \12113 , \403 );
and \U$11738 ( \12115 , \12112 , \12114 );
and \U$11739 ( \12116 , \12108 , \12115 );
and \U$11740 ( \12117 , \11029 , \422 );
and \U$11741 ( \12118 , \10409 , \420 );
nor \U$11742 ( \12119 , \12117 , \12118 );
xnor \U$11743 ( \12120 , \12119 , \403 );
and \U$11744 ( \12121 , \12115 , \12120 );
and \U$11745 ( \12122 , \12108 , \12120 );
or \U$11746 ( \12123 , \12116 , \12121 , \12122 );
xor \U$11747 ( \12124 , \11709 , \11713 );
xor \U$11748 ( \12125 , \12124 , \11718 );
xor \U$11749 ( \12126 , \11745 , \11749 );
xor \U$11750 ( \12127 , \12126 , \11754 );
and \U$11751 ( \12128 , \12125 , \12127 );
xor \U$11752 ( \12129 , \11762 , \11766 );
xor \U$11753 ( \12130 , \12129 , \11771 );
and \U$11754 ( \12131 , \12127 , \12130 );
and \U$11755 ( \12132 , \12125 , \12130 );
or \U$11756 ( \12133 , \12128 , \12131 , \12132 );
and \U$11757 ( \12134 , \12123 , \12133 );
xor \U$11758 ( \12135 , \11676 , \11680 );
xor \U$11759 ( \12136 , \12135 , \11685 );
xor \U$11760 ( \12137 , \11692 , \11696 );
xor \U$11761 ( \12138 , \12137 , \11701 );
and \U$11762 ( \12139 , \12136 , \12138 );
xor \U$11763 ( \12140 , \11794 , \11798 );
xor \U$11764 ( \12141 , \12140 , \11803 );
and \U$11765 ( \12142 , \12138 , \12141 );
and \U$11766 ( \12143 , \12136 , \12141 );
or \U$11767 ( \12144 , \12139 , \12142 , \12143 );
and \U$11768 ( \12145 , \12133 , \12144 );
and \U$11769 ( \12146 , \12123 , \12144 );
or \U$11770 ( \12147 , \12134 , \12145 , \12146 );
and \U$11771 ( \12148 , \12092 , \12147 );
xor \U$11772 ( \12149 , \11624 , \11628 );
xor \U$11773 ( \12150 , \12149 , \11633 );
xor \U$11774 ( \12151 , \11729 , \11733 );
xor \U$11775 ( \12152 , \12151 , \11738 );
and \U$11776 ( \12153 , \12150 , \12152 );
xor \U$11777 ( \12154 , \11657 , \11661 );
xor \U$11778 ( \12155 , \12154 , \11666 );
and \U$11779 ( \12156 , \12152 , \12155 );
and \U$11780 ( \12157 , \12150 , \12155 );
or \U$11781 ( \12158 , \12153 , \12156 , \12157 );
xor \U$11782 ( \12159 , \11831 , \11833 );
xor \U$11783 ( \12160 , \12159 , \11836 );
and \U$11784 ( \12161 , \12158 , \12160 );
xor \U$11785 ( \12162 , \11782 , \11784 );
xor \U$11786 ( \12163 , \12162 , \11787 );
and \U$11787 ( \12164 , \12160 , \12163 );
and \U$11788 ( \12165 , \12158 , \12163 );
or \U$11789 ( \12166 , \12161 , \12164 , \12165 );
and \U$11790 ( \12167 , \12147 , \12166 );
and \U$11791 ( \12168 , \12092 , \12166 );
or \U$11792 ( \12169 , \12148 , \12167 , \12168 );
xor \U$11793 ( \12170 , \11688 , \11704 );
xor \U$11794 ( \12171 , \12170 , \11721 );
xor \U$11795 ( \12172 , \11806 , \11808 );
xor \U$11796 ( \12173 , \12172 , \11811 );
and \U$11797 ( \12174 , \12171 , \12173 );
xor \U$11798 ( \12175 , \11817 , \11819 );
xor \U$11799 ( \12176 , \12175 , \11822 );
and \U$11800 ( \12177 , \12173 , \12176 );
and \U$11801 ( \12178 , \12171 , \12176 );
or \U$11802 ( \12179 , \12174 , \12177 , \12178 );
xor \U$11803 ( \12180 , \11851 , \11853 );
xor \U$11804 ( \12181 , \12180 , \11856 );
and \U$11805 ( \12182 , \12179 , \12181 );
xor \U$11806 ( \12183 , \11861 , \11863 );
xor \U$11807 ( \12184 , \12183 , \11866 );
and \U$11808 ( \12185 , \12181 , \12184 );
and \U$11809 ( \12186 , \12179 , \12184 );
or \U$11810 ( \12187 , \12182 , \12185 , \12186 );
and \U$11811 ( \12188 , \12169 , \12187 );
xor \U$11812 ( \12189 , \11672 , \11724 );
xor \U$11813 ( \12190 , \12189 , \11777 );
xor \U$11814 ( \12191 , \11790 , \11814 );
xor \U$11815 ( \12192 , \12191 , \11825 );
and \U$11816 ( \12193 , \12190 , \12192 );
xor \U$11817 ( \12194 , \11839 , \11841 );
xor \U$11818 ( \12195 , \12194 , \11843 );
and \U$11819 ( \12196 , \12192 , \12195 );
and \U$11820 ( \12197 , \12190 , \12195 );
or \U$11821 ( \12198 , \12193 , \12196 , \12197 );
and \U$11822 ( \12199 , \12187 , \12198 );
and \U$11823 ( \12200 , \12169 , \12198 );
or \U$11824 ( \12201 , \12188 , \12199 , \12200 );
xor \U$11825 ( \12202 , \11340 , \11352 );
xor \U$11826 ( \12203 , \12202 , \11363 );
xor \U$11827 ( \12204 , \11418 , \11466 );
xor \U$11828 ( \12205 , \12204 , \11519 );
and \U$11829 ( \12206 , \12203 , \12205 );
xor \U$11830 ( \12207 , \11878 , \11880 );
xor \U$11831 ( \12208 , \12207 , \11883 );
and \U$11832 ( \12209 , \12205 , \12208 );
and \U$11833 ( \12210 , \12203 , \12208 );
or \U$11834 ( \12211 , \12206 , \12209 , \12210 );
and \U$11835 ( \12212 , \12201 , \12211 );
xor \U$11836 ( \12213 , \11366 , \11522 );
xor \U$11837 ( \12214 , \12213 , \11543 );
and \U$11838 ( \12215 , \12211 , \12214 );
and \U$11839 ( \12216 , \12201 , \12214 );
or \U$11840 ( \12217 , \12212 , \12215 , \12216 );
xor \U$11841 ( \12218 , \11889 , \11899 );
xor \U$11842 ( \12219 , \12218 , \11902 );
and \U$11843 ( \12220 , \12217 , \12219 );
xor \U$11844 ( \12221 , \11907 , \11909 );
xor \U$11845 ( \12222 , \12221 , \11912 );
and \U$11846 ( \12223 , \12219 , \12222 );
and \U$11847 ( \12224 , \12217 , \12222 );
or \U$11848 ( \12225 , \12220 , \12223 , \12224 );
xor \U$11849 ( \12226 , \11905 , \11915 );
xor \U$11850 ( \12227 , \12226 , \11918 );
and \U$11851 ( \12228 , \12225 , \12227 );
xor \U$11852 ( \12229 , \11923 , \11925 );
and \U$11853 ( \12230 , \12227 , \12229 );
and \U$11854 ( \12231 , \12225 , \12229 );
or \U$11855 ( \12232 , \12228 , \12230 , \12231 );
and \U$11856 ( \12233 , \11936 , \12232 );
xor \U$11857 ( \12234 , \11936 , \12232 );
xor \U$11858 ( \12235 , \12225 , \12227 );
xor \U$11859 ( \12236 , \12235 , \12229 );
xor \U$11860 ( \12237 , \11940 , \11944 );
xor \U$11861 ( \12238 , \12237 , \11949 );
xor \U$11862 ( \12239 , \11956 , \11960 );
xor \U$11863 ( \12240 , \12239 , \11965 );
and \U$11864 ( \12241 , \12238 , \12240 );
xor \U$11865 ( \12242 , \11973 , \11977 );
xor \U$11866 ( \12243 , \12242 , \11982 );
and \U$11867 ( \12244 , \12240 , \12243 );
and \U$11868 ( \12245 , \12238 , \12243 );
or \U$11869 ( \12246 , \12241 , \12244 , \12245 );
xor \U$11870 ( \12247 , \12041 , \12045 );
xor \U$11871 ( \12248 , \12247 , \12050 );
xor \U$11872 ( \12249 , \12057 , \12061 );
xor \U$11873 ( \12250 , \12249 , \12066 );
and \U$11874 ( \12251 , \12248 , \12250 );
xor \U$11875 ( \12252 , \12074 , \12078 );
xor \U$11876 ( \12253 , \12252 , \12083 );
and \U$11877 ( \12254 , \12250 , \12253 );
and \U$11878 ( \12255 , \12248 , \12253 );
or \U$11879 ( \12256 , \12251 , \12254 , \12255 );
and \U$11880 ( \12257 , \12246 , \12256 );
and \U$11881 ( \12258 , \9620 , \641 );
and \U$11882 ( \12259 , \9612 , \639 );
nor \U$11883 ( \12260 , \12258 , \12259 );
xnor \U$11884 ( \12261 , \12260 , \592 );
and \U$11885 ( \12262 , \10228 , \540 );
and \U$11886 ( \12263 , \10223 , \538 );
nor \U$11887 ( \12264 , \12262 , \12263 );
xnor \U$11888 ( \12265 , \12264 , \499 );
and \U$11889 ( \12266 , \12261 , \12265 );
and \U$11890 ( \12267 , \11029 , \470 );
and \U$11891 ( \12268 , \10409 , \468 );
nor \U$11892 ( \12269 , \12267 , \12268 );
xnor \U$11893 ( \12270 , \12269 , \440 );
and \U$11894 ( \12271 , \12265 , \12270 );
and \U$11895 ( \12272 , \12261 , \12270 );
or \U$11896 ( \12273 , \12266 , \12271 , \12272 );
xor \U$11897 ( \12274 , \12096 , \12100 );
xor \U$11898 ( \12275 , \12274 , \12105 );
and \U$11899 ( \12276 , \12273 , \12275 );
xor \U$11900 ( \12277 , \12112 , \12114 );
and \U$11901 ( \12278 , \12275 , \12277 );
and \U$11902 ( \12279 , \12273 , \12277 );
or \U$11903 ( \12280 , \12276 , \12278 , \12279 );
and \U$11904 ( \12281 , \12256 , \12280 );
and \U$11905 ( \12282 , \12246 , \12280 );
or \U$11906 ( \12283 , \12257 , \12281 , \12282 );
and \U$11907 ( \12284 , \3951 , \3386 );
and \U$11908 ( \12285 , \3743 , \3384 );
nor \U$11909 ( \12286 , \12284 , \12285 );
xnor \U$11910 ( \12287 , \12286 , \3181 );
and \U$11911 ( \12288 , \4078 , \2980 );
and \U$11912 ( \12289 , \4073 , \2978 );
nor \U$11913 ( \12290 , \12288 , \12289 );
xnor \U$11914 ( \12291 , \12290 , \2831 );
and \U$11915 ( \12292 , \12287 , \12291 );
and \U$11916 ( \12293 , \4531 , \2658 );
and \U$11917 ( \12294 , \4334 , \2656 );
nor \U$11918 ( \12295 , \12293 , \12294 );
xnor \U$11919 ( \12296 , \12295 , \2516 );
and \U$11920 ( \12297 , \12291 , \12296 );
and \U$11921 ( \12298 , \12287 , \12296 );
or \U$11922 ( \12299 , \12292 , \12297 , \12298 );
and \U$11923 ( \12300 , \1861 , \5708 );
and \U$11924 ( \12301 , \1853 , \5706 );
nor \U$11925 ( \12302 , \12300 , \12301 );
xnor \U$11926 ( \12303 , \12302 , \5467 );
and \U$11927 ( \12304 , \2109 , \5242 );
and \U$11928 ( \12305 , \2104 , \5240 );
nor \U$11929 ( \12306 , \12304 , \12305 );
xnor \U$11930 ( \12307 , \12306 , \5054 );
and \U$11931 ( \12308 , \12303 , \12307 );
and \U$11932 ( \12309 , \2439 , \4868 );
and \U$11933 ( \12310 , \2295 , \4866 );
nor \U$11934 ( \12311 , \12309 , \12310 );
xnor \U$11935 ( \12312 , \12311 , \4636 );
and \U$11936 ( \12313 , \12307 , \12312 );
and \U$11937 ( \12314 , \12303 , \12312 );
or \U$11938 ( \12315 , \12308 , \12313 , \12314 );
and \U$11939 ( \12316 , \12299 , \12315 );
and \U$11940 ( \12317 , \2728 , \4417 );
and \U$11941 ( \12318 , \2703 , \4415 );
nor \U$11942 ( \12319 , \12317 , \12318 );
xnor \U$11943 ( \12320 , \12319 , \4274 );
and \U$11944 ( \12321 , \3069 , \4094 );
and \U$11945 ( \12322 , \2902 , \4092 );
nor \U$11946 ( \12323 , \12321 , \12322 );
xnor \U$11947 ( \12324 , \12323 , \3848 );
and \U$11948 ( \12325 , \12320 , \12324 );
and \U$11949 ( \12326 , \3326 , \3699 );
and \U$11950 ( \12327 , \3207 , \3697 );
nor \U$11951 ( \12328 , \12326 , \12327 );
xnor \U$11952 ( \12329 , \12328 , \3512 );
and \U$11953 ( \12330 , \12324 , \12329 );
and \U$11954 ( \12331 , \12320 , \12329 );
or \U$11955 ( \12332 , \12325 , \12330 , \12331 );
and \U$11956 ( \12333 , \12315 , \12332 );
and \U$11957 ( \12334 , \12299 , \12332 );
or \U$11958 ( \12335 , \12316 , \12333 , \12334 );
and \U$11959 ( \12336 , \1336 , \7300 );
and \U$11960 ( \12337 , \1248 , \7298 );
nor \U$11961 ( \12338 , \12336 , \12337 );
xnor \U$11962 ( \12339 , \12338 , \7040 );
and \U$11963 ( \12340 , \1446 , \6806 );
and \U$11964 ( \12341 , \1441 , \6804 );
nor \U$11965 ( \12342 , \12340 , \12341 );
xnor \U$11966 ( \12343 , \12342 , \6491 );
and \U$11967 ( \12344 , \12339 , \12343 );
and \U$11968 ( \12345 , \1677 , \6297 );
and \U$11969 ( \12346 , \1562 , \6295 );
nor \U$11970 ( \12347 , \12345 , \12346 );
xnor \U$11971 ( \12348 , \12347 , \5957 );
and \U$11972 ( \12349 , \12343 , \12348 );
and \U$11973 ( \12350 , \12339 , \12348 );
or \U$11974 ( \12351 , \12344 , \12349 , \12350 );
and \U$11975 ( \12352 , \487 , \10876 );
and \U$11976 ( \12353 , \479 , \10873 );
nor \U$11977 ( \12354 , \12352 , \12353 );
xnor \U$11978 ( \12355 , \12354 , \9821 );
and \U$11979 ( \12356 , \561 , \10063 );
and \U$11980 ( \12357 , \556 , \10061 );
nor \U$11981 ( \12358 , \12356 , \12357 );
xnor \U$11982 ( \12359 , \12358 , \9824 );
and \U$11983 ( \12360 , \12355 , \12359 );
and \U$11984 ( \12361 , \666 , \9495 );
and \U$11985 ( \12362 , \615 , \9493 );
nor \U$11986 ( \12363 , \12361 , \12362 );
xnor \U$11987 ( \12364 , \12363 , \9185 );
and \U$11988 ( \12365 , \12359 , \12364 );
and \U$11989 ( \12366 , \12355 , \12364 );
or \U$11990 ( \12367 , \12360 , \12365 , \12366 );
and \U$11991 ( \12368 , \12351 , \12367 );
and \U$11992 ( \12369 , \771 , \8958 );
and \U$11993 ( \12370 , \743 , \8956 );
nor \U$11994 ( \12371 , \12369 , \12370 );
xnor \U$11995 ( \12372 , \12371 , \8587 );
and \U$11996 ( \12373 , \925 , \8396 );
and \U$11997 ( \12374 , \851 , \8394 );
nor \U$11998 ( \12375 , \12373 , \12374 );
xnor \U$11999 ( \12376 , \12375 , \8078 );
and \U$12000 ( \12377 , \12372 , \12376 );
and \U$12001 ( \12378 , \1050 , \7829 );
and \U$12002 ( \12379 , \987 , \7827 );
nor \U$12003 ( \12380 , \12378 , \12379 );
xnor \U$12004 ( \12381 , \12380 , \7580 );
and \U$12005 ( \12382 , \12376 , \12381 );
and \U$12006 ( \12383 , \12372 , \12381 );
or \U$12007 ( \12384 , \12377 , \12382 , \12383 );
and \U$12008 ( \12385 , \12367 , \12384 );
and \U$12009 ( \12386 , \12351 , \12384 );
or \U$12010 ( \12387 , \12368 , \12385 , \12386 );
and \U$12011 ( \12388 , \12335 , \12387 );
and \U$12012 ( \12389 , \4841 , \2362 );
and \U$12013 ( \12390 , \4833 , \2360 );
nor \U$12014 ( \12391 , \12389 , \12390 );
xnor \U$12015 ( \12392 , \12391 , \2225 );
and \U$12016 ( \12393 , \5315 , \2156 );
and \U$12017 ( \12394 , \5310 , \2154 );
nor \U$12018 ( \12395 , \12393 , \12394 );
xnor \U$12019 ( \12396 , \12395 , \2004 );
and \U$12020 ( \12397 , \12392 , \12396 );
and \U$12021 ( \12398 , \5838 , \1888 );
and \U$12022 ( \12399 , \5579 , \1886 );
nor \U$12023 ( \12400 , \12398 , \12399 );
xnor \U$12024 ( \12401 , \12400 , \1732 );
and \U$12025 ( \12402 , \12396 , \12401 );
and \U$12026 ( \12403 , \12392 , \12401 );
or \U$12027 ( \12404 , \12397 , \12402 , \12403 );
and \U$12028 ( \12405 , \8189 , \1058 );
and \U$12029 ( \12406 , \7765 , \1056 );
nor \U$12030 ( \12407 , \12405 , \12406 );
xnor \U$12031 ( \12408 , \12407 , \964 );
and \U$12032 ( \12409 , \8440 , \888 );
and \U$12033 ( \12410 , \8435 , \886 );
nor \U$12034 ( \12411 , \12409 , \12410 );
xnor \U$12035 ( \12412 , \12411 , \816 );
and \U$12036 ( \12413 , \12408 , \12412 );
and \U$12037 ( \12414 , \9043 , \754 );
and \U$12038 ( \12415 , \8759 , \752 );
nor \U$12039 ( \12416 , \12414 , \12415 );
xnor \U$12040 ( \12417 , \12416 , \711 );
and \U$12041 ( \12418 , \12412 , \12417 );
and \U$12042 ( \12419 , \12408 , \12417 );
or \U$12043 ( \12420 , \12413 , \12418 , \12419 );
and \U$12044 ( \12421 , \12404 , \12420 );
and \U$12045 ( \12422 , \6219 , \1616 );
and \U$12046 ( \12423 , \6210 , \1614 );
nor \U$12047 ( \12424 , \12422 , \12423 );
xnor \U$12048 ( \12425 , \12424 , \1503 );
and \U$12049 ( \12426 , \6764 , \1422 );
and \U$12050 ( \12427 , \6562 , \1420 );
nor \U$12051 ( \12428 , \12426 , \12427 );
xnor \U$12052 ( \12429 , \12428 , \1286 );
and \U$12053 ( \12430 , \12425 , \12429 );
and \U$12054 ( \12431 , \7239 , \1222 );
and \U$12055 ( \12432 , \7067 , \1220 );
nor \U$12056 ( \12433 , \12431 , \12432 );
xnor \U$12057 ( \12434 , \12433 , \1144 );
and \U$12058 ( \12435 , \12429 , \12434 );
and \U$12059 ( \12436 , \12425 , \12434 );
or \U$12060 ( \12437 , \12430 , \12435 , \12436 );
and \U$12061 ( \12438 , \12420 , \12437 );
and \U$12062 ( \12439 , \12404 , \12437 );
or \U$12063 ( \12440 , \12421 , \12438 , \12439 );
and \U$12064 ( \12441 , \12387 , \12440 );
and \U$12065 ( \12442 , \12335 , \12440 );
or \U$12066 ( \12443 , \12388 , \12441 , \12442 );
and \U$12067 ( \12444 , \12283 , \12443 );
xor \U$12068 ( \12445 , \11992 , \11996 );
xor \U$12069 ( \12446 , \12445 , \12001 );
xor \U$12070 ( \12447 , \12008 , \12012 );
xor \U$12071 ( \12448 , \12447 , \12017 );
and \U$12072 ( \12449 , \12446 , \12448 );
xor \U$12073 ( \12450 , \12025 , \12029 );
xor \U$12074 ( \12451 , \12450 , \403 );
and \U$12075 ( \12452 , \12448 , \12451 );
and \U$12076 ( \12453 , \12446 , \12451 );
or \U$12077 ( \12454 , \12449 , \12452 , \12453 );
xor \U$12078 ( \12455 , \11640 , \11644 );
xor \U$12079 ( \12456 , \12455 , \11649 );
and \U$12080 ( \12457 , \12454 , \12456 );
xor \U$12081 ( \12458 , \12150 , \12152 );
xor \U$12082 ( \12459 , \12458 , \12155 );
and \U$12083 ( \12460 , \12456 , \12459 );
and \U$12084 ( \12461 , \12454 , \12459 );
or \U$12085 ( \12462 , \12457 , \12460 , \12461 );
and \U$12086 ( \12463 , \12443 , \12462 );
and \U$12087 ( \12464 , \12283 , \12462 );
or \U$12088 ( \12465 , \12444 , \12463 , \12464 );
xor \U$12089 ( \12466 , \11952 , \11968 );
xor \U$12090 ( \12467 , \12466 , \11985 );
xor \U$12091 ( \12468 , \12004 , \12020 );
xor \U$12092 ( \12469 , \12468 , \12033 );
and \U$12093 ( \12470 , \12467 , \12469 );
xor \U$12094 ( \12471 , \12053 , \12069 );
xor \U$12095 ( \12472 , \12471 , \12086 );
and \U$12096 ( \12473 , \12469 , \12472 );
and \U$12097 ( \12474 , \12467 , \12472 );
or \U$12098 ( \12475 , \12470 , \12473 , \12474 );
xor \U$12099 ( \12476 , \12108 , \12115 );
xor \U$12100 ( \12477 , \12476 , \12120 );
xor \U$12101 ( \12478 , \12125 , \12127 );
xor \U$12102 ( \12479 , \12478 , \12130 );
and \U$12103 ( \12480 , \12477 , \12479 );
xor \U$12104 ( \12481 , \12136 , \12138 );
xor \U$12105 ( \12482 , \12481 , \12141 );
and \U$12106 ( \12483 , \12479 , \12482 );
and \U$12107 ( \12484 , \12477 , \12482 );
or \U$12108 ( \12485 , \12480 , \12483 , \12484 );
and \U$12109 ( \12486 , \12475 , \12485 );
xor \U$12110 ( \12487 , \11741 , \11757 );
xor \U$12111 ( \12488 , \12487 , \11774 );
and \U$12112 ( \12489 , \12485 , \12488 );
and \U$12113 ( \12490 , \12475 , \12488 );
or \U$12114 ( \12491 , \12486 , \12489 , \12490 );
and \U$12115 ( \12492 , \12465 , \12491 );
xor \U$12116 ( \12493 , \11636 , \11652 );
xor \U$12117 ( \12494 , \12493 , \11669 );
xor \U$12118 ( \12495 , \12171 , \12173 );
xor \U$12119 ( \12496 , \12495 , \12176 );
and \U$12120 ( \12497 , \12494 , \12496 );
xor \U$12121 ( \12498 , \12158 , \12160 );
xor \U$12122 ( \12499 , \12498 , \12163 );
and \U$12123 ( \12500 , \12496 , \12499 );
and \U$12124 ( \12501 , \12494 , \12499 );
or \U$12125 ( \12502 , \12497 , \12500 , \12501 );
and \U$12126 ( \12503 , \12491 , \12502 );
and \U$12127 ( \12504 , \12465 , \12502 );
or \U$12128 ( \12505 , \12492 , \12503 , \12504 );
xor \U$12129 ( \12506 , \12092 , \12147 );
xor \U$12130 ( \12507 , \12506 , \12166 );
xor \U$12131 ( \12508 , \12179 , \12181 );
xor \U$12132 ( \12509 , \12508 , \12184 );
and \U$12133 ( \12510 , \12507 , \12509 );
xor \U$12134 ( \12511 , \12190 , \12192 );
xor \U$12135 ( \12512 , \12511 , \12195 );
and \U$12136 ( \12513 , \12509 , \12512 );
and \U$12137 ( \12514 , \12507 , \12512 );
or \U$12138 ( \12515 , \12510 , \12513 , \12514 );
and \U$12139 ( \12516 , \12505 , \12515 );
xor \U$12140 ( \12517 , \11859 , \11869 );
xor \U$12141 ( \12518 , \12517 , \11872 );
and \U$12142 ( \12519 , \12515 , \12518 );
and \U$12143 ( \12520 , \12505 , \12518 );
or \U$12144 ( \12521 , \12516 , \12519 , \12520 );
xor \U$12145 ( \12522 , \11780 , \11828 );
xor \U$12146 ( \12523 , \12522 , \11846 );
xor \U$12147 ( \12524 , \12169 , \12187 );
xor \U$12148 ( \12525 , \12524 , \12198 );
and \U$12149 ( \12526 , \12523 , \12525 );
xor \U$12150 ( \12527 , \12203 , \12205 );
xor \U$12151 ( \12528 , \12527 , \12208 );
and \U$12152 ( \12529 , \12525 , \12528 );
and \U$12153 ( \12530 , \12523 , \12528 );
or \U$12154 ( \12531 , \12526 , \12529 , \12530 );
and \U$12155 ( \12532 , \12521 , \12531 );
xor \U$12156 ( \12533 , \11891 , \11893 );
xor \U$12157 ( \12534 , \12533 , \11896 );
and \U$12158 ( \12535 , \12531 , \12534 );
and \U$12159 ( \12536 , \12521 , \12534 );
or \U$12160 ( \12537 , \12532 , \12535 , \12536 );
xor \U$12161 ( \12538 , \11849 , \11875 );
xor \U$12162 ( \12539 , \12538 , \11886 );
xor \U$12163 ( \12540 , \12201 , \12211 );
xor \U$12164 ( \12541 , \12540 , \12214 );
and \U$12165 ( \12542 , \12539 , \12541 );
and \U$12166 ( \12543 , \12537 , \12542 );
xor \U$12167 ( \12544 , \12217 , \12219 );
xor \U$12168 ( \12545 , \12544 , \12222 );
and \U$12169 ( \12546 , \12542 , \12545 );
and \U$12170 ( \12547 , \12537 , \12545 );
or \U$12171 ( \12548 , \12543 , \12546 , \12547 );
and \U$12172 ( \12549 , \12236 , \12548 );
xor \U$12173 ( \12550 , \12236 , \12548 );
xor \U$12174 ( \12551 , \12537 , \12542 );
xor \U$12175 ( \12552 , \12551 , \12545 );
xor \U$12176 ( \12553 , \12287 , \12291 );
xor \U$12177 ( \12554 , \12553 , \12296 );
xor \U$12178 ( \12555 , \12392 , \12396 );
xor \U$12179 ( \12556 , \12555 , \12401 );
and \U$12180 ( \12557 , \12554 , \12556 );
xor \U$12181 ( \12558 , \12425 , \12429 );
xor \U$12182 ( \12559 , \12558 , \12434 );
and \U$12183 ( \12560 , \12556 , \12559 );
and \U$12184 ( \12561 , \12554 , \12559 );
or \U$12185 ( \12562 , \12557 , \12560 , \12561 );
and \U$12186 ( \12563 , \9612 , \754 );
and \U$12187 ( \12564 , \9043 , \752 );
nor \U$12188 ( \12565 , \12563 , \12564 );
xnor \U$12189 ( \12566 , \12565 , \711 );
and \U$12190 ( \12567 , \10223 , \641 );
and \U$12191 ( \12568 , \9620 , \639 );
nor \U$12192 ( \12569 , \12567 , \12568 );
xnor \U$12193 ( \12570 , \12569 , \592 );
and \U$12194 ( \12571 , \12566 , \12570 );
and \U$12195 ( \12572 , \10409 , \540 );
and \U$12196 ( \12573 , \10228 , \538 );
nor \U$12197 ( \12574 , \12572 , \12573 );
xnor \U$12198 ( \12575 , \12574 , \499 );
and \U$12199 ( \12576 , \12570 , \12575 );
and \U$12200 ( \12577 , \12566 , \12575 );
or \U$12201 ( \12578 , \12571 , \12576 , \12577 );
xor \U$12202 ( \12579 , \12408 , \12412 );
xor \U$12203 ( \12580 , \12579 , \12417 );
and \U$12204 ( \12581 , \12578 , \12580 );
xor \U$12205 ( \12582 , \12261 , \12265 );
xor \U$12206 ( \12583 , \12582 , \12270 );
and \U$12207 ( \12584 , \12580 , \12583 );
and \U$12208 ( \12585 , \12578 , \12583 );
or \U$12209 ( \12586 , \12581 , \12584 , \12585 );
and \U$12210 ( \12587 , \12562 , \12586 );
xor \U$12211 ( \12588 , \12339 , \12343 );
xor \U$12212 ( \12589 , \12588 , \12348 );
xor \U$12213 ( \12590 , \12303 , \12307 );
xor \U$12214 ( \12591 , \12590 , \12312 );
and \U$12215 ( \12592 , \12589 , \12591 );
xor \U$12216 ( \12593 , \12320 , \12324 );
xor \U$12217 ( \12594 , \12593 , \12329 );
and \U$12218 ( \12595 , \12591 , \12594 );
and \U$12219 ( \12596 , \12589 , \12594 );
or \U$12220 ( \12597 , \12592 , \12595 , \12596 );
and \U$12221 ( \12598 , \12586 , \12597 );
and \U$12222 ( \12599 , \12562 , \12597 );
or \U$12223 ( \12600 , \12587 , \12598 , \12599 );
and \U$12224 ( \12601 , \1248 , \7829 );
and \U$12225 ( \12602 , \1050 , \7827 );
nor \U$12226 ( \12603 , \12601 , \12602 );
xnor \U$12227 ( \12604 , \12603 , \7580 );
and \U$12228 ( \12605 , \1441 , \7300 );
and \U$12229 ( \12606 , \1336 , \7298 );
nor \U$12230 ( \12607 , \12605 , \12606 );
xnor \U$12231 ( \12608 , \12607 , \7040 );
and \U$12232 ( \12609 , \12604 , \12608 );
and \U$12233 ( \12610 , \1562 , \6806 );
and \U$12234 ( \12611 , \1446 , \6804 );
nor \U$12235 ( \12612 , \12610 , \12611 );
xnor \U$12236 ( \12613 , \12612 , \6491 );
and \U$12237 ( \12614 , \12608 , \12613 );
and \U$12238 ( \12615 , \12604 , \12613 );
or \U$12239 ( \12616 , \12609 , \12614 , \12615 );
and \U$12240 ( \12617 , \556 , \10876 );
and \U$12241 ( \12618 , \487 , \10873 );
nor \U$12242 ( \12619 , \12617 , \12618 );
xnor \U$12243 ( \12620 , \12619 , \9821 );
and \U$12244 ( \12621 , \615 , \10063 );
and \U$12245 ( \12622 , \561 , \10061 );
nor \U$12246 ( \12623 , \12621 , \12622 );
xnor \U$12247 ( \12624 , \12623 , \9824 );
and \U$12248 ( \12625 , \12620 , \12624 );
and \U$12249 ( \12626 , \12624 , \440 );
and \U$12250 ( \12627 , \12620 , \440 );
or \U$12251 ( \12628 , \12625 , \12626 , \12627 );
and \U$12252 ( \12629 , \12616 , \12628 );
and \U$12253 ( \12630 , \743 , \9495 );
and \U$12254 ( \12631 , \666 , \9493 );
nor \U$12255 ( \12632 , \12630 , \12631 );
xnor \U$12256 ( \12633 , \12632 , \9185 );
and \U$12257 ( \12634 , \851 , \8958 );
and \U$12258 ( \12635 , \771 , \8956 );
nor \U$12259 ( \12636 , \12634 , \12635 );
xnor \U$12260 ( \12637 , \12636 , \8587 );
and \U$12261 ( \12638 , \12633 , \12637 );
and \U$12262 ( \12639 , \987 , \8396 );
and \U$12263 ( \12640 , \925 , \8394 );
nor \U$12264 ( \12641 , \12639 , \12640 );
xnor \U$12265 ( \12642 , \12641 , \8078 );
and \U$12266 ( \12643 , \12637 , \12642 );
and \U$12267 ( \12644 , \12633 , \12642 );
or \U$12268 ( \12645 , \12638 , \12643 , \12644 );
and \U$12269 ( \12646 , \12628 , \12645 );
and \U$12270 ( \12647 , \12616 , \12645 );
or \U$12271 ( \12648 , \12629 , \12646 , \12647 );
and \U$12272 ( \12649 , \3743 , \3699 );
and \U$12273 ( \12650 , \3326 , \3697 );
nor \U$12274 ( \12651 , \12649 , \12650 );
xnor \U$12275 ( \12652 , \12651 , \3512 );
and \U$12276 ( \12653 , \4073 , \3386 );
and \U$12277 ( \12654 , \3951 , \3384 );
nor \U$12278 ( \12655 , \12653 , \12654 );
xnor \U$12279 ( \12656 , \12655 , \3181 );
and \U$12280 ( \12657 , \12652 , \12656 );
and \U$12281 ( \12658 , \4334 , \2980 );
and \U$12282 ( \12659 , \4078 , \2978 );
nor \U$12283 ( \12660 , \12658 , \12659 );
xnor \U$12284 ( \12661 , \12660 , \2831 );
and \U$12285 ( \12662 , \12656 , \12661 );
and \U$12286 ( \12663 , \12652 , \12661 );
or \U$12287 ( \12664 , \12657 , \12662 , \12663 );
and \U$12288 ( \12665 , \2703 , \4868 );
and \U$12289 ( \12666 , \2439 , \4866 );
nor \U$12290 ( \12667 , \12665 , \12666 );
xnor \U$12291 ( \12668 , \12667 , \4636 );
and \U$12292 ( \12669 , \2902 , \4417 );
and \U$12293 ( \12670 , \2728 , \4415 );
nor \U$12294 ( \12671 , \12669 , \12670 );
xnor \U$12295 ( \12672 , \12671 , \4274 );
and \U$12296 ( \12673 , \12668 , \12672 );
and \U$12297 ( \12674 , \3207 , \4094 );
and \U$12298 ( \12675 , \3069 , \4092 );
nor \U$12299 ( \12676 , \12674 , \12675 );
xnor \U$12300 ( \12677 , \12676 , \3848 );
and \U$12301 ( \12678 , \12672 , \12677 );
and \U$12302 ( \12679 , \12668 , \12677 );
or \U$12303 ( \12680 , \12673 , \12678 , \12679 );
and \U$12304 ( \12681 , \12664 , \12680 );
and \U$12305 ( \12682 , \1853 , \6297 );
and \U$12306 ( \12683 , \1677 , \6295 );
nor \U$12307 ( \12684 , \12682 , \12683 );
xnor \U$12308 ( \12685 , \12684 , \5957 );
and \U$12309 ( \12686 , \2104 , \5708 );
and \U$12310 ( \12687 , \1861 , \5706 );
nor \U$12311 ( \12688 , \12686 , \12687 );
xnor \U$12312 ( \12689 , \12688 , \5467 );
and \U$12313 ( \12690 , \12685 , \12689 );
and \U$12314 ( \12691 , \2295 , \5242 );
and \U$12315 ( \12692 , \2109 , \5240 );
nor \U$12316 ( \12693 , \12691 , \12692 );
xnor \U$12317 ( \12694 , \12693 , \5054 );
and \U$12318 ( \12695 , \12689 , \12694 );
and \U$12319 ( \12696 , \12685 , \12694 );
or \U$12320 ( \12697 , \12690 , \12695 , \12696 );
and \U$12321 ( \12698 , \12680 , \12697 );
and \U$12322 ( \12699 , \12664 , \12697 );
or \U$12323 ( \12700 , \12681 , \12698 , \12699 );
and \U$12324 ( \12701 , \12648 , \12700 );
and \U$12325 ( \12702 , \4833 , \2658 );
and \U$12326 ( \12703 , \4531 , \2656 );
nor \U$12327 ( \12704 , \12702 , \12703 );
xnor \U$12328 ( \12705 , \12704 , \2516 );
and \U$12329 ( \12706 , \5310 , \2362 );
and \U$12330 ( \12707 , \4841 , \2360 );
nor \U$12331 ( \12708 , \12706 , \12707 );
xnor \U$12332 ( \12709 , \12708 , \2225 );
and \U$12333 ( \12710 , \12705 , \12709 );
and \U$12334 ( \12711 , \5579 , \2156 );
and \U$12335 ( \12712 , \5315 , \2154 );
nor \U$12336 ( \12713 , \12711 , \12712 );
xnor \U$12337 ( \12714 , \12713 , \2004 );
and \U$12338 ( \12715 , \12709 , \12714 );
and \U$12339 ( \12716 , \12705 , \12714 );
or \U$12340 ( \12717 , \12710 , \12715 , \12716 );
and \U$12341 ( \12718 , \6210 , \1888 );
and \U$12342 ( \12719 , \5838 , \1886 );
nor \U$12343 ( \12720 , \12718 , \12719 );
xnor \U$12344 ( \12721 , \12720 , \1732 );
and \U$12345 ( \12722 , \6562 , \1616 );
and \U$12346 ( \12723 , \6219 , \1614 );
nor \U$12347 ( \12724 , \12722 , \12723 );
xnor \U$12348 ( \12725 , \12724 , \1503 );
and \U$12349 ( \12726 , \12721 , \12725 );
and \U$12350 ( \12727 , \7067 , \1422 );
and \U$12351 ( \12728 , \6764 , \1420 );
nor \U$12352 ( \12729 , \12727 , \12728 );
xnor \U$12353 ( \12730 , \12729 , \1286 );
and \U$12354 ( \12731 , \12725 , \12730 );
and \U$12355 ( \12732 , \12721 , \12730 );
or \U$12356 ( \12733 , \12726 , \12731 , \12732 );
and \U$12357 ( \12734 , \12717 , \12733 );
and \U$12358 ( \12735 , \7765 , \1222 );
and \U$12359 ( \12736 , \7239 , \1220 );
nor \U$12360 ( \12737 , \12735 , \12736 );
xnor \U$12361 ( \12738 , \12737 , \1144 );
and \U$12362 ( \12739 , \8435 , \1058 );
and \U$12363 ( \12740 , \8189 , \1056 );
nor \U$12364 ( \12741 , \12739 , \12740 );
xnor \U$12365 ( \12742 , \12741 , \964 );
and \U$12366 ( \12743 , \12738 , \12742 );
and \U$12367 ( \12744 , \8759 , \888 );
and \U$12368 ( \12745 , \8440 , \886 );
nor \U$12369 ( \12746 , \12744 , \12745 );
xnor \U$12370 ( \12747 , \12746 , \816 );
and \U$12371 ( \12748 , \12742 , \12747 );
and \U$12372 ( \12749 , \12738 , \12747 );
or \U$12373 ( \12750 , \12743 , \12748 , \12749 );
and \U$12374 ( \12751 , \12733 , \12750 );
and \U$12375 ( \12752 , \12717 , \12750 );
or \U$12376 ( \12753 , \12734 , \12751 , \12752 );
and \U$12377 ( \12754 , \12700 , \12753 );
and \U$12378 ( \12755 , \12648 , \12753 );
or \U$12379 ( \12756 , \12701 , \12754 , \12755 );
and \U$12380 ( \12757 , \12600 , \12756 );
xor \U$12381 ( \12758 , \12446 , \12448 );
xor \U$12382 ( \12759 , \12758 , \12451 );
xor \U$12383 ( \12760 , \12238 , \12240 );
xor \U$12384 ( \12761 , \12760 , \12243 );
and \U$12385 ( \12762 , \12759 , \12761 );
xor \U$12386 ( \12763 , \12248 , \12250 );
xor \U$12387 ( \12764 , \12763 , \12253 );
and \U$12388 ( \12765 , \12761 , \12764 );
and \U$12389 ( \12766 , \12759 , \12764 );
or \U$12390 ( \12767 , \12762 , \12765 , \12766 );
and \U$12391 ( \12768 , \12756 , \12767 );
and \U$12392 ( \12769 , \12600 , \12767 );
or \U$12393 ( \12770 , \12757 , \12768 , \12769 );
xor \U$12394 ( \12771 , \12299 , \12315 );
xor \U$12395 ( \12772 , \12771 , \12332 );
xor \U$12396 ( \12773 , \12404 , \12420 );
xor \U$12397 ( \12774 , \12773 , \12437 );
and \U$12398 ( \12775 , \12772 , \12774 );
xor \U$12399 ( \12776 , \12273 , \12275 );
xor \U$12400 ( \12777 , \12776 , \12277 );
and \U$12401 ( \12778 , \12774 , \12777 );
and \U$12402 ( \12779 , \12772 , \12777 );
or \U$12403 ( \12780 , \12775 , \12778 , \12779 );
xor \U$12404 ( \12781 , \12467 , \12469 );
xor \U$12405 ( \12782 , \12781 , \12472 );
and \U$12406 ( \12783 , \12780 , \12782 );
xor \U$12407 ( \12784 , \12477 , \12479 );
xor \U$12408 ( \12785 , \12784 , \12482 );
and \U$12409 ( \12786 , \12782 , \12785 );
and \U$12410 ( \12787 , \12780 , \12785 );
or \U$12411 ( \12788 , \12783 , \12786 , \12787 );
and \U$12412 ( \12789 , \12770 , \12788 );
xor \U$12413 ( \12790 , \12246 , \12256 );
xor \U$12414 ( \12791 , \12790 , \12280 );
xor \U$12415 ( \12792 , \12335 , \12387 );
xor \U$12416 ( \12793 , \12792 , \12440 );
and \U$12417 ( \12794 , \12791 , \12793 );
xor \U$12418 ( \12795 , \12454 , \12456 );
xor \U$12419 ( \12796 , \12795 , \12459 );
and \U$12420 ( \12797 , \12793 , \12796 );
and \U$12421 ( \12798 , \12791 , \12796 );
or \U$12422 ( \12799 , \12794 , \12797 , \12798 );
and \U$12423 ( \12800 , \12788 , \12799 );
and \U$12424 ( \12801 , \12770 , \12799 );
or \U$12425 ( \12802 , \12789 , \12800 , \12801 );
xor \U$12426 ( \12803 , \11988 , \12036 );
xor \U$12427 ( \12804 , \12803 , \12089 );
xor \U$12428 ( \12805 , \12123 , \12133 );
xor \U$12429 ( \12806 , \12805 , \12144 );
and \U$12430 ( \12807 , \12804 , \12806 );
xor \U$12431 ( \12808 , \12494 , \12496 );
xor \U$12432 ( \12809 , \12808 , \12499 );
and \U$12433 ( \12810 , \12806 , \12809 );
and \U$12434 ( \12811 , \12804 , \12809 );
or \U$12435 ( \12812 , \12807 , \12810 , \12811 );
and \U$12436 ( \12813 , \12802 , \12812 );
xor \U$12437 ( \12814 , \12507 , \12509 );
xor \U$12438 ( \12815 , \12814 , \12512 );
and \U$12439 ( \12816 , \12812 , \12815 );
and \U$12440 ( \12817 , \12802 , \12815 );
or \U$12441 ( \12818 , \12813 , \12816 , \12817 );
xor \U$12442 ( \12819 , \12505 , \12515 );
xor \U$12443 ( \12820 , \12819 , \12518 );
and \U$12444 ( \12821 , \12818 , \12820 );
xor \U$12445 ( \12822 , \12523 , \12525 );
xor \U$12446 ( \12823 , \12822 , \12528 );
and \U$12447 ( \12824 , \12820 , \12823 );
and \U$12448 ( \12825 , \12818 , \12823 );
or \U$12449 ( \12826 , \12821 , \12824 , \12825 );
xor \U$12450 ( \12827 , \12521 , \12531 );
xor \U$12451 ( \12828 , \12827 , \12534 );
and \U$12452 ( \12829 , \12826 , \12828 );
xor \U$12453 ( \12830 , \12539 , \12541 );
and \U$12454 ( \12831 , \12828 , \12830 );
and \U$12455 ( \12832 , \12826 , \12830 );
or \U$12456 ( \12833 , \12829 , \12831 , \12832 );
and \U$12457 ( \12834 , \12552 , \12833 );
xor \U$12458 ( \12835 , \12552 , \12833 );
xor \U$12459 ( \12836 , \12826 , \12828 );
xor \U$12460 ( \12837 , \12836 , \12830 );
and \U$12461 ( \12838 , \3069 , \4417 );
and \U$12462 ( \12839 , \2902 , \4415 );
nor \U$12463 ( \12840 , \12838 , \12839 );
xnor \U$12464 ( \12841 , \12840 , \4274 );
and \U$12465 ( \12842 , \3326 , \4094 );
and \U$12466 ( \12843 , \3207 , \4092 );
nor \U$12467 ( \12844 , \12842 , \12843 );
xnor \U$12468 ( \12845 , \12844 , \3848 );
and \U$12469 ( \12846 , \12841 , \12845 );
and \U$12470 ( \12847 , \3951 , \3699 );
and \U$12471 ( \12848 , \3743 , \3697 );
nor \U$12472 ( \12849 , \12847 , \12848 );
xnor \U$12473 ( \12850 , \12849 , \3512 );
and \U$12474 ( \12851 , \12845 , \12850 );
and \U$12475 ( \12852 , \12841 , \12850 );
or \U$12476 ( \12853 , \12846 , \12851 , \12852 );
and \U$12477 ( \12854 , \4078 , \3386 );
and \U$12478 ( \12855 , \4073 , \3384 );
nor \U$12479 ( \12856 , \12854 , \12855 );
xnor \U$12480 ( \12857 , \12856 , \3181 );
and \U$12481 ( \12858 , \4531 , \2980 );
and \U$12482 ( \12859 , \4334 , \2978 );
nor \U$12483 ( \12860 , \12858 , \12859 );
xnor \U$12484 ( \12861 , \12860 , \2831 );
and \U$12485 ( \12862 , \12857 , \12861 );
and \U$12486 ( \12863 , \4841 , \2658 );
and \U$12487 ( \12864 , \4833 , \2656 );
nor \U$12488 ( \12865 , \12863 , \12864 );
xnor \U$12489 ( \12866 , \12865 , \2516 );
and \U$12490 ( \12867 , \12861 , \12866 );
and \U$12491 ( \12868 , \12857 , \12866 );
or \U$12492 ( \12869 , \12862 , \12867 , \12868 );
and \U$12493 ( \12870 , \12853 , \12869 );
and \U$12494 ( \12871 , \2109 , \5708 );
and \U$12495 ( \12872 , \2104 , \5706 );
nor \U$12496 ( \12873 , \12871 , \12872 );
xnor \U$12497 ( \12874 , \12873 , \5467 );
and \U$12498 ( \12875 , \2439 , \5242 );
and \U$12499 ( \12876 , \2295 , \5240 );
nor \U$12500 ( \12877 , \12875 , \12876 );
xnor \U$12501 ( \12878 , \12877 , \5054 );
and \U$12502 ( \12879 , \12874 , \12878 );
and \U$12503 ( \12880 , \2728 , \4868 );
and \U$12504 ( \12881 , \2703 , \4866 );
nor \U$12505 ( \12882 , \12880 , \12881 );
xnor \U$12506 ( \12883 , \12882 , \4636 );
and \U$12507 ( \12884 , \12878 , \12883 );
and \U$12508 ( \12885 , \12874 , \12883 );
or \U$12509 ( \12886 , \12879 , \12884 , \12885 );
and \U$12510 ( \12887 , \12869 , \12886 );
and \U$12511 ( \12888 , \12853 , \12886 );
or \U$12512 ( \12889 , \12870 , \12887 , \12888 );
and \U$12513 ( \12890 , \6764 , \1616 );
and \U$12514 ( \12891 , \6562 , \1614 );
nor \U$12515 ( \12892 , \12890 , \12891 );
xnor \U$12516 ( \12893 , \12892 , \1503 );
and \U$12517 ( \12894 , \7239 , \1422 );
and \U$12518 ( \12895 , \7067 , \1420 );
nor \U$12519 ( \12896 , \12894 , \12895 );
xnor \U$12520 ( \12897 , \12896 , \1286 );
and \U$12521 ( \12898 , \12893 , \12897 );
and \U$12522 ( \12899 , \8189 , \1222 );
and \U$12523 ( \12900 , \7765 , \1220 );
nor \U$12524 ( \12901 , \12899 , \12900 );
xnor \U$12525 ( \12902 , \12901 , \1144 );
and \U$12526 ( \12903 , \12897 , \12902 );
and \U$12527 ( \12904 , \12893 , \12902 );
or \U$12528 ( \12905 , \12898 , \12903 , \12904 );
and \U$12529 ( \12906 , \8440 , \1058 );
and \U$12530 ( \12907 , \8435 , \1056 );
nor \U$12531 ( \12908 , \12906 , \12907 );
xnor \U$12532 ( \12909 , \12908 , \964 );
and \U$12533 ( \12910 , \9043 , \888 );
and \U$12534 ( \12911 , \8759 , \886 );
nor \U$12535 ( \12912 , \12910 , \12911 );
xnor \U$12536 ( \12913 , \12912 , \816 );
and \U$12537 ( \12914 , \12909 , \12913 );
and \U$12538 ( \12915 , \9620 , \754 );
and \U$12539 ( \12916 , \9612 , \752 );
nor \U$12540 ( \12917 , \12915 , \12916 );
xnor \U$12541 ( \12918 , \12917 , \711 );
and \U$12542 ( \12919 , \12913 , \12918 );
and \U$12543 ( \12920 , \12909 , \12918 );
or \U$12544 ( \12921 , \12914 , \12919 , \12920 );
and \U$12545 ( \12922 , \12905 , \12921 );
and \U$12546 ( \12923 , \5315 , \2362 );
and \U$12547 ( \12924 , \5310 , \2360 );
nor \U$12548 ( \12925 , \12923 , \12924 );
xnor \U$12549 ( \12926 , \12925 , \2225 );
and \U$12550 ( \12927 , \5838 , \2156 );
and \U$12551 ( \12928 , \5579 , \2154 );
nor \U$12552 ( \12929 , \12927 , \12928 );
xnor \U$12553 ( \12930 , \12929 , \2004 );
and \U$12554 ( \12931 , \12926 , \12930 );
and \U$12555 ( \12932 , \6219 , \1888 );
and \U$12556 ( \12933 , \6210 , \1886 );
nor \U$12557 ( \12934 , \12932 , \12933 );
xnor \U$12558 ( \12935 , \12934 , \1732 );
and \U$12559 ( \12936 , \12930 , \12935 );
and \U$12560 ( \12937 , \12926 , \12935 );
or \U$12561 ( \12938 , \12931 , \12936 , \12937 );
and \U$12562 ( \12939 , \12921 , \12938 );
and \U$12563 ( \12940 , \12905 , \12938 );
or \U$12564 ( \12941 , \12922 , \12939 , \12940 );
and \U$12565 ( \12942 , \12889 , \12941 );
and \U$12566 ( \12943 , \561 , \10876 );
and \U$12567 ( \12944 , \556 , \10873 );
nor \U$12568 ( \12945 , \12943 , \12944 );
xnor \U$12569 ( \12946 , \12945 , \9821 );
and \U$12570 ( \12947 , \666 , \10063 );
and \U$12571 ( \12948 , \615 , \10061 );
nor \U$12572 ( \12949 , \12947 , \12948 );
xnor \U$12573 ( \12950 , \12949 , \9824 );
and \U$12574 ( \12951 , \12946 , \12950 );
and \U$12575 ( \12952 , \771 , \9495 );
and \U$12576 ( \12953 , \743 , \9493 );
nor \U$12577 ( \12954 , \12952 , \12953 );
xnor \U$12578 ( \12955 , \12954 , \9185 );
and \U$12579 ( \12956 , \12950 , \12955 );
and \U$12580 ( \12957 , \12946 , \12955 );
or \U$12581 ( \12958 , \12951 , \12956 , \12957 );
and \U$12582 ( \12959 , \925 , \8958 );
and \U$12583 ( \12960 , \851 , \8956 );
nor \U$12584 ( \12961 , \12959 , \12960 );
xnor \U$12585 ( \12962 , \12961 , \8587 );
and \U$12586 ( \12963 , \1050 , \8396 );
and \U$12587 ( \12964 , \987 , \8394 );
nor \U$12588 ( \12965 , \12963 , \12964 );
xnor \U$12589 ( \12966 , \12965 , \8078 );
and \U$12590 ( \12967 , \12962 , \12966 );
and \U$12591 ( \12968 , \1336 , \7829 );
and \U$12592 ( \12969 , \1248 , \7827 );
nor \U$12593 ( \12970 , \12968 , \12969 );
xnor \U$12594 ( \12971 , \12970 , \7580 );
and \U$12595 ( \12972 , \12966 , \12971 );
and \U$12596 ( \12973 , \12962 , \12971 );
or \U$12597 ( \12974 , \12967 , \12972 , \12973 );
and \U$12598 ( \12975 , \12958 , \12974 );
and \U$12599 ( \12976 , \1446 , \7300 );
and \U$12600 ( \12977 , \1441 , \7298 );
nor \U$12601 ( \12978 , \12976 , \12977 );
xnor \U$12602 ( \12979 , \12978 , \7040 );
and \U$12603 ( \12980 , \1677 , \6806 );
and \U$12604 ( \12981 , \1562 , \6804 );
nor \U$12605 ( \12982 , \12980 , \12981 );
xnor \U$12606 ( \12983 , \12982 , \6491 );
and \U$12607 ( \12984 , \12979 , \12983 );
and \U$12608 ( \12985 , \1861 , \6297 );
and \U$12609 ( \12986 , \1853 , \6295 );
nor \U$12610 ( \12987 , \12985 , \12986 );
xnor \U$12611 ( \12988 , \12987 , \5957 );
and \U$12612 ( \12989 , \12983 , \12988 );
and \U$12613 ( \12990 , \12979 , \12988 );
or \U$12614 ( \12991 , \12984 , \12989 , \12990 );
and \U$12615 ( \12992 , \12974 , \12991 );
and \U$12616 ( \12993 , \12958 , \12991 );
or \U$12617 ( \12994 , \12975 , \12992 , \12993 );
and \U$12618 ( \12995 , \12941 , \12994 );
and \U$12619 ( \12996 , \12889 , \12994 );
or \U$12620 ( \12997 , \12942 , \12995 , \12996 );
xor \U$12621 ( \12998 , \12604 , \12608 );
xor \U$12622 ( \12999 , \12998 , \12613 );
xor \U$12623 ( \13000 , \12668 , \12672 );
xor \U$12624 ( \13001 , \13000 , \12677 );
and \U$12625 ( \13002 , \12999 , \13001 );
xor \U$12626 ( \13003 , \12685 , \12689 );
xor \U$12627 ( \13004 , \13003 , \12694 );
and \U$12628 ( \13005 , \13001 , \13004 );
and \U$12629 ( \13006 , \12999 , \13004 );
or \U$12630 ( \13007 , \13002 , \13005 , \13006 );
xor \U$12631 ( \13008 , \12652 , \12656 );
xor \U$12632 ( \13009 , \13008 , \12661 );
xor \U$12633 ( \13010 , \12705 , \12709 );
xor \U$12634 ( \13011 , \13010 , \12714 );
and \U$12635 ( \13012 , \13009 , \13011 );
xor \U$12636 ( \13013 , \12721 , \12725 );
xor \U$12637 ( \13014 , \13013 , \12730 );
and \U$12638 ( \13015 , \13011 , \13014 );
and \U$12639 ( \13016 , \13009 , \13014 );
or \U$12640 ( \13017 , \13012 , \13015 , \13016 );
and \U$12641 ( \13018 , \13007 , \13017 );
nand \U$12642 ( \13019 , \11029 , \468 );
xnor \U$12643 ( \13020 , \13019 , \440 );
xor \U$12644 ( \13021 , \12738 , \12742 );
xor \U$12645 ( \13022 , \13021 , \12747 );
and \U$12646 ( \13023 , \13020 , \13022 );
xor \U$12647 ( \13024 , \12566 , \12570 );
xor \U$12648 ( \13025 , \13024 , \12575 );
and \U$12649 ( \13026 , \13022 , \13025 );
and \U$12650 ( \13027 , \13020 , \13025 );
or \U$12651 ( \13028 , \13023 , \13026 , \13027 );
and \U$12652 ( \13029 , \13017 , \13028 );
and \U$12653 ( \13030 , \13007 , \13028 );
or \U$12654 ( \13031 , \13018 , \13029 , \13030 );
and \U$12655 ( \13032 , \12997 , \13031 );
xor \U$12656 ( \13033 , \12355 , \12359 );
xor \U$12657 ( \13034 , \13033 , \12364 );
xor \U$12658 ( \13035 , \12372 , \12376 );
xor \U$12659 ( \13036 , \13035 , \12381 );
and \U$12660 ( \13037 , \13034 , \13036 );
xor \U$12661 ( \13038 , \12589 , \12591 );
xor \U$12662 ( \13039 , \13038 , \12594 );
and \U$12663 ( \13040 , \13036 , \13039 );
and \U$12664 ( \13041 , \13034 , \13039 );
or \U$12665 ( \13042 , \13037 , \13040 , \13041 );
and \U$12666 ( \13043 , \13031 , \13042 );
and \U$12667 ( \13044 , \12997 , \13042 );
or \U$12668 ( \13045 , \13032 , \13043 , \13044 );
xor \U$12669 ( \13046 , \12562 , \12586 );
xor \U$12670 ( \13047 , \13046 , \12597 );
xor \U$12671 ( \13048 , \12648 , \12700 );
xor \U$12672 ( \13049 , \13048 , \12753 );
and \U$12673 ( \13050 , \13047 , \13049 );
xor \U$12674 ( \13051 , \12759 , \12761 );
xor \U$12675 ( \13052 , \13051 , \12764 );
and \U$12676 ( \13053 , \13049 , \13052 );
and \U$12677 ( \13054 , \13047 , \13052 );
or \U$12678 ( \13055 , \13050 , \13053 , \13054 );
and \U$12679 ( \13056 , \13045 , \13055 );
xor \U$12680 ( \13057 , \12717 , \12733 );
xor \U$12681 ( \13058 , \13057 , \12750 );
xor \U$12682 ( \13059 , \12554 , \12556 );
xor \U$12683 ( \13060 , \13059 , \12559 );
and \U$12684 ( \13061 , \13058 , \13060 );
xor \U$12685 ( \13062 , \12578 , \12580 );
xor \U$12686 ( \13063 , \13062 , \12583 );
and \U$12687 ( \13064 , \13060 , \13063 );
and \U$12688 ( \13065 , \13058 , \13063 );
or \U$12689 ( \13066 , \13061 , \13064 , \13065 );
xor \U$12690 ( \13067 , \12351 , \12367 );
xor \U$12691 ( \13068 , \13067 , \12384 );
and \U$12692 ( \13069 , \13066 , \13068 );
xor \U$12693 ( \13070 , \12772 , \12774 );
xor \U$12694 ( \13071 , \13070 , \12777 );
and \U$12695 ( \13072 , \13068 , \13071 );
and \U$12696 ( \13073 , \13066 , \13071 );
or \U$12697 ( \13074 , \13069 , \13072 , \13073 );
and \U$12698 ( \13075 , \13055 , \13074 );
and \U$12699 ( \13076 , \13045 , \13074 );
or \U$12700 ( \13077 , \13056 , \13075 , \13076 );
xor \U$12701 ( \13078 , \12600 , \12756 );
xor \U$12702 ( \13079 , \13078 , \12767 );
xor \U$12703 ( \13080 , \12780 , \12782 );
xor \U$12704 ( \13081 , \13080 , \12785 );
and \U$12705 ( \13082 , \13079 , \13081 );
xor \U$12706 ( \13083 , \12791 , \12793 );
xor \U$12707 ( \13084 , \13083 , \12796 );
and \U$12708 ( \13085 , \13081 , \13084 );
and \U$12709 ( \13086 , \13079 , \13084 );
or \U$12710 ( \13087 , \13082 , \13085 , \13086 );
and \U$12711 ( \13088 , \13077 , \13087 );
xor \U$12712 ( \13089 , \12475 , \12485 );
xor \U$12713 ( \13090 , \13089 , \12488 );
and \U$12714 ( \13091 , \13087 , \13090 );
and \U$12715 ( \13092 , \13077 , \13090 );
or \U$12716 ( \13093 , \13088 , \13091 , \13092 );
xor \U$12717 ( \13094 , \12283 , \12443 );
xor \U$12718 ( \13095 , \13094 , \12462 );
xor \U$12719 ( \13096 , \12770 , \12788 );
xor \U$12720 ( \13097 , \13096 , \12799 );
and \U$12721 ( \13098 , \13095 , \13097 );
xor \U$12722 ( \13099 , \12804 , \12806 );
xor \U$12723 ( \13100 , \13099 , \12809 );
and \U$12724 ( \13101 , \13097 , \13100 );
and \U$12725 ( \13102 , \13095 , \13100 );
or \U$12726 ( \13103 , \13098 , \13101 , \13102 );
and \U$12727 ( \13104 , \13093 , \13103 );
xor \U$12728 ( \13105 , \12465 , \12491 );
xor \U$12729 ( \13106 , \13105 , \12502 );
and \U$12730 ( \13107 , \13103 , \13106 );
and \U$12731 ( \13108 , \13093 , \13106 );
or \U$12732 ( \13109 , \13104 , \13107 , \13108 );
xor \U$12733 ( \13110 , \12818 , \12820 );
xor \U$12734 ( \13111 , \13110 , \12823 );
and \U$12735 ( \13112 , \13109 , \13111 );
and \U$12736 ( \13113 , \12837 , \13112 );
xor \U$12737 ( \13114 , \12837 , \13112 );
xor \U$12738 ( \13115 , \13109 , \13111 );
and \U$12739 ( \13116 , \10223 , \754 );
and \U$12740 ( \13117 , \9620 , \752 );
nor \U$12741 ( \13118 , \13116 , \13117 );
xnor \U$12742 ( \13119 , \13118 , \711 );
and \U$12743 ( \13120 , \10409 , \641 );
and \U$12744 ( \13121 , \10228 , \639 );
nor \U$12745 ( \13122 , \13120 , \13121 );
xnor \U$12746 ( \13123 , \13122 , \592 );
and \U$12747 ( \13124 , \13119 , \13123 );
nand \U$12748 ( \13125 , \11029 , \538 );
xnor \U$12749 ( \13126 , \13125 , \499 );
and \U$12750 ( \13127 , \13123 , \13126 );
and \U$12751 ( \13128 , \13119 , \13126 );
or \U$12752 ( \13129 , \13124 , \13127 , \13128 );
and \U$12753 ( \13130 , \10228 , \641 );
and \U$12754 ( \13131 , \10223 , \639 );
nor \U$12755 ( \13132 , \13130 , \13131 );
xnor \U$12756 ( \13133 , \13132 , \592 );
and \U$12757 ( \13134 , \13129 , \13133 );
and \U$12758 ( \13135 , \11029 , \540 );
and \U$12759 ( \13136 , \10409 , \538 );
nor \U$12760 ( \13137 , \13135 , \13136 );
xnor \U$12761 ( \13138 , \13137 , \499 );
and \U$12762 ( \13139 , \13133 , \13138 );
and \U$12763 ( \13140 , \13129 , \13138 );
or \U$12764 ( \13141 , \13134 , \13139 , \13140 );
xor \U$12765 ( \13142 , \12893 , \12897 );
xor \U$12766 ( \13143 , \13142 , \12902 );
xor \U$12767 ( \13144 , \12909 , \12913 );
xor \U$12768 ( \13145 , \13144 , \12918 );
and \U$12769 ( \13146 , \13143 , \13145 );
xor \U$12770 ( \13147 , \12926 , \12930 );
xor \U$12771 ( \13148 , \13147 , \12935 );
and \U$12772 ( \13149 , \13145 , \13148 );
and \U$12773 ( \13150 , \13143 , \13148 );
or \U$12774 ( \13151 , \13146 , \13149 , \13150 );
and \U$12775 ( \13152 , \13141 , \13151 );
xor \U$12776 ( \13153 , \12841 , \12845 );
xor \U$12777 ( \13154 , \13153 , \12850 );
xor \U$12778 ( \13155 , \12857 , \12861 );
xor \U$12779 ( \13156 , \13155 , \12866 );
and \U$12780 ( \13157 , \13154 , \13156 );
xor \U$12781 ( \13158 , \12874 , \12878 );
xor \U$12782 ( \13159 , \13158 , \12883 );
and \U$12783 ( \13160 , \13156 , \13159 );
and \U$12784 ( \13161 , \13154 , \13159 );
or \U$12785 ( \13162 , \13157 , \13160 , \13161 );
and \U$12786 ( \13163 , \13151 , \13162 );
and \U$12787 ( \13164 , \13141 , \13162 );
or \U$12788 ( \13165 , \13152 , \13163 , \13164 );
and \U$12789 ( \13166 , \851 , \9495 );
and \U$12790 ( \13167 , \771 , \9493 );
nor \U$12791 ( \13168 , \13166 , \13167 );
xnor \U$12792 ( \13169 , \13168 , \9185 );
and \U$12793 ( \13170 , \987 , \8958 );
and \U$12794 ( \13171 , \925 , \8956 );
nor \U$12795 ( \13172 , \13170 , \13171 );
xnor \U$12796 ( \13173 , \13172 , \8587 );
and \U$12797 ( \13174 , \13169 , \13173 );
and \U$12798 ( \13175 , \1248 , \8396 );
and \U$12799 ( \13176 , \1050 , \8394 );
nor \U$12800 ( \13177 , \13175 , \13176 );
xnor \U$12801 ( \13178 , \13177 , \8078 );
and \U$12802 ( \13179 , \13173 , \13178 );
and \U$12803 ( \13180 , \13169 , \13178 );
or \U$12804 ( \13181 , \13174 , \13179 , \13180 );
and \U$12805 ( \13182 , \1441 , \7829 );
and \U$12806 ( \13183 , \1336 , \7827 );
nor \U$12807 ( \13184 , \13182 , \13183 );
xnor \U$12808 ( \13185 , \13184 , \7580 );
and \U$12809 ( \13186 , \1562 , \7300 );
and \U$12810 ( \13187 , \1446 , \7298 );
nor \U$12811 ( \13188 , \13186 , \13187 );
xnor \U$12812 ( \13189 , \13188 , \7040 );
and \U$12813 ( \13190 , \13185 , \13189 );
and \U$12814 ( \13191 , \1853 , \6806 );
and \U$12815 ( \13192 , \1677 , \6804 );
nor \U$12816 ( \13193 , \13191 , \13192 );
xnor \U$12817 ( \13194 , \13193 , \6491 );
and \U$12818 ( \13195 , \13189 , \13194 );
and \U$12819 ( \13196 , \13185 , \13194 );
or \U$12820 ( \13197 , \13190 , \13195 , \13196 );
and \U$12821 ( \13198 , \13181 , \13197 );
and \U$12822 ( \13199 , \615 , \10876 );
and \U$12823 ( \13200 , \561 , \10873 );
nor \U$12824 ( \13201 , \13199 , \13200 );
xnor \U$12825 ( \13202 , \13201 , \9821 );
and \U$12826 ( \13203 , \743 , \10063 );
and \U$12827 ( \13204 , \666 , \10061 );
nor \U$12828 ( \13205 , \13203 , \13204 );
xnor \U$12829 ( \13206 , \13205 , \9824 );
and \U$12830 ( \13207 , \13202 , \13206 );
and \U$12831 ( \13208 , \13206 , \499 );
and \U$12832 ( \13209 , \13202 , \499 );
or \U$12833 ( \13210 , \13207 , \13208 , \13209 );
and \U$12834 ( \13211 , \13197 , \13210 );
and \U$12835 ( \13212 , \13181 , \13210 );
or \U$12836 ( \13213 , \13198 , \13211 , \13212 );
and \U$12837 ( \13214 , \4073 , \3699 );
and \U$12838 ( \13215 , \3951 , \3697 );
nor \U$12839 ( \13216 , \13214 , \13215 );
xnor \U$12840 ( \13217 , \13216 , \3512 );
and \U$12841 ( \13218 , \4334 , \3386 );
and \U$12842 ( \13219 , \4078 , \3384 );
nor \U$12843 ( \13220 , \13218 , \13219 );
xnor \U$12844 ( \13221 , \13220 , \3181 );
and \U$12845 ( \13222 , \13217 , \13221 );
and \U$12846 ( \13223 , \4833 , \2980 );
and \U$12847 ( \13224 , \4531 , \2978 );
nor \U$12848 ( \13225 , \13223 , \13224 );
xnor \U$12849 ( \13226 , \13225 , \2831 );
and \U$12850 ( \13227 , \13221 , \13226 );
and \U$12851 ( \13228 , \13217 , \13226 );
or \U$12852 ( \13229 , \13222 , \13227 , \13228 );
and \U$12853 ( \13230 , \2104 , \6297 );
and \U$12854 ( \13231 , \1861 , \6295 );
nor \U$12855 ( \13232 , \13230 , \13231 );
xnor \U$12856 ( \13233 , \13232 , \5957 );
and \U$12857 ( \13234 , \2295 , \5708 );
and \U$12858 ( \13235 , \2109 , \5706 );
nor \U$12859 ( \13236 , \13234 , \13235 );
xnor \U$12860 ( \13237 , \13236 , \5467 );
and \U$12861 ( \13238 , \13233 , \13237 );
and \U$12862 ( \13239 , \2703 , \5242 );
and \U$12863 ( \13240 , \2439 , \5240 );
nor \U$12864 ( \13241 , \13239 , \13240 );
xnor \U$12865 ( \13242 , \13241 , \5054 );
and \U$12866 ( \13243 , \13237 , \13242 );
and \U$12867 ( \13244 , \13233 , \13242 );
or \U$12868 ( \13245 , \13238 , \13243 , \13244 );
and \U$12869 ( \13246 , \13229 , \13245 );
and \U$12870 ( \13247 , \2902 , \4868 );
and \U$12871 ( \13248 , \2728 , \4866 );
nor \U$12872 ( \13249 , \13247 , \13248 );
xnor \U$12873 ( \13250 , \13249 , \4636 );
and \U$12874 ( \13251 , \3207 , \4417 );
and \U$12875 ( \13252 , \3069 , \4415 );
nor \U$12876 ( \13253 , \13251 , \13252 );
xnor \U$12877 ( \13254 , \13253 , \4274 );
and \U$12878 ( \13255 , \13250 , \13254 );
and \U$12879 ( \13256 , \3743 , \4094 );
and \U$12880 ( \13257 , \3326 , \4092 );
nor \U$12881 ( \13258 , \13256 , \13257 );
xnor \U$12882 ( \13259 , \13258 , \3848 );
and \U$12883 ( \13260 , \13254 , \13259 );
and \U$12884 ( \13261 , \13250 , \13259 );
or \U$12885 ( \13262 , \13255 , \13260 , \13261 );
and \U$12886 ( \13263 , \13245 , \13262 );
and \U$12887 ( \13264 , \13229 , \13262 );
or \U$12888 ( \13265 , \13246 , \13263 , \13264 );
and \U$12889 ( \13266 , \13213 , \13265 );
and \U$12890 ( \13267 , \6562 , \1888 );
and \U$12891 ( \13268 , \6219 , \1886 );
nor \U$12892 ( \13269 , \13267 , \13268 );
xnor \U$12893 ( \13270 , \13269 , \1732 );
and \U$12894 ( \13271 , \7067 , \1616 );
and \U$12895 ( \13272 , \6764 , \1614 );
nor \U$12896 ( \13273 , \13271 , \13272 );
xnor \U$12897 ( \13274 , \13273 , \1503 );
and \U$12898 ( \13275 , \13270 , \13274 );
and \U$12899 ( \13276 , \7765 , \1422 );
and \U$12900 ( \13277 , \7239 , \1420 );
nor \U$12901 ( \13278 , \13276 , \13277 );
xnor \U$12902 ( \13279 , \13278 , \1286 );
and \U$12903 ( \13280 , \13274 , \13279 );
and \U$12904 ( \13281 , \13270 , \13279 );
or \U$12905 ( \13282 , \13275 , \13280 , \13281 );
and \U$12906 ( \13283 , \8435 , \1222 );
and \U$12907 ( \13284 , \8189 , \1220 );
nor \U$12908 ( \13285 , \13283 , \13284 );
xnor \U$12909 ( \13286 , \13285 , \1144 );
and \U$12910 ( \13287 , \8759 , \1058 );
and \U$12911 ( \13288 , \8440 , \1056 );
nor \U$12912 ( \13289 , \13287 , \13288 );
xnor \U$12913 ( \13290 , \13289 , \964 );
and \U$12914 ( \13291 , \13286 , \13290 );
and \U$12915 ( \13292 , \9612 , \888 );
and \U$12916 ( \13293 , \9043 , \886 );
nor \U$12917 ( \13294 , \13292 , \13293 );
xnor \U$12918 ( \13295 , \13294 , \816 );
and \U$12919 ( \13296 , \13290 , \13295 );
and \U$12920 ( \13297 , \13286 , \13295 );
or \U$12921 ( \13298 , \13291 , \13296 , \13297 );
and \U$12922 ( \13299 , \13282 , \13298 );
and \U$12923 ( \13300 , \5310 , \2658 );
and \U$12924 ( \13301 , \4841 , \2656 );
nor \U$12925 ( \13302 , \13300 , \13301 );
xnor \U$12926 ( \13303 , \13302 , \2516 );
and \U$12927 ( \13304 , \5579 , \2362 );
and \U$12928 ( \13305 , \5315 , \2360 );
nor \U$12929 ( \13306 , \13304 , \13305 );
xnor \U$12930 ( \13307 , \13306 , \2225 );
and \U$12931 ( \13308 , \13303 , \13307 );
and \U$12932 ( \13309 , \6210 , \2156 );
and \U$12933 ( \13310 , \5838 , \2154 );
nor \U$12934 ( \13311 , \13309 , \13310 );
xnor \U$12935 ( \13312 , \13311 , \2004 );
and \U$12936 ( \13313 , \13307 , \13312 );
and \U$12937 ( \13314 , \13303 , \13312 );
or \U$12938 ( \13315 , \13308 , \13313 , \13314 );
and \U$12939 ( \13316 , \13298 , \13315 );
and \U$12940 ( \13317 , \13282 , \13315 );
or \U$12941 ( \13318 , \13299 , \13316 , \13317 );
and \U$12942 ( \13319 , \13265 , \13318 );
and \U$12943 ( \13320 , \13213 , \13318 );
or \U$12944 ( \13321 , \13266 , \13319 , \13320 );
and \U$12945 ( \13322 , \13165 , \13321 );
xor \U$12946 ( \13323 , \12946 , \12950 );
xor \U$12947 ( \13324 , \13323 , \12955 );
xor \U$12948 ( \13325 , \12962 , \12966 );
xor \U$12949 ( \13326 , \13325 , \12971 );
and \U$12950 ( \13327 , \13324 , \13326 );
xor \U$12951 ( \13328 , \12979 , \12983 );
xor \U$12952 ( \13329 , \13328 , \12988 );
and \U$12953 ( \13330 , \13326 , \13329 );
and \U$12954 ( \13331 , \13324 , \13329 );
or \U$12955 ( \13332 , \13327 , \13330 , \13331 );
xor \U$12956 ( \13333 , \12620 , \12624 );
xor \U$12957 ( \13334 , \13333 , \440 );
and \U$12958 ( \13335 , \13332 , \13334 );
xor \U$12959 ( \13336 , \12633 , \12637 );
xor \U$12960 ( \13337 , \13336 , \12642 );
and \U$12961 ( \13338 , \13334 , \13337 );
and \U$12962 ( \13339 , \13332 , \13337 );
or \U$12963 ( \13340 , \13335 , \13338 , \13339 );
and \U$12964 ( \13341 , \13321 , \13340 );
and \U$12965 ( \13342 , \13165 , \13340 );
or \U$12966 ( \13343 , \13322 , \13341 , \13342 );
xor \U$12967 ( \13344 , \12853 , \12869 );
xor \U$12968 ( \13345 , \13344 , \12886 );
xor \U$12969 ( \13346 , \12905 , \12921 );
xor \U$12970 ( \13347 , \13346 , \12938 );
and \U$12971 ( \13348 , \13345 , \13347 );
xor \U$12972 ( \13349 , \12958 , \12974 );
xor \U$12973 ( \13350 , \13349 , \12991 );
and \U$12974 ( \13351 , \13347 , \13350 );
and \U$12975 ( \13352 , \13345 , \13350 );
or \U$12976 ( \13353 , \13348 , \13351 , \13352 );
xor \U$12977 ( \13354 , \12999 , \13001 );
xor \U$12978 ( \13355 , \13354 , \13004 );
xor \U$12979 ( \13356 , \13009 , \13011 );
xor \U$12980 ( \13357 , \13356 , \13014 );
and \U$12981 ( \13358 , \13355 , \13357 );
xor \U$12982 ( \13359 , \13020 , \13022 );
xor \U$12983 ( \13360 , \13359 , \13025 );
and \U$12984 ( \13361 , \13357 , \13360 );
and \U$12985 ( \13362 , \13355 , \13360 );
or \U$12986 ( \13363 , \13358 , \13361 , \13362 );
and \U$12987 ( \13364 , \13353 , \13363 );
xor \U$12988 ( \13365 , \12664 , \12680 );
xor \U$12989 ( \13366 , \13365 , \12697 );
and \U$12990 ( \13367 , \13363 , \13366 );
and \U$12991 ( \13368 , \13353 , \13366 );
or \U$12992 ( \13369 , \13364 , \13367 , \13368 );
and \U$12993 ( \13370 , \13343 , \13369 );
xor \U$12994 ( \13371 , \12616 , \12628 );
xor \U$12995 ( \13372 , \13371 , \12645 );
xor \U$12996 ( \13373 , \13034 , \13036 );
xor \U$12997 ( \13374 , \13373 , \13039 );
and \U$12998 ( \13375 , \13372 , \13374 );
xor \U$12999 ( \13376 , \13058 , \13060 );
xor \U$13000 ( \13377 , \13376 , \13063 );
and \U$13001 ( \13378 , \13374 , \13377 );
and \U$13002 ( \13379 , \13372 , \13377 );
or \U$13003 ( \13380 , \13375 , \13378 , \13379 );
and \U$13004 ( \13381 , \13369 , \13380 );
and \U$13005 ( \13382 , \13343 , \13380 );
or \U$13006 ( \13383 , \13370 , \13381 , \13382 );
xor \U$13007 ( \13384 , \12997 , \13031 );
xor \U$13008 ( \13385 , \13384 , \13042 );
xor \U$13009 ( \13386 , \13047 , \13049 );
xor \U$13010 ( \13387 , \13386 , \13052 );
and \U$13011 ( \13388 , \13385 , \13387 );
xor \U$13012 ( \13389 , \13066 , \13068 );
xor \U$13013 ( \13390 , \13389 , \13071 );
and \U$13014 ( \13391 , \13387 , \13390 );
and \U$13015 ( \13392 , \13385 , \13390 );
or \U$13016 ( \13393 , \13388 , \13391 , \13392 );
and \U$13017 ( \13394 , \13383 , \13393 );
xor \U$13018 ( \13395 , \13079 , \13081 );
xor \U$13019 ( \13396 , \13395 , \13084 );
and \U$13020 ( \13397 , \13393 , \13396 );
and \U$13021 ( \13398 , \13383 , \13396 );
or \U$13022 ( \13399 , \13394 , \13397 , \13398 );
xor \U$13023 ( \13400 , \13077 , \13087 );
xor \U$13024 ( \13401 , \13400 , \13090 );
and \U$13025 ( \13402 , \13399 , \13401 );
xor \U$13026 ( \13403 , \13095 , \13097 );
xor \U$13027 ( \13404 , \13403 , \13100 );
and \U$13028 ( \13405 , \13401 , \13404 );
and \U$13029 ( \13406 , \13399 , \13404 );
or \U$13030 ( \13407 , \13402 , \13405 , \13406 );
xor \U$13031 ( \13408 , \13093 , \13103 );
xor \U$13032 ( \13409 , \13408 , \13106 );
and \U$13033 ( \13410 , \13407 , \13409 );
xor \U$13034 ( \13411 , \12802 , \12812 );
xor \U$13035 ( \13412 , \13411 , \12815 );
and \U$13036 ( \13413 , \13409 , \13412 );
and \U$13037 ( \13414 , \13407 , \13412 );
or \U$13038 ( \13415 , \13410 , \13413 , \13414 );
and \U$13039 ( \13416 , \13115 , \13415 );
xor \U$13040 ( \13417 , \13115 , \13415 );
xor \U$13041 ( \13418 , \13407 , \13409 );
xor \U$13042 ( \13419 , \13418 , \13412 );
xor \U$13043 ( \13420 , \13169 , \13173 );
xor \U$13044 ( \13421 , \13420 , \13178 );
xor \U$13045 ( \13422 , \13185 , \13189 );
xor \U$13046 ( \13423 , \13422 , \13194 );
and \U$13047 ( \13424 , \13421 , \13423 );
xor \U$13048 ( \13425 , \13233 , \13237 );
xor \U$13049 ( \13426 , \13425 , \13242 );
and \U$13050 ( \13427 , \13423 , \13426 );
and \U$13051 ( \13428 , \13421 , \13426 );
or \U$13052 ( \13429 , \13424 , \13427 , \13428 );
xor \U$13053 ( \13430 , \13217 , \13221 );
xor \U$13054 ( \13431 , \13430 , \13226 );
xor \U$13055 ( \13432 , \13250 , \13254 );
xor \U$13056 ( \13433 , \13432 , \13259 );
and \U$13057 ( \13434 , \13431 , \13433 );
xor \U$13058 ( \13435 , \13303 , \13307 );
xor \U$13059 ( \13436 , \13435 , \13312 );
and \U$13060 ( \13437 , \13433 , \13436 );
and \U$13061 ( \13438 , \13431 , \13436 );
or \U$13062 ( \13439 , \13434 , \13437 , \13438 );
and \U$13063 ( \13440 , \13429 , \13439 );
xor \U$13064 ( \13441 , \13270 , \13274 );
xor \U$13065 ( \13442 , \13441 , \13279 );
xor \U$13066 ( \13443 , \13119 , \13123 );
xor \U$13067 ( \13444 , \13443 , \13126 );
and \U$13068 ( \13445 , \13442 , \13444 );
xor \U$13069 ( \13446 , \13286 , \13290 );
xor \U$13070 ( \13447 , \13446 , \13295 );
and \U$13071 ( \13448 , \13444 , \13447 );
and \U$13072 ( \13449 , \13442 , \13447 );
or \U$13073 ( \13450 , \13445 , \13448 , \13449 );
and \U$13074 ( \13451 , \13439 , \13450 );
and \U$13075 ( \13452 , \13429 , \13450 );
or \U$13076 ( \13453 , \13440 , \13451 , \13452 );
and \U$13077 ( \13454 , \2439 , \5708 );
and \U$13078 ( \13455 , \2295 , \5706 );
nor \U$13079 ( \13456 , \13454 , \13455 );
xnor \U$13080 ( \13457 , \13456 , \5467 );
and \U$13081 ( \13458 , \2728 , \5242 );
and \U$13082 ( \13459 , \2703 , \5240 );
nor \U$13083 ( \13460 , \13458 , \13459 );
xnor \U$13084 ( \13461 , \13460 , \5054 );
and \U$13085 ( \13462 , \13457 , \13461 );
and \U$13086 ( \13463 , \3069 , \4868 );
and \U$13087 ( \13464 , \2902 , \4866 );
nor \U$13088 ( \13465 , \13463 , \13464 );
xnor \U$13089 ( \13466 , \13465 , \4636 );
and \U$13090 ( \13467 , \13461 , \13466 );
and \U$13091 ( \13468 , \13457 , \13466 );
or \U$13092 ( \13469 , \13462 , \13467 , \13468 );
and \U$13093 ( \13470 , \4531 , \3386 );
and \U$13094 ( \13471 , \4334 , \3384 );
nor \U$13095 ( \13472 , \13470 , \13471 );
xnor \U$13096 ( \13473 , \13472 , \3181 );
and \U$13097 ( \13474 , \4841 , \2980 );
and \U$13098 ( \13475 , \4833 , \2978 );
nor \U$13099 ( \13476 , \13474 , \13475 );
xnor \U$13100 ( \13477 , \13476 , \2831 );
and \U$13101 ( \13478 , \13473 , \13477 );
and \U$13102 ( \13479 , \5315 , \2658 );
and \U$13103 ( \13480 , \5310 , \2656 );
nor \U$13104 ( \13481 , \13479 , \13480 );
xnor \U$13105 ( \13482 , \13481 , \2516 );
and \U$13106 ( \13483 , \13477 , \13482 );
and \U$13107 ( \13484 , \13473 , \13482 );
or \U$13108 ( \13485 , \13478 , \13483 , \13484 );
and \U$13109 ( \13486 , \13469 , \13485 );
and \U$13110 ( \13487 , \3326 , \4417 );
and \U$13111 ( \13488 , \3207 , \4415 );
nor \U$13112 ( \13489 , \13487 , \13488 );
xnor \U$13113 ( \13490 , \13489 , \4274 );
and \U$13114 ( \13491 , \3951 , \4094 );
and \U$13115 ( \13492 , \3743 , \4092 );
nor \U$13116 ( \13493 , \13491 , \13492 );
xnor \U$13117 ( \13494 , \13493 , \3848 );
and \U$13118 ( \13495 , \13490 , \13494 );
and \U$13119 ( \13496 , \4078 , \3699 );
and \U$13120 ( \13497 , \4073 , \3697 );
nor \U$13121 ( \13498 , \13496 , \13497 );
xnor \U$13122 ( \13499 , \13498 , \3512 );
and \U$13123 ( \13500 , \13494 , \13499 );
and \U$13124 ( \13501 , \13490 , \13499 );
or \U$13125 ( \13502 , \13495 , \13500 , \13501 );
and \U$13126 ( \13503 , \13485 , \13502 );
and \U$13127 ( \13504 , \13469 , \13502 );
or \U$13128 ( \13505 , \13486 , \13503 , \13504 );
and \U$13129 ( \13506 , \9043 , \1058 );
and \U$13130 ( \13507 , \8759 , \1056 );
nor \U$13131 ( \13508 , \13506 , \13507 );
xnor \U$13132 ( \13509 , \13508 , \964 );
and \U$13133 ( \13510 , \9620 , \888 );
and \U$13134 ( \13511 , \9612 , \886 );
nor \U$13135 ( \13512 , \13510 , \13511 );
xnor \U$13136 ( \13513 , \13512 , \816 );
and \U$13137 ( \13514 , \13509 , \13513 );
and \U$13138 ( \13515 , \10228 , \754 );
and \U$13139 ( \13516 , \10223 , \752 );
nor \U$13140 ( \13517 , \13515 , \13516 );
xnor \U$13141 ( \13518 , \13517 , \711 );
and \U$13142 ( \13519 , \13513 , \13518 );
and \U$13143 ( \13520 , \13509 , \13518 );
or \U$13144 ( \13521 , \13514 , \13519 , \13520 );
and \U$13145 ( \13522 , \7239 , \1616 );
and \U$13146 ( \13523 , \7067 , \1614 );
nor \U$13147 ( \13524 , \13522 , \13523 );
xnor \U$13148 ( \13525 , \13524 , \1503 );
and \U$13149 ( \13526 , \8189 , \1422 );
and \U$13150 ( \13527 , \7765 , \1420 );
nor \U$13151 ( \13528 , \13526 , \13527 );
xnor \U$13152 ( \13529 , \13528 , \1286 );
and \U$13153 ( \13530 , \13525 , \13529 );
and \U$13154 ( \13531 , \8440 , \1222 );
and \U$13155 ( \13532 , \8435 , \1220 );
nor \U$13156 ( \13533 , \13531 , \13532 );
xnor \U$13157 ( \13534 , \13533 , \1144 );
and \U$13158 ( \13535 , \13529 , \13534 );
and \U$13159 ( \13536 , \13525 , \13534 );
or \U$13160 ( \13537 , \13530 , \13535 , \13536 );
and \U$13161 ( \13538 , \13521 , \13537 );
and \U$13162 ( \13539 , \5838 , \2362 );
and \U$13163 ( \13540 , \5579 , \2360 );
nor \U$13164 ( \13541 , \13539 , \13540 );
xnor \U$13165 ( \13542 , \13541 , \2225 );
and \U$13166 ( \13543 , \6219 , \2156 );
and \U$13167 ( \13544 , \6210 , \2154 );
nor \U$13168 ( \13545 , \13543 , \13544 );
xnor \U$13169 ( \13546 , \13545 , \2004 );
and \U$13170 ( \13547 , \13542 , \13546 );
and \U$13171 ( \13548 , \6764 , \1888 );
and \U$13172 ( \13549 , \6562 , \1886 );
nor \U$13173 ( \13550 , \13548 , \13549 );
xnor \U$13174 ( \13551 , \13550 , \1732 );
and \U$13175 ( \13552 , \13546 , \13551 );
and \U$13176 ( \13553 , \13542 , \13551 );
or \U$13177 ( \13554 , \13547 , \13552 , \13553 );
and \U$13178 ( \13555 , \13537 , \13554 );
and \U$13179 ( \13556 , \13521 , \13554 );
or \U$13180 ( \13557 , \13538 , \13555 , \13556 );
and \U$13181 ( \13558 , \13505 , \13557 );
and \U$13182 ( \13559 , \1677 , \7300 );
and \U$13183 ( \13560 , \1562 , \7298 );
nor \U$13184 ( \13561 , \13559 , \13560 );
xnor \U$13185 ( \13562 , \13561 , \7040 );
and \U$13186 ( \13563 , \1861 , \6806 );
and \U$13187 ( \13564 , \1853 , \6804 );
nor \U$13188 ( \13565 , \13563 , \13564 );
xnor \U$13189 ( \13566 , \13565 , \6491 );
and \U$13190 ( \13567 , \13562 , \13566 );
and \U$13191 ( \13568 , \2109 , \6297 );
and \U$13192 ( \13569 , \2104 , \6295 );
nor \U$13193 ( \13570 , \13568 , \13569 );
xnor \U$13194 ( \13571 , \13570 , \5957 );
and \U$13195 ( \13572 , \13566 , \13571 );
and \U$13196 ( \13573 , \13562 , \13571 );
or \U$13197 ( \13574 , \13567 , \13572 , \13573 );
and \U$13198 ( \13575 , \666 , \10876 );
and \U$13199 ( \13576 , \615 , \10873 );
nor \U$13200 ( \13577 , \13575 , \13576 );
xnor \U$13201 ( \13578 , \13577 , \9821 );
and \U$13202 ( \13579 , \771 , \10063 );
and \U$13203 ( \13580 , \743 , \10061 );
nor \U$13204 ( \13581 , \13579 , \13580 );
xnor \U$13205 ( \13582 , \13581 , \9824 );
and \U$13206 ( \13583 , \13578 , \13582 );
and \U$13207 ( \13584 , \925 , \9495 );
and \U$13208 ( \13585 , \851 , \9493 );
nor \U$13209 ( \13586 , \13584 , \13585 );
xnor \U$13210 ( \13587 , \13586 , \9185 );
and \U$13211 ( \13588 , \13582 , \13587 );
and \U$13212 ( \13589 , \13578 , \13587 );
or \U$13213 ( \13590 , \13583 , \13588 , \13589 );
and \U$13214 ( \13591 , \13574 , \13590 );
and \U$13215 ( \13592 , \1050 , \8958 );
and \U$13216 ( \13593 , \987 , \8956 );
nor \U$13217 ( \13594 , \13592 , \13593 );
xnor \U$13218 ( \13595 , \13594 , \8587 );
and \U$13219 ( \13596 , \1336 , \8396 );
and \U$13220 ( \13597 , \1248 , \8394 );
nor \U$13221 ( \13598 , \13596 , \13597 );
xnor \U$13222 ( \13599 , \13598 , \8078 );
and \U$13223 ( \13600 , \13595 , \13599 );
and \U$13224 ( \13601 , \1446 , \7829 );
and \U$13225 ( \13602 , \1441 , \7827 );
nor \U$13226 ( \13603 , \13601 , \13602 );
xnor \U$13227 ( \13604 , \13603 , \7580 );
and \U$13228 ( \13605 , \13599 , \13604 );
and \U$13229 ( \13606 , \13595 , \13604 );
or \U$13230 ( \13607 , \13600 , \13605 , \13606 );
and \U$13231 ( \13608 , \13590 , \13607 );
and \U$13232 ( \13609 , \13574 , \13607 );
or \U$13233 ( \13610 , \13591 , \13608 , \13609 );
and \U$13234 ( \13611 , \13557 , \13610 );
and \U$13235 ( \13612 , \13505 , \13610 );
or \U$13236 ( \13613 , \13558 , \13611 , \13612 );
and \U$13237 ( \13614 , \13453 , \13613 );
xor \U$13238 ( \13615 , \13143 , \13145 );
xor \U$13239 ( \13616 , \13615 , \13148 );
xor \U$13240 ( \13617 , \13324 , \13326 );
xor \U$13241 ( \13618 , \13617 , \13329 );
and \U$13242 ( \13619 , \13616 , \13618 );
xor \U$13243 ( \13620 , \13154 , \13156 );
xor \U$13244 ( \13621 , \13620 , \13159 );
and \U$13245 ( \13622 , \13618 , \13621 );
and \U$13246 ( \13623 , \13616 , \13621 );
or \U$13247 ( \13624 , \13619 , \13622 , \13623 );
and \U$13248 ( \13625 , \13613 , \13624 );
and \U$13249 ( \13626 , \13453 , \13624 );
or \U$13250 ( \13627 , \13614 , \13625 , \13626 );
xor \U$13251 ( \13628 , \13141 , \13151 );
xor \U$13252 ( \13629 , \13628 , \13162 );
xor \U$13253 ( \13630 , \13213 , \13265 );
xor \U$13254 ( \13631 , \13630 , \13318 );
and \U$13255 ( \13632 , \13629 , \13631 );
xor \U$13256 ( \13633 , \13332 , \13334 );
xor \U$13257 ( \13634 , \13633 , \13337 );
and \U$13258 ( \13635 , \13631 , \13634 );
and \U$13259 ( \13636 , \13629 , \13634 );
or \U$13260 ( \13637 , \13632 , \13635 , \13636 );
and \U$13261 ( \13638 , \13627 , \13637 );
xor \U$13262 ( \13639 , \13129 , \13133 );
xor \U$13263 ( \13640 , \13639 , \13138 );
xor \U$13264 ( \13641 , \13229 , \13245 );
xor \U$13265 ( \13642 , \13641 , \13262 );
and \U$13266 ( \13643 , \13640 , \13642 );
xor \U$13267 ( \13644 , \13282 , \13298 );
xor \U$13268 ( \13645 , \13644 , \13315 );
and \U$13269 ( \13646 , \13642 , \13645 );
and \U$13270 ( \13647 , \13640 , \13645 );
or \U$13271 ( \13648 , \13643 , \13646 , \13647 );
xor \U$13272 ( \13649 , \13345 , \13347 );
xor \U$13273 ( \13650 , \13649 , \13350 );
and \U$13274 ( \13651 , \13648 , \13650 );
xor \U$13275 ( \13652 , \13355 , \13357 );
xor \U$13276 ( \13653 , \13652 , \13360 );
and \U$13277 ( \13654 , \13650 , \13653 );
and \U$13278 ( \13655 , \13648 , \13653 );
or \U$13279 ( \13656 , \13651 , \13654 , \13655 );
and \U$13280 ( \13657 , \13637 , \13656 );
and \U$13281 ( \13658 , \13627 , \13656 );
or \U$13282 ( \13659 , \13638 , \13657 , \13658 );
xor \U$13283 ( \13660 , \12889 , \12941 );
xor \U$13284 ( \13661 , \13660 , \12994 );
xor \U$13285 ( \13662 , \13007 , \13017 );
xor \U$13286 ( \13663 , \13662 , \13028 );
and \U$13287 ( \13664 , \13661 , \13663 );
xor \U$13288 ( \13665 , \13372 , \13374 );
xor \U$13289 ( \13666 , \13665 , \13377 );
and \U$13290 ( \13667 , \13663 , \13666 );
and \U$13291 ( \13668 , \13661 , \13666 );
or \U$13292 ( \13669 , \13664 , \13667 , \13668 );
and \U$13293 ( \13670 , \13659 , \13669 );
xor \U$13294 ( \13671 , \13385 , \13387 );
xor \U$13295 ( \13672 , \13671 , \13390 );
and \U$13296 ( \13673 , \13669 , \13672 );
and \U$13297 ( \13674 , \13659 , \13672 );
or \U$13298 ( \13675 , \13670 , \13673 , \13674 );
xor \U$13299 ( \13676 , \13045 , \13055 );
xor \U$13300 ( \13677 , \13676 , \13074 );
and \U$13301 ( \13678 , \13675 , \13677 );
xor \U$13302 ( \13679 , \13383 , \13393 );
xor \U$13303 ( \13680 , \13679 , \13396 );
and \U$13304 ( \13681 , \13677 , \13680 );
and \U$13305 ( \13682 , \13675 , \13680 );
or \U$13306 ( \13683 , \13678 , \13681 , \13682 );
xor \U$13307 ( \13684 , \13399 , \13401 );
xor \U$13308 ( \13685 , \13684 , \13404 );
and \U$13309 ( \13686 , \13683 , \13685 );
and \U$13310 ( \13687 , \13419 , \13686 );
xor \U$13311 ( \13688 , \13419 , \13686 );
xor \U$13312 ( \13689 , \13683 , \13685 );
xor \U$13313 ( \13690 , \13473 , \13477 );
xor \U$13314 ( \13691 , \13690 , \13482 );
xor \U$13315 ( \13692 , \13490 , \13494 );
xor \U$13316 ( \13693 , \13692 , \13499 );
and \U$13317 ( \13694 , \13691 , \13693 );
xor \U$13318 ( \13695 , \13542 , \13546 );
xor \U$13319 ( \13696 , \13695 , \13551 );
and \U$13320 ( \13697 , \13693 , \13696 );
and \U$13321 ( \13698 , \13691 , \13696 );
or \U$13322 ( \13699 , \13694 , \13697 , \13698 );
xor \U$13323 ( \13700 , \13457 , \13461 );
xor \U$13324 ( \13701 , \13700 , \13466 );
xor \U$13325 ( \13702 , \13562 , \13566 );
xor \U$13326 ( \13703 , \13702 , \13571 );
and \U$13327 ( \13704 , \13701 , \13703 );
xor \U$13328 ( \13705 , \13595 , \13599 );
xor \U$13329 ( \13706 , \13705 , \13604 );
and \U$13330 ( \13707 , \13703 , \13706 );
and \U$13331 ( \13708 , \13701 , \13706 );
or \U$13332 ( \13709 , \13704 , \13707 , \13708 );
and \U$13333 ( \13710 , \13699 , \13709 );
and \U$13334 ( \13711 , \11029 , \641 );
and \U$13335 ( \13712 , \10409 , \639 );
nor \U$13336 ( \13713 , \13711 , \13712 );
xnor \U$13337 ( \13714 , \13713 , \592 );
xor \U$13338 ( \13715 , \13509 , \13513 );
xor \U$13339 ( \13716 , \13715 , \13518 );
and \U$13340 ( \13717 , \13714 , \13716 );
xor \U$13341 ( \13718 , \13525 , \13529 );
xor \U$13342 ( \13719 , \13718 , \13534 );
and \U$13343 ( \13720 , \13716 , \13719 );
and \U$13344 ( \13721 , \13714 , \13719 );
or \U$13345 ( \13722 , \13717 , \13720 , \13721 );
and \U$13346 ( \13723 , \13709 , \13722 );
and \U$13347 ( \13724 , \13699 , \13722 );
or \U$13348 ( \13725 , \13710 , \13723 , \13724 );
and \U$13349 ( \13726 , \1562 , \7829 );
and \U$13350 ( \13727 , \1446 , \7827 );
nor \U$13351 ( \13728 , \13726 , \13727 );
xnor \U$13352 ( \13729 , \13728 , \7580 );
and \U$13353 ( \13730 , \1853 , \7300 );
and \U$13354 ( \13731 , \1677 , \7298 );
nor \U$13355 ( \13732 , \13730 , \13731 );
xnor \U$13356 ( \13733 , \13732 , \7040 );
and \U$13357 ( \13734 , \13729 , \13733 );
and \U$13358 ( \13735 , \2104 , \6806 );
and \U$13359 ( \13736 , \1861 , \6804 );
nor \U$13360 ( \13737 , \13735 , \13736 );
xnor \U$13361 ( \13738 , \13737 , \6491 );
and \U$13362 ( \13739 , \13733 , \13738 );
and \U$13363 ( \13740 , \13729 , \13738 );
or \U$13364 ( \13741 , \13734 , \13739 , \13740 );
and \U$13365 ( \13742 , \987 , \9495 );
and \U$13366 ( \13743 , \925 , \9493 );
nor \U$13367 ( \13744 , \13742 , \13743 );
xnor \U$13368 ( \13745 , \13744 , \9185 );
and \U$13369 ( \13746 , \1248 , \8958 );
and \U$13370 ( \13747 , \1050 , \8956 );
nor \U$13371 ( \13748 , \13746 , \13747 );
xnor \U$13372 ( \13749 , \13748 , \8587 );
and \U$13373 ( \13750 , \13745 , \13749 );
and \U$13374 ( \13751 , \1441 , \8396 );
and \U$13375 ( \13752 , \1336 , \8394 );
nor \U$13376 ( \13753 , \13751 , \13752 );
xnor \U$13377 ( \13754 , \13753 , \8078 );
and \U$13378 ( \13755 , \13749 , \13754 );
and \U$13379 ( \13756 , \13745 , \13754 );
or \U$13380 ( \13757 , \13750 , \13755 , \13756 );
and \U$13381 ( \13758 , \13741 , \13757 );
and \U$13382 ( \13759 , \743 , \10876 );
and \U$13383 ( \13760 , \666 , \10873 );
nor \U$13384 ( \13761 , \13759 , \13760 );
xnor \U$13385 ( \13762 , \13761 , \9821 );
and \U$13386 ( \13763 , \851 , \10063 );
and \U$13387 ( \13764 , \771 , \10061 );
nor \U$13388 ( \13765 , \13763 , \13764 );
xnor \U$13389 ( \13766 , \13765 , \9824 );
and \U$13390 ( \13767 , \13762 , \13766 );
and \U$13391 ( \13768 , \13766 , \592 );
and \U$13392 ( \13769 , \13762 , \592 );
or \U$13393 ( \13770 , \13767 , \13768 , \13769 );
and \U$13394 ( \13771 , \13757 , \13770 );
and \U$13395 ( \13772 , \13741 , \13770 );
or \U$13396 ( \13773 , \13758 , \13771 , \13772 );
and \U$13397 ( \13774 , \8759 , \1222 );
and \U$13398 ( \13775 , \8440 , \1220 );
nor \U$13399 ( \13776 , \13774 , \13775 );
xnor \U$13400 ( \13777 , \13776 , \1144 );
and \U$13401 ( \13778 , \9612 , \1058 );
and \U$13402 ( \13779 , \9043 , \1056 );
nor \U$13403 ( \13780 , \13778 , \13779 );
xnor \U$13404 ( \13781 , \13780 , \964 );
and \U$13405 ( \13782 , \13777 , \13781 );
and \U$13406 ( \13783 , \10223 , \888 );
and \U$13407 ( \13784 , \9620 , \886 );
nor \U$13408 ( \13785 , \13783 , \13784 );
xnor \U$13409 ( \13786 , \13785 , \816 );
and \U$13410 ( \13787 , \13781 , \13786 );
and \U$13411 ( \13788 , \13777 , \13786 );
or \U$13412 ( \13789 , \13782 , \13787 , \13788 );
and \U$13413 ( \13790 , \5579 , \2658 );
and \U$13414 ( \13791 , \5315 , \2656 );
nor \U$13415 ( \13792 , \13790 , \13791 );
xnor \U$13416 ( \13793 , \13792 , \2516 );
and \U$13417 ( \13794 , \6210 , \2362 );
and \U$13418 ( \13795 , \5838 , \2360 );
nor \U$13419 ( \13796 , \13794 , \13795 );
xnor \U$13420 ( \13797 , \13796 , \2225 );
and \U$13421 ( \13798 , \13793 , \13797 );
and \U$13422 ( \13799 , \6562 , \2156 );
and \U$13423 ( \13800 , \6219 , \2154 );
nor \U$13424 ( \13801 , \13799 , \13800 );
xnor \U$13425 ( \13802 , \13801 , \2004 );
and \U$13426 ( \13803 , \13797 , \13802 );
and \U$13427 ( \13804 , \13793 , \13802 );
or \U$13428 ( \13805 , \13798 , \13803 , \13804 );
and \U$13429 ( \13806 , \13789 , \13805 );
and \U$13430 ( \13807 , \7067 , \1888 );
and \U$13431 ( \13808 , \6764 , \1886 );
nor \U$13432 ( \13809 , \13807 , \13808 );
xnor \U$13433 ( \13810 , \13809 , \1732 );
and \U$13434 ( \13811 , \7765 , \1616 );
and \U$13435 ( \13812 , \7239 , \1614 );
nor \U$13436 ( \13813 , \13811 , \13812 );
xnor \U$13437 ( \13814 , \13813 , \1503 );
and \U$13438 ( \13815 , \13810 , \13814 );
and \U$13439 ( \13816 , \8435 , \1422 );
and \U$13440 ( \13817 , \8189 , \1420 );
nor \U$13441 ( \13818 , \13816 , \13817 );
xnor \U$13442 ( \13819 , \13818 , \1286 );
and \U$13443 ( \13820 , \13814 , \13819 );
and \U$13444 ( \13821 , \13810 , \13819 );
or \U$13445 ( \13822 , \13815 , \13820 , \13821 );
and \U$13446 ( \13823 , \13805 , \13822 );
and \U$13447 ( \13824 , \13789 , \13822 );
or \U$13448 ( \13825 , \13806 , \13823 , \13824 );
and \U$13449 ( \13826 , \13773 , \13825 );
and \U$13450 ( \13827 , \4334 , \3699 );
and \U$13451 ( \13828 , \4078 , \3697 );
nor \U$13452 ( \13829 , \13827 , \13828 );
xnor \U$13453 ( \13830 , \13829 , \3512 );
and \U$13454 ( \13831 , \4833 , \3386 );
and \U$13455 ( \13832 , \4531 , \3384 );
nor \U$13456 ( \13833 , \13831 , \13832 );
xnor \U$13457 ( \13834 , \13833 , \3181 );
and \U$13458 ( \13835 , \13830 , \13834 );
and \U$13459 ( \13836 , \5310 , \2980 );
and \U$13460 ( \13837 , \4841 , \2978 );
nor \U$13461 ( \13838 , \13836 , \13837 );
xnor \U$13462 ( \13839 , \13838 , \2831 );
and \U$13463 ( \13840 , \13834 , \13839 );
and \U$13464 ( \13841 , \13830 , \13839 );
or \U$13465 ( \13842 , \13835 , \13840 , \13841 );
and \U$13466 ( \13843 , \3207 , \4868 );
and \U$13467 ( \13844 , \3069 , \4866 );
nor \U$13468 ( \13845 , \13843 , \13844 );
xnor \U$13469 ( \13846 , \13845 , \4636 );
and \U$13470 ( \13847 , \3743 , \4417 );
and \U$13471 ( \13848 , \3326 , \4415 );
nor \U$13472 ( \13849 , \13847 , \13848 );
xnor \U$13473 ( \13850 , \13849 , \4274 );
and \U$13474 ( \13851 , \13846 , \13850 );
and \U$13475 ( \13852 , \4073 , \4094 );
and \U$13476 ( \13853 , \3951 , \4092 );
nor \U$13477 ( \13854 , \13852 , \13853 );
xnor \U$13478 ( \13855 , \13854 , \3848 );
and \U$13479 ( \13856 , \13850 , \13855 );
and \U$13480 ( \13857 , \13846 , \13855 );
or \U$13481 ( \13858 , \13851 , \13856 , \13857 );
and \U$13482 ( \13859 , \13842 , \13858 );
and \U$13483 ( \13860 , \2295 , \6297 );
and \U$13484 ( \13861 , \2109 , \6295 );
nor \U$13485 ( \13862 , \13860 , \13861 );
xnor \U$13486 ( \13863 , \13862 , \5957 );
and \U$13487 ( \13864 , \2703 , \5708 );
and \U$13488 ( \13865 , \2439 , \5706 );
nor \U$13489 ( \13866 , \13864 , \13865 );
xnor \U$13490 ( \13867 , \13866 , \5467 );
and \U$13491 ( \13868 , \13863 , \13867 );
and \U$13492 ( \13869 , \2902 , \5242 );
and \U$13493 ( \13870 , \2728 , \5240 );
nor \U$13494 ( \13871 , \13869 , \13870 );
xnor \U$13495 ( \13872 , \13871 , \5054 );
and \U$13496 ( \13873 , \13867 , \13872 );
and \U$13497 ( \13874 , \13863 , \13872 );
or \U$13498 ( \13875 , \13868 , \13873 , \13874 );
and \U$13499 ( \13876 , \13858 , \13875 );
and \U$13500 ( \13877 , \13842 , \13875 );
or \U$13501 ( \13878 , \13859 , \13876 , \13877 );
and \U$13502 ( \13879 , \13825 , \13878 );
and \U$13503 ( \13880 , \13773 , \13878 );
or \U$13504 ( \13881 , \13826 , \13879 , \13880 );
and \U$13505 ( \13882 , \13725 , \13881 );
xor \U$13506 ( \13883 , \13202 , \13206 );
xor \U$13507 ( \13884 , \13883 , \499 );
xor \U$13508 ( \13885 , \13421 , \13423 );
xor \U$13509 ( \13886 , \13885 , \13426 );
and \U$13510 ( \13887 , \13884 , \13886 );
xor \U$13511 ( \13888 , \13431 , \13433 );
xor \U$13512 ( \13889 , \13888 , \13436 );
and \U$13513 ( \13890 , \13886 , \13889 );
and \U$13514 ( \13891 , \13884 , \13889 );
or \U$13515 ( \13892 , \13887 , \13890 , \13891 );
and \U$13516 ( \13893 , \13881 , \13892 );
and \U$13517 ( \13894 , \13725 , \13892 );
or \U$13518 ( \13895 , \13882 , \13893 , \13894 );
xor \U$13519 ( \13896 , \13469 , \13485 );
xor \U$13520 ( \13897 , \13896 , \13502 );
xor \U$13521 ( \13898 , \13521 , \13537 );
xor \U$13522 ( \13899 , \13898 , \13554 );
and \U$13523 ( \13900 , \13897 , \13899 );
xor \U$13524 ( \13901 , \13442 , \13444 );
xor \U$13525 ( \13902 , \13901 , \13447 );
and \U$13526 ( \13903 , \13899 , \13902 );
and \U$13527 ( \13904 , \13897 , \13902 );
or \U$13528 ( \13905 , \13900 , \13903 , \13904 );
xor \U$13529 ( \13906 , \13181 , \13197 );
xor \U$13530 ( \13907 , \13906 , \13210 );
and \U$13531 ( \13908 , \13905 , \13907 );
xor \U$13532 ( \13909 , \13640 , \13642 );
xor \U$13533 ( \13910 , \13909 , \13645 );
and \U$13534 ( \13911 , \13907 , \13910 );
and \U$13535 ( \13912 , \13905 , \13910 );
or \U$13536 ( \13913 , \13908 , \13911 , \13912 );
and \U$13537 ( \13914 , \13895 , \13913 );
xor \U$13538 ( \13915 , \13429 , \13439 );
xor \U$13539 ( \13916 , \13915 , \13450 );
xor \U$13540 ( \13917 , \13505 , \13557 );
xor \U$13541 ( \13918 , \13917 , \13610 );
and \U$13542 ( \13919 , \13916 , \13918 );
xor \U$13543 ( \13920 , \13616 , \13618 );
xor \U$13544 ( \13921 , \13920 , \13621 );
and \U$13545 ( \13922 , \13918 , \13921 );
and \U$13546 ( \13923 , \13916 , \13921 );
or \U$13547 ( \13924 , \13919 , \13922 , \13923 );
and \U$13548 ( \13925 , \13913 , \13924 );
and \U$13549 ( \13926 , \13895 , \13924 );
or \U$13550 ( \13927 , \13914 , \13925 , \13926 );
xor \U$13551 ( \13928 , \13453 , \13613 );
xor \U$13552 ( \13929 , \13928 , \13624 );
xor \U$13553 ( \13930 , \13629 , \13631 );
xor \U$13554 ( \13931 , \13930 , \13634 );
and \U$13555 ( \13932 , \13929 , \13931 );
xor \U$13556 ( \13933 , \13648 , \13650 );
xor \U$13557 ( \13934 , \13933 , \13653 );
and \U$13558 ( \13935 , \13931 , \13934 );
and \U$13559 ( \13936 , \13929 , \13934 );
or \U$13560 ( \13937 , \13932 , \13935 , \13936 );
and \U$13561 ( \13938 , \13927 , \13937 );
xor \U$13562 ( \13939 , \13353 , \13363 );
xor \U$13563 ( \13940 , \13939 , \13366 );
and \U$13564 ( \13941 , \13937 , \13940 );
and \U$13565 ( \13942 , \13927 , \13940 );
or \U$13566 ( \13943 , \13938 , \13941 , \13942 );
xor \U$13567 ( \13944 , \13165 , \13321 );
xor \U$13568 ( \13945 , \13944 , \13340 );
xor \U$13569 ( \13946 , \13627 , \13637 );
xor \U$13570 ( \13947 , \13946 , \13656 );
and \U$13571 ( \13948 , \13945 , \13947 );
xor \U$13572 ( \13949 , \13661 , \13663 );
xor \U$13573 ( \13950 , \13949 , \13666 );
and \U$13574 ( \13951 , \13947 , \13950 );
and \U$13575 ( \13952 , \13945 , \13950 );
or \U$13576 ( \13953 , \13948 , \13951 , \13952 );
and \U$13577 ( \13954 , \13943 , \13953 );
xor \U$13578 ( \13955 , \13343 , \13369 );
xor \U$13579 ( \13956 , \13955 , \13380 );
and \U$13580 ( \13957 , \13953 , \13956 );
and \U$13581 ( \13958 , \13943 , \13956 );
or \U$13582 ( \13959 , \13954 , \13957 , \13958 );
xor \U$13583 ( \13960 , \13675 , \13677 );
xor \U$13584 ( \13961 , \13960 , \13680 );
and \U$13585 ( \13962 , \13959 , \13961 );
and \U$13586 ( \13963 , \13689 , \13962 );
xor \U$13587 ( \13964 , \13689 , \13962 );
xor \U$13588 ( \13965 , \13959 , \13961 );
xor \U$13589 ( \13966 , \13830 , \13834 );
xor \U$13590 ( \13967 , \13966 , \13839 );
xor \U$13591 ( \13968 , \13793 , \13797 );
xor \U$13592 ( \13969 , \13968 , \13802 );
and \U$13593 ( \13970 , \13967 , \13969 );
xor \U$13594 ( \13971 , \13810 , \13814 );
xor \U$13595 ( \13972 , \13971 , \13819 );
and \U$13596 ( \13973 , \13969 , \13972 );
and \U$13597 ( \13974 , \13967 , \13972 );
or \U$13598 ( \13975 , \13970 , \13973 , \13974 );
and \U$13599 ( \13976 , \10409 , \754 );
and \U$13600 ( \13977 , \10228 , \752 );
nor \U$13601 ( \13978 , \13976 , \13977 );
xnor \U$13602 ( \13979 , \13978 , \711 );
nand \U$13603 ( \13980 , \11029 , \639 );
xnor \U$13604 ( \13981 , \13980 , \592 );
and \U$13605 ( \13982 , \13979 , \13981 );
xor \U$13606 ( \13983 , \13777 , \13781 );
xor \U$13607 ( \13984 , \13983 , \13786 );
and \U$13608 ( \13985 , \13981 , \13984 );
and \U$13609 ( \13986 , \13979 , \13984 );
or \U$13610 ( \13987 , \13982 , \13985 , \13986 );
and \U$13611 ( \13988 , \13975 , \13987 );
xor \U$13612 ( \13989 , \13729 , \13733 );
xor \U$13613 ( \13990 , \13989 , \13738 );
xor \U$13614 ( \13991 , \13846 , \13850 );
xor \U$13615 ( \13992 , \13991 , \13855 );
and \U$13616 ( \13993 , \13990 , \13992 );
xor \U$13617 ( \13994 , \13863 , \13867 );
xor \U$13618 ( \13995 , \13994 , \13872 );
and \U$13619 ( \13996 , \13992 , \13995 );
and \U$13620 ( \13997 , \13990 , \13995 );
or \U$13621 ( \13998 , \13993 , \13996 , \13997 );
and \U$13622 ( \13999 , \13987 , \13998 );
and \U$13623 ( \14000 , \13975 , \13998 );
or \U$13624 ( \14001 , \13988 , \13999 , \14000 );
and \U$13625 ( \14002 , \9620 , \1058 );
and \U$13626 ( \14003 , \9612 , \1056 );
nor \U$13627 ( \14004 , \14002 , \14003 );
xnor \U$13628 ( \14005 , \14004 , \964 );
and \U$13629 ( \14006 , \10228 , \888 );
and \U$13630 ( \14007 , \10223 , \886 );
nor \U$13631 ( \14008 , \14006 , \14007 );
xnor \U$13632 ( \14009 , \14008 , \816 );
and \U$13633 ( \14010 , \14005 , \14009 );
and \U$13634 ( \14011 , \11029 , \754 );
and \U$13635 ( \14012 , \10409 , \752 );
nor \U$13636 ( \14013 , \14011 , \14012 );
xnor \U$13637 ( \14014 , \14013 , \711 );
and \U$13638 ( \14015 , \14009 , \14014 );
and \U$13639 ( \14016 , \14005 , \14014 );
or \U$13640 ( \14017 , \14010 , \14015 , \14016 );
and \U$13641 ( \14018 , \6219 , \2362 );
and \U$13642 ( \14019 , \6210 , \2360 );
nor \U$13643 ( \14020 , \14018 , \14019 );
xnor \U$13644 ( \14021 , \14020 , \2225 );
and \U$13645 ( \14022 , \6764 , \2156 );
and \U$13646 ( \14023 , \6562 , \2154 );
nor \U$13647 ( \14024 , \14022 , \14023 );
xnor \U$13648 ( \14025 , \14024 , \2004 );
and \U$13649 ( \14026 , \14021 , \14025 );
and \U$13650 ( \14027 , \7239 , \1888 );
and \U$13651 ( \14028 , \7067 , \1886 );
nor \U$13652 ( \14029 , \14027 , \14028 );
xnor \U$13653 ( \14030 , \14029 , \1732 );
and \U$13654 ( \14031 , \14025 , \14030 );
and \U$13655 ( \14032 , \14021 , \14030 );
or \U$13656 ( \14033 , \14026 , \14031 , \14032 );
and \U$13657 ( \14034 , \14017 , \14033 );
and \U$13658 ( \14035 , \8189 , \1616 );
and \U$13659 ( \14036 , \7765 , \1614 );
nor \U$13660 ( \14037 , \14035 , \14036 );
xnor \U$13661 ( \14038 , \14037 , \1503 );
and \U$13662 ( \14039 , \8440 , \1422 );
and \U$13663 ( \14040 , \8435 , \1420 );
nor \U$13664 ( \14041 , \14039 , \14040 );
xnor \U$13665 ( \14042 , \14041 , \1286 );
and \U$13666 ( \14043 , \14038 , \14042 );
and \U$13667 ( \14044 , \9043 , \1222 );
and \U$13668 ( \14045 , \8759 , \1220 );
nor \U$13669 ( \14046 , \14044 , \14045 );
xnor \U$13670 ( \14047 , \14046 , \1144 );
and \U$13671 ( \14048 , \14042 , \14047 );
and \U$13672 ( \14049 , \14038 , \14047 );
or \U$13673 ( \14050 , \14043 , \14048 , \14049 );
and \U$13674 ( \14051 , \14033 , \14050 );
and \U$13675 ( \14052 , \14017 , \14050 );
or \U$13676 ( \14053 , \14034 , \14051 , \14052 );
and \U$13677 ( \14054 , \1336 , \8958 );
and \U$13678 ( \14055 , \1248 , \8956 );
nor \U$13679 ( \14056 , \14054 , \14055 );
xnor \U$13680 ( \14057 , \14056 , \8587 );
and \U$13681 ( \14058 , \1446 , \8396 );
and \U$13682 ( \14059 , \1441 , \8394 );
nor \U$13683 ( \14060 , \14058 , \14059 );
xnor \U$13684 ( \14061 , \14060 , \8078 );
and \U$13685 ( \14062 , \14057 , \14061 );
and \U$13686 ( \14063 , \1677 , \7829 );
and \U$13687 ( \14064 , \1562 , \7827 );
nor \U$13688 ( \14065 , \14063 , \14064 );
xnor \U$13689 ( \14066 , \14065 , \7580 );
and \U$13690 ( \14067 , \14061 , \14066 );
and \U$13691 ( \14068 , \14057 , \14066 );
or \U$13692 ( \14069 , \14062 , \14067 , \14068 );
and \U$13693 ( \14070 , \1861 , \7300 );
and \U$13694 ( \14071 , \1853 , \7298 );
nor \U$13695 ( \14072 , \14070 , \14071 );
xnor \U$13696 ( \14073 , \14072 , \7040 );
and \U$13697 ( \14074 , \2109 , \6806 );
and \U$13698 ( \14075 , \2104 , \6804 );
nor \U$13699 ( \14076 , \14074 , \14075 );
xnor \U$13700 ( \14077 , \14076 , \6491 );
and \U$13701 ( \14078 , \14073 , \14077 );
and \U$13702 ( \14079 , \2439 , \6297 );
and \U$13703 ( \14080 , \2295 , \6295 );
nor \U$13704 ( \14081 , \14079 , \14080 );
xnor \U$13705 ( \14082 , \14081 , \5957 );
and \U$13706 ( \14083 , \14077 , \14082 );
and \U$13707 ( \14084 , \14073 , \14082 );
or \U$13708 ( \14085 , \14078 , \14083 , \14084 );
and \U$13709 ( \14086 , \14069 , \14085 );
and \U$13710 ( \14087 , \771 , \10876 );
and \U$13711 ( \14088 , \743 , \10873 );
nor \U$13712 ( \14089 , \14087 , \14088 );
xnor \U$13713 ( \14090 , \14089 , \9821 );
and \U$13714 ( \14091 , \925 , \10063 );
and \U$13715 ( \14092 , \851 , \10061 );
nor \U$13716 ( \14093 , \14091 , \14092 );
xnor \U$13717 ( \14094 , \14093 , \9824 );
and \U$13718 ( \14095 , \14090 , \14094 );
and \U$13719 ( \14096 , \1050 , \9495 );
and \U$13720 ( \14097 , \987 , \9493 );
nor \U$13721 ( \14098 , \14096 , \14097 );
xnor \U$13722 ( \14099 , \14098 , \9185 );
and \U$13723 ( \14100 , \14094 , \14099 );
and \U$13724 ( \14101 , \14090 , \14099 );
or \U$13725 ( \14102 , \14095 , \14100 , \14101 );
and \U$13726 ( \14103 , \14085 , \14102 );
and \U$13727 ( \14104 , \14069 , \14102 );
or \U$13728 ( \14105 , \14086 , \14103 , \14104 );
and \U$13729 ( \14106 , \14053 , \14105 );
and \U$13730 ( \14107 , \4841 , \3386 );
and \U$13731 ( \14108 , \4833 , \3384 );
nor \U$13732 ( \14109 , \14107 , \14108 );
xnor \U$13733 ( \14110 , \14109 , \3181 );
and \U$13734 ( \14111 , \5315 , \2980 );
and \U$13735 ( \14112 , \5310 , \2978 );
nor \U$13736 ( \14113 , \14111 , \14112 );
xnor \U$13737 ( \14114 , \14113 , \2831 );
and \U$13738 ( \14115 , \14110 , \14114 );
and \U$13739 ( \14116 , \5838 , \2658 );
and \U$13740 ( \14117 , \5579 , \2656 );
nor \U$13741 ( \14118 , \14116 , \14117 );
xnor \U$13742 ( \14119 , \14118 , \2516 );
and \U$13743 ( \14120 , \14114 , \14119 );
and \U$13744 ( \14121 , \14110 , \14119 );
or \U$13745 ( \14122 , \14115 , \14120 , \14121 );
and \U$13746 ( \14123 , \3951 , \4417 );
and \U$13747 ( \14124 , \3743 , \4415 );
nor \U$13748 ( \14125 , \14123 , \14124 );
xnor \U$13749 ( \14126 , \14125 , \4274 );
and \U$13750 ( \14127 , \4078 , \4094 );
and \U$13751 ( \14128 , \4073 , \4092 );
nor \U$13752 ( \14129 , \14127 , \14128 );
xnor \U$13753 ( \14130 , \14129 , \3848 );
and \U$13754 ( \14131 , \14126 , \14130 );
and \U$13755 ( \14132 , \4531 , \3699 );
and \U$13756 ( \14133 , \4334 , \3697 );
nor \U$13757 ( \14134 , \14132 , \14133 );
xnor \U$13758 ( \14135 , \14134 , \3512 );
and \U$13759 ( \14136 , \14130 , \14135 );
and \U$13760 ( \14137 , \14126 , \14135 );
or \U$13761 ( \14138 , \14131 , \14136 , \14137 );
and \U$13762 ( \14139 , \14122 , \14138 );
and \U$13763 ( \14140 , \2728 , \5708 );
and \U$13764 ( \14141 , \2703 , \5706 );
nor \U$13765 ( \14142 , \14140 , \14141 );
xnor \U$13766 ( \14143 , \14142 , \5467 );
and \U$13767 ( \14144 , \3069 , \5242 );
and \U$13768 ( \14145 , \2902 , \5240 );
nor \U$13769 ( \14146 , \14144 , \14145 );
xnor \U$13770 ( \14147 , \14146 , \5054 );
and \U$13771 ( \14148 , \14143 , \14147 );
and \U$13772 ( \14149 , \3326 , \4868 );
and \U$13773 ( \14150 , \3207 , \4866 );
nor \U$13774 ( \14151 , \14149 , \14150 );
xnor \U$13775 ( \14152 , \14151 , \4636 );
and \U$13776 ( \14153 , \14147 , \14152 );
and \U$13777 ( \14154 , \14143 , \14152 );
or \U$13778 ( \14155 , \14148 , \14153 , \14154 );
and \U$13779 ( \14156 , \14138 , \14155 );
and \U$13780 ( \14157 , \14122 , \14155 );
or \U$13781 ( \14158 , \14139 , \14156 , \14157 );
and \U$13782 ( \14159 , \14105 , \14158 );
and \U$13783 ( \14160 , \14053 , \14158 );
or \U$13784 ( \14161 , \14106 , \14159 , \14160 );
and \U$13785 ( \14162 , \14001 , \14161 );
xor \U$13786 ( \14163 , \13578 , \13582 );
xor \U$13787 ( \14164 , \14163 , \13587 );
xor \U$13788 ( \14165 , \13691 , \13693 );
xor \U$13789 ( \14166 , \14165 , \13696 );
and \U$13790 ( \14167 , \14164 , \14166 );
xor \U$13791 ( \14168 , \13701 , \13703 );
xor \U$13792 ( \14169 , \14168 , \13706 );
and \U$13793 ( \14170 , \14166 , \14169 );
and \U$13794 ( \14171 , \14164 , \14169 );
or \U$13795 ( \14172 , \14167 , \14170 , \14171 );
and \U$13796 ( \14173 , \14161 , \14172 );
and \U$13797 ( \14174 , \14001 , \14172 );
or \U$13798 ( \14175 , \14162 , \14173 , \14174 );
xor \U$13799 ( \14176 , \13789 , \13805 );
xor \U$13800 ( \14177 , \14176 , \13822 );
xor \U$13801 ( \14178 , \13842 , \13858 );
xor \U$13802 ( \14179 , \14178 , \13875 );
and \U$13803 ( \14180 , \14177 , \14179 );
xor \U$13804 ( \14181 , \13714 , \13716 );
xor \U$13805 ( \14182 , \14181 , \13719 );
and \U$13806 ( \14183 , \14179 , \14182 );
and \U$13807 ( \14184 , \14177 , \14182 );
or \U$13808 ( \14185 , \14180 , \14183 , \14184 );
xor \U$13809 ( \14186 , \13574 , \13590 );
xor \U$13810 ( \14187 , \14186 , \13607 );
and \U$13811 ( \14188 , \14185 , \14187 );
xor \U$13812 ( \14189 , \13897 , \13899 );
xor \U$13813 ( \14190 , \14189 , \13902 );
and \U$13814 ( \14191 , \14187 , \14190 );
and \U$13815 ( \14192 , \14185 , \14190 );
or \U$13816 ( \14193 , \14188 , \14191 , \14192 );
and \U$13817 ( \14194 , \14175 , \14193 );
xor \U$13818 ( \14195 , \13699 , \13709 );
xor \U$13819 ( \14196 , \14195 , \13722 );
xor \U$13820 ( \14197 , \13773 , \13825 );
xor \U$13821 ( \14198 , \14197 , \13878 );
and \U$13822 ( \14199 , \14196 , \14198 );
xor \U$13823 ( \14200 , \13884 , \13886 );
xor \U$13824 ( \14201 , \14200 , \13889 );
and \U$13825 ( \14202 , \14198 , \14201 );
and \U$13826 ( \14203 , \14196 , \14201 );
or \U$13827 ( \14204 , \14199 , \14202 , \14203 );
and \U$13828 ( \14205 , \14193 , \14204 );
and \U$13829 ( \14206 , \14175 , \14204 );
or \U$13830 ( \14207 , \14194 , \14205 , \14206 );
xor \U$13831 ( \14208 , \13725 , \13881 );
xor \U$13832 ( \14209 , \14208 , \13892 );
xor \U$13833 ( \14210 , \13905 , \13907 );
xor \U$13834 ( \14211 , \14210 , \13910 );
and \U$13835 ( \14212 , \14209 , \14211 );
xor \U$13836 ( \14213 , \13916 , \13918 );
xor \U$13837 ( \14214 , \14213 , \13921 );
and \U$13838 ( \14215 , \14211 , \14214 );
and \U$13839 ( \14216 , \14209 , \14214 );
or \U$13840 ( \14217 , \14212 , \14215 , \14216 );
and \U$13841 ( \14218 , \14207 , \14217 );
xor \U$13842 ( \14219 , \13929 , \13931 );
xor \U$13843 ( \14220 , \14219 , \13934 );
and \U$13844 ( \14221 , \14217 , \14220 );
and \U$13845 ( \14222 , \14207 , \14220 );
or \U$13846 ( \14223 , \14218 , \14221 , \14222 );
xor \U$13847 ( \14224 , \13927 , \13937 );
xor \U$13848 ( \14225 , \14224 , \13940 );
and \U$13849 ( \14226 , \14223 , \14225 );
xor \U$13850 ( \14227 , \13945 , \13947 );
xor \U$13851 ( \14228 , \14227 , \13950 );
and \U$13852 ( \14229 , \14225 , \14228 );
and \U$13853 ( \14230 , \14223 , \14228 );
or \U$13854 ( \14231 , \14226 , \14229 , \14230 );
xor \U$13855 ( \14232 , \13943 , \13953 );
xor \U$13856 ( \14233 , \14232 , \13956 );
and \U$13857 ( \14234 , \14231 , \14233 );
xor \U$13858 ( \14235 , \13659 , \13669 );
xor \U$13859 ( \14236 , \14235 , \13672 );
and \U$13860 ( \14237 , \14233 , \14236 );
and \U$13861 ( \14238 , \14231 , \14236 );
or \U$13862 ( \14239 , \14234 , \14237 , \14238 );
and \U$13863 ( \14240 , \13965 , \14239 );
xor \U$13864 ( \14241 , \13965 , \14239 );
xor \U$13865 ( \14242 , \14231 , \14233 );
xor \U$13866 ( \14243 , \14242 , \14236 );
xor \U$13867 ( \14244 , \14110 , \14114 );
xor \U$13868 ( \14245 , \14244 , \14119 );
xor \U$13869 ( \14246 , \14126 , \14130 );
xor \U$13870 ( \14247 , \14246 , \14135 );
and \U$13871 ( \14248 , \14245 , \14247 );
xor \U$13872 ( \14249 , \14143 , \14147 );
xor \U$13873 ( \14250 , \14249 , \14152 );
and \U$13874 ( \14251 , \14247 , \14250 );
and \U$13875 ( \14252 , \14245 , \14250 );
or \U$13876 ( \14253 , \14248 , \14251 , \14252 );
xor \U$13877 ( \14254 , \14005 , \14009 );
xor \U$13878 ( \14255 , \14254 , \14014 );
xor \U$13879 ( \14256 , \14021 , \14025 );
xor \U$13880 ( \14257 , \14256 , \14030 );
and \U$13881 ( \14258 , \14255 , \14257 );
xor \U$13882 ( \14259 , \14038 , \14042 );
xor \U$13883 ( \14260 , \14259 , \14047 );
and \U$13884 ( \14261 , \14257 , \14260 );
and \U$13885 ( \14262 , \14255 , \14260 );
or \U$13886 ( \14263 , \14258 , \14261 , \14262 );
and \U$13887 ( \14264 , \14253 , \14263 );
xor \U$13888 ( \14265 , \14057 , \14061 );
xor \U$13889 ( \14266 , \14265 , \14066 );
xor \U$13890 ( \14267 , \14073 , \14077 );
xor \U$13891 ( \14268 , \14267 , \14082 );
and \U$13892 ( \14269 , \14266 , \14268 );
xor \U$13893 ( \14270 , \14090 , \14094 );
xor \U$13894 ( \14271 , \14270 , \14099 );
and \U$13895 ( \14272 , \14268 , \14271 );
and \U$13896 ( \14273 , \14266 , \14271 );
or \U$13897 ( \14274 , \14269 , \14272 , \14273 );
and \U$13898 ( \14275 , \14263 , \14274 );
and \U$13899 ( \14276 , \14253 , \14274 );
or \U$13900 ( \14277 , \14264 , \14275 , \14276 );
and \U$13901 ( \14278 , \4833 , \3699 );
and \U$13902 ( \14279 , \4531 , \3697 );
nor \U$13903 ( \14280 , \14278 , \14279 );
xnor \U$13904 ( \14281 , \14280 , \3512 );
and \U$13905 ( \14282 , \5310 , \3386 );
and \U$13906 ( \14283 , \4841 , \3384 );
nor \U$13907 ( \14284 , \14282 , \14283 );
xnor \U$13908 ( \14285 , \14284 , \3181 );
and \U$13909 ( \14286 , \14281 , \14285 );
and \U$13910 ( \14287 , \5579 , \2980 );
and \U$13911 ( \14288 , \5315 , \2978 );
nor \U$13912 ( \14289 , \14287 , \14288 );
xnor \U$13913 ( \14290 , \14289 , \2831 );
and \U$13914 ( \14291 , \14285 , \14290 );
and \U$13915 ( \14292 , \14281 , \14290 );
or \U$13916 ( \14293 , \14286 , \14291 , \14292 );
and \U$13917 ( \14294 , \2703 , \6297 );
and \U$13918 ( \14295 , \2439 , \6295 );
nor \U$13919 ( \14296 , \14294 , \14295 );
xnor \U$13920 ( \14297 , \14296 , \5957 );
and \U$13921 ( \14298 , \2902 , \5708 );
and \U$13922 ( \14299 , \2728 , \5706 );
nor \U$13923 ( \14300 , \14298 , \14299 );
xnor \U$13924 ( \14301 , \14300 , \5467 );
and \U$13925 ( \14302 , \14297 , \14301 );
and \U$13926 ( \14303 , \3207 , \5242 );
and \U$13927 ( \14304 , \3069 , \5240 );
nor \U$13928 ( \14305 , \14303 , \14304 );
xnor \U$13929 ( \14306 , \14305 , \5054 );
and \U$13930 ( \14307 , \14301 , \14306 );
and \U$13931 ( \14308 , \14297 , \14306 );
or \U$13932 ( \14309 , \14302 , \14307 , \14308 );
and \U$13933 ( \14310 , \14293 , \14309 );
and \U$13934 ( \14311 , \3743 , \4868 );
and \U$13935 ( \14312 , \3326 , \4866 );
nor \U$13936 ( \14313 , \14311 , \14312 );
xnor \U$13937 ( \14314 , \14313 , \4636 );
and \U$13938 ( \14315 , \4073 , \4417 );
and \U$13939 ( \14316 , \3951 , \4415 );
nor \U$13940 ( \14317 , \14315 , \14316 );
xnor \U$13941 ( \14318 , \14317 , \4274 );
and \U$13942 ( \14319 , \14314 , \14318 );
and \U$13943 ( \14320 , \4334 , \4094 );
and \U$13944 ( \14321 , \4078 , \4092 );
nor \U$13945 ( \14322 , \14320 , \14321 );
xnor \U$13946 ( \14323 , \14322 , \3848 );
and \U$13947 ( \14324 , \14318 , \14323 );
and \U$13948 ( \14325 , \14314 , \14323 );
or \U$13949 ( \14326 , \14319 , \14324 , \14325 );
and \U$13950 ( \14327 , \14309 , \14326 );
and \U$13951 ( \14328 , \14293 , \14326 );
or \U$13952 ( \14329 , \14310 , \14327 , \14328 );
and \U$13953 ( \14330 , \1248 , \9495 );
and \U$13954 ( \14331 , \1050 , \9493 );
nor \U$13955 ( \14332 , \14330 , \14331 );
xnor \U$13956 ( \14333 , \14332 , \9185 );
and \U$13957 ( \14334 , \1441 , \8958 );
and \U$13958 ( \14335 , \1336 , \8956 );
nor \U$13959 ( \14336 , \14334 , \14335 );
xnor \U$13960 ( \14337 , \14336 , \8587 );
and \U$13961 ( \14338 , \14333 , \14337 );
and \U$13962 ( \14339 , \1562 , \8396 );
and \U$13963 ( \14340 , \1446 , \8394 );
nor \U$13964 ( \14341 , \14339 , \14340 );
xnor \U$13965 ( \14342 , \14341 , \8078 );
and \U$13966 ( \14343 , \14337 , \14342 );
and \U$13967 ( \14344 , \14333 , \14342 );
or \U$13968 ( \14345 , \14338 , \14343 , \14344 );
and \U$13969 ( \14346 , \851 , \10876 );
and \U$13970 ( \14347 , \771 , \10873 );
nor \U$13971 ( \14348 , \14346 , \14347 );
xnor \U$13972 ( \14349 , \14348 , \9821 );
and \U$13973 ( \14350 , \987 , \10063 );
and \U$13974 ( \14351 , \925 , \10061 );
nor \U$13975 ( \14352 , \14350 , \14351 );
xnor \U$13976 ( \14353 , \14352 , \9824 );
and \U$13977 ( \14354 , \14349 , \14353 );
and \U$13978 ( \14355 , \14353 , \711 );
and \U$13979 ( \14356 , \14349 , \711 );
or \U$13980 ( \14357 , \14354 , \14355 , \14356 );
and \U$13981 ( \14358 , \14345 , \14357 );
and \U$13982 ( \14359 , \1853 , \7829 );
and \U$13983 ( \14360 , \1677 , \7827 );
nor \U$13984 ( \14361 , \14359 , \14360 );
xnor \U$13985 ( \14362 , \14361 , \7580 );
and \U$13986 ( \14363 , \2104 , \7300 );
and \U$13987 ( \14364 , \1861 , \7298 );
nor \U$13988 ( \14365 , \14363 , \14364 );
xnor \U$13989 ( \14366 , \14365 , \7040 );
and \U$13990 ( \14367 , \14362 , \14366 );
and \U$13991 ( \14368 , \2295 , \6806 );
and \U$13992 ( \14369 , \2109 , \6804 );
nor \U$13993 ( \14370 , \14368 , \14369 );
xnor \U$13994 ( \14371 , \14370 , \6491 );
and \U$13995 ( \14372 , \14366 , \14371 );
and \U$13996 ( \14373 , \14362 , \14371 );
or \U$13997 ( \14374 , \14367 , \14372 , \14373 );
and \U$13998 ( \14375 , \14357 , \14374 );
and \U$13999 ( \14376 , \14345 , \14374 );
or \U$14000 ( \14377 , \14358 , \14375 , \14376 );
and \U$14001 ( \14378 , \14329 , \14377 );
and \U$14002 ( \14379 , \9612 , \1222 );
and \U$14003 ( \14380 , \9043 , \1220 );
nor \U$14004 ( \14381 , \14379 , \14380 );
xnor \U$14005 ( \14382 , \14381 , \1144 );
and \U$14006 ( \14383 , \10223 , \1058 );
and \U$14007 ( \14384 , \9620 , \1056 );
nor \U$14008 ( \14385 , \14383 , \14384 );
xnor \U$14009 ( \14386 , \14385 , \964 );
and \U$14010 ( \14387 , \14382 , \14386 );
and \U$14011 ( \14388 , \10409 , \888 );
and \U$14012 ( \14389 , \10228 , \886 );
nor \U$14013 ( \14390 , \14388 , \14389 );
xnor \U$14014 ( \14391 , \14390 , \816 );
and \U$14015 ( \14392 , \14386 , \14391 );
and \U$14016 ( \14393 , \14382 , \14391 );
or \U$14017 ( \14394 , \14387 , \14392 , \14393 );
and \U$14018 ( \14395 , \6210 , \2658 );
and \U$14019 ( \14396 , \5838 , \2656 );
nor \U$14020 ( \14397 , \14395 , \14396 );
xnor \U$14021 ( \14398 , \14397 , \2516 );
and \U$14022 ( \14399 , \6562 , \2362 );
and \U$14023 ( \14400 , \6219 , \2360 );
nor \U$14024 ( \14401 , \14399 , \14400 );
xnor \U$14025 ( \14402 , \14401 , \2225 );
and \U$14026 ( \14403 , \14398 , \14402 );
and \U$14027 ( \14404 , \7067 , \2156 );
and \U$14028 ( \14405 , \6764 , \2154 );
nor \U$14029 ( \14406 , \14404 , \14405 );
xnor \U$14030 ( \14407 , \14406 , \2004 );
and \U$14031 ( \14408 , \14402 , \14407 );
and \U$14032 ( \14409 , \14398 , \14407 );
or \U$14033 ( \14410 , \14403 , \14408 , \14409 );
and \U$14034 ( \14411 , \14394 , \14410 );
and \U$14035 ( \14412 , \7765 , \1888 );
and \U$14036 ( \14413 , \7239 , \1886 );
nor \U$14037 ( \14414 , \14412 , \14413 );
xnor \U$14038 ( \14415 , \14414 , \1732 );
and \U$14039 ( \14416 , \8435 , \1616 );
and \U$14040 ( \14417 , \8189 , \1614 );
nor \U$14041 ( \14418 , \14416 , \14417 );
xnor \U$14042 ( \14419 , \14418 , \1503 );
and \U$14043 ( \14420 , \14415 , \14419 );
and \U$14044 ( \14421 , \8759 , \1422 );
and \U$14045 ( \14422 , \8440 , \1420 );
nor \U$14046 ( \14423 , \14421 , \14422 );
xnor \U$14047 ( \14424 , \14423 , \1286 );
and \U$14048 ( \14425 , \14419 , \14424 );
and \U$14049 ( \14426 , \14415 , \14424 );
or \U$14050 ( \14427 , \14420 , \14425 , \14426 );
and \U$14051 ( \14428 , \14410 , \14427 );
and \U$14052 ( \14429 , \14394 , \14427 );
or \U$14053 ( \14430 , \14411 , \14428 , \14429 );
and \U$14054 ( \14431 , \14377 , \14430 );
and \U$14055 ( \14432 , \14329 , \14430 );
or \U$14056 ( \14433 , \14378 , \14431 , \14432 );
and \U$14057 ( \14434 , \14277 , \14433 );
xor \U$14058 ( \14435 , \13745 , \13749 );
xor \U$14059 ( \14436 , \14435 , \13754 );
xor \U$14060 ( \14437 , \13762 , \13766 );
xor \U$14061 ( \14438 , \14437 , \592 );
and \U$14062 ( \14439 , \14436 , \14438 );
xor \U$14063 ( \14440 , \13990 , \13992 );
xor \U$14064 ( \14441 , \14440 , \13995 );
and \U$14065 ( \14442 , \14438 , \14441 );
and \U$14066 ( \14443 , \14436 , \14441 );
or \U$14067 ( \14444 , \14439 , \14442 , \14443 );
and \U$14068 ( \14445 , \14433 , \14444 );
and \U$14069 ( \14446 , \14277 , \14444 );
or \U$14070 ( \14447 , \14434 , \14445 , \14446 );
xor \U$14071 ( \14448 , \14017 , \14033 );
xor \U$14072 ( \14449 , \14448 , \14050 );
xor \U$14073 ( \14450 , \13967 , \13969 );
xor \U$14074 ( \14451 , \14450 , \13972 );
and \U$14075 ( \14452 , \14449 , \14451 );
xor \U$14076 ( \14453 , \13979 , \13981 );
xor \U$14077 ( \14454 , \14453 , \13984 );
and \U$14078 ( \14455 , \14451 , \14454 );
and \U$14079 ( \14456 , \14449 , \14454 );
or \U$14080 ( \14457 , \14452 , \14455 , \14456 );
xor \U$14081 ( \14458 , \14069 , \14085 );
xor \U$14082 ( \14459 , \14458 , \14102 );
xor \U$14083 ( \14460 , \14122 , \14138 );
xor \U$14084 ( \14461 , \14460 , \14155 );
and \U$14085 ( \14462 , \14459 , \14461 );
and \U$14086 ( \14463 , \14457 , \14462 );
xor \U$14087 ( \14464 , \13741 , \13757 );
xor \U$14088 ( \14465 , \14464 , \13770 );
and \U$14089 ( \14466 , \14462 , \14465 );
and \U$14090 ( \14467 , \14457 , \14465 );
or \U$14091 ( \14468 , \14463 , \14466 , \14467 );
and \U$14092 ( \14469 , \14447 , \14468 );
xor \U$14093 ( \14470 , \13975 , \13987 );
xor \U$14094 ( \14471 , \14470 , \13998 );
xor \U$14095 ( \14472 , \14177 , \14179 );
xor \U$14096 ( \14473 , \14472 , \14182 );
and \U$14097 ( \14474 , \14471 , \14473 );
xor \U$14098 ( \14475 , \14164 , \14166 );
xor \U$14099 ( \14476 , \14475 , \14169 );
and \U$14100 ( \14477 , \14473 , \14476 );
and \U$14101 ( \14478 , \14471 , \14476 );
or \U$14102 ( \14479 , \14474 , \14477 , \14478 );
and \U$14103 ( \14480 , \14468 , \14479 );
and \U$14104 ( \14481 , \14447 , \14479 );
or \U$14105 ( \14482 , \14469 , \14480 , \14481 );
xor \U$14106 ( \14483 , \14001 , \14161 );
xor \U$14107 ( \14484 , \14483 , \14172 );
xor \U$14108 ( \14485 , \14185 , \14187 );
xor \U$14109 ( \14486 , \14485 , \14190 );
and \U$14110 ( \14487 , \14484 , \14486 );
xor \U$14111 ( \14488 , \14196 , \14198 );
xor \U$14112 ( \14489 , \14488 , \14201 );
and \U$14113 ( \14490 , \14486 , \14489 );
and \U$14114 ( \14491 , \14484 , \14489 );
or \U$14115 ( \14492 , \14487 , \14490 , \14491 );
and \U$14116 ( \14493 , \14482 , \14492 );
xor \U$14117 ( \14494 , \14209 , \14211 );
xor \U$14118 ( \14495 , \14494 , \14214 );
and \U$14119 ( \14496 , \14492 , \14495 );
and \U$14120 ( \14497 , \14482 , \14495 );
or \U$14121 ( \14498 , \14493 , \14496 , \14497 );
xor \U$14122 ( \14499 , \13895 , \13913 );
xor \U$14123 ( \14500 , \14499 , \13924 );
and \U$14124 ( \14501 , \14498 , \14500 );
xor \U$14125 ( \14502 , \14207 , \14217 );
xor \U$14126 ( \14503 , \14502 , \14220 );
and \U$14127 ( \14504 , \14500 , \14503 );
and \U$14128 ( \14505 , \14498 , \14503 );
or \U$14129 ( \14506 , \14501 , \14504 , \14505 );
xor \U$14130 ( \14507 , \14223 , \14225 );
xor \U$14131 ( \14508 , \14507 , \14228 );
and \U$14132 ( \14509 , \14506 , \14508 );
and \U$14133 ( \14510 , \14243 , \14509 );
xor \U$14134 ( \14511 , \14243 , \14509 );
xor \U$14135 ( \14512 , \14506 , \14508 );
and \U$14136 ( \14513 , \4078 , \4417 );
and \U$14137 ( \14514 , \4073 , \4415 );
nor \U$14138 ( \14515 , \14513 , \14514 );
xnor \U$14139 ( \14516 , \14515 , \4274 );
and \U$14140 ( \14517 , \4531 , \4094 );
and \U$14141 ( \14518 , \4334 , \4092 );
nor \U$14142 ( \14519 , \14517 , \14518 );
xnor \U$14143 ( \14520 , \14519 , \3848 );
and \U$14144 ( \14521 , \14516 , \14520 );
and \U$14145 ( \14522 , \4841 , \3699 );
and \U$14146 ( \14523 , \4833 , \3697 );
nor \U$14147 ( \14524 , \14522 , \14523 );
xnor \U$14148 ( \14525 , \14524 , \3512 );
and \U$14149 ( \14526 , \14520 , \14525 );
and \U$14150 ( \14527 , \14516 , \14525 );
or \U$14151 ( \14528 , \14521 , \14526 , \14527 );
and \U$14152 ( \14529 , \3069 , \5708 );
and \U$14153 ( \14530 , \2902 , \5706 );
nor \U$14154 ( \14531 , \14529 , \14530 );
xnor \U$14155 ( \14532 , \14531 , \5467 );
and \U$14156 ( \14533 , \3326 , \5242 );
and \U$14157 ( \14534 , \3207 , \5240 );
nor \U$14158 ( \14535 , \14533 , \14534 );
xnor \U$14159 ( \14536 , \14535 , \5054 );
and \U$14160 ( \14537 , \14532 , \14536 );
and \U$14161 ( \14538 , \3951 , \4868 );
and \U$14162 ( \14539 , \3743 , \4866 );
nor \U$14163 ( \14540 , \14538 , \14539 );
xnor \U$14164 ( \14541 , \14540 , \4636 );
and \U$14165 ( \14542 , \14536 , \14541 );
and \U$14166 ( \14543 , \14532 , \14541 );
or \U$14167 ( \14544 , \14537 , \14542 , \14543 );
and \U$14168 ( \14545 , \14528 , \14544 );
and \U$14169 ( \14546 , \5315 , \3386 );
and \U$14170 ( \14547 , \5310 , \3384 );
nor \U$14171 ( \14548 , \14546 , \14547 );
xnor \U$14172 ( \14549 , \14548 , \3181 );
and \U$14173 ( \14550 , \5838 , \2980 );
and \U$14174 ( \14551 , \5579 , \2978 );
nor \U$14175 ( \14552 , \14550 , \14551 );
xnor \U$14176 ( \14553 , \14552 , \2831 );
and \U$14177 ( \14554 , \14549 , \14553 );
and \U$14178 ( \14555 , \6219 , \2658 );
and \U$14179 ( \14556 , \6210 , \2656 );
nor \U$14180 ( \14557 , \14555 , \14556 );
xnor \U$14181 ( \14558 , \14557 , \2516 );
and \U$14182 ( \14559 , \14553 , \14558 );
and \U$14183 ( \14560 , \14549 , \14558 );
or \U$14184 ( \14561 , \14554 , \14559 , \14560 );
and \U$14185 ( \14562 , \14544 , \14561 );
and \U$14186 ( \14563 , \14528 , \14561 );
or \U$14187 ( \14564 , \14545 , \14562 , \14563 );
and \U$14188 ( \14565 , \8440 , \1616 );
and \U$14189 ( \14566 , \8435 , \1614 );
nor \U$14190 ( \14567 , \14565 , \14566 );
xnor \U$14191 ( \14568 , \14567 , \1503 );
and \U$14192 ( \14569 , \9043 , \1422 );
and \U$14193 ( \14570 , \8759 , \1420 );
nor \U$14194 ( \14571 , \14569 , \14570 );
xnor \U$14195 ( \14572 , \14571 , \1286 );
and \U$14196 ( \14573 , \14568 , \14572 );
and \U$14197 ( \14574 , \9620 , \1222 );
and \U$14198 ( \14575 , \9612 , \1220 );
nor \U$14199 ( \14576 , \14574 , \14575 );
xnor \U$14200 ( \14577 , \14576 , \1144 );
and \U$14201 ( \14578 , \14572 , \14577 );
and \U$14202 ( \14579 , \14568 , \14577 );
or \U$14203 ( \14580 , \14573 , \14578 , \14579 );
and \U$14204 ( \14581 , \6764 , \2362 );
and \U$14205 ( \14582 , \6562 , \2360 );
nor \U$14206 ( \14583 , \14581 , \14582 );
xnor \U$14207 ( \14584 , \14583 , \2225 );
and \U$14208 ( \14585 , \7239 , \2156 );
and \U$14209 ( \14586 , \7067 , \2154 );
nor \U$14210 ( \14587 , \14585 , \14586 );
xnor \U$14211 ( \14588 , \14587 , \2004 );
and \U$14212 ( \14589 , \14584 , \14588 );
and \U$14213 ( \14590 , \8189 , \1888 );
and \U$14214 ( \14591 , \7765 , \1886 );
nor \U$14215 ( \14592 , \14590 , \14591 );
xnor \U$14216 ( \14593 , \14592 , \1732 );
and \U$14217 ( \14594 , \14588 , \14593 );
and \U$14218 ( \14595 , \14584 , \14593 );
or \U$14219 ( \14596 , \14589 , \14594 , \14595 );
and \U$14220 ( \14597 , \14580 , \14596 );
and \U$14221 ( \14598 , \10228 , \1058 );
and \U$14222 ( \14599 , \10223 , \1056 );
nor \U$14223 ( \14600 , \14598 , \14599 );
xnor \U$14224 ( \14601 , \14600 , \964 );
and \U$14225 ( \14602 , \11029 , \888 );
and \U$14226 ( \14603 , \10409 , \886 );
nor \U$14227 ( \14604 , \14602 , \14603 );
xnor \U$14228 ( \14605 , \14604 , \816 );
and \U$14229 ( \14606 , \14601 , \14605 );
and \U$14230 ( \14607 , \14596 , \14606 );
and \U$14231 ( \14608 , \14580 , \14606 );
or \U$14232 ( \14609 , \14597 , \14607 , \14608 );
and \U$14233 ( \14610 , \14564 , \14609 );
and \U$14234 ( \14611 , \2109 , \7300 );
and \U$14235 ( \14612 , \2104 , \7298 );
nor \U$14236 ( \14613 , \14611 , \14612 );
xnor \U$14237 ( \14614 , \14613 , \7040 );
and \U$14238 ( \14615 , \2439 , \6806 );
and \U$14239 ( \14616 , \2295 , \6804 );
nor \U$14240 ( \14617 , \14615 , \14616 );
xnor \U$14241 ( \14618 , \14617 , \6491 );
and \U$14242 ( \14619 , \14614 , \14618 );
and \U$14243 ( \14620 , \2728 , \6297 );
and \U$14244 ( \14621 , \2703 , \6295 );
nor \U$14245 ( \14622 , \14620 , \14621 );
xnor \U$14246 ( \14623 , \14622 , \5957 );
and \U$14247 ( \14624 , \14618 , \14623 );
and \U$14248 ( \14625 , \14614 , \14623 );
or \U$14249 ( \14626 , \14619 , \14624 , \14625 );
and \U$14250 ( \14627 , \925 , \10876 );
and \U$14251 ( \14628 , \851 , \10873 );
nor \U$14252 ( \14629 , \14627 , \14628 );
xnor \U$14253 ( \14630 , \14629 , \9821 );
and \U$14254 ( \14631 , \1050 , \10063 );
and \U$14255 ( \14632 , \987 , \10061 );
nor \U$14256 ( \14633 , \14631 , \14632 );
xnor \U$14257 ( \14634 , \14633 , \9824 );
and \U$14258 ( \14635 , \14630 , \14634 );
and \U$14259 ( \14636 , \1336 , \9495 );
and \U$14260 ( \14637 , \1248 , \9493 );
nor \U$14261 ( \14638 , \14636 , \14637 );
xnor \U$14262 ( \14639 , \14638 , \9185 );
and \U$14263 ( \14640 , \14634 , \14639 );
and \U$14264 ( \14641 , \14630 , \14639 );
or \U$14265 ( \14642 , \14635 , \14640 , \14641 );
and \U$14266 ( \14643 , \14626 , \14642 );
and \U$14267 ( \14644 , \1446 , \8958 );
and \U$14268 ( \14645 , \1441 , \8956 );
nor \U$14269 ( \14646 , \14644 , \14645 );
xnor \U$14270 ( \14647 , \14646 , \8587 );
and \U$14271 ( \14648 , \1677 , \8396 );
and \U$14272 ( \14649 , \1562 , \8394 );
nor \U$14273 ( \14650 , \14648 , \14649 );
xnor \U$14274 ( \14651 , \14650 , \8078 );
and \U$14275 ( \14652 , \14647 , \14651 );
and \U$14276 ( \14653 , \1861 , \7829 );
and \U$14277 ( \14654 , \1853 , \7827 );
nor \U$14278 ( \14655 , \14653 , \14654 );
xnor \U$14279 ( \14656 , \14655 , \7580 );
and \U$14280 ( \14657 , \14651 , \14656 );
and \U$14281 ( \14658 , \14647 , \14656 );
or \U$14282 ( \14659 , \14652 , \14657 , \14658 );
and \U$14283 ( \14660 , \14642 , \14659 );
and \U$14284 ( \14661 , \14626 , \14659 );
or \U$14285 ( \14662 , \14643 , \14660 , \14661 );
and \U$14286 ( \14663 , \14609 , \14662 );
and \U$14287 ( \14664 , \14564 , \14662 );
or \U$14288 ( \14665 , \14610 , \14663 , \14664 );
xor \U$14289 ( \14666 , \14333 , \14337 );
xor \U$14290 ( \14667 , \14666 , \14342 );
xor \U$14291 ( \14668 , \14362 , \14366 );
xor \U$14292 ( \14669 , \14668 , \14371 );
and \U$14293 ( \14670 , \14667 , \14669 );
xor \U$14294 ( \14671 , \14297 , \14301 );
xor \U$14295 ( \14672 , \14671 , \14306 );
and \U$14296 ( \14673 , \14669 , \14672 );
and \U$14297 ( \14674 , \14667 , \14672 );
or \U$14298 ( \14675 , \14670 , \14673 , \14674 );
nand \U$14299 ( \14676 , \11029 , \752 );
xnor \U$14300 ( \14677 , \14676 , \711 );
xor \U$14301 ( \14678 , \14382 , \14386 );
xor \U$14302 ( \14679 , \14678 , \14391 );
and \U$14303 ( \14680 , \14677 , \14679 );
xor \U$14304 ( \14681 , \14415 , \14419 );
xor \U$14305 ( \14682 , \14681 , \14424 );
and \U$14306 ( \14683 , \14679 , \14682 );
and \U$14307 ( \14684 , \14677 , \14682 );
or \U$14308 ( \14685 , \14680 , \14683 , \14684 );
and \U$14309 ( \14686 , \14675 , \14685 );
xor \U$14310 ( \14687 , \14398 , \14402 );
xor \U$14311 ( \14688 , \14687 , \14407 );
xor \U$14312 ( \14689 , \14281 , \14285 );
xor \U$14313 ( \14690 , \14689 , \14290 );
and \U$14314 ( \14691 , \14688 , \14690 );
xor \U$14315 ( \14692 , \14314 , \14318 );
xor \U$14316 ( \14693 , \14692 , \14323 );
and \U$14317 ( \14694 , \14690 , \14693 );
and \U$14318 ( \14695 , \14688 , \14693 );
or \U$14319 ( \14696 , \14691 , \14694 , \14695 );
and \U$14320 ( \14697 , \14685 , \14696 );
and \U$14321 ( \14698 , \14675 , \14696 );
or \U$14322 ( \14699 , \14686 , \14697 , \14698 );
and \U$14323 ( \14700 , \14665 , \14699 );
xor \U$14324 ( \14701 , \14245 , \14247 );
xor \U$14325 ( \14702 , \14701 , \14250 );
xor \U$14326 ( \14703 , \14255 , \14257 );
xor \U$14327 ( \14704 , \14703 , \14260 );
and \U$14328 ( \14705 , \14702 , \14704 );
xor \U$14329 ( \14706 , \14266 , \14268 );
xor \U$14330 ( \14707 , \14706 , \14271 );
and \U$14331 ( \14708 , \14704 , \14707 );
and \U$14332 ( \14709 , \14702 , \14707 );
or \U$14333 ( \14710 , \14705 , \14708 , \14709 );
and \U$14334 ( \14711 , \14699 , \14710 );
and \U$14335 ( \14712 , \14665 , \14710 );
or \U$14336 ( \14713 , \14700 , \14711 , \14712 );
xor \U$14337 ( \14714 , \14253 , \14263 );
xor \U$14338 ( \14715 , \14714 , \14274 );
xor \U$14339 ( \14716 , \14329 , \14377 );
xor \U$14340 ( \14717 , \14716 , \14430 );
and \U$14341 ( \14718 , \14715 , \14717 );
xor \U$14342 ( \14719 , \14436 , \14438 );
xor \U$14343 ( \14720 , \14719 , \14441 );
and \U$14344 ( \14721 , \14717 , \14720 );
and \U$14345 ( \14722 , \14715 , \14720 );
or \U$14346 ( \14723 , \14718 , \14721 , \14722 );
and \U$14347 ( \14724 , \14713 , \14723 );
xor \U$14348 ( \14725 , \14293 , \14309 );
xor \U$14349 ( \14726 , \14725 , \14326 );
xor \U$14350 ( \14727 , \14345 , \14357 );
xor \U$14351 ( \14728 , \14727 , \14374 );
and \U$14352 ( \14729 , \14726 , \14728 );
xor \U$14353 ( \14730 , \14394 , \14410 );
xor \U$14354 ( \14731 , \14730 , \14427 );
and \U$14355 ( \14732 , \14728 , \14731 );
and \U$14356 ( \14733 , \14726 , \14731 );
or \U$14357 ( \14734 , \14729 , \14732 , \14733 );
xor \U$14358 ( \14735 , \14449 , \14451 );
xor \U$14359 ( \14736 , \14735 , \14454 );
and \U$14360 ( \14737 , \14734 , \14736 );
xor \U$14361 ( \14738 , \14459 , \14461 );
and \U$14362 ( \14739 , \14736 , \14738 );
and \U$14363 ( \14740 , \14734 , \14738 );
or \U$14364 ( \14741 , \14737 , \14739 , \14740 );
and \U$14365 ( \14742 , \14723 , \14741 );
and \U$14366 ( \14743 , \14713 , \14741 );
or \U$14367 ( \14744 , \14724 , \14742 , \14743 );
xor \U$14368 ( \14745 , \14053 , \14105 );
xor \U$14369 ( \14746 , \14745 , \14158 );
xor \U$14370 ( \14747 , \14457 , \14462 );
xor \U$14371 ( \14748 , \14747 , \14465 );
and \U$14372 ( \14749 , \14746 , \14748 );
xor \U$14373 ( \14750 , \14471 , \14473 );
xor \U$14374 ( \14751 , \14750 , \14476 );
and \U$14375 ( \14752 , \14748 , \14751 );
and \U$14376 ( \14753 , \14746 , \14751 );
or \U$14377 ( \14754 , \14749 , \14752 , \14753 );
and \U$14378 ( \14755 , \14744 , \14754 );
xor \U$14379 ( \14756 , \14484 , \14486 );
xor \U$14380 ( \14757 , \14756 , \14489 );
and \U$14381 ( \14758 , \14754 , \14757 );
and \U$14382 ( \14759 , \14744 , \14757 );
or \U$14383 ( \14760 , \14755 , \14758 , \14759 );
xor \U$14384 ( \14761 , \14175 , \14193 );
xor \U$14385 ( \14762 , \14761 , \14204 );
and \U$14386 ( \14763 , \14760 , \14762 );
xor \U$14387 ( \14764 , \14482 , \14492 );
xor \U$14388 ( \14765 , \14764 , \14495 );
and \U$14389 ( \14766 , \14762 , \14765 );
and \U$14390 ( \14767 , \14760 , \14765 );
or \U$14391 ( \14768 , \14763 , \14766 , \14767 );
xor \U$14392 ( \14769 , \14498 , \14500 );
xor \U$14393 ( \14770 , \14769 , \14503 );
and \U$14394 ( \14771 , \14768 , \14770 );
and \U$14395 ( \14772 , \14512 , \14771 );
xor \U$14396 ( \14773 , \14512 , \14771 );
xor \U$14397 ( \14774 , \14768 , \14770 );
and \U$14398 ( \14775 , \4073 , \4868 );
and \U$14399 ( \14776 , \3951 , \4866 );
nor \U$14400 ( \14777 , \14775 , \14776 );
xnor \U$14401 ( \14778 , \14777 , \4636 );
and \U$14402 ( \14779 , \4334 , \4417 );
and \U$14403 ( \14780 , \4078 , \4415 );
nor \U$14404 ( \14781 , \14779 , \14780 );
xnor \U$14405 ( \14782 , \14781 , \4274 );
and \U$14406 ( \14783 , \14778 , \14782 );
and \U$14407 ( \14784 , \4833 , \4094 );
and \U$14408 ( \14785 , \4531 , \4092 );
nor \U$14409 ( \14786 , \14784 , \14785 );
xnor \U$14410 ( \14787 , \14786 , \3848 );
and \U$14411 ( \14788 , \14782 , \14787 );
and \U$14412 ( \14789 , \14778 , \14787 );
or \U$14413 ( \14790 , \14783 , \14788 , \14789 );
and \U$14414 ( \14791 , \2902 , \6297 );
and \U$14415 ( \14792 , \2728 , \6295 );
nor \U$14416 ( \14793 , \14791 , \14792 );
xnor \U$14417 ( \14794 , \14793 , \5957 );
and \U$14418 ( \14795 , \3207 , \5708 );
and \U$14419 ( \14796 , \3069 , \5706 );
nor \U$14420 ( \14797 , \14795 , \14796 );
xnor \U$14421 ( \14798 , \14797 , \5467 );
and \U$14422 ( \14799 , \14794 , \14798 );
and \U$14423 ( \14800 , \3743 , \5242 );
and \U$14424 ( \14801 , \3326 , \5240 );
nor \U$14425 ( \14802 , \14800 , \14801 );
xnor \U$14426 ( \14803 , \14802 , \5054 );
and \U$14427 ( \14804 , \14798 , \14803 );
and \U$14428 ( \14805 , \14794 , \14803 );
or \U$14429 ( \14806 , \14799 , \14804 , \14805 );
and \U$14430 ( \14807 , \14790 , \14806 );
and \U$14431 ( \14808 , \5310 , \3699 );
and \U$14432 ( \14809 , \4841 , \3697 );
nor \U$14433 ( \14810 , \14808 , \14809 );
xnor \U$14434 ( \14811 , \14810 , \3512 );
and \U$14435 ( \14812 , \5579 , \3386 );
and \U$14436 ( \14813 , \5315 , \3384 );
nor \U$14437 ( \14814 , \14812 , \14813 );
xnor \U$14438 ( \14815 , \14814 , \3181 );
and \U$14439 ( \14816 , \14811 , \14815 );
and \U$14440 ( \14817 , \6210 , \2980 );
and \U$14441 ( \14818 , \5838 , \2978 );
nor \U$14442 ( \14819 , \14817 , \14818 );
xnor \U$14443 ( \14820 , \14819 , \2831 );
and \U$14444 ( \14821 , \14815 , \14820 );
and \U$14445 ( \14822 , \14811 , \14820 );
or \U$14446 ( \14823 , \14816 , \14821 , \14822 );
and \U$14447 ( \14824 , \14806 , \14823 );
and \U$14448 ( \14825 , \14790 , \14823 );
or \U$14449 ( \14826 , \14807 , \14824 , \14825 );
and \U$14450 ( \14827 , \2104 , \7829 );
and \U$14451 ( \14828 , \1861 , \7827 );
nor \U$14452 ( \14829 , \14827 , \14828 );
xnor \U$14453 ( \14830 , \14829 , \7580 );
and \U$14454 ( \14831 , \2295 , \7300 );
and \U$14455 ( \14832 , \2109 , \7298 );
nor \U$14456 ( \14833 , \14831 , \14832 );
xnor \U$14457 ( \14834 , \14833 , \7040 );
and \U$14458 ( \14835 , \14830 , \14834 );
and \U$14459 ( \14836 , \2703 , \6806 );
and \U$14460 ( \14837 , \2439 , \6804 );
nor \U$14461 ( \14838 , \14836 , \14837 );
xnor \U$14462 ( \14839 , \14838 , \6491 );
and \U$14463 ( \14840 , \14834 , \14839 );
and \U$14464 ( \14841 , \14830 , \14839 );
or \U$14465 ( \14842 , \14835 , \14840 , \14841 );
and \U$14466 ( \14843 , \1441 , \9495 );
and \U$14467 ( \14844 , \1336 , \9493 );
nor \U$14468 ( \14845 , \14843 , \14844 );
xnor \U$14469 ( \14846 , \14845 , \9185 );
and \U$14470 ( \14847 , \1562 , \8958 );
and \U$14471 ( \14848 , \1446 , \8956 );
nor \U$14472 ( \14849 , \14847 , \14848 );
xnor \U$14473 ( \14850 , \14849 , \8587 );
and \U$14474 ( \14851 , \14846 , \14850 );
and \U$14475 ( \14852 , \1853 , \8396 );
and \U$14476 ( \14853 , \1677 , \8394 );
nor \U$14477 ( \14854 , \14852 , \14853 );
xnor \U$14478 ( \14855 , \14854 , \8078 );
and \U$14479 ( \14856 , \14850 , \14855 );
and \U$14480 ( \14857 , \14846 , \14855 );
or \U$14481 ( \14858 , \14851 , \14856 , \14857 );
and \U$14482 ( \14859 , \14842 , \14858 );
and \U$14483 ( \14860 , \987 , \10876 );
and \U$14484 ( \14861 , \925 , \10873 );
nor \U$14485 ( \14862 , \14860 , \14861 );
xnor \U$14486 ( \14863 , \14862 , \9821 );
and \U$14487 ( \14864 , \1248 , \10063 );
and \U$14488 ( \14865 , \1050 , \10061 );
nor \U$14489 ( \14866 , \14864 , \14865 );
xnor \U$14490 ( \14867 , \14866 , \9824 );
and \U$14491 ( \14868 , \14863 , \14867 );
and \U$14492 ( \14869 , \14867 , \816 );
and \U$14493 ( \14870 , \14863 , \816 );
or \U$14494 ( \14871 , \14868 , \14869 , \14870 );
and \U$14495 ( \14872 , \14858 , \14871 );
and \U$14496 ( \14873 , \14842 , \14871 );
or \U$14497 ( \14874 , \14859 , \14872 , \14873 );
and \U$14498 ( \14875 , \14826 , \14874 );
and \U$14499 ( \14876 , \6562 , \2658 );
and \U$14500 ( \14877 , \6219 , \2656 );
nor \U$14501 ( \14878 , \14876 , \14877 );
xnor \U$14502 ( \14879 , \14878 , \2516 );
and \U$14503 ( \14880 , \7067 , \2362 );
and \U$14504 ( \14881 , \6764 , \2360 );
nor \U$14505 ( \14882 , \14880 , \14881 );
xnor \U$14506 ( \14883 , \14882 , \2225 );
and \U$14507 ( \14884 , \14879 , \14883 );
and \U$14508 ( \14885 , \7765 , \2156 );
and \U$14509 ( \14886 , \7239 , \2154 );
nor \U$14510 ( \14887 , \14885 , \14886 );
xnor \U$14511 ( \14888 , \14887 , \2004 );
and \U$14512 ( \14889 , \14883 , \14888 );
and \U$14513 ( \14890 , \14879 , \14888 );
or \U$14514 ( \14891 , \14884 , \14889 , \14890 );
and \U$14515 ( \14892 , \10223 , \1222 );
and \U$14516 ( \14893 , \9620 , \1220 );
nor \U$14517 ( \14894 , \14892 , \14893 );
xnor \U$14518 ( \14895 , \14894 , \1144 );
and \U$14519 ( \14896 , \10409 , \1058 );
and \U$14520 ( \14897 , \10228 , \1056 );
nor \U$14521 ( \14898 , \14896 , \14897 );
xnor \U$14522 ( \14899 , \14898 , \964 );
and \U$14523 ( \14900 , \14895 , \14899 );
nand \U$14524 ( \14901 , \11029 , \886 );
xnor \U$14525 ( \14902 , \14901 , \816 );
and \U$14526 ( \14903 , \14899 , \14902 );
and \U$14527 ( \14904 , \14895 , \14902 );
or \U$14528 ( \14905 , \14900 , \14903 , \14904 );
and \U$14529 ( \14906 , \14891 , \14905 );
and \U$14530 ( \14907 , \8435 , \1888 );
and \U$14531 ( \14908 , \8189 , \1886 );
nor \U$14532 ( \14909 , \14907 , \14908 );
xnor \U$14533 ( \14910 , \14909 , \1732 );
and \U$14534 ( \14911 , \8759 , \1616 );
and \U$14535 ( \14912 , \8440 , \1614 );
nor \U$14536 ( \14913 , \14911 , \14912 );
xnor \U$14537 ( \14914 , \14913 , \1503 );
and \U$14538 ( \14915 , \14910 , \14914 );
and \U$14539 ( \14916 , \9612 , \1422 );
and \U$14540 ( \14917 , \9043 , \1420 );
nor \U$14541 ( \14918 , \14916 , \14917 );
xnor \U$14542 ( \14919 , \14918 , \1286 );
and \U$14543 ( \14920 , \14914 , \14919 );
and \U$14544 ( \14921 , \14910 , \14919 );
or \U$14545 ( \14922 , \14915 , \14920 , \14921 );
and \U$14546 ( \14923 , \14905 , \14922 );
and \U$14547 ( \14924 , \14891 , \14922 );
or \U$14548 ( \14925 , \14906 , \14923 , \14924 );
and \U$14549 ( \14926 , \14874 , \14925 );
and \U$14550 ( \14927 , \14826 , \14925 );
or \U$14551 ( \14928 , \14875 , \14926 , \14927 );
xor \U$14552 ( \14929 , \14614 , \14618 );
xor \U$14553 ( \14930 , \14929 , \14623 );
xor \U$14554 ( \14931 , \14630 , \14634 );
xor \U$14555 ( \14932 , \14931 , \14639 );
and \U$14556 ( \14933 , \14930 , \14932 );
xor \U$14557 ( \14934 , \14647 , \14651 );
xor \U$14558 ( \14935 , \14934 , \14656 );
and \U$14559 ( \14936 , \14932 , \14935 );
and \U$14560 ( \14937 , \14930 , \14935 );
or \U$14561 ( \14938 , \14933 , \14936 , \14937 );
xor \U$14562 ( \14939 , \14516 , \14520 );
xor \U$14563 ( \14940 , \14939 , \14525 );
xor \U$14564 ( \14941 , \14532 , \14536 );
xor \U$14565 ( \14942 , \14941 , \14541 );
and \U$14566 ( \14943 , \14940 , \14942 );
xor \U$14567 ( \14944 , \14549 , \14553 );
xor \U$14568 ( \14945 , \14944 , \14558 );
and \U$14569 ( \14946 , \14942 , \14945 );
and \U$14570 ( \14947 , \14940 , \14945 );
or \U$14571 ( \14948 , \14943 , \14946 , \14947 );
and \U$14572 ( \14949 , \14938 , \14948 );
xor \U$14573 ( \14950 , \14568 , \14572 );
xor \U$14574 ( \14951 , \14950 , \14577 );
xor \U$14575 ( \14952 , \14584 , \14588 );
xor \U$14576 ( \14953 , \14952 , \14593 );
and \U$14577 ( \14954 , \14951 , \14953 );
xor \U$14578 ( \14955 , \14601 , \14605 );
and \U$14579 ( \14956 , \14953 , \14955 );
and \U$14580 ( \14957 , \14951 , \14955 );
or \U$14581 ( \14958 , \14954 , \14956 , \14957 );
and \U$14582 ( \14959 , \14948 , \14958 );
and \U$14583 ( \14960 , \14938 , \14958 );
or \U$14584 ( \14961 , \14949 , \14959 , \14960 );
and \U$14585 ( \14962 , \14928 , \14961 );
xor \U$14586 ( \14963 , \14349 , \14353 );
xor \U$14587 ( \14964 , \14963 , \711 );
xor \U$14588 ( \14965 , \14667 , \14669 );
xor \U$14589 ( \14966 , \14965 , \14672 );
and \U$14590 ( \14967 , \14964 , \14966 );
xor \U$14591 ( \14968 , \14688 , \14690 );
xor \U$14592 ( \14969 , \14968 , \14693 );
and \U$14593 ( \14970 , \14966 , \14969 );
and \U$14594 ( \14971 , \14964 , \14969 );
or \U$14595 ( \14972 , \14967 , \14970 , \14971 );
and \U$14596 ( \14973 , \14961 , \14972 );
and \U$14597 ( \14974 , \14928 , \14972 );
or \U$14598 ( \14975 , \14962 , \14973 , \14974 );
xor \U$14599 ( \14976 , \14528 , \14544 );
xor \U$14600 ( \14977 , \14976 , \14561 );
xor \U$14601 ( \14978 , \14580 , \14596 );
xor \U$14602 ( \14979 , \14978 , \14606 );
and \U$14603 ( \14980 , \14977 , \14979 );
xor \U$14604 ( \14981 , \14677 , \14679 );
xor \U$14605 ( \14982 , \14981 , \14682 );
and \U$14606 ( \14983 , \14979 , \14982 );
and \U$14607 ( \14984 , \14977 , \14982 );
or \U$14608 ( \14985 , \14980 , \14983 , \14984 );
xor \U$14609 ( \14986 , \14726 , \14728 );
xor \U$14610 ( \14987 , \14986 , \14731 );
and \U$14611 ( \14988 , \14985 , \14987 );
xor \U$14612 ( \14989 , \14702 , \14704 );
xor \U$14613 ( \14990 , \14989 , \14707 );
and \U$14614 ( \14991 , \14987 , \14990 );
and \U$14615 ( \14992 , \14985 , \14990 );
or \U$14616 ( \14993 , \14988 , \14991 , \14992 );
and \U$14617 ( \14994 , \14975 , \14993 );
xor \U$14618 ( \14995 , \14564 , \14609 );
xor \U$14619 ( \14996 , \14995 , \14662 );
xor \U$14620 ( \14997 , \14675 , \14685 );
xor \U$14621 ( \14998 , \14997 , \14696 );
and \U$14622 ( \14999 , \14996 , \14998 );
and \U$14623 ( \15000 , \14993 , \14999 );
and \U$14624 ( \15001 , \14975 , \14999 );
or \U$14625 ( \15002 , \14994 , \15000 , \15001 );
xor \U$14626 ( \15003 , \14665 , \14699 );
xor \U$14627 ( \15004 , \15003 , \14710 );
xor \U$14628 ( \15005 , \14715 , \14717 );
xor \U$14629 ( \15006 , \15005 , \14720 );
and \U$14630 ( \15007 , \15004 , \15006 );
xor \U$14631 ( \15008 , \14734 , \14736 );
xor \U$14632 ( \15009 , \15008 , \14738 );
and \U$14633 ( \15010 , \15006 , \15009 );
and \U$14634 ( \15011 , \15004 , \15009 );
or \U$14635 ( \15012 , \15007 , \15010 , \15011 );
and \U$14636 ( \15013 , \15002 , \15012 );
xor \U$14637 ( \15014 , \14277 , \14433 );
xor \U$14638 ( \15015 , \15014 , \14444 );
and \U$14639 ( \15016 , \15012 , \15015 );
and \U$14640 ( \15017 , \15002 , \15015 );
or \U$14641 ( \15018 , \15013 , \15016 , \15017 );
xor \U$14642 ( \15019 , \14713 , \14723 );
xor \U$14643 ( \15020 , \15019 , \14741 );
xor \U$14644 ( \15021 , \14746 , \14748 );
xor \U$14645 ( \15022 , \15021 , \14751 );
and \U$14646 ( \15023 , \15020 , \15022 );
and \U$14647 ( \15024 , \15018 , \15023 );
xor \U$14648 ( \15025 , \14447 , \14468 );
xor \U$14649 ( \15026 , \15025 , \14479 );
and \U$14650 ( \15027 , \15023 , \15026 );
and \U$14651 ( \15028 , \15018 , \15026 );
or \U$14652 ( \15029 , \15024 , \15027 , \15028 );
xor \U$14653 ( \15030 , \14760 , \14762 );
xor \U$14654 ( \15031 , \15030 , \14765 );
and \U$14655 ( \15032 , \15029 , \15031 );
and \U$14656 ( \15033 , \14774 , \15032 );
xor \U$14657 ( \15034 , \14774 , \15032 );
xor \U$14658 ( \15035 , \15029 , \15031 );
xor \U$14659 ( \15036 , \15018 , \15023 );
xor \U$14660 ( \15037 , \15036 , \15026 );
xor \U$14661 ( \15038 , \14744 , \14754 );
xor \U$14662 ( \15039 , \15038 , \14757 );
and \U$14663 ( \15040 , \15037 , \15039 );
and \U$14664 ( \15041 , \15035 , \15040 );
xor \U$14665 ( \15042 , \15035 , \15040 );
xor \U$14666 ( \15043 , \15037 , \15039 );
and \U$14667 ( \15044 , \2439 , \7300 );
and \U$14668 ( \15045 , \2295 , \7298 );
nor \U$14669 ( \15046 , \15044 , \15045 );
xnor \U$14670 ( \15047 , \15046 , \7040 );
and \U$14671 ( \15048 , \2728 , \6806 );
and \U$14672 ( \15049 , \2703 , \6804 );
nor \U$14673 ( \15050 , \15048 , \15049 );
xnor \U$14674 ( \15051 , \15050 , \6491 );
and \U$14675 ( \15052 , \15047 , \15051 );
and \U$14676 ( \15053 , \3069 , \6297 );
and \U$14677 ( \15054 , \2902 , \6295 );
nor \U$14678 ( \15055 , \15053 , \15054 );
xnor \U$14679 ( \15056 , \15055 , \5957 );
and \U$14680 ( \15057 , \15051 , \15056 );
and \U$14681 ( \15058 , \15047 , \15056 );
or \U$14682 ( \15059 , \15052 , \15057 , \15058 );
and \U$14683 ( \15060 , \1050 , \10876 );
and \U$14684 ( \15061 , \987 , \10873 );
nor \U$14685 ( \15062 , \15060 , \15061 );
xnor \U$14686 ( \15063 , \15062 , \9821 );
and \U$14687 ( \15064 , \1336 , \10063 );
and \U$14688 ( \15065 , \1248 , \10061 );
nor \U$14689 ( \15066 , \15064 , \15065 );
xnor \U$14690 ( \15067 , \15066 , \9824 );
and \U$14691 ( \15068 , \15063 , \15067 );
and \U$14692 ( \15069 , \1446 , \9495 );
and \U$14693 ( \15070 , \1441 , \9493 );
nor \U$14694 ( \15071 , \15069 , \15070 );
xnor \U$14695 ( \15072 , \15071 , \9185 );
and \U$14696 ( \15073 , \15067 , \15072 );
and \U$14697 ( \15074 , \15063 , \15072 );
or \U$14698 ( \15075 , \15068 , \15073 , \15074 );
and \U$14699 ( \15076 , \15059 , \15075 );
and \U$14700 ( \15077 , \1677 , \8958 );
and \U$14701 ( \15078 , \1562 , \8956 );
nor \U$14702 ( \15079 , \15077 , \15078 );
xnor \U$14703 ( \15080 , \15079 , \8587 );
and \U$14704 ( \15081 , \1861 , \8396 );
and \U$14705 ( \15082 , \1853 , \8394 );
nor \U$14706 ( \15083 , \15081 , \15082 );
xnor \U$14707 ( \15084 , \15083 , \8078 );
and \U$14708 ( \15085 , \15080 , \15084 );
and \U$14709 ( \15086 , \2109 , \7829 );
and \U$14710 ( \15087 , \2104 , \7827 );
nor \U$14711 ( \15088 , \15086 , \15087 );
xnor \U$14712 ( \15089 , \15088 , \7580 );
and \U$14713 ( \15090 , \15084 , \15089 );
and \U$14714 ( \15091 , \15080 , \15089 );
or \U$14715 ( \15092 , \15085 , \15090 , \15091 );
and \U$14716 ( \15093 , \15075 , \15092 );
and \U$14717 ( \15094 , \15059 , \15092 );
or \U$14718 ( \15095 , \15076 , \15093 , \15094 );
and \U$14719 ( \15096 , \4531 , \4417 );
and \U$14720 ( \15097 , \4334 , \4415 );
nor \U$14721 ( \15098 , \15096 , \15097 );
xnor \U$14722 ( \15099 , \15098 , \4274 );
and \U$14723 ( \15100 , \4841 , \4094 );
and \U$14724 ( \15101 , \4833 , \4092 );
nor \U$14725 ( \15102 , \15100 , \15101 );
xnor \U$14726 ( \15103 , \15102 , \3848 );
and \U$14727 ( \15104 , \15099 , \15103 );
and \U$14728 ( \15105 , \5315 , \3699 );
and \U$14729 ( \15106 , \5310 , \3697 );
nor \U$14730 ( \15107 , \15105 , \15106 );
xnor \U$14731 ( \15108 , \15107 , \3512 );
and \U$14732 ( \15109 , \15103 , \15108 );
and \U$14733 ( \15110 , \15099 , \15108 );
or \U$14734 ( \15111 , \15104 , \15109 , \15110 );
and \U$14735 ( \15112 , \3326 , \5708 );
and \U$14736 ( \15113 , \3207 , \5706 );
nor \U$14737 ( \15114 , \15112 , \15113 );
xnor \U$14738 ( \15115 , \15114 , \5467 );
and \U$14739 ( \15116 , \3951 , \5242 );
and \U$14740 ( \15117 , \3743 , \5240 );
nor \U$14741 ( \15118 , \15116 , \15117 );
xnor \U$14742 ( \15119 , \15118 , \5054 );
and \U$14743 ( \15120 , \15115 , \15119 );
and \U$14744 ( \15121 , \4078 , \4868 );
and \U$14745 ( \15122 , \4073 , \4866 );
nor \U$14746 ( \15123 , \15121 , \15122 );
xnor \U$14747 ( \15124 , \15123 , \4636 );
and \U$14748 ( \15125 , \15119 , \15124 );
and \U$14749 ( \15126 , \15115 , \15124 );
or \U$14750 ( \15127 , \15120 , \15125 , \15126 );
and \U$14751 ( \15128 , \15111 , \15127 );
and \U$14752 ( \15129 , \5838 , \3386 );
and \U$14753 ( \15130 , \5579 , \3384 );
nor \U$14754 ( \15131 , \15129 , \15130 );
xnor \U$14755 ( \15132 , \15131 , \3181 );
and \U$14756 ( \15133 , \6219 , \2980 );
and \U$14757 ( \15134 , \6210 , \2978 );
nor \U$14758 ( \15135 , \15133 , \15134 );
xnor \U$14759 ( \15136 , \15135 , \2831 );
and \U$14760 ( \15137 , \15132 , \15136 );
and \U$14761 ( \15138 , \6764 , \2658 );
and \U$14762 ( \15139 , \6562 , \2656 );
nor \U$14763 ( \15140 , \15138 , \15139 );
xnor \U$14764 ( \15141 , \15140 , \2516 );
and \U$14765 ( \15142 , \15136 , \15141 );
and \U$14766 ( \15143 , \15132 , \15141 );
or \U$14767 ( \15144 , \15137 , \15142 , \15143 );
and \U$14768 ( \15145 , \15127 , \15144 );
and \U$14769 ( \15146 , \15111 , \15144 );
or \U$14770 ( \15147 , \15128 , \15145 , \15146 );
and \U$14771 ( \15148 , \15095 , \15147 );
and \U$14772 ( \15149 , \9043 , \1616 );
and \U$14773 ( \15150 , \8759 , \1614 );
nor \U$14774 ( \15151 , \15149 , \15150 );
xnor \U$14775 ( \15152 , \15151 , \1503 );
and \U$14776 ( \15153 , \9620 , \1422 );
and \U$14777 ( \15154 , \9612 , \1420 );
nor \U$14778 ( \15155 , \15153 , \15154 );
xnor \U$14779 ( \15156 , \15155 , \1286 );
and \U$14780 ( \15157 , \15152 , \15156 );
and \U$14781 ( \15158 , \10228 , \1222 );
and \U$14782 ( \15159 , \10223 , \1220 );
nor \U$14783 ( \15160 , \15158 , \15159 );
xnor \U$14784 ( \15161 , \15160 , \1144 );
and \U$14785 ( \15162 , \15156 , \15161 );
and \U$14786 ( \15163 , \15152 , \15161 );
or \U$14787 ( \15164 , \15157 , \15162 , \15163 );
and \U$14788 ( \15165 , \7239 , \2362 );
and \U$14789 ( \15166 , \7067 , \2360 );
nor \U$14790 ( \15167 , \15165 , \15166 );
xnor \U$14791 ( \15168 , \15167 , \2225 );
and \U$14792 ( \15169 , \8189 , \2156 );
and \U$14793 ( \15170 , \7765 , \2154 );
nor \U$14794 ( \15171 , \15169 , \15170 );
xnor \U$14795 ( \15172 , \15171 , \2004 );
and \U$14796 ( \15173 , \15168 , \15172 );
and \U$14797 ( \15174 , \8440 , \1888 );
and \U$14798 ( \15175 , \8435 , \1886 );
nor \U$14799 ( \15176 , \15174 , \15175 );
xnor \U$14800 ( \15177 , \15176 , \1732 );
and \U$14801 ( \15178 , \15172 , \15177 );
and \U$14802 ( \15179 , \15168 , \15177 );
or \U$14803 ( \15180 , \15173 , \15178 , \15179 );
and \U$14804 ( \15181 , \15164 , \15180 );
xor \U$14805 ( \15182 , \14895 , \14899 );
xor \U$14806 ( \15183 , \15182 , \14902 );
and \U$14807 ( \15184 , \15180 , \15183 );
and \U$14808 ( \15185 , \15164 , \15183 );
or \U$14809 ( \15186 , \15181 , \15184 , \15185 );
and \U$14810 ( \15187 , \15147 , \15186 );
and \U$14811 ( \15188 , \15095 , \15186 );
or \U$14812 ( \15189 , \15148 , \15187 , \15188 );
xor \U$14813 ( \15190 , \14879 , \14883 );
xor \U$14814 ( \15191 , \15190 , \14888 );
xor \U$14815 ( \15192 , \14811 , \14815 );
xor \U$14816 ( \15193 , \15192 , \14820 );
and \U$14817 ( \15194 , \15191 , \15193 );
xor \U$14818 ( \15195 , \14910 , \14914 );
xor \U$14819 ( \15196 , \15195 , \14919 );
and \U$14820 ( \15197 , \15193 , \15196 );
and \U$14821 ( \15198 , \15191 , \15196 );
or \U$14822 ( \15199 , \15194 , \15197 , \15198 );
xor \U$14823 ( \15200 , \14778 , \14782 );
xor \U$14824 ( \15201 , \15200 , \14787 );
xor \U$14825 ( \15202 , \14794 , \14798 );
xor \U$14826 ( \15203 , \15202 , \14803 );
and \U$14827 ( \15204 , \15201 , \15203 );
xor \U$14828 ( \15205 , \14830 , \14834 );
xor \U$14829 ( \15206 , \15205 , \14839 );
and \U$14830 ( \15207 , \15203 , \15206 );
and \U$14831 ( \15208 , \15201 , \15206 );
or \U$14832 ( \15209 , \15204 , \15207 , \15208 );
and \U$14833 ( \15210 , \15199 , \15209 );
xor \U$14834 ( \15211 , \14846 , \14850 );
xor \U$14835 ( \15212 , \15211 , \14855 );
xor \U$14836 ( \15213 , \14863 , \14867 );
xor \U$14837 ( \15214 , \15213 , \816 );
and \U$14838 ( \15215 , \15212 , \15214 );
and \U$14839 ( \15216 , \15209 , \15215 );
and \U$14840 ( \15217 , \15199 , \15215 );
or \U$14841 ( \15218 , \15210 , \15216 , \15217 );
and \U$14842 ( \15219 , \15189 , \15218 );
xor \U$14843 ( \15220 , \14930 , \14932 );
xor \U$14844 ( \15221 , \15220 , \14935 );
xor \U$14845 ( \15222 , \14940 , \14942 );
xor \U$14846 ( \15223 , \15222 , \14945 );
and \U$14847 ( \15224 , \15221 , \15223 );
xor \U$14848 ( \15225 , \14951 , \14953 );
xor \U$14849 ( \15226 , \15225 , \14955 );
and \U$14850 ( \15227 , \15223 , \15226 );
and \U$14851 ( \15228 , \15221 , \15226 );
or \U$14852 ( \15229 , \15224 , \15227 , \15228 );
and \U$14853 ( \15230 , \15218 , \15229 );
and \U$14854 ( \15231 , \15189 , \15229 );
or \U$14855 ( \15232 , \15219 , \15230 , \15231 );
xor \U$14856 ( \15233 , \14790 , \14806 );
xor \U$14857 ( \15234 , \15233 , \14823 );
xor \U$14858 ( \15235 , \14842 , \14858 );
xor \U$14859 ( \15236 , \15235 , \14871 );
and \U$14860 ( \15237 , \15234 , \15236 );
xor \U$14861 ( \15238 , \14891 , \14905 );
xor \U$14862 ( \15239 , \15238 , \14922 );
and \U$14863 ( \15240 , \15236 , \15239 );
and \U$14864 ( \15241 , \15234 , \15239 );
or \U$14865 ( \15242 , \15237 , \15240 , \15241 );
xor \U$14866 ( \15243 , \14626 , \14642 );
xor \U$14867 ( \15244 , \15243 , \14659 );
and \U$14868 ( \15245 , \15242 , \15244 );
xor \U$14869 ( \15246 , \14977 , \14979 );
xor \U$14870 ( \15247 , \15246 , \14982 );
and \U$14871 ( \15248 , \15244 , \15247 );
and \U$14872 ( \15249 , \15242 , \15247 );
or \U$14873 ( \15250 , \15245 , \15248 , \15249 );
and \U$14874 ( \15251 , \15232 , \15250 );
xor \U$14875 ( \15252 , \14826 , \14874 );
xor \U$14876 ( \15253 , \15252 , \14925 );
xor \U$14877 ( \15254 , \14938 , \14948 );
xor \U$14878 ( \15255 , \15254 , \14958 );
and \U$14879 ( \15256 , \15253 , \15255 );
xor \U$14880 ( \15257 , \14964 , \14966 );
xor \U$14881 ( \15258 , \15257 , \14969 );
and \U$14882 ( \15259 , \15255 , \15258 );
and \U$14883 ( \15260 , \15253 , \15258 );
or \U$14884 ( \15261 , \15256 , \15259 , \15260 );
and \U$14885 ( \15262 , \15250 , \15261 );
and \U$14886 ( \15263 , \15232 , \15261 );
or \U$14887 ( \15264 , \15251 , \15262 , \15263 );
xor \U$14888 ( \15265 , \14928 , \14961 );
xor \U$14889 ( \15266 , \15265 , \14972 );
xor \U$14890 ( \15267 , \14985 , \14987 );
xor \U$14891 ( \15268 , \15267 , \14990 );
and \U$14892 ( \15269 , \15266 , \15268 );
xor \U$14893 ( \15270 , \14996 , \14998 );
and \U$14894 ( \15271 , \15268 , \15270 );
and \U$14895 ( \15272 , \15266 , \15270 );
or \U$14896 ( \15273 , \15269 , \15271 , \15272 );
and \U$14897 ( \15274 , \15264 , \15273 );
xor \U$14898 ( \15275 , \15004 , \15006 );
xor \U$14899 ( \15276 , \15275 , \15009 );
and \U$14900 ( \15277 , \15273 , \15276 );
and \U$14901 ( \15278 , \15264 , \15276 );
or \U$14902 ( \15279 , \15274 , \15277 , \15278 );
xor \U$14903 ( \15280 , \15002 , \15012 );
xor \U$14904 ( \15281 , \15280 , \15015 );
and \U$14905 ( \15282 , \15279 , \15281 );
xor \U$14906 ( \15283 , \15020 , \15022 );
and \U$14907 ( \15284 , \15281 , \15283 );
and \U$14908 ( \15285 , \15279 , \15283 );
or \U$14909 ( \15286 , \15282 , \15284 , \15285 );
and \U$14910 ( \15287 , \15043 , \15286 );
xor \U$14911 ( \15288 , \15043 , \15286 );
xor \U$14912 ( \15289 , \15279 , \15281 );
xor \U$14913 ( \15290 , \15289 , \15283 );
and \U$14914 ( \15291 , \2295 , \7829 );
and \U$14915 ( \15292 , \2109 , \7827 );
nor \U$14916 ( \15293 , \15291 , \15292 );
xnor \U$14917 ( \15294 , \15293 , \7580 );
and \U$14918 ( \15295 , \2703 , \7300 );
and \U$14919 ( \15296 , \2439 , \7298 );
nor \U$14920 ( \15297 , \15295 , \15296 );
xnor \U$14921 ( \15298 , \15297 , \7040 );
and \U$14922 ( \15299 , \15294 , \15298 );
and \U$14923 ( \15300 , \2902 , \6806 );
and \U$14924 ( \15301 , \2728 , \6804 );
nor \U$14925 ( \15302 , \15300 , \15301 );
xnor \U$14926 ( \15303 , \15302 , \6491 );
and \U$14927 ( \15304 , \15298 , \15303 );
and \U$14928 ( \15305 , \15294 , \15303 );
or \U$14929 ( \15306 , \15299 , \15304 , \15305 );
and \U$14930 ( \15307 , \1562 , \9495 );
and \U$14931 ( \15308 , \1446 , \9493 );
nor \U$14932 ( \15309 , \15307 , \15308 );
xnor \U$14933 ( \15310 , \15309 , \9185 );
and \U$14934 ( \15311 , \1853 , \8958 );
and \U$14935 ( \15312 , \1677 , \8956 );
nor \U$14936 ( \15313 , \15311 , \15312 );
xnor \U$14937 ( \15314 , \15313 , \8587 );
and \U$14938 ( \15315 , \15310 , \15314 );
and \U$14939 ( \15316 , \2104 , \8396 );
and \U$14940 ( \15317 , \1861 , \8394 );
nor \U$14941 ( \15318 , \15316 , \15317 );
xnor \U$14942 ( \15319 , \15318 , \8078 );
and \U$14943 ( \15320 , \15314 , \15319 );
and \U$14944 ( \15321 , \15310 , \15319 );
or \U$14945 ( \15322 , \15315 , \15320 , \15321 );
and \U$14946 ( \15323 , \15306 , \15322 );
and \U$14947 ( \15324 , \1248 , \10876 );
and \U$14948 ( \15325 , \1050 , \10873 );
nor \U$14949 ( \15326 , \15324 , \15325 );
xnor \U$14950 ( \15327 , \15326 , \9821 );
and \U$14951 ( \15328 , \1441 , \10063 );
and \U$14952 ( \15329 , \1336 , \10061 );
nor \U$14953 ( \15330 , \15328 , \15329 );
xnor \U$14954 ( \15331 , \15330 , \9824 );
and \U$14955 ( \15332 , \15327 , \15331 );
and \U$14956 ( \15333 , \15331 , \964 );
and \U$14957 ( \15334 , \15327 , \964 );
or \U$14958 ( \15335 , \15332 , \15333 , \15334 );
and \U$14959 ( \15336 , \15322 , \15335 );
and \U$14960 ( \15337 , \15306 , \15335 );
or \U$14961 ( \15338 , \15323 , \15336 , \15337 );
and \U$14962 ( \15339 , \7067 , \2658 );
and \U$14963 ( \15340 , \6764 , \2656 );
nor \U$14964 ( \15341 , \15339 , \15340 );
xnor \U$14965 ( \15342 , \15341 , \2516 );
and \U$14966 ( \15343 , \7765 , \2362 );
and \U$14967 ( \15344 , \7239 , \2360 );
nor \U$14968 ( \15345 , \15343 , \15344 );
xnor \U$14969 ( \15346 , \15345 , \2225 );
and \U$14970 ( \15347 , \15342 , \15346 );
and \U$14971 ( \15348 , \8435 , \2156 );
and \U$14972 ( \15349 , \8189 , \2154 );
nor \U$14973 ( \15350 , \15348 , \15349 );
xnor \U$14974 ( \15351 , \15350 , \2004 );
and \U$14975 ( \15352 , \15346 , \15351 );
and \U$14976 ( \15353 , \15342 , \15351 );
or \U$14977 ( \15354 , \15347 , \15352 , \15353 );
and \U$14978 ( \15355 , \8759 , \1888 );
and \U$14979 ( \15356 , \8440 , \1886 );
nor \U$14980 ( \15357 , \15355 , \15356 );
xnor \U$14981 ( \15358 , \15357 , \1732 );
and \U$14982 ( \15359 , \9612 , \1616 );
and \U$14983 ( \15360 , \9043 , \1614 );
nor \U$14984 ( \15361 , \15359 , \15360 );
xnor \U$14985 ( \15362 , \15361 , \1503 );
and \U$14986 ( \15363 , \15358 , \15362 );
and \U$14987 ( \15364 , \10223 , \1422 );
and \U$14988 ( \15365 , \9620 , \1420 );
nor \U$14989 ( \15366 , \15364 , \15365 );
xnor \U$14990 ( \15367 , \15366 , \1286 );
and \U$14991 ( \15368 , \15362 , \15367 );
and \U$14992 ( \15369 , \15358 , \15367 );
or \U$14993 ( \15370 , \15363 , \15368 , \15369 );
and \U$14994 ( \15371 , \15354 , \15370 );
and \U$14995 ( \15372 , \11029 , \1058 );
and \U$14996 ( \15373 , \10409 , \1056 );
nor \U$14997 ( \15374 , \15372 , \15373 );
xnor \U$14998 ( \15375 , \15374 , \964 );
and \U$14999 ( \15376 , \15370 , \15375 );
and \U$15000 ( \15377 , \15354 , \15375 );
or \U$15001 ( \15378 , \15371 , \15376 , \15377 );
and \U$15002 ( \15379 , \15338 , \15378 );
and \U$15003 ( \15380 , \4334 , \4868 );
and \U$15004 ( \15381 , \4078 , \4866 );
nor \U$15005 ( \15382 , \15380 , \15381 );
xnor \U$15006 ( \15383 , \15382 , \4636 );
and \U$15007 ( \15384 , \4833 , \4417 );
and \U$15008 ( \15385 , \4531 , \4415 );
nor \U$15009 ( \15386 , \15384 , \15385 );
xnor \U$15010 ( \15387 , \15386 , \4274 );
and \U$15011 ( \15388 , \15383 , \15387 );
and \U$15012 ( \15389 , \5310 , \4094 );
and \U$15013 ( \15390 , \4841 , \4092 );
nor \U$15014 ( \15391 , \15389 , \15390 );
xnor \U$15015 ( \15392 , \15391 , \3848 );
and \U$15016 ( \15393 , \15387 , \15392 );
and \U$15017 ( \15394 , \15383 , \15392 );
or \U$15018 ( \15395 , \15388 , \15393 , \15394 );
and \U$15019 ( \15396 , \3207 , \6297 );
and \U$15020 ( \15397 , \3069 , \6295 );
nor \U$15021 ( \15398 , \15396 , \15397 );
xnor \U$15022 ( \15399 , \15398 , \5957 );
and \U$15023 ( \15400 , \3743 , \5708 );
and \U$15024 ( \15401 , \3326 , \5706 );
nor \U$15025 ( \15402 , \15400 , \15401 );
xnor \U$15026 ( \15403 , \15402 , \5467 );
and \U$15027 ( \15404 , \15399 , \15403 );
and \U$15028 ( \15405 , \4073 , \5242 );
and \U$15029 ( \15406 , \3951 , \5240 );
nor \U$15030 ( \15407 , \15405 , \15406 );
xnor \U$15031 ( \15408 , \15407 , \5054 );
and \U$15032 ( \15409 , \15403 , \15408 );
and \U$15033 ( \15410 , \15399 , \15408 );
or \U$15034 ( \15411 , \15404 , \15409 , \15410 );
and \U$15035 ( \15412 , \15395 , \15411 );
and \U$15036 ( \15413 , \5579 , \3699 );
and \U$15037 ( \15414 , \5315 , \3697 );
nor \U$15038 ( \15415 , \15413 , \15414 );
xnor \U$15039 ( \15416 , \15415 , \3512 );
and \U$15040 ( \15417 , \6210 , \3386 );
and \U$15041 ( \15418 , \5838 , \3384 );
nor \U$15042 ( \15419 , \15417 , \15418 );
xnor \U$15043 ( \15420 , \15419 , \3181 );
and \U$15044 ( \15421 , \15416 , \15420 );
and \U$15045 ( \15422 , \6562 , \2980 );
and \U$15046 ( \15423 , \6219 , \2978 );
nor \U$15047 ( \15424 , \15422 , \15423 );
xnor \U$15048 ( \15425 , \15424 , \2831 );
and \U$15049 ( \15426 , \15420 , \15425 );
and \U$15050 ( \15427 , \15416 , \15425 );
or \U$15051 ( \15428 , \15421 , \15426 , \15427 );
and \U$15052 ( \15429 , \15411 , \15428 );
and \U$15053 ( \15430 , \15395 , \15428 );
or \U$15054 ( \15431 , \15412 , \15429 , \15430 );
and \U$15055 ( \15432 , \15378 , \15431 );
and \U$15056 ( \15433 , \15338 , \15431 );
or \U$15057 ( \15434 , \15379 , \15432 , \15433 );
xor \U$15058 ( \15435 , \15152 , \15156 );
xor \U$15059 ( \15436 , \15435 , \15161 );
xor \U$15060 ( \15437 , \15132 , \15136 );
xor \U$15061 ( \15438 , \15437 , \15141 );
and \U$15062 ( \15439 , \15436 , \15438 );
xor \U$15063 ( \15440 , \15168 , \15172 );
xor \U$15064 ( \15441 , \15440 , \15177 );
and \U$15065 ( \15442 , \15438 , \15441 );
and \U$15066 ( \15443 , \15436 , \15441 );
or \U$15067 ( \15444 , \15439 , \15442 , \15443 );
xor \U$15068 ( \15445 , \15099 , \15103 );
xor \U$15069 ( \15446 , \15445 , \15108 );
xor \U$15070 ( \15447 , \15115 , \15119 );
xor \U$15071 ( \15448 , \15447 , \15124 );
and \U$15072 ( \15449 , \15446 , \15448 );
xor \U$15073 ( \15450 , \15047 , \15051 );
xor \U$15074 ( \15451 , \15450 , \15056 );
and \U$15075 ( \15452 , \15448 , \15451 );
and \U$15076 ( \15453 , \15446 , \15451 );
or \U$15077 ( \15454 , \15449 , \15452 , \15453 );
and \U$15078 ( \15455 , \15444 , \15454 );
xor \U$15079 ( \15456 , \15063 , \15067 );
xor \U$15080 ( \15457 , \15456 , \15072 );
xor \U$15081 ( \15458 , \15080 , \15084 );
xor \U$15082 ( \15459 , \15458 , \15089 );
and \U$15083 ( \15460 , \15457 , \15459 );
and \U$15084 ( \15461 , \15454 , \15460 );
and \U$15085 ( \15462 , \15444 , \15460 );
or \U$15086 ( \15463 , \15455 , \15461 , \15462 );
and \U$15087 ( \15464 , \15434 , \15463 );
xor \U$15088 ( \15465 , \15191 , \15193 );
xor \U$15089 ( \15466 , \15465 , \15196 );
xor \U$15090 ( \15467 , \15201 , \15203 );
xor \U$15091 ( \15468 , \15467 , \15206 );
and \U$15092 ( \15469 , \15466 , \15468 );
xor \U$15093 ( \15470 , \15212 , \15214 );
and \U$15094 ( \15471 , \15468 , \15470 );
and \U$15095 ( \15472 , \15466 , \15470 );
or \U$15096 ( \15473 , \15469 , \15471 , \15472 );
and \U$15097 ( \15474 , \15463 , \15473 );
and \U$15098 ( \15475 , \15434 , \15473 );
or \U$15099 ( \15476 , \15464 , \15474 , \15475 );
xor \U$15100 ( \15477 , \15059 , \15075 );
xor \U$15101 ( \15478 , \15477 , \15092 );
xor \U$15102 ( \15479 , \15111 , \15127 );
xor \U$15103 ( \15480 , \15479 , \15144 );
and \U$15104 ( \15481 , \15478 , \15480 );
xor \U$15105 ( \15482 , \15164 , \15180 );
xor \U$15106 ( \15483 , \15482 , \15183 );
and \U$15107 ( \15484 , \15480 , \15483 );
and \U$15108 ( \15485 , \15478 , \15483 );
or \U$15109 ( \15486 , \15481 , \15484 , \15485 );
xor \U$15110 ( \15487 , \15234 , \15236 );
xor \U$15111 ( \15488 , \15487 , \15239 );
and \U$15112 ( \15489 , \15486 , \15488 );
xor \U$15113 ( \15490 , \15221 , \15223 );
xor \U$15114 ( \15491 , \15490 , \15226 );
and \U$15115 ( \15492 , \15488 , \15491 );
and \U$15116 ( \15493 , \15486 , \15491 );
or \U$15117 ( \15494 , \15489 , \15492 , \15493 );
and \U$15118 ( \15495 , \15476 , \15494 );
xor \U$15119 ( \15496 , \15253 , \15255 );
xor \U$15120 ( \15497 , \15496 , \15258 );
and \U$15121 ( \15498 , \15494 , \15497 );
and \U$15122 ( \15499 , \15476 , \15497 );
or \U$15123 ( \15500 , \15495 , \15498 , \15499 );
xor \U$15124 ( \15501 , \15232 , \15250 );
xor \U$15125 ( \15502 , \15501 , \15261 );
and \U$15126 ( \15503 , \15500 , \15502 );
xor \U$15127 ( \15504 , \15266 , \15268 );
xor \U$15128 ( \15505 , \15504 , \15270 );
and \U$15129 ( \15506 , \15502 , \15505 );
and \U$15130 ( \15507 , \15500 , \15505 );
or \U$15131 ( \15508 , \15503 , \15506 , \15507 );
xor \U$15132 ( \15509 , \14975 , \14993 );
xor \U$15133 ( \15510 , \15509 , \14999 );
and \U$15134 ( \15511 , \15508 , \15510 );
xor \U$15135 ( \15512 , \15264 , \15273 );
xor \U$15136 ( \15513 , \15512 , \15276 );
and \U$15137 ( \15514 , \15510 , \15513 );
and \U$15138 ( \15515 , \15508 , \15513 );
or \U$15139 ( \15516 , \15511 , \15514 , \15515 );
and \U$15140 ( \15517 , \15290 , \15516 );
xor \U$15141 ( \15518 , \15290 , \15516 );
xor \U$15142 ( \15519 , \15508 , \15510 );
xor \U$15143 ( \15520 , \15519 , \15513 );
xor \U$15144 ( \15521 , \15294 , \15298 );
xor \U$15145 ( \15522 , \15521 , \15303 );
xor \U$15146 ( \15523 , \15310 , \15314 );
xor \U$15147 ( \15524 , \15523 , \15319 );
and \U$15148 ( \15525 , \15522 , \15524 );
xor \U$15149 ( \15526 , \15327 , \15331 );
xor \U$15150 ( \15527 , \15526 , \964 );
and \U$15151 ( \15528 , \15524 , \15527 );
and \U$15152 ( \15529 , \15522 , \15527 );
or \U$15153 ( \15530 , \15525 , \15528 , \15529 );
nand \U$15154 ( \15531 , \11029 , \1056 );
xnor \U$15155 ( \15532 , \15531 , \964 );
xor \U$15156 ( \15533 , \15342 , \15346 );
xor \U$15157 ( \15534 , \15533 , \15351 );
and \U$15158 ( \15535 , \15532 , \15534 );
xor \U$15159 ( \15536 , \15358 , \15362 );
xor \U$15160 ( \15537 , \15536 , \15367 );
and \U$15161 ( \15538 , \15534 , \15537 );
and \U$15162 ( \15539 , \15532 , \15537 );
or \U$15163 ( \15540 , \15535 , \15538 , \15539 );
and \U$15164 ( \15541 , \15530 , \15540 );
xor \U$15165 ( \15542 , \15383 , \15387 );
xor \U$15166 ( \15543 , \15542 , \15392 );
xor \U$15167 ( \15544 , \15399 , \15403 );
xor \U$15168 ( \15545 , \15544 , \15408 );
and \U$15169 ( \15546 , \15543 , \15545 );
xor \U$15170 ( \15547 , \15416 , \15420 );
xor \U$15171 ( \15548 , \15547 , \15425 );
and \U$15172 ( \15549 , \15545 , \15548 );
and \U$15173 ( \15550 , \15543 , \15548 );
or \U$15174 ( \15551 , \15546 , \15549 , \15550 );
and \U$15175 ( \15552 , \15540 , \15551 );
and \U$15176 ( \15553 , \15530 , \15551 );
or \U$15177 ( \15554 , \15541 , \15552 , \15553 );
and \U$15178 ( \15555 , \8189 , \2362 );
and \U$15179 ( \15556 , \7765 , \2360 );
nor \U$15180 ( \15557 , \15555 , \15556 );
xnor \U$15181 ( \15558 , \15557 , \2225 );
and \U$15182 ( \15559 , \8440 , \2156 );
and \U$15183 ( \15560 , \8435 , \2154 );
nor \U$15184 ( \15561 , \15559 , \15560 );
xnor \U$15185 ( \15562 , \15561 , \2004 );
and \U$15186 ( \15563 , \15558 , \15562 );
and \U$15187 ( \15564 , \9043 , \1888 );
and \U$15188 ( \15565 , \8759 , \1886 );
nor \U$15189 ( \15566 , \15564 , \15565 );
xnor \U$15190 ( \15567 , \15566 , \1732 );
and \U$15191 ( \15568 , \15562 , \15567 );
and \U$15192 ( \15569 , \15558 , \15567 );
or \U$15193 ( \15570 , \15563 , \15568 , \15569 );
and \U$15194 ( \15571 , \9620 , \1616 );
and \U$15195 ( \15572 , \9612 , \1614 );
nor \U$15196 ( \15573 , \15571 , \15572 );
xnor \U$15197 ( \15574 , \15573 , \1503 );
and \U$15198 ( \15575 , \10228 , \1422 );
and \U$15199 ( \15576 , \10223 , \1420 );
nor \U$15200 ( \15577 , \15575 , \15576 );
xnor \U$15201 ( \15578 , \15577 , \1286 );
and \U$15202 ( \15579 , \15574 , \15578 );
and \U$15203 ( \15580 , \11029 , \1222 );
and \U$15204 ( \15581 , \10409 , \1220 );
nor \U$15205 ( \15582 , \15580 , \15581 );
xnor \U$15206 ( \15583 , \15582 , \1144 );
and \U$15207 ( \15584 , \15578 , \15583 );
and \U$15208 ( \15585 , \15574 , \15583 );
or \U$15209 ( \15586 , \15579 , \15584 , \15585 );
and \U$15210 ( \15587 , \15570 , \15586 );
and \U$15211 ( \15588 , \10409 , \1222 );
and \U$15212 ( \15589 , \10228 , \1220 );
nor \U$15213 ( \15590 , \15588 , \15589 );
xnor \U$15214 ( \15591 , \15590 , \1144 );
and \U$15215 ( \15592 , \15586 , \15591 );
and \U$15216 ( \15593 , \15570 , \15591 );
or \U$15217 ( \15594 , \15587 , \15592 , \15593 );
and \U$15218 ( \15595 , \1336 , \10876 );
and \U$15219 ( \15596 , \1248 , \10873 );
nor \U$15220 ( \15597 , \15595 , \15596 );
xnor \U$15221 ( \15598 , \15597 , \9821 );
and \U$15222 ( \15599 , \1446 , \10063 );
and \U$15223 ( \15600 , \1441 , \10061 );
nor \U$15224 ( \15601 , \15599 , \15600 );
xnor \U$15225 ( \15602 , \15601 , \9824 );
and \U$15226 ( \15603 , \15598 , \15602 );
and \U$15227 ( \15604 , \1677 , \9495 );
and \U$15228 ( \15605 , \1562 , \9493 );
nor \U$15229 ( \15606 , \15604 , \15605 );
xnor \U$15230 ( \15607 , \15606 , \9185 );
and \U$15231 ( \15608 , \15602 , \15607 );
and \U$15232 ( \15609 , \15598 , \15607 );
or \U$15233 ( \15610 , \15603 , \15608 , \15609 );
and \U$15234 ( \15611 , \1861 , \8958 );
and \U$15235 ( \15612 , \1853 , \8956 );
nor \U$15236 ( \15613 , \15611 , \15612 );
xnor \U$15237 ( \15614 , \15613 , \8587 );
and \U$15238 ( \15615 , \2109 , \8396 );
and \U$15239 ( \15616 , \2104 , \8394 );
nor \U$15240 ( \15617 , \15615 , \15616 );
xnor \U$15241 ( \15618 , \15617 , \8078 );
and \U$15242 ( \15619 , \15614 , \15618 );
and \U$15243 ( \15620 , \2439 , \7829 );
and \U$15244 ( \15621 , \2295 , \7827 );
nor \U$15245 ( \15622 , \15620 , \15621 );
xnor \U$15246 ( \15623 , \15622 , \7580 );
and \U$15247 ( \15624 , \15618 , \15623 );
and \U$15248 ( \15625 , \15614 , \15623 );
or \U$15249 ( \15626 , \15619 , \15624 , \15625 );
and \U$15250 ( \15627 , \15610 , \15626 );
and \U$15251 ( \15628 , \2728 , \7300 );
and \U$15252 ( \15629 , \2703 , \7298 );
nor \U$15253 ( \15630 , \15628 , \15629 );
xnor \U$15254 ( \15631 , \15630 , \7040 );
and \U$15255 ( \15632 , \3069 , \6806 );
and \U$15256 ( \15633 , \2902 , \6804 );
nor \U$15257 ( \15634 , \15632 , \15633 );
xnor \U$15258 ( \15635 , \15634 , \6491 );
and \U$15259 ( \15636 , \15631 , \15635 );
and \U$15260 ( \15637 , \3326 , \6297 );
and \U$15261 ( \15638 , \3207 , \6295 );
nor \U$15262 ( \15639 , \15637 , \15638 );
xnor \U$15263 ( \15640 , \15639 , \5957 );
and \U$15264 ( \15641 , \15635 , \15640 );
and \U$15265 ( \15642 , \15631 , \15640 );
or \U$15266 ( \15643 , \15636 , \15641 , \15642 );
and \U$15267 ( \15644 , \15626 , \15643 );
and \U$15268 ( \15645 , \15610 , \15643 );
or \U$15269 ( \15646 , \15627 , \15644 , \15645 );
and \U$15270 ( \15647 , \15594 , \15646 );
and \U$15271 ( \15648 , \4841 , \4417 );
and \U$15272 ( \15649 , \4833 , \4415 );
nor \U$15273 ( \15650 , \15648 , \15649 );
xnor \U$15274 ( \15651 , \15650 , \4274 );
and \U$15275 ( \15652 , \5315 , \4094 );
and \U$15276 ( \15653 , \5310 , \4092 );
nor \U$15277 ( \15654 , \15652 , \15653 );
xnor \U$15278 ( \15655 , \15654 , \3848 );
and \U$15279 ( \15656 , \15651 , \15655 );
and \U$15280 ( \15657 , \5838 , \3699 );
and \U$15281 ( \15658 , \5579 , \3697 );
nor \U$15282 ( \15659 , \15657 , \15658 );
xnor \U$15283 ( \15660 , \15659 , \3512 );
and \U$15284 ( \15661 , \15655 , \15660 );
and \U$15285 ( \15662 , \15651 , \15660 );
or \U$15286 ( \15663 , \15656 , \15661 , \15662 );
and \U$15287 ( \15664 , \6219 , \3386 );
and \U$15288 ( \15665 , \6210 , \3384 );
nor \U$15289 ( \15666 , \15664 , \15665 );
xnor \U$15290 ( \15667 , \15666 , \3181 );
and \U$15291 ( \15668 , \6764 , \2980 );
and \U$15292 ( \15669 , \6562 , \2978 );
nor \U$15293 ( \15670 , \15668 , \15669 );
xnor \U$15294 ( \15671 , \15670 , \2831 );
and \U$15295 ( \15672 , \15667 , \15671 );
and \U$15296 ( \15673 , \7239 , \2658 );
and \U$15297 ( \15674 , \7067 , \2656 );
nor \U$15298 ( \15675 , \15673 , \15674 );
xnor \U$15299 ( \15676 , \15675 , \2516 );
and \U$15300 ( \15677 , \15671 , \15676 );
and \U$15301 ( \15678 , \15667 , \15676 );
or \U$15302 ( \15679 , \15672 , \15677 , \15678 );
and \U$15303 ( \15680 , \15663 , \15679 );
and \U$15304 ( \15681 , \3951 , \5708 );
and \U$15305 ( \15682 , \3743 , \5706 );
nor \U$15306 ( \15683 , \15681 , \15682 );
xnor \U$15307 ( \15684 , \15683 , \5467 );
and \U$15308 ( \15685 , \4078 , \5242 );
and \U$15309 ( \15686 , \4073 , \5240 );
nor \U$15310 ( \15687 , \15685 , \15686 );
xnor \U$15311 ( \15688 , \15687 , \5054 );
and \U$15312 ( \15689 , \15684 , \15688 );
and \U$15313 ( \15690 , \4531 , \4868 );
and \U$15314 ( \15691 , \4334 , \4866 );
nor \U$15315 ( \15692 , \15690 , \15691 );
xnor \U$15316 ( \15693 , \15692 , \4636 );
and \U$15317 ( \15694 , \15688 , \15693 );
and \U$15318 ( \15695 , \15684 , \15693 );
or \U$15319 ( \15696 , \15689 , \15694 , \15695 );
and \U$15320 ( \15697 , \15679 , \15696 );
and \U$15321 ( \15698 , \15663 , \15696 );
or \U$15322 ( \15699 , \15680 , \15697 , \15698 );
and \U$15323 ( \15700 , \15646 , \15699 );
and \U$15324 ( \15701 , \15594 , \15699 );
or \U$15325 ( \15702 , \15647 , \15700 , \15701 );
and \U$15326 ( \15703 , \15554 , \15702 );
xor \U$15327 ( \15704 , \15436 , \15438 );
xor \U$15328 ( \15705 , \15704 , \15441 );
xor \U$15329 ( \15706 , \15446 , \15448 );
xor \U$15330 ( \15707 , \15706 , \15451 );
and \U$15331 ( \15708 , \15705 , \15707 );
xor \U$15332 ( \15709 , \15457 , \15459 );
and \U$15333 ( \15710 , \15707 , \15709 );
and \U$15334 ( \15711 , \15705 , \15709 );
or \U$15335 ( \15712 , \15708 , \15710 , \15711 );
and \U$15336 ( \15713 , \15702 , \15712 );
and \U$15337 ( \15714 , \15554 , \15712 );
or \U$15338 ( \15715 , \15703 , \15713 , \15714 );
xor \U$15339 ( \15716 , \15306 , \15322 );
xor \U$15340 ( \15717 , \15716 , \15335 );
xor \U$15341 ( \15718 , \15354 , \15370 );
xor \U$15342 ( \15719 , \15718 , \15375 );
and \U$15343 ( \15720 , \15717 , \15719 );
xor \U$15344 ( \15721 , \15395 , \15411 );
xor \U$15345 ( \15722 , \15721 , \15428 );
and \U$15346 ( \15723 , \15719 , \15722 );
and \U$15347 ( \15724 , \15717 , \15722 );
or \U$15348 ( \15725 , \15720 , \15723 , \15724 );
xor \U$15349 ( \15726 , \15478 , \15480 );
xor \U$15350 ( \15727 , \15726 , \15483 );
and \U$15351 ( \15728 , \15725 , \15727 );
xor \U$15352 ( \15729 , \15466 , \15468 );
xor \U$15353 ( \15730 , \15729 , \15470 );
and \U$15354 ( \15731 , \15727 , \15730 );
and \U$15355 ( \15732 , \15725 , \15730 );
or \U$15356 ( \15733 , \15728 , \15731 , \15732 );
and \U$15357 ( \15734 , \15715 , \15733 );
xor \U$15358 ( \15735 , \15199 , \15209 );
xor \U$15359 ( \15736 , \15735 , \15215 );
and \U$15360 ( \15737 , \15733 , \15736 );
and \U$15361 ( \15738 , \15715 , \15736 );
or \U$15362 ( \15739 , \15734 , \15737 , \15738 );
xor \U$15363 ( \15740 , \15095 , \15147 );
xor \U$15364 ( \15741 , \15740 , \15186 );
xor \U$15365 ( \15742 , \15434 , \15463 );
xor \U$15366 ( \15743 , \15742 , \15473 );
and \U$15367 ( \15744 , \15741 , \15743 );
xor \U$15368 ( \15745 , \15486 , \15488 );
xor \U$15369 ( \15746 , \15745 , \15491 );
and \U$15370 ( \15747 , \15743 , \15746 );
and \U$15371 ( \15748 , \15741 , \15746 );
or \U$15372 ( \15749 , \15744 , \15747 , \15748 );
and \U$15373 ( \15750 , \15739 , \15749 );
xor \U$15374 ( \15751 , \15242 , \15244 );
xor \U$15375 ( \15752 , \15751 , \15247 );
and \U$15376 ( \15753 , \15749 , \15752 );
and \U$15377 ( \15754 , \15739 , \15752 );
or \U$15378 ( \15755 , \15750 , \15753 , \15754 );
xor \U$15379 ( \15756 , \15189 , \15218 );
xor \U$15380 ( \15757 , \15756 , \15229 );
xor \U$15381 ( \15758 , \15476 , \15494 );
xor \U$15382 ( \15759 , \15758 , \15497 );
and \U$15383 ( \15760 , \15757 , \15759 );
and \U$15384 ( \15761 , \15755 , \15760 );
xor \U$15385 ( \15762 , \15500 , \15502 );
xor \U$15386 ( \15763 , \15762 , \15505 );
and \U$15387 ( \15764 , \15760 , \15763 );
and \U$15388 ( \15765 , \15755 , \15763 );
or \U$15389 ( \15766 , \15761 , \15764 , \15765 );
and \U$15390 ( \15767 , \15520 , \15766 );
xor \U$15391 ( \15768 , \15520 , \15766 );
xor \U$15392 ( \15769 , \15755 , \15760 );
xor \U$15393 ( \15770 , \15769 , \15763 );
and \U$15394 ( \15771 , \6210 , \3699 );
and \U$15395 ( \15772 , \5838 , \3697 );
nor \U$15396 ( \15773 , \15771 , \15772 );
xnor \U$15397 ( \15774 , \15773 , \3512 );
and \U$15398 ( \15775 , \6562 , \3386 );
and \U$15399 ( \15776 , \6219 , \3384 );
nor \U$15400 ( \15777 , \15775 , \15776 );
xnor \U$15401 ( \15778 , \15777 , \3181 );
and \U$15402 ( \15779 , \15774 , \15778 );
and \U$15403 ( \15780 , \7067 , \2980 );
and \U$15404 ( \15781 , \6764 , \2978 );
nor \U$15405 ( \15782 , \15780 , \15781 );
xnor \U$15406 ( \15783 , \15782 , \2831 );
and \U$15407 ( \15784 , \15778 , \15783 );
and \U$15408 ( \15785 , \15774 , \15783 );
or \U$15409 ( \15786 , \15779 , \15784 , \15785 );
and \U$15410 ( \15787 , \4833 , \4868 );
and \U$15411 ( \15788 , \4531 , \4866 );
nor \U$15412 ( \15789 , \15787 , \15788 );
xnor \U$15413 ( \15790 , \15789 , \4636 );
and \U$15414 ( \15791 , \5310 , \4417 );
and \U$15415 ( \15792 , \4841 , \4415 );
nor \U$15416 ( \15793 , \15791 , \15792 );
xnor \U$15417 ( \15794 , \15793 , \4274 );
and \U$15418 ( \15795 , \15790 , \15794 );
and \U$15419 ( \15796 , \5579 , \4094 );
and \U$15420 ( \15797 , \5315 , \4092 );
nor \U$15421 ( \15798 , \15796 , \15797 );
xnor \U$15422 ( \15799 , \15798 , \3848 );
and \U$15423 ( \15800 , \15794 , \15799 );
and \U$15424 ( \15801 , \15790 , \15799 );
or \U$15425 ( \15802 , \15795 , \15800 , \15801 );
and \U$15426 ( \15803 , \15786 , \15802 );
and \U$15427 ( \15804 , \3743 , \6297 );
and \U$15428 ( \15805 , \3326 , \6295 );
nor \U$15429 ( \15806 , \15804 , \15805 );
xnor \U$15430 ( \15807 , \15806 , \5957 );
and \U$15431 ( \15808 , \4073 , \5708 );
and \U$15432 ( \15809 , \3951 , \5706 );
nor \U$15433 ( \15810 , \15808 , \15809 );
xnor \U$15434 ( \15811 , \15810 , \5467 );
and \U$15435 ( \15812 , \15807 , \15811 );
and \U$15436 ( \15813 , \4334 , \5242 );
and \U$15437 ( \15814 , \4078 , \5240 );
nor \U$15438 ( \15815 , \15813 , \15814 );
xnor \U$15439 ( \15816 , \15815 , \5054 );
and \U$15440 ( \15817 , \15811 , \15816 );
and \U$15441 ( \15818 , \15807 , \15816 );
or \U$15442 ( \15819 , \15812 , \15817 , \15818 );
and \U$15443 ( \15820 , \15802 , \15819 );
and \U$15444 ( \15821 , \15786 , \15819 );
or \U$15445 ( \15822 , \15803 , \15820 , \15821 );
and \U$15446 ( \15823 , \1853 , \9495 );
and \U$15447 ( \15824 , \1677 , \9493 );
nor \U$15448 ( \15825 , \15823 , \15824 );
xnor \U$15449 ( \15826 , \15825 , \9185 );
and \U$15450 ( \15827 , \2104 , \8958 );
and \U$15451 ( \15828 , \1861 , \8956 );
nor \U$15452 ( \15829 , \15827 , \15828 );
xnor \U$15453 ( \15830 , \15829 , \8587 );
and \U$15454 ( \15831 , \15826 , \15830 );
and \U$15455 ( \15832 , \2295 , \8396 );
and \U$15456 ( \15833 , \2109 , \8394 );
nor \U$15457 ( \15834 , \15832 , \15833 );
xnor \U$15458 ( \15835 , \15834 , \8078 );
and \U$15459 ( \15836 , \15830 , \15835 );
and \U$15460 ( \15837 , \15826 , \15835 );
or \U$15461 ( \15838 , \15831 , \15836 , \15837 );
and \U$15462 ( \15839 , \1441 , \10876 );
and \U$15463 ( \15840 , \1336 , \10873 );
nor \U$15464 ( \15841 , \15839 , \15840 );
xnor \U$15465 ( \15842 , \15841 , \9821 );
and \U$15466 ( \15843 , \1562 , \10063 );
and \U$15467 ( \15844 , \1446 , \10061 );
nor \U$15468 ( \15845 , \15843 , \15844 );
xnor \U$15469 ( \15846 , \15845 , \9824 );
and \U$15470 ( \15847 , \15842 , \15846 );
and \U$15471 ( \15848 , \15846 , \1144 );
and \U$15472 ( \15849 , \15842 , \1144 );
or \U$15473 ( \15850 , \15847 , \15848 , \15849 );
and \U$15474 ( \15851 , \15838 , \15850 );
and \U$15475 ( \15852 , \2703 , \7829 );
and \U$15476 ( \15853 , \2439 , \7827 );
nor \U$15477 ( \15854 , \15852 , \15853 );
xnor \U$15478 ( \15855 , \15854 , \7580 );
and \U$15479 ( \15856 , \2902 , \7300 );
and \U$15480 ( \15857 , \2728 , \7298 );
nor \U$15481 ( \15858 , \15856 , \15857 );
xnor \U$15482 ( \15859 , \15858 , \7040 );
and \U$15483 ( \15860 , \15855 , \15859 );
and \U$15484 ( \15861 , \3207 , \6806 );
and \U$15485 ( \15862 , \3069 , \6804 );
nor \U$15486 ( \15863 , \15861 , \15862 );
xnor \U$15487 ( \15864 , \15863 , \6491 );
and \U$15488 ( \15865 , \15859 , \15864 );
and \U$15489 ( \15866 , \15855 , \15864 );
or \U$15490 ( \15867 , \15860 , \15865 , \15866 );
and \U$15491 ( \15868 , \15850 , \15867 );
and \U$15492 ( \15869 , \15838 , \15867 );
or \U$15493 ( \15870 , \15851 , \15868 , \15869 );
and \U$15494 ( \15871 , \15822 , \15870 );
and \U$15495 ( \15872 , \7765 , \2658 );
and \U$15496 ( \15873 , \7239 , \2656 );
nor \U$15497 ( \15874 , \15872 , \15873 );
xnor \U$15498 ( \15875 , \15874 , \2516 );
and \U$15499 ( \15876 , \8435 , \2362 );
and \U$15500 ( \15877 , \8189 , \2360 );
nor \U$15501 ( \15878 , \15876 , \15877 );
xnor \U$15502 ( \15879 , \15878 , \2225 );
and \U$15503 ( \15880 , \15875 , \15879 );
and \U$15504 ( \15881 , \8759 , \2156 );
and \U$15505 ( \15882 , \8440 , \2154 );
nor \U$15506 ( \15883 , \15881 , \15882 );
xnor \U$15507 ( \15884 , \15883 , \2004 );
and \U$15508 ( \15885 , \15879 , \15884 );
and \U$15509 ( \15886 , \15875 , \15884 );
or \U$15510 ( \15887 , \15880 , \15885 , \15886 );
and \U$15511 ( \15888 , \9612 , \1888 );
and \U$15512 ( \15889 , \9043 , \1886 );
nor \U$15513 ( \15890 , \15888 , \15889 );
xnor \U$15514 ( \15891 , \15890 , \1732 );
and \U$15515 ( \15892 , \10223 , \1616 );
and \U$15516 ( \15893 , \9620 , \1614 );
nor \U$15517 ( \15894 , \15892 , \15893 );
xnor \U$15518 ( \15895 , \15894 , \1503 );
and \U$15519 ( \15896 , \15891 , \15895 );
and \U$15520 ( \15897 , \10409 , \1422 );
and \U$15521 ( \15898 , \10228 , \1420 );
nor \U$15522 ( \15899 , \15897 , \15898 );
xnor \U$15523 ( \15900 , \15899 , \1286 );
and \U$15524 ( \15901 , \15895 , \15900 );
and \U$15525 ( \15902 , \15891 , \15900 );
or \U$15526 ( \15903 , \15896 , \15901 , \15902 );
and \U$15527 ( \15904 , \15887 , \15903 );
xor \U$15528 ( \15905 , \15574 , \15578 );
xor \U$15529 ( \15906 , \15905 , \15583 );
and \U$15530 ( \15907 , \15903 , \15906 );
and \U$15531 ( \15908 , \15887 , \15906 );
or \U$15532 ( \15909 , \15904 , \15907 , \15908 );
and \U$15533 ( \15910 , \15870 , \15909 );
and \U$15534 ( \15911 , \15822 , \15909 );
or \U$15535 ( \15912 , \15871 , \15910 , \15911 );
xor \U$15536 ( \15913 , \15558 , \15562 );
xor \U$15537 ( \15914 , \15913 , \15567 );
xor \U$15538 ( \15915 , \15651 , \15655 );
xor \U$15539 ( \15916 , \15915 , \15660 );
and \U$15540 ( \15917 , \15914 , \15916 );
xor \U$15541 ( \15918 , \15667 , \15671 );
xor \U$15542 ( \15919 , \15918 , \15676 );
and \U$15543 ( \15920 , \15916 , \15919 );
and \U$15544 ( \15921 , \15914 , \15919 );
or \U$15545 ( \15922 , \15917 , \15920 , \15921 );
xor \U$15546 ( \15923 , \15614 , \15618 );
xor \U$15547 ( \15924 , \15923 , \15623 );
xor \U$15548 ( \15925 , \15684 , \15688 );
xor \U$15549 ( \15926 , \15925 , \15693 );
and \U$15550 ( \15927 , \15924 , \15926 );
xor \U$15551 ( \15928 , \15631 , \15635 );
xor \U$15552 ( \15929 , \15928 , \15640 );
and \U$15553 ( \15930 , \15926 , \15929 );
and \U$15554 ( \15931 , \15924 , \15929 );
or \U$15555 ( \15932 , \15927 , \15930 , \15931 );
and \U$15556 ( \15933 , \15922 , \15932 );
xor \U$15557 ( \15934 , \15522 , \15524 );
xor \U$15558 ( \15935 , \15934 , \15527 );
and \U$15559 ( \15936 , \15932 , \15935 );
and \U$15560 ( \15937 , \15922 , \15935 );
or \U$15561 ( \15938 , \15933 , \15936 , \15937 );
and \U$15562 ( \15939 , \15912 , \15938 );
xor \U$15563 ( \15940 , \15570 , \15586 );
xor \U$15564 ( \15941 , \15940 , \15591 );
xor \U$15565 ( \15942 , \15532 , \15534 );
xor \U$15566 ( \15943 , \15942 , \15537 );
and \U$15567 ( \15944 , \15941 , \15943 );
xor \U$15568 ( \15945 , \15543 , \15545 );
xor \U$15569 ( \15946 , \15945 , \15548 );
and \U$15570 ( \15947 , \15943 , \15946 );
and \U$15571 ( \15948 , \15941 , \15946 );
or \U$15572 ( \15949 , \15944 , \15947 , \15948 );
and \U$15573 ( \15950 , \15938 , \15949 );
and \U$15574 ( \15951 , \15912 , \15949 );
or \U$15575 ( \15952 , \15939 , \15950 , \15951 );
xor \U$15576 ( \15953 , \15530 , \15540 );
xor \U$15577 ( \15954 , \15953 , \15551 );
xor \U$15578 ( \15955 , \15717 , \15719 );
xor \U$15579 ( \15956 , \15955 , \15722 );
and \U$15580 ( \15957 , \15954 , \15956 );
xor \U$15581 ( \15958 , \15705 , \15707 );
xor \U$15582 ( \15959 , \15958 , \15709 );
and \U$15583 ( \15960 , \15956 , \15959 );
and \U$15584 ( \15961 , \15954 , \15959 );
or \U$15585 ( \15962 , \15957 , \15960 , \15961 );
and \U$15586 ( \15963 , \15952 , \15962 );
xor \U$15587 ( \15964 , \15444 , \15454 );
xor \U$15588 ( \15965 , \15964 , \15460 );
and \U$15589 ( \15966 , \15962 , \15965 );
and \U$15590 ( \15967 , \15952 , \15965 );
or \U$15591 ( \15968 , \15963 , \15966 , \15967 );
xor \U$15592 ( \15969 , \15338 , \15378 );
xor \U$15593 ( \15970 , \15969 , \15431 );
xor \U$15594 ( \15971 , \15554 , \15702 );
xor \U$15595 ( \15972 , \15971 , \15712 );
and \U$15596 ( \15973 , \15970 , \15972 );
xor \U$15597 ( \15974 , \15725 , \15727 );
xor \U$15598 ( \15975 , \15974 , \15730 );
and \U$15599 ( \15976 , \15972 , \15975 );
and \U$15600 ( \15977 , \15970 , \15975 );
or \U$15601 ( \15978 , \15973 , \15976 , \15977 );
and \U$15602 ( \15979 , \15968 , \15978 );
xor \U$15603 ( \15980 , \15741 , \15743 );
xor \U$15604 ( \15981 , \15980 , \15746 );
and \U$15605 ( \15982 , \15978 , \15981 );
and \U$15606 ( \15983 , \15968 , \15981 );
or \U$15607 ( \15984 , \15979 , \15982 , \15983 );
xor \U$15608 ( \15985 , \15739 , \15749 );
xor \U$15609 ( \15986 , \15985 , \15752 );
and \U$15610 ( \15987 , \15984 , \15986 );
xor \U$15611 ( \15988 , \15757 , \15759 );
and \U$15612 ( \15989 , \15986 , \15988 );
and \U$15613 ( \15990 , \15984 , \15988 );
or \U$15614 ( \15991 , \15987 , \15989 , \15990 );
and \U$15615 ( \15992 , \15770 , \15991 );
xor \U$15616 ( \15993 , \15770 , \15991 );
xor \U$15617 ( \15994 , \15984 , \15986 );
xor \U$15618 ( \15995 , \15994 , \15988 );
and \U$15619 ( \15996 , \4078 , \5708 );
and \U$15620 ( \15997 , \4073 , \5706 );
nor \U$15621 ( \15998 , \15996 , \15997 );
xnor \U$15622 ( \15999 , \15998 , \5467 );
and \U$15623 ( \16000 , \4531 , \5242 );
and \U$15624 ( \16001 , \4334 , \5240 );
nor \U$15625 ( \16002 , \16000 , \16001 );
xnor \U$15626 ( \16003 , \16002 , \5054 );
and \U$15627 ( \16004 , \15999 , \16003 );
and \U$15628 ( \16005 , \4841 , \4868 );
and \U$15629 ( \16006 , \4833 , \4866 );
nor \U$15630 ( \16007 , \16005 , \16006 );
xnor \U$15631 ( \16008 , \16007 , \4636 );
and \U$15632 ( \16009 , \16003 , \16008 );
and \U$15633 ( \16010 , \15999 , \16008 );
or \U$15634 ( \16011 , \16004 , \16009 , \16010 );
and \U$15635 ( \16012 , \5315 , \4417 );
and \U$15636 ( \16013 , \5310 , \4415 );
nor \U$15637 ( \16014 , \16012 , \16013 );
xnor \U$15638 ( \16015 , \16014 , \4274 );
and \U$15639 ( \16016 , \5838 , \4094 );
and \U$15640 ( \16017 , \5579 , \4092 );
nor \U$15641 ( \16018 , \16016 , \16017 );
xnor \U$15642 ( \16019 , \16018 , \3848 );
and \U$15643 ( \16020 , \16015 , \16019 );
and \U$15644 ( \16021 , \6219 , \3699 );
and \U$15645 ( \16022 , \6210 , \3697 );
nor \U$15646 ( \16023 , \16021 , \16022 );
xnor \U$15647 ( \16024 , \16023 , \3512 );
and \U$15648 ( \16025 , \16019 , \16024 );
and \U$15649 ( \16026 , \16015 , \16024 );
or \U$15650 ( \16027 , \16020 , \16025 , \16026 );
and \U$15651 ( \16028 , \16011 , \16027 );
and \U$15652 ( \16029 , \6764 , \3386 );
and \U$15653 ( \16030 , \6562 , \3384 );
nor \U$15654 ( \16031 , \16029 , \16030 );
xnor \U$15655 ( \16032 , \16031 , \3181 );
and \U$15656 ( \16033 , \7239 , \2980 );
and \U$15657 ( \16034 , \7067 , \2978 );
nor \U$15658 ( \16035 , \16033 , \16034 );
xnor \U$15659 ( \16036 , \16035 , \2831 );
and \U$15660 ( \16037 , \16032 , \16036 );
and \U$15661 ( \16038 , \8189 , \2658 );
and \U$15662 ( \16039 , \7765 , \2656 );
nor \U$15663 ( \16040 , \16038 , \16039 );
xnor \U$15664 ( \16041 , \16040 , \2516 );
and \U$15665 ( \16042 , \16036 , \16041 );
and \U$15666 ( \16043 , \16032 , \16041 );
or \U$15667 ( \16044 , \16037 , \16042 , \16043 );
and \U$15668 ( \16045 , \16027 , \16044 );
and \U$15669 ( \16046 , \16011 , \16044 );
or \U$15670 ( \16047 , \16028 , \16045 , \16046 );
and \U$15671 ( \16048 , \2109 , \8958 );
and \U$15672 ( \16049 , \2104 , \8956 );
nor \U$15673 ( \16050 , \16048 , \16049 );
xnor \U$15674 ( \16051 , \16050 , \8587 );
and \U$15675 ( \16052 , \2439 , \8396 );
and \U$15676 ( \16053 , \2295 , \8394 );
nor \U$15677 ( \16054 , \16052 , \16053 );
xnor \U$15678 ( \16055 , \16054 , \8078 );
and \U$15679 ( \16056 , \16051 , \16055 );
and \U$15680 ( \16057 , \2728 , \7829 );
and \U$15681 ( \16058 , \2703 , \7827 );
nor \U$15682 ( \16059 , \16057 , \16058 );
xnor \U$15683 ( \16060 , \16059 , \7580 );
and \U$15684 ( \16061 , \16055 , \16060 );
and \U$15685 ( \16062 , \16051 , \16060 );
or \U$15686 ( \16063 , \16056 , \16061 , \16062 );
and \U$15687 ( \16064 , \3069 , \7300 );
and \U$15688 ( \16065 , \2902 , \7298 );
nor \U$15689 ( \16066 , \16064 , \16065 );
xnor \U$15690 ( \16067 , \16066 , \7040 );
and \U$15691 ( \16068 , \3326 , \6806 );
and \U$15692 ( \16069 , \3207 , \6804 );
nor \U$15693 ( \16070 , \16068 , \16069 );
xnor \U$15694 ( \16071 , \16070 , \6491 );
and \U$15695 ( \16072 , \16067 , \16071 );
and \U$15696 ( \16073 , \3951 , \6297 );
and \U$15697 ( \16074 , \3743 , \6295 );
nor \U$15698 ( \16075 , \16073 , \16074 );
xnor \U$15699 ( \16076 , \16075 , \5957 );
and \U$15700 ( \16077 , \16071 , \16076 );
and \U$15701 ( \16078 , \16067 , \16076 );
or \U$15702 ( \16079 , \16072 , \16077 , \16078 );
and \U$15703 ( \16080 , \16063 , \16079 );
and \U$15704 ( \16081 , \1446 , \10876 );
and \U$15705 ( \16082 , \1441 , \10873 );
nor \U$15706 ( \16083 , \16081 , \16082 );
xnor \U$15707 ( \16084 , \16083 , \9821 );
and \U$15708 ( \16085 , \1677 , \10063 );
and \U$15709 ( \16086 , \1562 , \10061 );
nor \U$15710 ( \16087 , \16085 , \16086 );
xnor \U$15711 ( \16088 , \16087 , \9824 );
and \U$15712 ( \16089 , \16084 , \16088 );
and \U$15713 ( \16090 , \1861 , \9495 );
and \U$15714 ( \16091 , \1853 , \9493 );
nor \U$15715 ( \16092 , \16090 , \16091 );
xnor \U$15716 ( \16093 , \16092 , \9185 );
and \U$15717 ( \16094 , \16088 , \16093 );
and \U$15718 ( \16095 , \16084 , \16093 );
or \U$15719 ( \16096 , \16089 , \16094 , \16095 );
and \U$15720 ( \16097 , \16079 , \16096 );
and \U$15721 ( \16098 , \16063 , \16096 );
or \U$15722 ( \16099 , \16080 , \16097 , \16098 );
and \U$15723 ( \16100 , \16047 , \16099 );
and \U$15724 ( \16101 , \8440 , \2362 );
and \U$15725 ( \16102 , \8435 , \2360 );
nor \U$15726 ( \16103 , \16101 , \16102 );
xnor \U$15727 ( \16104 , \16103 , \2225 );
and \U$15728 ( \16105 , \9043 , \2156 );
and \U$15729 ( \16106 , \8759 , \2154 );
nor \U$15730 ( \16107 , \16105 , \16106 );
xnor \U$15731 ( \16108 , \16107 , \2004 );
and \U$15732 ( \16109 , \16104 , \16108 );
and \U$15733 ( \16110 , \9620 , \1888 );
and \U$15734 ( \16111 , \9612 , \1886 );
nor \U$15735 ( \16112 , \16110 , \16111 );
xnor \U$15736 ( \16113 , \16112 , \1732 );
and \U$15737 ( \16114 , \16108 , \16113 );
and \U$15738 ( \16115 , \16104 , \16113 );
or \U$15739 ( \16116 , \16109 , \16114 , \16115 );
nand \U$15740 ( \16117 , \11029 , \1220 );
xnor \U$15741 ( \16118 , \16117 , \1144 );
and \U$15742 ( \16119 , \16116 , \16118 );
xor \U$15743 ( \16120 , \15891 , \15895 );
xor \U$15744 ( \16121 , \16120 , \15900 );
and \U$15745 ( \16122 , \16118 , \16121 );
and \U$15746 ( \16123 , \16116 , \16121 );
or \U$15747 ( \16124 , \16119 , \16122 , \16123 );
and \U$15748 ( \16125 , \16099 , \16124 );
and \U$15749 ( \16126 , \16047 , \16124 );
or \U$15750 ( \16127 , \16100 , \16125 , \16126 );
xor \U$15751 ( \16128 , \15774 , \15778 );
xor \U$15752 ( \16129 , \16128 , \15783 );
xor \U$15753 ( \16130 , \15875 , \15879 );
xor \U$15754 ( \16131 , \16130 , \15884 );
and \U$15755 ( \16132 , \16129 , \16131 );
xor \U$15756 ( \16133 , \15790 , \15794 );
xor \U$15757 ( \16134 , \16133 , \15799 );
and \U$15758 ( \16135 , \16131 , \16134 );
and \U$15759 ( \16136 , \16129 , \16134 );
or \U$15760 ( \16137 , \16132 , \16135 , \16136 );
xor \U$15761 ( \16138 , \15826 , \15830 );
xor \U$15762 ( \16139 , \16138 , \15835 );
xor \U$15763 ( \16140 , \15807 , \15811 );
xor \U$15764 ( \16141 , \16140 , \15816 );
and \U$15765 ( \16142 , \16139 , \16141 );
xor \U$15766 ( \16143 , \15855 , \15859 );
xor \U$15767 ( \16144 , \16143 , \15864 );
and \U$15768 ( \16145 , \16141 , \16144 );
and \U$15769 ( \16146 , \16139 , \16144 );
or \U$15770 ( \16147 , \16142 , \16145 , \16146 );
and \U$15771 ( \16148 , \16137 , \16147 );
xor \U$15772 ( \16149 , \15598 , \15602 );
xor \U$15773 ( \16150 , \16149 , \15607 );
and \U$15774 ( \16151 , \16147 , \16150 );
and \U$15775 ( \16152 , \16137 , \16150 );
or \U$15776 ( \16153 , \16148 , \16151 , \16152 );
and \U$15777 ( \16154 , \16127 , \16153 );
xor \U$15778 ( \16155 , \15914 , \15916 );
xor \U$15779 ( \16156 , \16155 , \15919 );
xor \U$15780 ( \16157 , \15924 , \15926 );
xor \U$15781 ( \16158 , \16157 , \15929 );
and \U$15782 ( \16159 , \16156 , \16158 );
xor \U$15783 ( \16160 , \15887 , \15903 );
xor \U$15784 ( \16161 , \16160 , \15906 );
and \U$15785 ( \16162 , \16158 , \16161 );
and \U$15786 ( \16163 , \16156 , \16161 );
or \U$15787 ( \16164 , \16159 , \16162 , \16163 );
and \U$15788 ( \16165 , \16153 , \16164 );
and \U$15789 ( \16166 , \16127 , \16164 );
or \U$15790 ( \16167 , \16154 , \16165 , \16166 );
xor \U$15791 ( \16168 , \15610 , \15626 );
xor \U$15792 ( \16169 , \16168 , \15643 );
xor \U$15793 ( \16170 , \15663 , \15679 );
xor \U$15794 ( \16171 , \16170 , \15696 );
and \U$15795 ( \16172 , \16169 , \16171 );
xor \U$15796 ( \16173 , \15941 , \15943 );
xor \U$15797 ( \16174 , \16173 , \15946 );
and \U$15798 ( \16175 , \16171 , \16174 );
and \U$15799 ( \16176 , \16169 , \16174 );
or \U$15800 ( \16177 , \16172 , \16175 , \16176 );
and \U$15801 ( \16178 , \16167 , \16177 );
xor \U$15802 ( \16179 , \15822 , \15870 );
xor \U$15803 ( \16180 , \16179 , \15909 );
xor \U$15804 ( \16181 , \15922 , \15932 );
xor \U$15805 ( \16182 , \16181 , \15935 );
and \U$15806 ( \16183 , \16180 , \16182 );
and \U$15807 ( \16184 , \16177 , \16183 );
and \U$15808 ( \16185 , \16167 , \16183 );
or \U$15809 ( \16186 , \16178 , \16184 , \16185 );
xor \U$15810 ( \16187 , \15594 , \15646 );
xor \U$15811 ( \16188 , \16187 , \15699 );
xor \U$15812 ( \16189 , \15912 , \15938 );
xor \U$15813 ( \16190 , \16189 , \15949 );
and \U$15814 ( \16191 , \16188 , \16190 );
xor \U$15815 ( \16192 , \15954 , \15956 );
xor \U$15816 ( \16193 , \16192 , \15959 );
and \U$15817 ( \16194 , \16190 , \16193 );
and \U$15818 ( \16195 , \16188 , \16193 );
or \U$15819 ( \16196 , \16191 , \16194 , \16195 );
and \U$15820 ( \16197 , \16186 , \16196 );
xor \U$15821 ( \16198 , \15970 , \15972 );
xor \U$15822 ( \16199 , \16198 , \15975 );
and \U$15823 ( \16200 , \16196 , \16199 );
and \U$15824 ( \16201 , \16186 , \16199 );
or \U$15825 ( \16202 , \16197 , \16200 , \16201 );
xor \U$15826 ( \16203 , \15715 , \15733 );
xor \U$15827 ( \16204 , \16203 , \15736 );
and \U$15828 ( \16205 , \16202 , \16204 );
xor \U$15829 ( \16206 , \15968 , \15978 );
xor \U$15830 ( \16207 , \16206 , \15981 );
and \U$15831 ( \16208 , \16204 , \16207 );
and \U$15832 ( \16209 , \16202 , \16207 );
or \U$15833 ( \16210 , \16205 , \16208 , \16209 );
and \U$15834 ( \16211 , \15995 , \16210 );
xor \U$15835 ( \16212 , \15995 , \16210 );
xor \U$15836 ( \16213 , \16202 , \16204 );
xor \U$15837 ( \16214 , \16213 , \16207 );
and \U$15838 ( \16215 , \1562 , \10876 );
and \U$15839 ( \16216 , \1446 , \10873 );
nor \U$15840 ( \16217 , \16215 , \16216 );
xnor \U$15841 ( \16218 , \16217 , \9821 );
and \U$15842 ( \16219 , \1853 , \10063 );
and \U$15843 ( \16220 , \1677 , \10061 );
nor \U$15844 ( \16221 , \16219 , \16220 );
xnor \U$15845 ( \16222 , \16221 , \9824 );
and \U$15846 ( \16223 , \16218 , \16222 );
and \U$15847 ( \16224 , \16222 , \1286 );
and \U$15848 ( \16225 , \16218 , \1286 );
or \U$15849 ( \16226 , \16223 , \16224 , \16225 );
and \U$15850 ( \16227 , \2902 , \7829 );
and \U$15851 ( \16228 , \2728 , \7827 );
nor \U$15852 ( \16229 , \16227 , \16228 );
xnor \U$15853 ( \16230 , \16229 , \7580 );
and \U$15854 ( \16231 , \3207 , \7300 );
and \U$15855 ( \16232 , \3069 , \7298 );
nor \U$15856 ( \16233 , \16231 , \16232 );
xnor \U$15857 ( \16234 , \16233 , \7040 );
and \U$15858 ( \16235 , \16230 , \16234 );
and \U$15859 ( \16236 , \3743 , \6806 );
and \U$15860 ( \16237 , \3326 , \6804 );
nor \U$15861 ( \16238 , \16236 , \16237 );
xnor \U$15862 ( \16239 , \16238 , \6491 );
and \U$15863 ( \16240 , \16234 , \16239 );
and \U$15864 ( \16241 , \16230 , \16239 );
or \U$15865 ( \16242 , \16235 , \16240 , \16241 );
and \U$15866 ( \16243 , \16226 , \16242 );
and \U$15867 ( \16244 , \2104 , \9495 );
and \U$15868 ( \16245 , \1861 , \9493 );
nor \U$15869 ( \16246 , \16244 , \16245 );
xnor \U$15870 ( \16247 , \16246 , \9185 );
and \U$15871 ( \16248 , \2295 , \8958 );
and \U$15872 ( \16249 , \2109 , \8956 );
nor \U$15873 ( \16250 , \16248 , \16249 );
xnor \U$15874 ( \16251 , \16250 , \8587 );
and \U$15875 ( \16252 , \16247 , \16251 );
and \U$15876 ( \16253 , \2703 , \8396 );
and \U$15877 ( \16254 , \2439 , \8394 );
nor \U$15878 ( \16255 , \16253 , \16254 );
xnor \U$15879 ( \16256 , \16255 , \8078 );
and \U$15880 ( \16257 , \16251 , \16256 );
and \U$15881 ( \16258 , \16247 , \16256 );
or \U$15882 ( \16259 , \16252 , \16257 , \16258 );
and \U$15883 ( \16260 , \16242 , \16259 );
and \U$15884 ( \16261 , \16226 , \16259 );
or \U$15885 ( \16262 , \16243 , \16260 , \16261 );
and \U$15886 ( \16263 , \4073 , \6297 );
and \U$15887 ( \16264 , \3951 , \6295 );
nor \U$15888 ( \16265 , \16263 , \16264 );
xnor \U$15889 ( \16266 , \16265 , \5957 );
and \U$15890 ( \16267 , \4334 , \5708 );
and \U$15891 ( \16268 , \4078 , \5706 );
nor \U$15892 ( \16269 , \16267 , \16268 );
xnor \U$15893 ( \16270 , \16269 , \5467 );
and \U$15894 ( \16271 , \16266 , \16270 );
and \U$15895 ( \16272 , \4833 , \5242 );
and \U$15896 ( \16273 , \4531 , \5240 );
nor \U$15897 ( \16274 , \16272 , \16273 );
xnor \U$15898 ( \16275 , \16274 , \5054 );
and \U$15899 ( \16276 , \16270 , \16275 );
and \U$15900 ( \16277 , \16266 , \16275 );
or \U$15901 ( \16278 , \16271 , \16276 , \16277 );
and \U$15902 ( \16279 , \5310 , \4868 );
and \U$15903 ( \16280 , \4841 , \4866 );
nor \U$15904 ( \16281 , \16279 , \16280 );
xnor \U$15905 ( \16282 , \16281 , \4636 );
and \U$15906 ( \16283 , \5579 , \4417 );
and \U$15907 ( \16284 , \5315 , \4415 );
nor \U$15908 ( \16285 , \16283 , \16284 );
xnor \U$15909 ( \16286 , \16285 , \4274 );
and \U$15910 ( \16287 , \16282 , \16286 );
and \U$15911 ( \16288 , \6210 , \4094 );
and \U$15912 ( \16289 , \5838 , \4092 );
nor \U$15913 ( \16290 , \16288 , \16289 );
xnor \U$15914 ( \16291 , \16290 , \3848 );
and \U$15915 ( \16292 , \16286 , \16291 );
and \U$15916 ( \16293 , \16282 , \16291 );
or \U$15917 ( \16294 , \16287 , \16292 , \16293 );
and \U$15918 ( \16295 , \16278 , \16294 );
and \U$15919 ( \16296 , \6562 , \3699 );
and \U$15920 ( \16297 , \6219 , \3697 );
nor \U$15921 ( \16298 , \16296 , \16297 );
xnor \U$15922 ( \16299 , \16298 , \3512 );
and \U$15923 ( \16300 , \7067 , \3386 );
and \U$15924 ( \16301 , \6764 , \3384 );
nor \U$15925 ( \16302 , \16300 , \16301 );
xnor \U$15926 ( \16303 , \16302 , \3181 );
and \U$15927 ( \16304 , \16299 , \16303 );
and \U$15928 ( \16305 , \7765 , \2980 );
and \U$15929 ( \16306 , \7239 , \2978 );
nor \U$15930 ( \16307 , \16305 , \16306 );
xnor \U$15931 ( \16308 , \16307 , \2831 );
and \U$15932 ( \16309 , \16303 , \16308 );
and \U$15933 ( \16310 , \16299 , \16308 );
or \U$15934 ( \16311 , \16304 , \16309 , \16310 );
and \U$15935 ( \16312 , \16294 , \16311 );
and \U$15936 ( \16313 , \16278 , \16311 );
or \U$15937 ( \16314 , \16295 , \16312 , \16313 );
and \U$15938 ( \16315 , \16262 , \16314 );
and \U$15939 ( \16316 , \10223 , \1888 );
and \U$15940 ( \16317 , \9620 , \1886 );
nor \U$15941 ( \16318 , \16316 , \16317 );
xnor \U$15942 ( \16319 , \16318 , \1732 );
and \U$15943 ( \16320 , \10409 , \1616 );
and \U$15944 ( \16321 , \10228 , \1614 );
nor \U$15945 ( \16322 , \16320 , \16321 );
xnor \U$15946 ( \16323 , \16322 , \1503 );
and \U$15947 ( \16324 , \16319 , \16323 );
nand \U$15948 ( \16325 , \11029 , \1420 );
xnor \U$15949 ( \16326 , \16325 , \1286 );
and \U$15950 ( \16327 , \16323 , \16326 );
and \U$15951 ( \16328 , \16319 , \16326 );
or \U$15952 ( \16329 , \16324 , \16327 , \16328 );
and \U$15953 ( \16330 , \8435 , \2658 );
and \U$15954 ( \16331 , \8189 , \2656 );
nor \U$15955 ( \16332 , \16330 , \16331 );
xnor \U$15956 ( \16333 , \16332 , \2516 );
and \U$15957 ( \16334 , \8759 , \2362 );
and \U$15958 ( \16335 , \8440 , \2360 );
nor \U$15959 ( \16336 , \16334 , \16335 );
xnor \U$15960 ( \16337 , \16336 , \2225 );
and \U$15961 ( \16338 , \16333 , \16337 );
and \U$15962 ( \16339 , \9612 , \2156 );
and \U$15963 ( \16340 , \9043 , \2154 );
nor \U$15964 ( \16341 , \16339 , \16340 );
xnor \U$15965 ( \16342 , \16341 , \2004 );
and \U$15966 ( \16343 , \16337 , \16342 );
and \U$15967 ( \16344 , \16333 , \16342 );
or \U$15968 ( \16345 , \16338 , \16343 , \16344 );
and \U$15969 ( \16346 , \16329 , \16345 );
and \U$15970 ( \16347 , \10228 , \1616 );
and \U$15971 ( \16348 , \10223 , \1614 );
nor \U$15972 ( \16349 , \16347 , \16348 );
xnor \U$15973 ( \16350 , \16349 , \1503 );
and \U$15974 ( \16351 , \16345 , \16350 );
and \U$15975 ( \16352 , \16329 , \16350 );
or \U$15976 ( \16353 , \16346 , \16351 , \16352 );
and \U$15977 ( \16354 , \16314 , \16353 );
and \U$15978 ( \16355 , \16262 , \16353 );
or \U$15979 ( \16356 , \16315 , \16354 , \16355 );
and \U$15980 ( \16357 , \11029 , \1422 );
and \U$15981 ( \16358 , \10409 , \1420 );
nor \U$15982 ( \16359 , \16357 , \16358 );
xnor \U$15983 ( \16360 , \16359 , \1286 );
xor \U$15984 ( \16361 , \16032 , \16036 );
xor \U$15985 ( \16362 , \16361 , \16041 );
and \U$15986 ( \16363 , \16360 , \16362 );
xor \U$15987 ( \16364 , \16104 , \16108 );
xor \U$15988 ( \16365 , \16364 , \16113 );
and \U$15989 ( \16366 , \16362 , \16365 );
and \U$15990 ( \16367 , \16360 , \16365 );
or \U$15991 ( \16368 , \16363 , \16366 , \16367 );
xor \U$15992 ( \16369 , \15999 , \16003 );
xor \U$15993 ( \16370 , \16369 , \16008 );
xor \U$15994 ( \16371 , \16015 , \16019 );
xor \U$15995 ( \16372 , \16371 , \16024 );
and \U$15996 ( \16373 , \16370 , \16372 );
xor \U$15997 ( \16374 , \16067 , \16071 );
xor \U$15998 ( \16375 , \16374 , \16076 );
and \U$15999 ( \16376 , \16372 , \16375 );
and \U$16000 ( \16377 , \16370 , \16375 );
or \U$16001 ( \16378 , \16373 , \16376 , \16377 );
and \U$16002 ( \16379 , \16368 , \16378 );
xor \U$16003 ( \16380 , \15842 , \15846 );
xor \U$16004 ( \16381 , \16380 , \1144 );
and \U$16005 ( \16382 , \16378 , \16381 );
and \U$16006 ( \16383 , \16368 , \16381 );
or \U$16007 ( \16384 , \16379 , \16382 , \16383 );
and \U$16008 ( \16385 , \16356 , \16384 );
xor \U$16009 ( \16386 , \16116 , \16118 );
xor \U$16010 ( \16387 , \16386 , \16121 );
xor \U$16011 ( \16388 , \16129 , \16131 );
xor \U$16012 ( \16389 , \16388 , \16134 );
and \U$16013 ( \16390 , \16387 , \16389 );
xor \U$16014 ( \16391 , \16139 , \16141 );
xor \U$16015 ( \16392 , \16391 , \16144 );
and \U$16016 ( \16393 , \16389 , \16392 );
and \U$16017 ( \16394 , \16387 , \16392 );
or \U$16018 ( \16395 , \16390 , \16393 , \16394 );
and \U$16019 ( \16396 , \16384 , \16395 );
and \U$16020 ( \16397 , \16356 , \16395 );
or \U$16021 ( \16398 , \16385 , \16396 , \16397 );
xor \U$16022 ( \16399 , \15786 , \15802 );
xor \U$16023 ( \16400 , \16399 , \15819 );
xor \U$16024 ( \16401 , \15838 , \15850 );
xor \U$16025 ( \16402 , \16401 , \15867 );
and \U$16026 ( \16403 , \16400 , \16402 );
xor \U$16027 ( \16404 , \16156 , \16158 );
xor \U$16028 ( \16405 , \16404 , \16161 );
and \U$16029 ( \16406 , \16402 , \16405 );
and \U$16030 ( \16407 , \16400 , \16405 );
or \U$16031 ( \16408 , \16403 , \16406 , \16407 );
and \U$16032 ( \16409 , \16398 , \16408 );
xor \U$16033 ( \16410 , \16047 , \16099 );
xor \U$16034 ( \16411 , \16410 , \16124 );
xor \U$16035 ( \16412 , \16137 , \16147 );
xor \U$16036 ( \16413 , \16412 , \16150 );
and \U$16037 ( \16414 , \16411 , \16413 );
and \U$16038 ( \16415 , \16408 , \16414 );
and \U$16039 ( \16416 , \16398 , \16414 );
or \U$16040 ( \16417 , \16409 , \16415 , \16416 );
xor \U$16041 ( \16418 , \16127 , \16153 );
xor \U$16042 ( \16419 , \16418 , \16164 );
xor \U$16043 ( \16420 , \16169 , \16171 );
xor \U$16044 ( \16421 , \16420 , \16174 );
and \U$16045 ( \16422 , \16419 , \16421 );
xor \U$16046 ( \16423 , \16180 , \16182 );
and \U$16047 ( \16424 , \16421 , \16423 );
and \U$16048 ( \16425 , \16419 , \16423 );
or \U$16049 ( \16426 , \16422 , \16424 , \16425 );
and \U$16050 ( \16427 , \16417 , \16426 );
xor \U$16051 ( \16428 , \16188 , \16190 );
xor \U$16052 ( \16429 , \16428 , \16193 );
and \U$16053 ( \16430 , \16426 , \16429 );
and \U$16054 ( \16431 , \16417 , \16429 );
or \U$16055 ( \16432 , \16427 , \16430 , \16431 );
xor \U$16056 ( \16433 , \15952 , \15962 );
xor \U$16057 ( \16434 , \16433 , \15965 );
and \U$16058 ( \16435 , \16432 , \16434 );
xor \U$16059 ( \16436 , \16186 , \16196 );
xor \U$16060 ( \16437 , \16436 , \16199 );
and \U$16061 ( \16438 , \16434 , \16437 );
and \U$16062 ( \16439 , \16432 , \16437 );
or \U$16063 ( \16440 , \16435 , \16438 , \16439 );
and \U$16064 ( \16441 , \16214 , \16440 );
xor \U$16065 ( \16442 , \16214 , \16440 );
xor \U$16066 ( \16443 , \16432 , \16434 );
xor \U$16067 ( \16444 , \16443 , \16437 );
and \U$16068 ( \16445 , \1677 , \10876 );
and \U$16069 ( \16446 , \1562 , \10873 );
nor \U$16070 ( \16447 , \16445 , \16446 );
xnor \U$16071 ( \16448 , \16447 , \9821 );
and \U$16072 ( \16449 , \1861 , \10063 );
and \U$16073 ( \16450 , \1853 , \10061 );
nor \U$16074 ( \16451 , \16449 , \16450 );
xnor \U$16075 ( \16452 , \16451 , \9824 );
and \U$16076 ( \16453 , \16448 , \16452 );
and \U$16077 ( \16454 , \2109 , \9495 );
and \U$16078 ( \16455 , \2104 , \9493 );
nor \U$16079 ( \16456 , \16454 , \16455 );
xnor \U$16080 ( \16457 , \16456 , \9185 );
and \U$16081 ( \16458 , \16452 , \16457 );
and \U$16082 ( \16459 , \16448 , \16457 );
or \U$16083 ( \16460 , \16453 , \16458 , \16459 );
and \U$16084 ( \16461 , \2439 , \8958 );
and \U$16085 ( \16462 , \2295 , \8956 );
nor \U$16086 ( \16463 , \16461 , \16462 );
xnor \U$16087 ( \16464 , \16463 , \8587 );
and \U$16088 ( \16465 , \2728 , \8396 );
and \U$16089 ( \16466 , \2703 , \8394 );
nor \U$16090 ( \16467 , \16465 , \16466 );
xnor \U$16091 ( \16468 , \16467 , \8078 );
and \U$16092 ( \16469 , \16464 , \16468 );
and \U$16093 ( \16470 , \3069 , \7829 );
and \U$16094 ( \16471 , \2902 , \7827 );
nor \U$16095 ( \16472 , \16470 , \16471 );
xnor \U$16096 ( \16473 , \16472 , \7580 );
and \U$16097 ( \16474 , \16468 , \16473 );
and \U$16098 ( \16475 , \16464 , \16473 );
or \U$16099 ( \16476 , \16469 , \16474 , \16475 );
and \U$16100 ( \16477 , \16460 , \16476 );
and \U$16101 ( \16478 , \3326 , \7300 );
and \U$16102 ( \16479 , \3207 , \7298 );
nor \U$16103 ( \16480 , \16478 , \16479 );
xnor \U$16104 ( \16481 , \16480 , \7040 );
and \U$16105 ( \16482 , \3951 , \6806 );
and \U$16106 ( \16483 , \3743 , \6804 );
nor \U$16107 ( \16484 , \16482 , \16483 );
xnor \U$16108 ( \16485 , \16484 , \6491 );
and \U$16109 ( \16486 , \16481 , \16485 );
and \U$16110 ( \16487 , \4078 , \6297 );
and \U$16111 ( \16488 , \4073 , \6295 );
nor \U$16112 ( \16489 , \16487 , \16488 );
xnor \U$16113 ( \16490 , \16489 , \5957 );
and \U$16114 ( \16491 , \16485 , \16490 );
and \U$16115 ( \16492 , \16481 , \16490 );
or \U$16116 ( \16493 , \16486 , \16491 , \16492 );
and \U$16117 ( \16494 , \16476 , \16493 );
and \U$16118 ( \16495 , \16460 , \16493 );
or \U$16119 ( \16496 , \16477 , \16494 , \16495 );
and \U$16120 ( \16497 , \5838 , \4417 );
and \U$16121 ( \16498 , \5579 , \4415 );
nor \U$16122 ( \16499 , \16497 , \16498 );
xnor \U$16123 ( \16500 , \16499 , \4274 );
and \U$16124 ( \16501 , \6219 , \4094 );
and \U$16125 ( \16502 , \6210 , \4092 );
nor \U$16126 ( \16503 , \16501 , \16502 );
xnor \U$16127 ( \16504 , \16503 , \3848 );
and \U$16128 ( \16505 , \16500 , \16504 );
and \U$16129 ( \16506 , \6764 , \3699 );
and \U$16130 ( \16507 , \6562 , \3697 );
nor \U$16131 ( \16508 , \16506 , \16507 );
xnor \U$16132 ( \16509 , \16508 , \3512 );
and \U$16133 ( \16510 , \16504 , \16509 );
and \U$16134 ( \16511 , \16500 , \16509 );
or \U$16135 ( \16512 , \16505 , \16510 , \16511 );
and \U$16136 ( \16513 , \7239 , \3386 );
and \U$16137 ( \16514 , \7067 , \3384 );
nor \U$16138 ( \16515 , \16513 , \16514 );
xnor \U$16139 ( \16516 , \16515 , \3181 );
and \U$16140 ( \16517 , \8189 , \2980 );
and \U$16141 ( \16518 , \7765 , \2978 );
nor \U$16142 ( \16519 , \16517 , \16518 );
xnor \U$16143 ( \16520 , \16519 , \2831 );
and \U$16144 ( \16521 , \16516 , \16520 );
and \U$16145 ( \16522 , \8440 , \2658 );
and \U$16146 ( \16523 , \8435 , \2656 );
nor \U$16147 ( \16524 , \16522 , \16523 );
xnor \U$16148 ( \16525 , \16524 , \2516 );
and \U$16149 ( \16526 , \16520 , \16525 );
and \U$16150 ( \16527 , \16516 , \16525 );
or \U$16151 ( \16528 , \16521 , \16526 , \16527 );
and \U$16152 ( \16529 , \16512 , \16528 );
and \U$16153 ( \16530 , \4531 , \5708 );
and \U$16154 ( \16531 , \4334 , \5706 );
nor \U$16155 ( \16532 , \16530 , \16531 );
xnor \U$16156 ( \16533 , \16532 , \5467 );
and \U$16157 ( \16534 , \4841 , \5242 );
and \U$16158 ( \16535 , \4833 , \5240 );
nor \U$16159 ( \16536 , \16534 , \16535 );
xnor \U$16160 ( \16537 , \16536 , \5054 );
and \U$16161 ( \16538 , \16533 , \16537 );
and \U$16162 ( \16539 , \5315 , \4868 );
and \U$16163 ( \16540 , \5310 , \4866 );
nor \U$16164 ( \16541 , \16539 , \16540 );
xnor \U$16165 ( \16542 , \16541 , \4636 );
and \U$16166 ( \16543 , \16537 , \16542 );
and \U$16167 ( \16544 , \16533 , \16542 );
or \U$16168 ( \16545 , \16538 , \16543 , \16544 );
and \U$16169 ( \16546 , \16528 , \16545 );
and \U$16170 ( \16547 , \16512 , \16545 );
or \U$16171 ( \16548 , \16529 , \16546 , \16547 );
and \U$16172 ( \16549 , \16496 , \16548 );
and \U$16173 ( \16550 , \9043 , \2362 );
and \U$16174 ( \16551 , \8759 , \2360 );
nor \U$16175 ( \16552 , \16550 , \16551 );
xnor \U$16176 ( \16553 , \16552 , \2225 );
and \U$16177 ( \16554 , \9620 , \2156 );
and \U$16178 ( \16555 , \9612 , \2154 );
nor \U$16179 ( \16556 , \16554 , \16555 );
xnor \U$16180 ( \16557 , \16556 , \2004 );
and \U$16181 ( \16558 , \16553 , \16557 );
and \U$16182 ( \16559 , \10228 , \1888 );
and \U$16183 ( \16560 , \10223 , \1886 );
nor \U$16184 ( \16561 , \16559 , \16560 );
xnor \U$16185 ( \16562 , \16561 , \1732 );
and \U$16186 ( \16563 , \16557 , \16562 );
and \U$16187 ( \16564 , \16553 , \16562 );
or \U$16188 ( \16565 , \16558 , \16563 , \16564 );
xor \U$16189 ( \16566 , \16319 , \16323 );
xor \U$16190 ( \16567 , \16566 , \16326 );
and \U$16191 ( \16568 , \16565 , \16567 );
xor \U$16192 ( \16569 , \16333 , \16337 );
xor \U$16193 ( \16570 , \16569 , \16342 );
and \U$16194 ( \16571 , \16567 , \16570 );
and \U$16195 ( \16572 , \16565 , \16570 );
or \U$16196 ( \16573 , \16568 , \16571 , \16572 );
and \U$16197 ( \16574 , \16548 , \16573 );
and \U$16198 ( \16575 , \16496 , \16573 );
or \U$16199 ( \16576 , \16549 , \16574 , \16575 );
xor \U$16200 ( \16577 , \16266 , \16270 );
xor \U$16201 ( \16578 , \16577 , \16275 );
xor \U$16202 ( \16579 , \16282 , \16286 );
xor \U$16203 ( \16580 , \16579 , \16291 );
and \U$16204 ( \16581 , \16578 , \16580 );
xor \U$16205 ( \16582 , \16299 , \16303 );
xor \U$16206 ( \16583 , \16582 , \16308 );
and \U$16207 ( \16584 , \16580 , \16583 );
and \U$16208 ( \16585 , \16578 , \16583 );
or \U$16209 ( \16586 , \16581 , \16584 , \16585 );
xor \U$16210 ( \16587 , \16218 , \16222 );
xor \U$16211 ( \16588 , \16587 , \1286 );
xor \U$16212 ( \16589 , \16230 , \16234 );
xor \U$16213 ( \16590 , \16589 , \16239 );
and \U$16214 ( \16591 , \16588 , \16590 );
xor \U$16215 ( \16592 , \16247 , \16251 );
xor \U$16216 ( \16593 , \16592 , \16256 );
and \U$16217 ( \16594 , \16590 , \16593 );
and \U$16218 ( \16595 , \16588 , \16593 );
or \U$16219 ( \16596 , \16591 , \16594 , \16595 );
and \U$16220 ( \16597 , \16586 , \16596 );
xor \U$16221 ( \16598 , \16051 , \16055 );
xor \U$16222 ( \16599 , \16598 , \16060 );
and \U$16223 ( \16600 , \16596 , \16599 );
and \U$16224 ( \16601 , \16586 , \16599 );
or \U$16225 ( \16602 , \16597 , \16600 , \16601 );
and \U$16226 ( \16603 , \16576 , \16602 );
xor \U$16227 ( \16604 , \16084 , \16088 );
xor \U$16228 ( \16605 , \16604 , \16093 );
xor \U$16229 ( \16606 , \16360 , \16362 );
xor \U$16230 ( \16607 , \16606 , \16365 );
and \U$16231 ( \16608 , \16605 , \16607 );
xor \U$16232 ( \16609 , \16370 , \16372 );
xor \U$16233 ( \16610 , \16609 , \16375 );
and \U$16234 ( \16611 , \16607 , \16610 );
and \U$16235 ( \16612 , \16605 , \16610 );
or \U$16236 ( \16613 , \16608 , \16611 , \16612 );
and \U$16237 ( \16614 , \16602 , \16613 );
and \U$16238 ( \16615 , \16576 , \16613 );
or \U$16239 ( \16616 , \16603 , \16614 , \16615 );
xor \U$16240 ( \16617 , \16226 , \16242 );
xor \U$16241 ( \16618 , \16617 , \16259 );
xor \U$16242 ( \16619 , \16278 , \16294 );
xor \U$16243 ( \16620 , \16619 , \16311 );
and \U$16244 ( \16621 , \16618 , \16620 );
xor \U$16245 ( \16622 , \16329 , \16345 );
xor \U$16246 ( \16623 , \16622 , \16350 );
and \U$16247 ( \16624 , \16620 , \16623 );
and \U$16248 ( \16625 , \16618 , \16623 );
or \U$16249 ( \16626 , \16621 , \16624 , \16625 );
xor \U$16250 ( \16627 , \16011 , \16027 );
xor \U$16251 ( \16628 , \16627 , \16044 );
and \U$16252 ( \16629 , \16626 , \16628 );
xor \U$16253 ( \16630 , \16063 , \16079 );
xor \U$16254 ( \16631 , \16630 , \16096 );
and \U$16255 ( \16632 , \16628 , \16631 );
and \U$16256 ( \16633 , \16626 , \16631 );
or \U$16257 ( \16634 , \16629 , \16632 , \16633 );
and \U$16258 ( \16635 , \16616 , \16634 );
xor \U$16259 ( \16636 , \16262 , \16314 );
xor \U$16260 ( \16637 , \16636 , \16353 );
xor \U$16261 ( \16638 , \16368 , \16378 );
xor \U$16262 ( \16639 , \16638 , \16381 );
and \U$16263 ( \16640 , \16637 , \16639 );
xor \U$16264 ( \16641 , \16387 , \16389 );
xor \U$16265 ( \16642 , \16641 , \16392 );
and \U$16266 ( \16643 , \16639 , \16642 );
and \U$16267 ( \16644 , \16637 , \16642 );
or \U$16268 ( \16645 , \16640 , \16643 , \16644 );
and \U$16269 ( \16646 , \16634 , \16645 );
and \U$16270 ( \16647 , \16616 , \16645 );
or \U$16271 ( \16648 , \16635 , \16646 , \16647 );
xor \U$16272 ( \16649 , \16356 , \16384 );
xor \U$16273 ( \16650 , \16649 , \16395 );
xor \U$16274 ( \16651 , \16400 , \16402 );
xor \U$16275 ( \16652 , \16651 , \16405 );
and \U$16276 ( \16653 , \16650 , \16652 );
xor \U$16277 ( \16654 , \16411 , \16413 );
and \U$16278 ( \16655 , \16652 , \16654 );
and \U$16279 ( \16656 , \16650 , \16654 );
or \U$16280 ( \16657 , \16653 , \16655 , \16656 );
and \U$16281 ( \16658 , \16648 , \16657 );
xor \U$16282 ( \16659 , \16419 , \16421 );
xor \U$16283 ( \16660 , \16659 , \16423 );
and \U$16284 ( \16661 , \16657 , \16660 );
and \U$16285 ( \16662 , \16648 , \16660 );
or \U$16286 ( \16663 , \16658 , \16661 , \16662 );
xor \U$16287 ( \16664 , \16167 , \16177 );
xor \U$16288 ( \16665 , \16664 , \16183 );
and \U$16289 ( \16666 , \16663 , \16665 );
xor \U$16290 ( \16667 , \16417 , \16426 );
xor \U$16291 ( \16668 , \16667 , \16429 );
and \U$16292 ( \16669 , \16665 , \16668 );
and \U$16293 ( \16670 , \16663 , \16668 );
or \U$16294 ( \16671 , \16666 , \16669 , \16670 );
and \U$16295 ( \16672 , \16444 , \16671 );
xor \U$16296 ( \16673 , \16444 , \16671 );
xor \U$16297 ( \16674 , \16663 , \16665 );
xor \U$16298 ( \16675 , \16674 , \16668 );
and \U$16299 ( \16676 , \7067 , \3699 );
and \U$16300 ( \16677 , \6764 , \3697 );
nor \U$16301 ( \16678 , \16676 , \16677 );
xnor \U$16302 ( \16679 , \16678 , \3512 );
and \U$16303 ( \16680 , \7765 , \3386 );
and \U$16304 ( \16681 , \7239 , \3384 );
nor \U$16305 ( \16682 , \16680 , \16681 );
xnor \U$16306 ( \16683 , \16682 , \3181 );
and \U$16307 ( \16684 , \16679 , \16683 );
and \U$16308 ( \16685 , \8435 , \2980 );
and \U$16309 ( \16686 , \8189 , \2978 );
nor \U$16310 ( \16687 , \16685 , \16686 );
xnor \U$16311 ( \16688 , \16687 , \2831 );
and \U$16312 ( \16689 , \16683 , \16688 );
and \U$16313 ( \16690 , \16679 , \16688 );
or \U$16314 ( \16691 , \16684 , \16689 , \16690 );
and \U$16315 ( \16692 , \4334 , \6297 );
and \U$16316 ( \16693 , \4078 , \6295 );
nor \U$16317 ( \16694 , \16692 , \16693 );
xnor \U$16318 ( \16695 , \16694 , \5957 );
and \U$16319 ( \16696 , \4833 , \5708 );
and \U$16320 ( \16697 , \4531 , \5706 );
nor \U$16321 ( \16698 , \16696 , \16697 );
xnor \U$16322 ( \16699 , \16698 , \5467 );
and \U$16323 ( \16700 , \16695 , \16699 );
and \U$16324 ( \16701 , \5310 , \5242 );
and \U$16325 ( \16702 , \4841 , \5240 );
nor \U$16326 ( \16703 , \16701 , \16702 );
xnor \U$16327 ( \16704 , \16703 , \5054 );
and \U$16328 ( \16705 , \16699 , \16704 );
and \U$16329 ( \16706 , \16695 , \16704 );
or \U$16330 ( \16707 , \16700 , \16705 , \16706 );
and \U$16331 ( \16708 , \16691 , \16707 );
and \U$16332 ( \16709 , \5579 , \4868 );
and \U$16333 ( \16710 , \5315 , \4866 );
nor \U$16334 ( \16711 , \16709 , \16710 );
xnor \U$16335 ( \16712 , \16711 , \4636 );
and \U$16336 ( \16713 , \6210 , \4417 );
and \U$16337 ( \16714 , \5838 , \4415 );
nor \U$16338 ( \16715 , \16713 , \16714 );
xnor \U$16339 ( \16716 , \16715 , \4274 );
and \U$16340 ( \16717 , \16712 , \16716 );
and \U$16341 ( \16718 , \6562 , \4094 );
and \U$16342 ( \16719 , \6219 , \4092 );
nor \U$16343 ( \16720 , \16718 , \16719 );
xnor \U$16344 ( \16721 , \16720 , \3848 );
and \U$16345 ( \16722 , \16716 , \16721 );
and \U$16346 ( \16723 , \16712 , \16721 );
or \U$16347 ( \16724 , \16717 , \16722 , \16723 );
and \U$16348 ( \16725 , \16707 , \16724 );
and \U$16349 ( \16726 , \16691 , \16724 );
or \U$16350 ( \16727 , \16708 , \16725 , \16726 );
and \U$16351 ( \16728 , \1853 , \10876 );
and \U$16352 ( \16729 , \1677 , \10873 );
nor \U$16353 ( \16730 , \16728 , \16729 );
xnor \U$16354 ( \16731 , \16730 , \9821 );
and \U$16355 ( \16732 , \2104 , \10063 );
and \U$16356 ( \16733 , \1861 , \10061 );
nor \U$16357 ( \16734 , \16732 , \16733 );
xnor \U$16358 ( \16735 , \16734 , \9824 );
and \U$16359 ( \16736 , \16731 , \16735 );
and \U$16360 ( \16737 , \16735 , \1503 );
and \U$16361 ( \16738 , \16731 , \1503 );
or \U$16362 ( \16739 , \16736 , \16737 , \16738 );
and \U$16363 ( \16740 , \3207 , \7829 );
and \U$16364 ( \16741 , \3069 , \7827 );
nor \U$16365 ( \16742 , \16740 , \16741 );
xnor \U$16366 ( \16743 , \16742 , \7580 );
and \U$16367 ( \16744 , \3743 , \7300 );
and \U$16368 ( \16745 , \3326 , \7298 );
nor \U$16369 ( \16746 , \16744 , \16745 );
xnor \U$16370 ( \16747 , \16746 , \7040 );
and \U$16371 ( \16748 , \16743 , \16747 );
and \U$16372 ( \16749 , \4073 , \6806 );
and \U$16373 ( \16750 , \3951 , \6804 );
nor \U$16374 ( \16751 , \16749 , \16750 );
xnor \U$16375 ( \16752 , \16751 , \6491 );
and \U$16376 ( \16753 , \16747 , \16752 );
and \U$16377 ( \16754 , \16743 , \16752 );
or \U$16378 ( \16755 , \16748 , \16753 , \16754 );
and \U$16379 ( \16756 , \16739 , \16755 );
and \U$16380 ( \16757 , \2295 , \9495 );
and \U$16381 ( \16758 , \2109 , \9493 );
nor \U$16382 ( \16759 , \16757 , \16758 );
xnor \U$16383 ( \16760 , \16759 , \9185 );
and \U$16384 ( \16761 , \2703 , \8958 );
and \U$16385 ( \16762 , \2439 , \8956 );
nor \U$16386 ( \16763 , \16761 , \16762 );
xnor \U$16387 ( \16764 , \16763 , \8587 );
and \U$16388 ( \16765 , \16760 , \16764 );
and \U$16389 ( \16766 , \2902 , \8396 );
and \U$16390 ( \16767 , \2728 , \8394 );
nor \U$16391 ( \16768 , \16766 , \16767 );
xnor \U$16392 ( \16769 , \16768 , \8078 );
and \U$16393 ( \16770 , \16764 , \16769 );
and \U$16394 ( \16771 , \16760 , \16769 );
or \U$16395 ( \16772 , \16765 , \16770 , \16771 );
and \U$16396 ( \16773 , \16755 , \16772 );
and \U$16397 ( \16774 , \16739 , \16772 );
or \U$16398 ( \16775 , \16756 , \16773 , \16774 );
and \U$16399 ( \16776 , \16727 , \16775 );
and \U$16400 ( \16777 , \8759 , \2658 );
and \U$16401 ( \16778 , \8440 , \2656 );
nor \U$16402 ( \16779 , \16777 , \16778 );
xnor \U$16403 ( \16780 , \16779 , \2516 );
and \U$16404 ( \16781 , \9612 , \2362 );
and \U$16405 ( \16782 , \9043 , \2360 );
nor \U$16406 ( \16783 , \16781 , \16782 );
xnor \U$16407 ( \16784 , \16783 , \2225 );
and \U$16408 ( \16785 , \16780 , \16784 );
and \U$16409 ( \16786 , \10223 , \2156 );
and \U$16410 ( \16787 , \9620 , \2154 );
nor \U$16411 ( \16788 , \16786 , \16787 );
xnor \U$16412 ( \16789 , \16788 , \2004 );
and \U$16413 ( \16790 , \16784 , \16789 );
and \U$16414 ( \16791 , \16780 , \16789 );
or \U$16415 ( \16792 , \16785 , \16790 , \16791 );
and \U$16416 ( \16793 , \10409 , \1888 );
and \U$16417 ( \16794 , \10228 , \1886 );
nor \U$16418 ( \16795 , \16793 , \16794 );
xnor \U$16419 ( \16796 , \16795 , \1732 );
nand \U$16420 ( \16797 , \11029 , \1614 );
xnor \U$16421 ( \16798 , \16797 , \1503 );
and \U$16422 ( \16799 , \16796 , \16798 );
and \U$16423 ( \16800 , \16792 , \16799 );
and \U$16424 ( \16801 , \11029 , \1616 );
and \U$16425 ( \16802 , \10409 , \1614 );
nor \U$16426 ( \16803 , \16801 , \16802 );
xnor \U$16427 ( \16804 , \16803 , \1503 );
and \U$16428 ( \16805 , \16799 , \16804 );
and \U$16429 ( \16806 , \16792 , \16804 );
or \U$16430 ( \16807 , \16800 , \16805 , \16806 );
and \U$16431 ( \16808 , \16775 , \16807 );
and \U$16432 ( \16809 , \16727 , \16807 );
or \U$16433 ( \16810 , \16776 , \16808 , \16809 );
xor \U$16434 ( \16811 , \16464 , \16468 );
xor \U$16435 ( \16812 , \16811 , \16473 );
xor \U$16436 ( \16813 , \16533 , \16537 );
xor \U$16437 ( \16814 , \16813 , \16542 );
and \U$16438 ( \16815 , \16812 , \16814 );
xor \U$16439 ( \16816 , \16481 , \16485 );
xor \U$16440 ( \16817 , \16816 , \16490 );
and \U$16441 ( \16818 , \16814 , \16817 );
and \U$16442 ( \16819 , \16812 , \16817 );
or \U$16443 ( \16820 , \16815 , \16818 , \16819 );
xor \U$16444 ( \16821 , \16500 , \16504 );
xor \U$16445 ( \16822 , \16821 , \16509 );
xor \U$16446 ( \16823 , \16553 , \16557 );
xor \U$16447 ( \16824 , \16823 , \16562 );
and \U$16448 ( \16825 , \16822 , \16824 );
xor \U$16449 ( \16826 , \16516 , \16520 );
xor \U$16450 ( \16827 , \16826 , \16525 );
and \U$16451 ( \16828 , \16824 , \16827 );
and \U$16452 ( \16829 , \16822 , \16827 );
or \U$16453 ( \16830 , \16825 , \16828 , \16829 );
and \U$16454 ( \16831 , \16820 , \16830 );
xor \U$16455 ( \16832 , \16588 , \16590 );
xor \U$16456 ( \16833 , \16832 , \16593 );
and \U$16457 ( \16834 , \16830 , \16833 );
and \U$16458 ( \16835 , \16820 , \16833 );
or \U$16459 ( \16836 , \16831 , \16834 , \16835 );
and \U$16460 ( \16837 , \16810 , \16836 );
xor \U$16461 ( \16838 , \16512 , \16528 );
xor \U$16462 ( \16839 , \16838 , \16545 );
xor \U$16463 ( \16840 , \16578 , \16580 );
xor \U$16464 ( \16841 , \16840 , \16583 );
and \U$16465 ( \16842 , \16839 , \16841 );
xor \U$16466 ( \16843 , \16565 , \16567 );
xor \U$16467 ( \16844 , \16843 , \16570 );
and \U$16468 ( \16845 , \16841 , \16844 );
and \U$16469 ( \16846 , \16839 , \16844 );
or \U$16470 ( \16847 , \16842 , \16845 , \16846 );
and \U$16471 ( \16848 , \16836 , \16847 );
and \U$16472 ( \16849 , \16810 , \16847 );
or \U$16473 ( \16850 , \16837 , \16848 , \16849 );
xor \U$16474 ( \16851 , \16618 , \16620 );
xor \U$16475 ( \16852 , \16851 , \16623 );
xor \U$16476 ( \16853 , \16586 , \16596 );
xor \U$16477 ( \16854 , \16853 , \16599 );
and \U$16478 ( \16855 , \16852 , \16854 );
xor \U$16479 ( \16856 , \16605 , \16607 );
xor \U$16480 ( \16857 , \16856 , \16610 );
and \U$16481 ( \16858 , \16854 , \16857 );
and \U$16482 ( \16859 , \16852 , \16857 );
or \U$16483 ( \16860 , \16855 , \16858 , \16859 );
and \U$16484 ( \16861 , \16850 , \16860 );
xor \U$16485 ( \16862 , \16637 , \16639 );
xor \U$16486 ( \16863 , \16862 , \16642 );
and \U$16487 ( \16864 , \16860 , \16863 );
and \U$16488 ( \16865 , \16850 , \16863 );
or \U$16489 ( \16866 , \16861 , \16864 , \16865 );
xor \U$16490 ( \16867 , \16616 , \16634 );
xor \U$16491 ( \16868 , \16867 , \16645 );
and \U$16492 ( \16869 , \16866 , \16868 );
xor \U$16493 ( \16870 , \16650 , \16652 );
xor \U$16494 ( \16871 , \16870 , \16654 );
and \U$16495 ( \16872 , \16868 , \16871 );
and \U$16496 ( \16873 , \16866 , \16871 );
or \U$16497 ( \16874 , \16869 , \16872 , \16873 );
xor \U$16498 ( \16875 , \16398 , \16408 );
xor \U$16499 ( \16876 , \16875 , \16414 );
and \U$16500 ( \16877 , \16874 , \16876 );
xor \U$16501 ( \16878 , \16648 , \16657 );
xor \U$16502 ( \16879 , \16878 , \16660 );
and \U$16503 ( \16880 , \16876 , \16879 );
and \U$16504 ( \16881 , \16874 , \16879 );
or \U$16505 ( \16882 , \16877 , \16880 , \16881 );
and \U$16506 ( \16883 , \16675 , \16882 );
xor \U$16507 ( \16884 , \16675 , \16882 );
xor \U$16508 ( \16885 , \16874 , \16876 );
xor \U$16509 ( \16886 , \16885 , \16879 );
and \U$16510 ( \16887 , \6219 , \4417 );
and \U$16511 ( \16888 , \6210 , \4415 );
nor \U$16512 ( \16889 , \16887 , \16888 );
xnor \U$16513 ( \16890 , \16889 , \4274 );
and \U$16514 ( \16891 , \6764 , \4094 );
and \U$16515 ( \16892 , \6562 , \4092 );
nor \U$16516 ( \16893 , \16891 , \16892 );
xnor \U$16517 ( \16894 , \16893 , \3848 );
and \U$16518 ( \16895 , \16890 , \16894 );
and \U$16519 ( \16896 , \7239 , \3699 );
and \U$16520 ( \16897 , \7067 , \3697 );
nor \U$16521 ( \16898 , \16896 , \16897 );
xnor \U$16522 ( \16899 , \16898 , \3512 );
and \U$16523 ( \16900 , \16894 , \16899 );
and \U$16524 ( \16901 , \16890 , \16899 );
or \U$16525 ( \16902 , \16895 , \16900 , \16901 );
and \U$16526 ( \16903 , \8189 , \3386 );
and \U$16527 ( \16904 , \7765 , \3384 );
nor \U$16528 ( \16905 , \16903 , \16904 );
xnor \U$16529 ( \16906 , \16905 , \3181 );
and \U$16530 ( \16907 , \8440 , \2980 );
and \U$16531 ( \16908 , \8435 , \2978 );
nor \U$16532 ( \16909 , \16907 , \16908 );
xnor \U$16533 ( \16910 , \16909 , \2831 );
and \U$16534 ( \16911 , \16906 , \16910 );
and \U$16535 ( \16912 , \9043 , \2658 );
and \U$16536 ( \16913 , \8759 , \2656 );
nor \U$16537 ( \16914 , \16912 , \16913 );
xnor \U$16538 ( \16915 , \16914 , \2516 );
and \U$16539 ( \16916 , \16910 , \16915 );
and \U$16540 ( \16917 , \16906 , \16915 );
or \U$16541 ( \16918 , \16911 , \16916 , \16917 );
and \U$16542 ( \16919 , \16902 , \16918 );
and \U$16543 ( \16920 , \4841 , \5708 );
and \U$16544 ( \16921 , \4833 , \5706 );
nor \U$16545 ( \16922 , \16920 , \16921 );
xnor \U$16546 ( \16923 , \16922 , \5467 );
and \U$16547 ( \16924 , \5315 , \5242 );
and \U$16548 ( \16925 , \5310 , \5240 );
nor \U$16549 ( \16926 , \16924 , \16925 );
xnor \U$16550 ( \16927 , \16926 , \5054 );
and \U$16551 ( \16928 , \16923 , \16927 );
and \U$16552 ( \16929 , \5838 , \4868 );
and \U$16553 ( \16930 , \5579 , \4866 );
nor \U$16554 ( \16931 , \16929 , \16930 );
xnor \U$16555 ( \16932 , \16931 , \4636 );
and \U$16556 ( \16933 , \16927 , \16932 );
and \U$16557 ( \16934 , \16923 , \16932 );
or \U$16558 ( \16935 , \16928 , \16933 , \16934 );
and \U$16559 ( \16936 , \16918 , \16935 );
and \U$16560 ( \16937 , \16902 , \16935 );
or \U$16561 ( \16938 , \16919 , \16936 , \16937 );
and \U$16562 ( \16939 , \3951 , \7300 );
and \U$16563 ( \16940 , \3743 , \7298 );
nor \U$16564 ( \16941 , \16939 , \16940 );
xnor \U$16565 ( \16942 , \16941 , \7040 );
and \U$16566 ( \16943 , \4078 , \6806 );
and \U$16567 ( \16944 , \4073 , \6804 );
nor \U$16568 ( \16945 , \16943 , \16944 );
xnor \U$16569 ( \16946 , \16945 , \6491 );
and \U$16570 ( \16947 , \16942 , \16946 );
and \U$16571 ( \16948 , \4531 , \6297 );
and \U$16572 ( \16949 , \4334 , \6295 );
nor \U$16573 ( \16950 , \16948 , \16949 );
xnor \U$16574 ( \16951 , \16950 , \5957 );
and \U$16575 ( \16952 , \16946 , \16951 );
and \U$16576 ( \16953 , \16942 , \16951 );
or \U$16577 ( \16954 , \16947 , \16952 , \16953 );
and \U$16578 ( \16955 , \2728 , \8958 );
and \U$16579 ( \16956 , \2703 , \8956 );
nor \U$16580 ( \16957 , \16955 , \16956 );
xnor \U$16581 ( \16958 , \16957 , \8587 );
and \U$16582 ( \16959 , \3069 , \8396 );
and \U$16583 ( \16960 , \2902 , \8394 );
nor \U$16584 ( \16961 , \16959 , \16960 );
xnor \U$16585 ( \16962 , \16961 , \8078 );
and \U$16586 ( \16963 , \16958 , \16962 );
and \U$16587 ( \16964 , \3326 , \7829 );
and \U$16588 ( \16965 , \3207 , \7827 );
nor \U$16589 ( \16966 , \16964 , \16965 );
xnor \U$16590 ( \16967 , \16966 , \7580 );
and \U$16591 ( \16968 , \16962 , \16967 );
and \U$16592 ( \16969 , \16958 , \16967 );
or \U$16593 ( \16970 , \16963 , \16968 , \16969 );
and \U$16594 ( \16971 , \16954 , \16970 );
and \U$16595 ( \16972 , \1861 , \10876 );
and \U$16596 ( \16973 , \1853 , \10873 );
nor \U$16597 ( \16974 , \16972 , \16973 );
xnor \U$16598 ( \16975 , \16974 , \9821 );
and \U$16599 ( \16976 , \2109 , \10063 );
and \U$16600 ( \16977 , \2104 , \10061 );
nor \U$16601 ( \16978 , \16976 , \16977 );
xnor \U$16602 ( \16979 , \16978 , \9824 );
and \U$16603 ( \16980 , \16975 , \16979 );
and \U$16604 ( \16981 , \2439 , \9495 );
and \U$16605 ( \16982 , \2295 , \9493 );
nor \U$16606 ( \16983 , \16981 , \16982 );
xnor \U$16607 ( \16984 , \16983 , \9185 );
and \U$16608 ( \16985 , \16979 , \16984 );
and \U$16609 ( \16986 , \16975 , \16984 );
or \U$16610 ( \16987 , \16980 , \16985 , \16986 );
and \U$16611 ( \16988 , \16970 , \16987 );
and \U$16612 ( \16989 , \16954 , \16987 );
or \U$16613 ( \16990 , \16971 , \16988 , \16989 );
and \U$16614 ( \16991 , \16938 , \16990 );
and \U$16615 ( \16992 , \9620 , \2362 );
and \U$16616 ( \16993 , \9612 , \2360 );
nor \U$16617 ( \16994 , \16992 , \16993 );
xnor \U$16618 ( \16995 , \16994 , \2225 );
and \U$16619 ( \16996 , \10228 , \2156 );
and \U$16620 ( \16997 , \10223 , \2154 );
nor \U$16621 ( \16998 , \16996 , \16997 );
xnor \U$16622 ( \16999 , \16998 , \2004 );
and \U$16623 ( \17000 , \16995 , \16999 );
and \U$16624 ( \17001 , \11029 , \1888 );
and \U$16625 ( \17002 , \10409 , \1886 );
nor \U$16626 ( \17003 , \17001 , \17002 );
xnor \U$16627 ( \17004 , \17003 , \1732 );
and \U$16628 ( \17005 , \16999 , \17004 );
and \U$16629 ( \17006 , \16995 , \17004 );
or \U$16630 ( \17007 , \17000 , \17005 , \17006 );
xor \U$16631 ( \17008 , \16780 , \16784 );
xor \U$16632 ( \17009 , \17008 , \16789 );
and \U$16633 ( \17010 , \17007 , \17009 );
xor \U$16634 ( \17011 , \16796 , \16798 );
and \U$16635 ( \17012 , \17009 , \17011 );
and \U$16636 ( \17013 , \17007 , \17011 );
or \U$16637 ( \17014 , \17010 , \17012 , \17013 );
and \U$16638 ( \17015 , \16990 , \17014 );
and \U$16639 ( \17016 , \16938 , \17014 );
or \U$16640 ( \17017 , \16991 , \17015 , \17016 );
xor \U$16641 ( \17018 , \16731 , \16735 );
xor \U$16642 ( \17019 , \17018 , \1503 );
xor \U$16643 ( \17020 , \16743 , \16747 );
xor \U$16644 ( \17021 , \17020 , \16752 );
and \U$16645 ( \17022 , \17019 , \17021 );
xor \U$16646 ( \17023 , \16760 , \16764 );
xor \U$16647 ( \17024 , \17023 , \16769 );
and \U$16648 ( \17025 , \17021 , \17024 );
and \U$16649 ( \17026 , \17019 , \17024 );
or \U$16650 ( \17027 , \17022 , \17025 , \17026 );
xor \U$16651 ( \17028 , \16679 , \16683 );
xor \U$16652 ( \17029 , \17028 , \16688 );
xor \U$16653 ( \17030 , \16695 , \16699 );
xor \U$16654 ( \17031 , \17030 , \16704 );
and \U$16655 ( \17032 , \17029 , \17031 );
xor \U$16656 ( \17033 , \16712 , \16716 );
xor \U$16657 ( \17034 , \17033 , \16721 );
and \U$16658 ( \17035 , \17031 , \17034 );
and \U$16659 ( \17036 , \17029 , \17034 );
or \U$16660 ( \17037 , \17032 , \17035 , \17036 );
and \U$16661 ( \17038 , \17027 , \17037 );
xor \U$16662 ( \17039 , \16448 , \16452 );
xor \U$16663 ( \17040 , \17039 , \16457 );
and \U$16664 ( \17041 , \17037 , \17040 );
and \U$16665 ( \17042 , \17027 , \17040 );
or \U$16666 ( \17043 , \17038 , \17041 , \17042 );
and \U$16667 ( \17044 , \17017 , \17043 );
xor \U$16668 ( \17045 , \16792 , \16799 );
xor \U$16669 ( \17046 , \17045 , \16804 );
xor \U$16670 ( \17047 , \16812 , \16814 );
xor \U$16671 ( \17048 , \17047 , \16817 );
and \U$16672 ( \17049 , \17046 , \17048 );
xor \U$16673 ( \17050 , \16822 , \16824 );
xor \U$16674 ( \17051 , \17050 , \16827 );
and \U$16675 ( \17052 , \17048 , \17051 );
and \U$16676 ( \17053 , \17046 , \17051 );
or \U$16677 ( \17054 , \17049 , \17052 , \17053 );
and \U$16678 ( \17055 , \17043 , \17054 );
and \U$16679 ( \17056 , \17017 , \17054 );
or \U$16680 ( \17057 , \17044 , \17055 , \17056 );
xor \U$16681 ( \17058 , \16460 , \16476 );
xor \U$16682 ( \17059 , \17058 , \16493 );
xor \U$16683 ( \17060 , \16820 , \16830 );
xor \U$16684 ( \17061 , \17060 , \16833 );
and \U$16685 ( \17062 , \17059 , \17061 );
xor \U$16686 ( \17063 , \16839 , \16841 );
xor \U$16687 ( \17064 , \17063 , \16844 );
and \U$16688 ( \17065 , \17061 , \17064 );
and \U$16689 ( \17066 , \17059 , \17064 );
or \U$16690 ( \17067 , \17062 , \17065 , \17066 );
and \U$16691 ( \17068 , \17057 , \17067 );
xor \U$16692 ( \17069 , \16496 , \16548 );
xor \U$16693 ( \17070 , \17069 , \16573 );
and \U$16694 ( \17071 , \17067 , \17070 );
and \U$16695 ( \17072 , \17057 , \17070 );
or \U$16696 ( \17073 , \17068 , \17071 , \17072 );
xor \U$16697 ( \17074 , \16810 , \16836 );
xor \U$16698 ( \17075 , \17074 , \16847 );
xor \U$16699 ( \17076 , \16852 , \16854 );
xor \U$16700 ( \17077 , \17076 , \16857 );
and \U$16701 ( \17078 , \17075 , \17077 );
and \U$16702 ( \17079 , \17073 , \17078 );
xor \U$16703 ( \17080 , \16626 , \16628 );
xor \U$16704 ( \17081 , \17080 , \16631 );
and \U$16705 ( \17082 , \17078 , \17081 );
and \U$16706 ( \17083 , \17073 , \17081 );
or \U$16707 ( \17084 , \17079 , \17082 , \17083 );
xor \U$16708 ( \17085 , \16576 , \16602 );
xor \U$16709 ( \17086 , \17085 , \16613 );
xor \U$16710 ( \17087 , \16850 , \16860 );
xor \U$16711 ( \17088 , \17087 , \16863 );
and \U$16712 ( \17089 , \17086 , \17088 );
and \U$16713 ( \17090 , \17084 , \17089 );
xor \U$16714 ( \17091 , \16866 , \16868 );
xor \U$16715 ( \17092 , \17091 , \16871 );
and \U$16716 ( \17093 , \17089 , \17092 );
and \U$16717 ( \17094 , \17084 , \17092 );
or \U$16718 ( \17095 , \17090 , \17093 , \17094 );
and \U$16719 ( \17096 , \16886 , \17095 );
xor \U$16720 ( \17097 , \16886 , \17095 );
xor \U$16721 ( \17098 , \17084 , \17089 );
xor \U$16722 ( \17099 , \17098 , \17092 );
and \U$16723 ( \17100 , \3743 , \7829 );
and \U$16724 ( \17101 , \3326 , \7827 );
nor \U$16725 ( \17102 , \17100 , \17101 );
xnor \U$16726 ( \17103 , \17102 , \7580 );
and \U$16727 ( \17104 , \4073 , \7300 );
and \U$16728 ( \17105 , \3951 , \7298 );
nor \U$16729 ( \17106 , \17104 , \17105 );
xnor \U$16730 ( \17107 , \17106 , \7040 );
and \U$16731 ( \17108 , \17103 , \17107 );
and \U$16732 ( \17109 , \4334 , \6806 );
and \U$16733 ( \17110 , \4078 , \6804 );
nor \U$16734 ( \17111 , \17109 , \17110 );
xnor \U$16735 ( \17112 , \17111 , \6491 );
and \U$16736 ( \17113 , \17107 , \17112 );
and \U$16737 ( \17114 , \17103 , \17112 );
or \U$16738 ( \17115 , \17108 , \17113 , \17114 );
and \U$16739 ( \17116 , \2703 , \9495 );
and \U$16740 ( \17117 , \2439 , \9493 );
nor \U$16741 ( \17118 , \17116 , \17117 );
xnor \U$16742 ( \17119 , \17118 , \9185 );
and \U$16743 ( \17120 , \2902 , \8958 );
and \U$16744 ( \17121 , \2728 , \8956 );
nor \U$16745 ( \17122 , \17120 , \17121 );
xnor \U$16746 ( \17123 , \17122 , \8587 );
and \U$16747 ( \17124 , \17119 , \17123 );
and \U$16748 ( \17125 , \3207 , \8396 );
and \U$16749 ( \17126 , \3069 , \8394 );
nor \U$16750 ( \17127 , \17125 , \17126 );
xnor \U$16751 ( \17128 , \17127 , \8078 );
and \U$16752 ( \17129 , \17123 , \17128 );
and \U$16753 ( \17130 , \17119 , \17128 );
or \U$16754 ( \17131 , \17124 , \17129 , \17130 );
and \U$16755 ( \17132 , \17115 , \17131 );
and \U$16756 ( \17133 , \2104 , \10876 );
and \U$16757 ( \17134 , \1861 , \10873 );
nor \U$16758 ( \17135 , \17133 , \17134 );
xnor \U$16759 ( \17136 , \17135 , \9821 );
and \U$16760 ( \17137 , \2295 , \10063 );
and \U$16761 ( \17138 , \2109 , \10061 );
nor \U$16762 ( \17139 , \17137 , \17138 );
xnor \U$16763 ( \17140 , \17139 , \9824 );
and \U$16764 ( \17141 , \17136 , \17140 );
and \U$16765 ( \17142 , \17140 , \1732 );
and \U$16766 ( \17143 , \17136 , \1732 );
or \U$16767 ( \17144 , \17141 , \17142 , \17143 );
and \U$16768 ( \17145 , \17131 , \17144 );
and \U$16769 ( \17146 , \17115 , \17144 );
or \U$16770 ( \17147 , \17132 , \17145 , \17146 );
and \U$16771 ( \17148 , \7765 , \3699 );
and \U$16772 ( \17149 , \7239 , \3697 );
nor \U$16773 ( \17150 , \17148 , \17149 );
xnor \U$16774 ( \17151 , \17150 , \3512 );
and \U$16775 ( \17152 , \8435 , \3386 );
and \U$16776 ( \17153 , \8189 , \3384 );
nor \U$16777 ( \17154 , \17152 , \17153 );
xnor \U$16778 ( \17155 , \17154 , \3181 );
and \U$16779 ( \17156 , \17151 , \17155 );
and \U$16780 ( \17157 , \8759 , \2980 );
and \U$16781 ( \17158 , \8440 , \2978 );
nor \U$16782 ( \17159 , \17157 , \17158 );
xnor \U$16783 ( \17160 , \17159 , \2831 );
and \U$16784 ( \17161 , \17155 , \17160 );
and \U$16785 ( \17162 , \17151 , \17160 );
or \U$16786 ( \17163 , \17156 , \17161 , \17162 );
and \U$16787 ( \17164 , \4833 , \6297 );
and \U$16788 ( \17165 , \4531 , \6295 );
nor \U$16789 ( \17166 , \17164 , \17165 );
xnor \U$16790 ( \17167 , \17166 , \5957 );
and \U$16791 ( \17168 , \5310 , \5708 );
and \U$16792 ( \17169 , \4841 , \5706 );
nor \U$16793 ( \17170 , \17168 , \17169 );
xnor \U$16794 ( \17171 , \17170 , \5467 );
and \U$16795 ( \17172 , \17167 , \17171 );
and \U$16796 ( \17173 , \5579 , \5242 );
and \U$16797 ( \17174 , \5315 , \5240 );
nor \U$16798 ( \17175 , \17173 , \17174 );
xnor \U$16799 ( \17176 , \17175 , \5054 );
and \U$16800 ( \17177 , \17171 , \17176 );
and \U$16801 ( \17178 , \17167 , \17176 );
or \U$16802 ( \17179 , \17172 , \17177 , \17178 );
and \U$16803 ( \17180 , \17163 , \17179 );
and \U$16804 ( \17181 , \6210 , \4868 );
and \U$16805 ( \17182 , \5838 , \4866 );
nor \U$16806 ( \17183 , \17181 , \17182 );
xnor \U$16807 ( \17184 , \17183 , \4636 );
and \U$16808 ( \17185 , \6562 , \4417 );
and \U$16809 ( \17186 , \6219 , \4415 );
nor \U$16810 ( \17187 , \17185 , \17186 );
xnor \U$16811 ( \17188 , \17187 , \4274 );
and \U$16812 ( \17189 , \17184 , \17188 );
and \U$16813 ( \17190 , \7067 , \4094 );
and \U$16814 ( \17191 , \6764 , \4092 );
nor \U$16815 ( \17192 , \17190 , \17191 );
xnor \U$16816 ( \17193 , \17192 , \3848 );
and \U$16817 ( \17194 , \17188 , \17193 );
and \U$16818 ( \17195 , \17184 , \17193 );
or \U$16819 ( \17196 , \17189 , \17194 , \17195 );
and \U$16820 ( \17197 , \17179 , \17196 );
and \U$16821 ( \17198 , \17163 , \17196 );
or \U$16822 ( \17199 , \17180 , \17197 , \17198 );
and \U$16823 ( \17200 , \17147 , \17199 );
and \U$16824 ( \17201 , \9612 , \2658 );
and \U$16825 ( \17202 , \9043 , \2656 );
nor \U$16826 ( \17203 , \17201 , \17202 );
xnor \U$16827 ( \17204 , \17203 , \2516 );
and \U$16828 ( \17205 , \10223 , \2362 );
and \U$16829 ( \17206 , \9620 , \2360 );
nor \U$16830 ( \17207 , \17205 , \17206 );
xnor \U$16831 ( \17208 , \17207 , \2225 );
and \U$16832 ( \17209 , \17204 , \17208 );
and \U$16833 ( \17210 , \10409 , \2156 );
and \U$16834 ( \17211 , \10228 , \2154 );
nor \U$16835 ( \17212 , \17210 , \17211 );
xnor \U$16836 ( \17213 , \17212 , \2004 );
and \U$16837 ( \17214 , \17208 , \17213 );
and \U$16838 ( \17215 , \17204 , \17213 );
or \U$16839 ( \17216 , \17209 , \17214 , \17215 );
xor \U$16840 ( \17217 , \16906 , \16910 );
xor \U$16841 ( \17218 , \17217 , \16915 );
and \U$16842 ( \17219 , \17216 , \17218 );
xor \U$16843 ( \17220 , \16995 , \16999 );
xor \U$16844 ( \17221 , \17220 , \17004 );
and \U$16845 ( \17222 , \17218 , \17221 );
and \U$16846 ( \17223 , \17216 , \17221 );
or \U$16847 ( \17224 , \17219 , \17222 , \17223 );
and \U$16848 ( \17225 , \17199 , \17224 );
and \U$16849 ( \17226 , \17147 , \17224 );
or \U$16850 ( \17227 , \17200 , \17225 , \17226 );
xor \U$16851 ( \17228 , \16890 , \16894 );
xor \U$16852 ( \17229 , \17228 , \16899 );
xor \U$16853 ( \17230 , \16942 , \16946 );
xor \U$16854 ( \17231 , \17230 , \16951 );
and \U$16855 ( \17232 , \17229 , \17231 );
xor \U$16856 ( \17233 , \16923 , \16927 );
xor \U$16857 ( \17234 , \17233 , \16932 );
and \U$16858 ( \17235 , \17231 , \17234 );
and \U$16859 ( \17236 , \17229 , \17234 );
or \U$16860 ( \17237 , \17232 , \17235 , \17236 );
xor \U$16861 ( \17238 , \16958 , \16962 );
xor \U$16862 ( \17239 , \17238 , \16967 );
xor \U$16863 ( \17240 , \16975 , \16979 );
xor \U$16864 ( \17241 , \17240 , \16984 );
and \U$16865 ( \17242 , \17239 , \17241 );
and \U$16866 ( \17243 , \17237 , \17242 );
xor \U$16867 ( \17244 , \17019 , \17021 );
xor \U$16868 ( \17245 , \17244 , \17024 );
and \U$16869 ( \17246 , \17242 , \17245 );
and \U$16870 ( \17247 , \17237 , \17245 );
or \U$16871 ( \17248 , \17243 , \17246 , \17247 );
and \U$16872 ( \17249 , \17227 , \17248 );
xor \U$16873 ( \17250 , \16902 , \16918 );
xor \U$16874 ( \17251 , \17250 , \16935 );
xor \U$16875 ( \17252 , \17029 , \17031 );
xor \U$16876 ( \17253 , \17252 , \17034 );
and \U$16877 ( \17254 , \17251 , \17253 );
xor \U$16878 ( \17255 , \17007 , \17009 );
xor \U$16879 ( \17256 , \17255 , \17011 );
and \U$16880 ( \17257 , \17253 , \17256 );
and \U$16881 ( \17258 , \17251 , \17256 );
or \U$16882 ( \17259 , \17254 , \17257 , \17258 );
and \U$16883 ( \17260 , \17248 , \17259 );
and \U$16884 ( \17261 , \17227 , \17259 );
or \U$16885 ( \17262 , \17249 , \17260 , \17261 );
xor \U$16886 ( \17263 , \16691 , \16707 );
xor \U$16887 ( \17264 , \17263 , \16724 );
xor \U$16888 ( \17265 , \16739 , \16755 );
xor \U$16889 ( \17266 , \17265 , \16772 );
and \U$16890 ( \17267 , \17264 , \17266 );
xor \U$16891 ( \17268 , \17046 , \17048 );
xor \U$16892 ( \17269 , \17268 , \17051 );
and \U$16893 ( \17270 , \17266 , \17269 );
and \U$16894 ( \17271 , \17264 , \17269 );
or \U$16895 ( \17272 , \17267 , \17270 , \17271 );
and \U$16896 ( \17273 , \17262 , \17272 );
xor \U$16897 ( \17274 , \16727 , \16775 );
xor \U$16898 ( \17275 , \17274 , \16807 );
and \U$16899 ( \17276 , \17272 , \17275 );
and \U$16900 ( \17277 , \17262 , \17275 );
or \U$16901 ( \17278 , \17273 , \17276 , \17277 );
xor \U$16902 ( \17279 , \17057 , \17067 );
xor \U$16903 ( \17280 , \17279 , \17070 );
and \U$16904 ( \17281 , \17278 , \17280 );
xor \U$16905 ( \17282 , \17075 , \17077 );
and \U$16906 ( \17283 , \17280 , \17282 );
and \U$16907 ( \17284 , \17278 , \17282 );
or \U$16908 ( \17285 , \17281 , \17283 , \17284 );
xor \U$16909 ( \17286 , \17073 , \17078 );
xor \U$16910 ( \17287 , \17286 , \17081 );
and \U$16911 ( \17288 , \17285 , \17287 );
xor \U$16912 ( \17289 , \17086 , \17088 );
and \U$16913 ( \17290 , \17287 , \17289 );
and \U$16914 ( \17291 , \17285 , \17289 );
or \U$16915 ( \17292 , \17288 , \17290 , \17291 );
and \U$16916 ( \17293 , \17099 , \17292 );
xor \U$16917 ( \17294 , \17099 , \17292 );
xor \U$16918 ( \17295 , \17285 , \17287 );
xor \U$16919 ( \17296 , \17295 , \17289 );
and \U$16920 ( \17297 , \2109 , \10876 );
and \U$16921 ( \17298 , \2104 , \10873 );
nor \U$16922 ( \17299 , \17297 , \17298 );
xnor \U$16923 ( \17300 , \17299 , \9821 );
and \U$16924 ( \17301 , \2439 , \10063 );
and \U$16925 ( \17302 , \2295 , \10061 );
nor \U$16926 ( \17303 , \17301 , \17302 );
xnor \U$16927 ( \17304 , \17303 , \9824 );
and \U$16928 ( \17305 , \17300 , \17304 );
and \U$16929 ( \17306 , \2728 , \9495 );
and \U$16930 ( \17307 , \2703 , \9493 );
nor \U$16931 ( \17308 , \17306 , \17307 );
xnor \U$16932 ( \17309 , \17308 , \9185 );
and \U$16933 ( \17310 , \17304 , \17309 );
and \U$16934 ( \17311 , \17300 , \17309 );
or \U$16935 ( \17312 , \17305 , \17310 , \17311 );
and \U$16936 ( \17313 , \3069 , \8958 );
and \U$16937 ( \17314 , \2902 , \8956 );
nor \U$16938 ( \17315 , \17313 , \17314 );
xnor \U$16939 ( \17316 , \17315 , \8587 );
and \U$16940 ( \17317 , \3326 , \8396 );
and \U$16941 ( \17318 , \3207 , \8394 );
nor \U$16942 ( \17319 , \17317 , \17318 );
xnor \U$16943 ( \17320 , \17319 , \8078 );
and \U$16944 ( \17321 , \17316 , \17320 );
and \U$16945 ( \17322 , \3951 , \7829 );
and \U$16946 ( \17323 , \3743 , \7827 );
nor \U$16947 ( \17324 , \17322 , \17323 );
xnor \U$16948 ( \17325 , \17324 , \7580 );
and \U$16949 ( \17326 , \17320 , \17325 );
and \U$16950 ( \17327 , \17316 , \17325 );
or \U$16951 ( \17328 , \17321 , \17326 , \17327 );
and \U$16952 ( \17329 , \17312 , \17328 );
and \U$16953 ( \17330 , \4078 , \7300 );
and \U$16954 ( \17331 , \4073 , \7298 );
nor \U$16955 ( \17332 , \17330 , \17331 );
xnor \U$16956 ( \17333 , \17332 , \7040 );
and \U$16957 ( \17334 , \4531 , \6806 );
and \U$16958 ( \17335 , \4334 , \6804 );
nor \U$16959 ( \17336 , \17334 , \17335 );
xnor \U$16960 ( \17337 , \17336 , \6491 );
and \U$16961 ( \17338 , \17333 , \17337 );
and \U$16962 ( \17339 , \4841 , \6297 );
and \U$16963 ( \17340 , \4833 , \6295 );
nor \U$16964 ( \17341 , \17339 , \17340 );
xnor \U$16965 ( \17342 , \17341 , \5957 );
and \U$16966 ( \17343 , \17337 , \17342 );
and \U$16967 ( \17344 , \17333 , \17342 );
or \U$16968 ( \17345 , \17338 , \17343 , \17344 );
and \U$16969 ( \17346 , \17328 , \17345 );
and \U$16970 ( \17347 , \17312 , \17345 );
or \U$16971 ( \17348 , \17329 , \17346 , \17347 );
and \U$16972 ( \17349 , \6764 , \4417 );
and \U$16973 ( \17350 , \6562 , \4415 );
nor \U$16974 ( \17351 , \17349 , \17350 );
xnor \U$16975 ( \17352 , \17351 , \4274 );
and \U$16976 ( \17353 , \7239 , \4094 );
and \U$16977 ( \17354 , \7067 , \4092 );
nor \U$16978 ( \17355 , \17353 , \17354 );
xnor \U$16979 ( \17356 , \17355 , \3848 );
and \U$16980 ( \17357 , \17352 , \17356 );
and \U$16981 ( \17358 , \8189 , \3699 );
and \U$16982 ( \17359 , \7765 , \3697 );
nor \U$16983 ( \17360 , \17358 , \17359 );
xnor \U$16984 ( \17361 , \17360 , \3512 );
and \U$16985 ( \17362 , \17356 , \17361 );
and \U$16986 ( \17363 , \17352 , \17361 );
or \U$16987 ( \17364 , \17357 , \17362 , \17363 );
and \U$16988 ( \17365 , \5315 , \5708 );
and \U$16989 ( \17366 , \5310 , \5706 );
nor \U$16990 ( \17367 , \17365 , \17366 );
xnor \U$16991 ( \17368 , \17367 , \5467 );
and \U$16992 ( \17369 , \5838 , \5242 );
and \U$16993 ( \17370 , \5579 , \5240 );
nor \U$16994 ( \17371 , \17369 , \17370 );
xnor \U$16995 ( \17372 , \17371 , \5054 );
and \U$16996 ( \17373 , \17368 , \17372 );
and \U$16997 ( \17374 , \6219 , \4868 );
and \U$16998 ( \17375 , \6210 , \4866 );
nor \U$16999 ( \17376 , \17374 , \17375 );
xnor \U$17000 ( \17377 , \17376 , \4636 );
and \U$17001 ( \17378 , \17372 , \17377 );
and \U$17002 ( \17379 , \17368 , \17377 );
or \U$17003 ( \17380 , \17373 , \17378 , \17379 );
and \U$17004 ( \17381 , \17364 , \17380 );
and \U$17005 ( \17382 , \8440 , \3386 );
and \U$17006 ( \17383 , \8435 , \3384 );
nor \U$17007 ( \17384 , \17382 , \17383 );
xnor \U$17008 ( \17385 , \17384 , \3181 );
and \U$17009 ( \17386 , \9043 , \2980 );
and \U$17010 ( \17387 , \8759 , \2978 );
nor \U$17011 ( \17388 , \17386 , \17387 );
xnor \U$17012 ( \17389 , \17388 , \2831 );
and \U$17013 ( \17390 , \17385 , \17389 );
and \U$17014 ( \17391 , \9620 , \2658 );
and \U$17015 ( \17392 , \9612 , \2656 );
nor \U$17016 ( \17393 , \17391 , \17392 );
xnor \U$17017 ( \17394 , \17393 , \2516 );
and \U$17018 ( \17395 , \17389 , \17394 );
and \U$17019 ( \17396 , \17385 , \17394 );
or \U$17020 ( \17397 , \17390 , \17395 , \17396 );
and \U$17021 ( \17398 , \17380 , \17397 );
and \U$17022 ( \17399 , \17364 , \17397 );
or \U$17023 ( \17400 , \17381 , \17398 , \17399 );
and \U$17024 ( \17401 , \17348 , \17400 );
nand \U$17025 ( \17402 , \11029 , \1886 );
xnor \U$17026 ( \17403 , \17402 , \1732 );
xor \U$17027 ( \17404 , \17151 , \17155 );
xor \U$17028 ( \17405 , \17404 , \17160 );
and \U$17029 ( \17406 , \17403 , \17405 );
xor \U$17030 ( \17407 , \17204 , \17208 );
xor \U$17031 ( \17408 , \17407 , \17213 );
and \U$17032 ( \17409 , \17405 , \17408 );
and \U$17033 ( \17410 , \17403 , \17408 );
or \U$17034 ( \17411 , \17406 , \17409 , \17410 );
and \U$17035 ( \17412 , \17400 , \17411 );
and \U$17036 ( \17413 , \17348 , \17411 );
or \U$17037 ( \17414 , \17401 , \17412 , \17413 );
xor \U$17038 ( \17415 , \17115 , \17131 );
xor \U$17039 ( \17416 , \17415 , \17144 );
xor \U$17040 ( \17417 , \17163 , \17179 );
xor \U$17041 ( \17418 , \17417 , \17196 );
and \U$17042 ( \17419 , \17416 , \17418 );
xor \U$17043 ( \17420 , \17216 , \17218 );
xor \U$17044 ( \17421 , \17420 , \17221 );
and \U$17045 ( \17422 , \17418 , \17421 );
and \U$17046 ( \17423 , \17416 , \17421 );
or \U$17047 ( \17424 , \17419 , \17422 , \17423 );
and \U$17048 ( \17425 , \17414 , \17424 );
xor \U$17049 ( \17426 , \17103 , \17107 );
xor \U$17050 ( \17427 , \17426 , \17112 );
xor \U$17051 ( \17428 , \17167 , \17171 );
xor \U$17052 ( \17429 , \17428 , \17176 );
and \U$17053 ( \17430 , \17427 , \17429 );
xor \U$17054 ( \17431 , \17184 , \17188 );
xor \U$17055 ( \17432 , \17431 , \17193 );
and \U$17056 ( \17433 , \17429 , \17432 );
and \U$17057 ( \17434 , \17427 , \17432 );
or \U$17058 ( \17435 , \17430 , \17433 , \17434 );
xor \U$17059 ( \17436 , \17229 , \17231 );
xor \U$17060 ( \17437 , \17436 , \17234 );
and \U$17061 ( \17438 , \17435 , \17437 );
xor \U$17062 ( \17439 , \17239 , \17241 );
and \U$17063 ( \17440 , \17437 , \17439 );
and \U$17064 ( \17441 , \17435 , \17439 );
or \U$17065 ( \17442 , \17438 , \17440 , \17441 );
and \U$17066 ( \17443 , \17424 , \17442 );
and \U$17067 ( \17444 , \17414 , \17442 );
or \U$17068 ( \17445 , \17425 , \17443 , \17444 );
xor \U$17069 ( \17446 , \16954 , \16970 );
xor \U$17070 ( \17447 , \17446 , \16987 );
xor \U$17071 ( \17448 , \17237 , \17242 );
xor \U$17072 ( \17449 , \17448 , \17245 );
and \U$17073 ( \17450 , \17447 , \17449 );
xor \U$17074 ( \17451 , \17251 , \17253 );
xor \U$17075 ( \17452 , \17451 , \17256 );
and \U$17076 ( \17453 , \17449 , \17452 );
and \U$17077 ( \17454 , \17447 , \17452 );
or \U$17078 ( \17455 , \17450 , \17453 , \17454 );
and \U$17079 ( \17456 , \17445 , \17455 );
xor \U$17080 ( \17457 , \17027 , \17037 );
xor \U$17081 ( \17458 , \17457 , \17040 );
and \U$17082 ( \17459 , \17455 , \17458 );
and \U$17083 ( \17460 , \17445 , \17458 );
or \U$17084 ( \17461 , \17456 , \17459 , \17460 );
xor \U$17085 ( \17462 , \16938 , \16990 );
xor \U$17086 ( \17463 , \17462 , \17014 );
xor \U$17087 ( \17464 , \17227 , \17248 );
xor \U$17088 ( \17465 , \17464 , \17259 );
and \U$17089 ( \17466 , \17463 , \17465 );
xor \U$17090 ( \17467 , \17264 , \17266 );
xor \U$17091 ( \17468 , \17467 , \17269 );
and \U$17092 ( \17469 , \17465 , \17468 );
and \U$17093 ( \17470 , \17463 , \17468 );
or \U$17094 ( \17471 , \17466 , \17469 , \17470 );
and \U$17095 ( \17472 , \17461 , \17471 );
xor \U$17096 ( \17473 , \17059 , \17061 );
xor \U$17097 ( \17474 , \17473 , \17064 );
and \U$17098 ( \17475 , \17471 , \17474 );
and \U$17099 ( \17476 , \17461 , \17474 );
or \U$17100 ( \17477 , \17472 , \17475 , \17476 );
xor \U$17101 ( \17478 , \17017 , \17043 );
xor \U$17102 ( \17479 , \17478 , \17054 );
xor \U$17103 ( \17480 , \17262 , \17272 );
xor \U$17104 ( \17481 , \17480 , \17275 );
and \U$17105 ( \17482 , \17479 , \17481 );
and \U$17106 ( \17483 , \17477 , \17482 );
xor \U$17107 ( \17484 , \17278 , \17280 );
xor \U$17108 ( \17485 , \17484 , \17282 );
and \U$17109 ( \17486 , \17482 , \17485 );
and \U$17110 ( \17487 , \17477 , \17485 );
or \U$17111 ( \17488 , \17483 , \17486 , \17487 );
and \U$17112 ( \17489 , \17296 , \17488 );
xor \U$17113 ( \17490 , \17296 , \17488 );
xor \U$17114 ( \17491 , \17477 , \17482 );
xor \U$17115 ( \17492 , \17491 , \17485 );
and \U$17116 ( \17493 , \2295 , \10876 );
and \U$17117 ( \17494 , \2109 , \10873 );
nor \U$17118 ( \17495 , \17493 , \17494 );
xnor \U$17119 ( \17496 , \17495 , \9821 );
and \U$17120 ( \17497 , \2703 , \10063 );
and \U$17121 ( \17498 , \2439 , \10061 );
nor \U$17122 ( \17499 , \17497 , \17498 );
xnor \U$17123 ( \17500 , \17499 , \9824 );
and \U$17124 ( \17501 , \17496 , \17500 );
and \U$17125 ( \17502 , \17500 , \2004 );
and \U$17126 ( \17503 , \17496 , \2004 );
or \U$17127 ( \17504 , \17501 , \17502 , \17503 );
and \U$17128 ( \17505 , \4073 , \7829 );
and \U$17129 ( \17506 , \3951 , \7827 );
nor \U$17130 ( \17507 , \17505 , \17506 );
xnor \U$17131 ( \17508 , \17507 , \7580 );
and \U$17132 ( \17509 , \4334 , \7300 );
and \U$17133 ( \17510 , \4078 , \7298 );
nor \U$17134 ( \17511 , \17509 , \17510 );
xnor \U$17135 ( \17512 , \17511 , \7040 );
and \U$17136 ( \17513 , \17508 , \17512 );
and \U$17137 ( \17514 , \4833 , \6806 );
and \U$17138 ( \17515 , \4531 , \6804 );
nor \U$17139 ( \17516 , \17514 , \17515 );
xnor \U$17140 ( \17517 , \17516 , \6491 );
and \U$17141 ( \17518 , \17512 , \17517 );
and \U$17142 ( \17519 , \17508 , \17517 );
or \U$17143 ( \17520 , \17513 , \17518 , \17519 );
and \U$17144 ( \17521 , \17504 , \17520 );
and \U$17145 ( \17522 , \2902 , \9495 );
and \U$17146 ( \17523 , \2728 , \9493 );
nor \U$17147 ( \17524 , \17522 , \17523 );
xnor \U$17148 ( \17525 , \17524 , \9185 );
and \U$17149 ( \17526 , \3207 , \8958 );
and \U$17150 ( \17527 , \3069 , \8956 );
nor \U$17151 ( \17528 , \17526 , \17527 );
xnor \U$17152 ( \17529 , \17528 , \8587 );
and \U$17153 ( \17530 , \17525 , \17529 );
and \U$17154 ( \17531 , \3743 , \8396 );
and \U$17155 ( \17532 , \3326 , \8394 );
nor \U$17156 ( \17533 , \17531 , \17532 );
xnor \U$17157 ( \17534 , \17533 , \8078 );
and \U$17158 ( \17535 , \17529 , \17534 );
and \U$17159 ( \17536 , \17525 , \17534 );
or \U$17160 ( \17537 , \17530 , \17535 , \17536 );
and \U$17161 ( \17538 , \17520 , \17537 );
and \U$17162 ( \17539 , \17504 , \17537 );
or \U$17163 ( \17540 , \17521 , \17538 , \17539 );
and \U$17164 ( \17541 , \10223 , \2658 );
and \U$17165 ( \17542 , \9620 , \2656 );
nor \U$17166 ( \17543 , \17541 , \17542 );
xnor \U$17167 ( \17544 , \17543 , \2516 );
and \U$17168 ( \17545 , \10409 , \2362 );
and \U$17169 ( \17546 , \10228 , \2360 );
nor \U$17170 ( \17547 , \17545 , \17546 );
xnor \U$17171 ( \17548 , \17547 , \2225 );
and \U$17172 ( \17549 , \17544 , \17548 );
nand \U$17173 ( \17550 , \11029 , \2154 );
xnor \U$17174 ( \17551 , \17550 , \2004 );
and \U$17175 ( \17552 , \17548 , \17551 );
and \U$17176 ( \17553 , \17544 , \17551 );
or \U$17177 ( \17554 , \17549 , \17552 , \17553 );
and \U$17178 ( \17555 , \10228 , \2362 );
and \U$17179 ( \17556 , \10223 , \2360 );
nor \U$17180 ( \17557 , \17555 , \17556 );
xnor \U$17181 ( \17558 , \17557 , \2225 );
and \U$17182 ( \17559 , \17554 , \17558 );
and \U$17183 ( \17560 , \11029 , \2156 );
and \U$17184 ( \17561 , \10409 , \2154 );
nor \U$17185 ( \17562 , \17560 , \17561 );
xnor \U$17186 ( \17563 , \17562 , \2004 );
and \U$17187 ( \17564 , \17558 , \17563 );
and \U$17188 ( \17565 , \17554 , \17563 );
or \U$17189 ( \17566 , \17559 , \17564 , \17565 );
and \U$17190 ( \17567 , \17540 , \17566 );
and \U$17191 ( \17568 , \5310 , \6297 );
and \U$17192 ( \17569 , \4841 , \6295 );
nor \U$17193 ( \17570 , \17568 , \17569 );
xnor \U$17194 ( \17571 , \17570 , \5957 );
and \U$17195 ( \17572 , \5579 , \5708 );
and \U$17196 ( \17573 , \5315 , \5706 );
nor \U$17197 ( \17574 , \17572 , \17573 );
xnor \U$17198 ( \17575 , \17574 , \5467 );
and \U$17199 ( \17576 , \17571 , \17575 );
and \U$17200 ( \17577 , \6210 , \5242 );
and \U$17201 ( \17578 , \5838 , \5240 );
nor \U$17202 ( \17579 , \17577 , \17578 );
xnor \U$17203 ( \17580 , \17579 , \5054 );
and \U$17204 ( \17581 , \17575 , \17580 );
and \U$17205 ( \17582 , \17571 , \17580 );
or \U$17206 ( \17583 , \17576 , \17581 , \17582 );
and \U$17207 ( \17584 , \8435 , \3699 );
and \U$17208 ( \17585 , \8189 , \3697 );
nor \U$17209 ( \17586 , \17584 , \17585 );
xnor \U$17210 ( \17587 , \17586 , \3512 );
and \U$17211 ( \17588 , \8759 , \3386 );
and \U$17212 ( \17589 , \8440 , \3384 );
nor \U$17213 ( \17590 , \17588 , \17589 );
xnor \U$17214 ( \17591 , \17590 , \3181 );
and \U$17215 ( \17592 , \17587 , \17591 );
and \U$17216 ( \17593 , \9612 , \2980 );
and \U$17217 ( \17594 , \9043 , \2978 );
nor \U$17218 ( \17595 , \17593 , \17594 );
xnor \U$17219 ( \17596 , \17595 , \2831 );
and \U$17220 ( \17597 , \17591 , \17596 );
and \U$17221 ( \17598 , \17587 , \17596 );
or \U$17222 ( \17599 , \17592 , \17597 , \17598 );
and \U$17223 ( \17600 , \17583 , \17599 );
and \U$17224 ( \17601 , \6562 , \4868 );
and \U$17225 ( \17602 , \6219 , \4866 );
nor \U$17226 ( \17603 , \17601 , \17602 );
xnor \U$17227 ( \17604 , \17603 , \4636 );
and \U$17228 ( \17605 , \7067 , \4417 );
and \U$17229 ( \17606 , \6764 , \4415 );
nor \U$17230 ( \17607 , \17605 , \17606 );
xnor \U$17231 ( \17608 , \17607 , \4274 );
and \U$17232 ( \17609 , \17604 , \17608 );
and \U$17233 ( \17610 , \7765 , \4094 );
and \U$17234 ( \17611 , \7239 , \4092 );
nor \U$17235 ( \17612 , \17610 , \17611 );
xnor \U$17236 ( \17613 , \17612 , \3848 );
and \U$17237 ( \17614 , \17608 , \17613 );
and \U$17238 ( \17615 , \17604 , \17613 );
or \U$17239 ( \17616 , \17609 , \17614 , \17615 );
and \U$17240 ( \17617 , \17599 , \17616 );
and \U$17241 ( \17618 , \17583 , \17616 );
or \U$17242 ( \17619 , \17600 , \17617 , \17618 );
and \U$17243 ( \17620 , \17566 , \17619 );
and \U$17244 ( \17621 , \17540 , \17619 );
or \U$17245 ( \17622 , \17567 , \17620 , \17621 );
xor \U$17246 ( \17623 , \17300 , \17304 );
xor \U$17247 ( \17624 , \17623 , \17309 );
xor \U$17248 ( \17625 , \17316 , \17320 );
xor \U$17249 ( \17626 , \17625 , \17325 );
and \U$17250 ( \17627 , \17624 , \17626 );
xor \U$17251 ( \17628 , \17333 , \17337 );
xor \U$17252 ( \17629 , \17628 , \17342 );
and \U$17253 ( \17630 , \17626 , \17629 );
and \U$17254 ( \17631 , \17624 , \17629 );
or \U$17255 ( \17632 , \17627 , \17630 , \17631 );
xor \U$17256 ( \17633 , \17352 , \17356 );
xor \U$17257 ( \17634 , \17633 , \17361 );
xor \U$17258 ( \17635 , \17368 , \17372 );
xor \U$17259 ( \17636 , \17635 , \17377 );
and \U$17260 ( \17637 , \17634 , \17636 );
xor \U$17261 ( \17638 , \17385 , \17389 );
xor \U$17262 ( \17639 , \17638 , \17394 );
and \U$17263 ( \17640 , \17636 , \17639 );
and \U$17264 ( \17641 , \17634 , \17639 );
or \U$17265 ( \17642 , \17637 , \17640 , \17641 );
and \U$17266 ( \17643 , \17632 , \17642 );
xor \U$17267 ( \17644 , \17119 , \17123 );
xor \U$17268 ( \17645 , \17644 , \17128 );
and \U$17269 ( \17646 , \17642 , \17645 );
and \U$17270 ( \17647 , \17632 , \17645 );
or \U$17271 ( \17648 , \17643 , \17646 , \17647 );
and \U$17272 ( \17649 , \17622 , \17648 );
xor \U$17273 ( \17650 , \17136 , \17140 );
xor \U$17274 ( \17651 , \17650 , \1732 );
xor \U$17275 ( \17652 , \17427 , \17429 );
xor \U$17276 ( \17653 , \17652 , \17432 );
and \U$17277 ( \17654 , \17651 , \17653 );
xor \U$17278 ( \17655 , \17403 , \17405 );
xor \U$17279 ( \17656 , \17655 , \17408 );
and \U$17280 ( \17657 , \17653 , \17656 );
and \U$17281 ( \17658 , \17651 , \17656 );
or \U$17282 ( \17659 , \17654 , \17657 , \17658 );
and \U$17283 ( \17660 , \17648 , \17659 );
and \U$17284 ( \17661 , \17622 , \17659 );
or \U$17285 ( \17662 , \17649 , \17660 , \17661 );
xor \U$17286 ( \17663 , \17348 , \17400 );
xor \U$17287 ( \17664 , \17663 , \17411 );
xor \U$17288 ( \17665 , \17416 , \17418 );
xor \U$17289 ( \17666 , \17665 , \17421 );
and \U$17290 ( \17667 , \17664 , \17666 );
xor \U$17291 ( \17668 , \17435 , \17437 );
xor \U$17292 ( \17669 , \17668 , \17439 );
and \U$17293 ( \17670 , \17666 , \17669 );
and \U$17294 ( \17671 , \17664 , \17669 );
or \U$17295 ( \17672 , \17667 , \17670 , \17671 );
and \U$17296 ( \17673 , \17662 , \17672 );
xor \U$17297 ( \17674 , \17147 , \17199 );
xor \U$17298 ( \17675 , \17674 , \17224 );
and \U$17299 ( \17676 , \17672 , \17675 );
and \U$17300 ( \17677 , \17662 , \17675 );
or \U$17301 ( \17678 , \17673 , \17676 , \17677 );
xor \U$17302 ( \17679 , \17414 , \17424 );
xor \U$17303 ( \17680 , \17679 , \17442 );
xor \U$17304 ( \17681 , \17447 , \17449 );
xor \U$17305 ( \17682 , \17681 , \17452 );
and \U$17306 ( \17683 , \17680 , \17682 );
and \U$17307 ( \17684 , \17678 , \17683 );
xor \U$17308 ( \17685 , \17463 , \17465 );
xor \U$17309 ( \17686 , \17685 , \17468 );
and \U$17310 ( \17687 , \17683 , \17686 );
and \U$17311 ( \17688 , \17678 , \17686 );
or \U$17312 ( \17689 , \17684 , \17687 , \17688 );
xor \U$17313 ( \17690 , \17461 , \17471 );
xor \U$17314 ( \17691 , \17690 , \17474 );
and \U$17315 ( \17692 , \17689 , \17691 );
xor \U$17316 ( \17693 , \17479 , \17481 );
and \U$17317 ( \17694 , \17691 , \17693 );
and \U$17318 ( \17695 , \17689 , \17693 );
or \U$17319 ( \17696 , \17692 , \17694 , \17695 );
and \U$17320 ( \17697 , \17492 , \17696 );
xor \U$17321 ( \17698 , \17492 , \17696 );
xor \U$17322 ( \17699 , \17689 , \17691 );
xor \U$17323 ( \17700 , \17699 , \17693 );
and \U$17324 ( \17701 , \9043 , \3386 );
and \U$17325 ( \17702 , \8759 , \3384 );
nor \U$17326 ( \17703 , \17701 , \17702 );
xnor \U$17327 ( \17704 , \17703 , \3181 );
and \U$17328 ( \17705 , \9620 , \2980 );
and \U$17329 ( \17706 , \9612 , \2978 );
nor \U$17330 ( \17707 , \17705 , \17706 );
xnor \U$17331 ( \17708 , \17707 , \2831 );
and \U$17332 ( \17709 , \17704 , \17708 );
and \U$17333 ( \17710 , \10228 , \2658 );
and \U$17334 ( \17711 , \10223 , \2656 );
nor \U$17335 ( \17712 , \17710 , \17711 );
xnor \U$17336 ( \17713 , \17712 , \2516 );
and \U$17337 ( \17714 , \17708 , \17713 );
and \U$17338 ( \17715 , \17704 , \17713 );
or \U$17339 ( \17716 , \17709 , \17714 , \17715 );
and \U$17340 ( \17717 , \5838 , \5708 );
and \U$17341 ( \17718 , \5579 , \5706 );
nor \U$17342 ( \17719 , \17717 , \17718 );
xnor \U$17343 ( \17720 , \17719 , \5467 );
and \U$17344 ( \17721 , \6219 , \5242 );
and \U$17345 ( \17722 , \6210 , \5240 );
nor \U$17346 ( \17723 , \17721 , \17722 );
xnor \U$17347 ( \17724 , \17723 , \5054 );
and \U$17348 ( \17725 , \17720 , \17724 );
and \U$17349 ( \17726 , \6764 , \4868 );
and \U$17350 ( \17727 , \6562 , \4866 );
nor \U$17351 ( \17728 , \17726 , \17727 );
xnor \U$17352 ( \17729 , \17728 , \4636 );
and \U$17353 ( \17730 , \17724 , \17729 );
and \U$17354 ( \17731 , \17720 , \17729 );
or \U$17355 ( \17732 , \17725 , \17730 , \17731 );
and \U$17356 ( \17733 , \17716 , \17732 );
and \U$17357 ( \17734 , \7239 , \4417 );
and \U$17358 ( \17735 , \7067 , \4415 );
nor \U$17359 ( \17736 , \17734 , \17735 );
xnor \U$17360 ( \17737 , \17736 , \4274 );
and \U$17361 ( \17738 , \8189 , \4094 );
and \U$17362 ( \17739 , \7765 , \4092 );
nor \U$17363 ( \17740 , \17738 , \17739 );
xnor \U$17364 ( \17741 , \17740 , \3848 );
and \U$17365 ( \17742 , \17737 , \17741 );
and \U$17366 ( \17743 , \8440 , \3699 );
and \U$17367 ( \17744 , \8435 , \3697 );
nor \U$17368 ( \17745 , \17743 , \17744 );
xnor \U$17369 ( \17746 , \17745 , \3512 );
and \U$17370 ( \17747 , \17741 , \17746 );
and \U$17371 ( \17748 , \17737 , \17746 );
or \U$17372 ( \17749 , \17742 , \17747 , \17748 );
and \U$17373 ( \17750 , \17732 , \17749 );
and \U$17374 ( \17751 , \17716 , \17749 );
or \U$17375 ( \17752 , \17733 , \17750 , \17751 );
and \U$17376 ( \17753 , \4531 , \7300 );
and \U$17377 ( \17754 , \4334 , \7298 );
nor \U$17378 ( \17755 , \17753 , \17754 );
xnor \U$17379 ( \17756 , \17755 , \7040 );
and \U$17380 ( \17757 , \4841 , \6806 );
and \U$17381 ( \17758 , \4833 , \6804 );
nor \U$17382 ( \17759 , \17757 , \17758 );
xnor \U$17383 ( \17760 , \17759 , \6491 );
and \U$17384 ( \17761 , \17756 , \17760 );
and \U$17385 ( \17762 , \5315 , \6297 );
and \U$17386 ( \17763 , \5310 , \6295 );
nor \U$17387 ( \17764 , \17762 , \17763 );
xnor \U$17388 ( \17765 , \17764 , \5957 );
and \U$17389 ( \17766 , \17760 , \17765 );
and \U$17390 ( \17767 , \17756 , \17765 );
or \U$17391 ( \17768 , \17761 , \17766 , \17767 );
and \U$17392 ( \17769 , \3326 , \8958 );
and \U$17393 ( \17770 , \3207 , \8956 );
nor \U$17394 ( \17771 , \17769 , \17770 );
xnor \U$17395 ( \17772 , \17771 , \8587 );
and \U$17396 ( \17773 , \3951 , \8396 );
and \U$17397 ( \17774 , \3743 , \8394 );
nor \U$17398 ( \17775 , \17773 , \17774 );
xnor \U$17399 ( \17776 , \17775 , \8078 );
and \U$17400 ( \17777 , \17772 , \17776 );
and \U$17401 ( \17778 , \4078 , \7829 );
and \U$17402 ( \17779 , \4073 , \7827 );
nor \U$17403 ( \17780 , \17778 , \17779 );
xnor \U$17404 ( \17781 , \17780 , \7580 );
and \U$17405 ( \17782 , \17776 , \17781 );
and \U$17406 ( \17783 , \17772 , \17781 );
or \U$17407 ( \17784 , \17777 , \17782 , \17783 );
and \U$17408 ( \17785 , \17768 , \17784 );
and \U$17409 ( \17786 , \2439 , \10876 );
and \U$17410 ( \17787 , \2295 , \10873 );
nor \U$17411 ( \17788 , \17786 , \17787 );
xnor \U$17412 ( \17789 , \17788 , \9821 );
and \U$17413 ( \17790 , \2728 , \10063 );
and \U$17414 ( \17791 , \2703 , \10061 );
nor \U$17415 ( \17792 , \17790 , \17791 );
xnor \U$17416 ( \17793 , \17792 , \9824 );
and \U$17417 ( \17794 , \17789 , \17793 );
and \U$17418 ( \17795 , \3069 , \9495 );
and \U$17419 ( \17796 , \2902 , \9493 );
nor \U$17420 ( \17797 , \17795 , \17796 );
xnor \U$17421 ( \17798 , \17797 , \9185 );
and \U$17422 ( \17799 , \17793 , \17798 );
and \U$17423 ( \17800 , \17789 , \17798 );
or \U$17424 ( \17801 , \17794 , \17799 , \17800 );
and \U$17425 ( \17802 , \17784 , \17801 );
and \U$17426 ( \17803 , \17768 , \17801 );
or \U$17427 ( \17804 , \17785 , \17802 , \17803 );
and \U$17428 ( \17805 , \17752 , \17804 );
xor \U$17429 ( \17806 , \17544 , \17548 );
xor \U$17430 ( \17807 , \17806 , \17551 );
xor \U$17431 ( \17808 , \17587 , \17591 );
xor \U$17432 ( \17809 , \17808 , \17596 );
and \U$17433 ( \17810 , \17807 , \17809 );
xor \U$17434 ( \17811 , \17604 , \17608 );
xor \U$17435 ( \17812 , \17811 , \17613 );
and \U$17436 ( \17813 , \17809 , \17812 );
and \U$17437 ( \17814 , \17807 , \17812 );
or \U$17438 ( \17815 , \17810 , \17813 , \17814 );
and \U$17439 ( \17816 , \17804 , \17815 );
and \U$17440 ( \17817 , \17752 , \17815 );
or \U$17441 ( \17818 , \17805 , \17816 , \17817 );
xor \U$17442 ( \17819 , \17504 , \17520 );
xor \U$17443 ( \17820 , \17819 , \17537 );
xor \U$17444 ( \17821 , \17554 , \17558 );
xor \U$17445 ( \17822 , \17821 , \17563 );
and \U$17446 ( \17823 , \17820 , \17822 );
xor \U$17447 ( \17824 , \17583 , \17599 );
xor \U$17448 ( \17825 , \17824 , \17616 );
and \U$17449 ( \17826 , \17822 , \17825 );
and \U$17450 ( \17827 , \17820 , \17825 );
or \U$17451 ( \17828 , \17823 , \17826 , \17827 );
and \U$17452 ( \17829 , \17818 , \17828 );
xor \U$17453 ( \17830 , \17571 , \17575 );
xor \U$17454 ( \17831 , \17830 , \17580 );
xor \U$17455 ( \17832 , \17508 , \17512 );
xor \U$17456 ( \17833 , \17832 , \17517 );
and \U$17457 ( \17834 , \17831 , \17833 );
xor \U$17458 ( \17835 , \17525 , \17529 );
xor \U$17459 ( \17836 , \17835 , \17534 );
and \U$17460 ( \17837 , \17833 , \17836 );
and \U$17461 ( \17838 , \17831 , \17836 );
or \U$17462 ( \17839 , \17834 , \17837 , \17838 );
xor \U$17463 ( \17840 , \17624 , \17626 );
xor \U$17464 ( \17841 , \17840 , \17629 );
and \U$17465 ( \17842 , \17839 , \17841 );
xor \U$17466 ( \17843 , \17634 , \17636 );
xor \U$17467 ( \17844 , \17843 , \17639 );
and \U$17468 ( \17845 , \17841 , \17844 );
and \U$17469 ( \17846 , \17839 , \17844 );
or \U$17470 ( \17847 , \17842 , \17845 , \17846 );
and \U$17471 ( \17848 , \17828 , \17847 );
and \U$17472 ( \17849 , \17818 , \17847 );
or \U$17473 ( \17850 , \17829 , \17848 , \17849 );
xor \U$17474 ( \17851 , \17312 , \17328 );
xor \U$17475 ( \17852 , \17851 , \17345 );
xor \U$17476 ( \17853 , \17364 , \17380 );
xor \U$17477 ( \17854 , \17853 , \17397 );
and \U$17478 ( \17855 , \17852 , \17854 );
xor \U$17479 ( \17856 , \17651 , \17653 );
xor \U$17480 ( \17857 , \17856 , \17656 );
and \U$17481 ( \17858 , \17854 , \17857 );
and \U$17482 ( \17859 , \17852 , \17857 );
or \U$17483 ( \17860 , \17855 , \17858 , \17859 );
and \U$17484 ( \17861 , \17850 , \17860 );
xor \U$17485 ( \17862 , \17664 , \17666 );
xor \U$17486 ( \17863 , \17862 , \17669 );
and \U$17487 ( \17864 , \17860 , \17863 );
and \U$17488 ( \17865 , \17850 , \17863 );
or \U$17489 ( \17866 , \17861 , \17864 , \17865 );
xor \U$17490 ( \17867 , \17662 , \17672 );
xor \U$17491 ( \17868 , \17867 , \17675 );
and \U$17492 ( \17869 , \17866 , \17868 );
xor \U$17493 ( \17870 , \17680 , \17682 );
and \U$17494 ( \17871 , \17868 , \17870 );
and \U$17495 ( \17872 , \17866 , \17870 );
or \U$17496 ( \17873 , \17869 , \17871 , \17872 );
xor \U$17497 ( \17874 , \17445 , \17455 );
xor \U$17498 ( \17875 , \17874 , \17458 );
and \U$17499 ( \17876 , \17873 , \17875 );
xor \U$17500 ( \17877 , \17678 , \17683 );
xor \U$17501 ( \17878 , \17877 , \17686 );
and \U$17502 ( \17879 , \17875 , \17878 );
and \U$17503 ( \17880 , \17873 , \17878 );
or \U$17504 ( \17881 , \17876 , \17879 , \17880 );
and \U$17505 ( \17882 , \17700 , \17881 );
xor \U$17506 ( \17883 , \17700 , \17881 );
xor \U$17507 ( \17884 , \17873 , \17875 );
xor \U$17508 ( \17885 , \17884 , \17878 );
and \U$17509 ( \17886 , \4334 , \7829 );
and \U$17510 ( \17887 , \4078 , \7827 );
nor \U$17511 ( \17888 , \17886 , \17887 );
xnor \U$17512 ( \17889 , \17888 , \7580 );
and \U$17513 ( \17890 , \4833 , \7300 );
and \U$17514 ( \17891 , \4531 , \7298 );
nor \U$17515 ( \17892 , \17890 , \17891 );
xnor \U$17516 ( \17893 , \17892 , \7040 );
and \U$17517 ( \17894 , \17889 , \17893 );
and \U$17518 ( \17895 , \5310 , \6806 );
and \U$17519 ( \17896 , \4841 , \6804 );
nor \U$17520 ( \17897 , \17895 , \17896 );
xnor \U$17521 ( \17898 , \17897 , \6491 );
and \U$17522 ( \17899 , \17893 , \17898 );
and \U$17523 ( \17900 , \17889 , \17898 );
or \U$17524 ( \17901 , \17894 , \17899 , \17900 );
and \U$17525 ( \17902 , \3207 , \9495 );
and \U$17526 ( \17903 , \3069 , \9493 );
nor \U$17527 ( \17904 , \17902 , \17903 );
xnor \U$17528 ( \17905 , \17904 , \9185 );
and \U$17529 ( \17906 , \3743 , \8958 );
and \U$17530 ( \17907 , \3326 , \8956 );
nor \U$17531 ( \17908 , \17906 , \17907 );
xnor \U$17532 ( \17909 , \17908 , \8587 );
and \U$17533 ( \17910 , \17905 , \17909 );
and \U$17534 ( \17911 , \4073 , \8396 );
and \U$17535 ( \17912 , \3951 , \8394 );
nor \U$17536 ( \17913 , \17911 , \17912 );
xnor \U$17537 ( \17914 , \17913 , \8078 );
and \U$17538 ( \17915 , \17909 , \17914 );
and \U$17539 ( \17916 , \17905 , \17914 );
or \U$17540 ( \17917 , \17910 , \17915 , \17916 );
and \U$17541 ( \17918 , \17901 , \17917 );
and \U$17542 ( \17919 , \2703 , \10876 );
and \U$17543 ( \17920 , \2439 , \10873 );
nor \U$17544 ( \17921 , \17919 , \17920 );
xnor \U$17545 ( \17922 , \17921 , \9821 );
and \U$17546 ( \17923 , \2902 , \10063 );
and \U$17547 ( \17924 , \2728 , \10061 );
nor \U$17548 ( \17925 , \17923 , \17924 );
xnor \U$17549 ( \17926 , \17925 , \9824 );
and \U$17550 ( \17927 , \17922 , \17926 );
and \U$17551 ( \17928 , \17926 , \2225 );
and \U$17552 ( \17929 , \17922 , \2225 );
or \U$17553 ( \17930 , \17927 , \17928 , \17929 );
and \U$17554 ( \17931 , \17917 , \17930 );
and \U$17555 ( \17932 , \17901 , \17930 );
or \U$17556 ( \17933 , \17918 , \17931 , \17932 );
and \U$17557 ( \17934 , \8759 , \3699 );
and \U$17558 ( \17935 , \8440 , \3697 );
nor \U$17559 ( \17936 , \17934 , \17935 );
xnor \U$17560 ( \17937 , \17936 , \3512 );
and \U$17561 ( \17938 , \9612 , \3386 );
and \U$17562 ( \17939 , \9043 , \3384 );
nor \U$17563 ( \17940 , \17938 , \17939 );
xnor \U$17564 ( \17941 , \17940 , \3181 );
and \U$17565 ( \17942 , \17937 , \17941 );
and \U$17566 ( \17943 , \10223 , \2980 );
and \U$17567 ( \17944 , \9620 , \2978 );
nor \U$17568 ( \17945 , \17943 , \17944 );
xnor \U$17569 ( \17946 , \17945 , \2831 );
and \U$17570 ( \17947 , \17941 , \17946 );
and \U$17571 ( \17948 , \17937 , \17946 );
or \U$17572 ( \17949 , \17942 , \17947 , \17948 );
and \U$17573 ( \17950 , \5579 , \6297 );
and \U$17574 ( \17951 , \5315 , \6295 );
nor \U$17575 ( \17952 , \17950 , \17951 );
xnor \U$17576 ( \17953 , \17952 , \5957 );
and \U$17577 ( \17954 , \6210 , \5708 );
and \U$17578 ( \17955 , \5838 , \5706 );
nor \U$17579 ( \17956 , \17954 , \17955 );
xnor \U$17580 ( \17957 , \17956 , \5467 );
and \U$17581 ( \17958 , \17953 , \17957 );
and \U$17582 ( \17959 , \6562 , \5242 );
and \U$17583 ( \17960 , \6219 , \5240 );
nor \U$17584 ( \17961 , \17959 , \17960 );
xnor \U$17585 ( \17962 , \17961 , \5054 );
and \U$17586 ( \17963 , \17957 , \17962 );
and \U$17587 ( \17964 , \17953 , \17962 );
or \U$17588 ( \17965 , \17958 , \17963 , \17964 );
and \U$17589 ( \17966 , \17949 , \17965 );
and \U$17590 ( \17967 , \7067 , \4868 );
and \U$17591 ( \17968 , \6764 , \4866 );
nor \U$17592 ( \17969 , \17967 , \17968 );
xnor \U$17593 ( \17970 , \17969 , \4636 );
and \U$17594 ( \17971 , \7765 , \4417 );
and \U$17595 ( \17972 , \7239 , \4415 );
nor \U$17596 ( \17973 , \17971 , \17972 );
xnor \U$17597 ( \17974 , \17973 , \4274 );
and \U$17598 ( \17975 , \17970 , \17974 );
and \U$17599 ( \17976 , \8435 , \4094 );
and \U$17600 ( \17977 , \8189 , \4092 );
nor \U$17601 ( \17978 , \17976 , \17977 );
xnor \U$17602 ( \17979 , \17978 , \3848 );
and \U$17603 ( \17980 , \17974 , \17979 );
and \U$17604 ( \17981 , \17970 , \17979 );
or \U$17605 ( \17982 , \17975 , \17980 , \17981 );
and \U$17606 ( \17983 , \17965 , \17982 );
and \U$17607 ( \17984 , \17949 , \17982 );
or \U$17608 ( \17985 , \17966 , \17983 , \17984 );
and \U$17609 ( \17986 , \17933 , \17985 );
and \U$17610 ( \17987 , \11029 , \2362 );
and \U$17611 ( \17988 , \10409 , \2360 );
nor \U$17612 ( \17989 , \17987 , \17988 );
xnor \U$17613 ( \17990 , \17989 , \2225 );
xor \U$17614 ( \17991 , \17704 , \17708 );
xor \U$17615 ( \17992 , \17991 , \17713 );
and \U$17616 ( \17993 , \17990 , \17992 );
xor \U$17617 ( \17994 , \17737 , \17741 );
xor \U$17618 ( \17995 , \17994 , \17746 );
and \U$17619 ( \17996 , \17992 , \17995 );
and \U$17620 ( \17997 , \17990 , \17995 );
or \U$17621 ( \17998 , \17993 , \17996 , \17997 );
and \U$17622 ( \17999 , \17985 , \17998 );
and \U$17623 ( \18000 , \17933 , \17998 );
or \U$17624 ( \18001 , \17986 , \17999 , \18000 );
xor \U$17625 ( \18002 , \17756 , \17760 );
xor \U$17626 ( \18003 , \18002 , \17765 );
xor \U$17627 ( \18004 , \17720 , \17724 );
xor \U$17628 ( \18005 , \18004 , \17729 );
and \U$17629 ( \18006 , \18003 , \18005 );
xor \U$17630 ( \18007 , \17772 , \17776 );
xor \U$17631 ( \18008 , \18007 , \17781 );
and \U$17632 ( \18009 , \18005 , \18008 );
and \U$17633 ( \18010 , \18003 , \18008 );
or \U$17634 ( \18011 , \18006 , \18009 , \18010 );
xor \U$17635 ( \18012 , \17496 , \17500 );
xor \U$17636 ( \18013 , \18012 , \2004 );
and \U$17637 ( \18014 , \18011 , \18013 );
xor \U$17638 ( \18015 , \17831 , \17833 );
xor \U$17639 ( \18016 , \18015 , \17836 );
and \U$17640 ( \18017 , \18013 , \18016 );
and \U$17641 ( \18018 , \18011 , \18016 );
or \U$17642 ( \18019 , \18014 , \18017 , \18018 );
and \U$17643 ( \18020 , \18001 , \18019 );
xor \U$17644 ( \18021 , \17716 , \17732 );
xor \U$17645 ( \18022 , \18021 , \17749 );
xor \U$17646 ( \18023 , \17768 , \17784 );
xor \U$17647 ( \18024 , \18023 , \17801 );
and \U$17648 ( \18025 , \18022 , \18024 );
xor \U$17649 ( \18026 , \17807 , \17809 );
xor \U$17650 ( \18027 , \18026 , \17812 );
and \U$17651 ( \18028 , \18024 , \18027 );
and \U$17652 ( \18029 , \18022 , \18027 );
or \U$17653 ( \18030 , \18025 , \18028 , \18029 );
and \U$17654 ( \18031 , \18019 , \18030 );
and \U$17655 ( \18032 , \18001 , \18030 );
or \U$17656 ( \18033 , \18020 , \18031 , \18032 );
xor \U$17657 ( \18034 , \17752 , \17804 );
xor \U$17658 ( \18035 , \18034 , \17815 );
xor \U$17659 ( \18036 , \17820 , \17822 );
xor \U$17660 ( \18037 , \18036 , \17825 );
and \U$17661 ( \18038 , \18035 , \18037 );
xor \U$17662 ( \18039 , \17839 , \17841 );
xor \U$17663 ( \18040 , \18039 , \17844 );
and \U$17664 ( \18041 , \18037 , \18040 );
and \U$17665 ( \18042 , \18035 , \18040 );
or \U$17666 ( \18043 , \18038 , \18041 , \18042 );
and \U$17667 ( \18044 , \18033 , \18043 );
xor \U$17668 ( \18045 , \17632 , \17642 );
xor \U$17669 ( \18046 , \18045 , \17645 );
and \U$17670 ( \18047 , \18043 , \18046 );
and \U$17671 ( \18048 , \18033 , \18046 );
or \U$17672 ( \18049 , \18044 , \18047 , \18048 );
xor \U$17673 ( \18050 , \17540 , \17566 );
xor \U$17674 ( \18051 , \18050 , \17619 );
xor \U$17675 ( \18052 , \17818 , \17828 );
xor \U$17676 ( \18053 , \18052 , \17847 );
and \U$17677 ( \18054 , \18051 , \18053 );
xor \U$17678 ( \18055 , \17852 , \17854 );
xor \U$17679 ( \18056 , \18055 , \17857 );
and \U$17680 ( \18057 , \18053 , \18056 );
and \U$17681 ( \18058 , \18051 , \18056 );
or \U$17682 ( \18059 , \18054 , \18057 , \18058 );
and \U$17683 ( \18060 , \18049 , \18059 );
xor \U$17684 ( \18061 , \17622 , \17648 );
xor \U$17685 ( \18062 , \18061 , \17659 );
and \U$17686 ( \18063 , \18059 , \18062 );
and \U$17687 ( \18064 , \18049 , \18062 );
or \U$17688 ( \18065 , \18060 , \18063 , \18064 );
xor \U$17689 ( \18066 , \17866 , \17868 );
xor \U$17690 ( \18067 , \18066 , \17870 );
and \U$17691 ( \18068 , \18065 , \18067 );
and \U$17692 ( \18069 , \17885 , \18068 );
xor \U$17693 ( \18070 , \17885 , \18068 );
xor \U$17694 ( \18071 , \18065 , \18067 );
and \U$17695 ( \18072 , \2728 , \10876 );
and \U$17696 ( \18073 , \2703 , \10873 );
nor \U$17697 ( \18074 , \18072 , \18073 );
xnor \U$17698 ( \18075 , \18074 , \9821 );
and \U$17699 ( \18076 , \3069 , \10063 );
and \U$17700 ( \18077 , \2902 , \10061 );
nor \U$17701 ( \18078 , \18076 , \18077 );
xnor \U$17702 ( \18079 , \18078 , \9824 );
and \U$17703 ( \18080 , \18075 , \18079 );
and \U$17704 ( \18081 , \3326 , \9495 );
and \U$17705 ( \18082 , \3207 , \9493 );
nor \U$17706 ( \18083 , \18081 , \18082 );
xnor \U$17707 ( \18084 , \18083 , \9185 );
and \U$17708 ( \18085 , \18079 , \18084 );
and \U$17709 ( \18086 , \18075 , \18084 );
or \U$17710 ( \18087 , \18080 , \18085 , \18086 );
and \U$17711 ( \18088 , \3951 , \8958 );
and \U$17712 ( \18089 , \3743 , \8956 );
nor \U$17713 ( \18090 , \18088 , \18089 );
xnor \U$17714 ( \18091 , \18090 , \8587 );
and \U$17715 ( \18092 , \4078 , \8396 );
and \U$17716 ( \18093 , \4073 , \8394 );
nor \U$17717 ( \18094 , \18092 , \18093 );
xnor \U$17718 ( \18095 , \18094 , \8078 );
and \U$17719 ( \18096 , \18091 , \18095 );
and \U$17720 ( \18097 , \4531 , \7829 );
and \U$17721 ( \18098 , \4334 , \7827 );
nor \U$17722 ( \18099 , \18097 , \18098 );
xnor \U$17723 ( \18100 , \18099 , \7580 );
and \U$17724 ( \18101 , \18095 , \18100 );
and \U$17725 ( \18102 , \18091 , \18100 );
or \U$17726 ( \18103 , \18096 , \18101 , \18102 );
and \U$17727 ( \18104 , \18087 , \18103 );
and \U$17728 ( \18105 , \4841 , \7300 );
and \U$17729 ( \18106 , \4833 , \7298 );
nor \U$17730 ( \18107 , \18105 , \18106 );
xnor \U$17731 ( \18108 , \18107 , \7040 );
and \U$17732 ( \18109 , \5315 , \6806 );
and \U$17733 ( \18110 , \5310 , \6804 );
nor \U$17734 ( \18111 , \18109 , \18110 );
xnor \U$17735 ( \18112 , \18111 , \6491 );
and \U$17736 ( \18113 , \18108 , \18112 );
and \U$17737 ( \18114 , \5838 , \6297 );
and \U$17738 ( \18115 , \5579 , \6295 );
nor \U$17739 ( \18116 , \18114 , \18115 );
xnor \U$17740 ( \18117 , \18116 , \5957 );
and \U$17741 ( \18118 , \18112 , \18117 );
and \U$17742 ( \18119 , \18108 , \18117 );
or \U$17743 ( \18120 , \18113 , \18118 , \18119 );
and \U$17744 ( \18121 , \18103 , \18120 );
and \U$17745 ( \18122 , \18087 , \18120 );
or \U$17746 ( \18123 , \18104 , \18121 , \18122 );
and \U$17747 ( \18124 , \9620 , \3386 );
and \U$17748 ( \18125 , \9612 , \3384 );
nor \U$17749 ( \18126 , \18124 , \18125 );
xnor \U$17750 ( \18127 , \18126 , \3181 );
and \U$17751 ( \18128 , \10228 , \2980 );
and \U$17752 ( \18129 , \10223 , \2978 );
nor \U$17753 ( \18130 , \18128 , \18129 );
xnor \U$17754 ( \18131 , \18130 , \2831 );
and \U$17755 ( \18132 , \18127 , \18131 );
and \U$17756 ( \18133 , \11029 , \2658 );
and \U$17757 ( \18134 , \10409 , \2656 );
nor \U$17758 ( \18135 , \18133 , \18134 );
xnor \U$17759 ( \18136 , \18135 , \2516 );
and \U$17760 ( \18137 , \18131 , \18136 );
and \U$17761 ( \18138 , \18127 , \18136 );
or \U$17762 ( \18139 , \18132 , \18137 , \18138 );
and \U$17763 ( \18140 , \8189 , \4417 );
and \U$17764 ( \18141 , \7765 , \4415 );
nor \U$17765 ( \18142 , \18140 , \18141 );
xnor \U$17766 ( \18143 , \18142 , \4274 );
and \U$17767 ( \18144 , \8440 , \4094 );
and \U$17768 ( \18145 , \8435 , \4092 );
nor \U$17769 ( \18146 , \18144 , \18145 );
xnor \U$17770 ( \18147 , \18146 , \3848 );
and \U$17771 ( \18148 , \18143 , \18147 );
and \U$17772 ( \18149 , \9043 , \3699 );
and \U$17773 ( \18150 , \8759 , \3697 );
nor \U$17774 ( \18151 , \18149 , \18150 );
xnor \U$17775 ( \18152 , \18151 , \3512 );
and \U$17776 ( \18153 , \18147 , \18152 );
and \U$17777 ( \18154 , \18143 , \18152 );
or \U$17778 ( \18155 , \18148 , \18153 , \18154 );
and \U$17779 ( \18156 , \18139 , \18155 );
and \U$17780 ( \18157 , \6219 , \5708 );
and \U$17781 ( \18158 , \6210 , \5706 );
nor \U$17782 ( \18159 , \18157 , \18158 );
xnor \U$17783 ( \18160 , \18159 , \5467 );
and \U$17784 ( \18161 , \6764 , \5242 );
and \U$17785 ( \18162 , \6562 , \5240 );
nor \U$17786 ( \18163 , \18161 , \18162 );
xnor \U$17787 ( \18164 , \18163 , \5054 );
and \U$17788 ( \18165 , \18160 , \18164 );
and \U$17789 ( \18166 , \7239 , \4868 );
and \U$17790 ( \18167 , \7067 , \4866 );
nor \U$17791 ( \18168 , \18166 , \18167 );
xnor \U$17792 ( \18169 , \18168 , \4636 );
and \U$17793 ( \18170 , \18164 , \18169 );
and \U$17794 ( \18171 , \18160 , \18169 );
or \U$17795 ( \18172 , \18165 , \18170 , \18171 );
and \U$17796 ( \18173 , \18155 , \18172 );
and \U$17797 ( \18174 , \18139 , \18172 );
or \U$17798 ( \18175 , \18156 , \18173 , \18174 );
and \U$17799 ( \18176 , \18123 , \18175 );
and \U$17800 ( \18177 , \10409 , \2658 );
and \U$17801 ( \18178 , \10228 , \2656 );
nor \U$17802 ( \18179 , \18177 , \18178 );
xnor \U$17803 ( \18180 , \18179 , \2516 );
nand \U$17804 ( \18181 , \11029 , \2360 );
xnor \U$17805 ( \18182 , \18181 , \2225 );
and \U$17806 ( \18183 , \18180 , \18182 );
xor \U$17807 ( \18184 , \17937 , \17941 );
xor \U$17808 ( \18185 , \18184 , \17946 );
and \U$17809 ( \18186 , \18182 , \18185 );
and \U$17810 ( \18187 , \18180 , \18185 );
or \U$17811 ( \18188 , \18183 , \18186 , \18187 );
and \U$17812 ( \18189 , \18175 , \18188 );
and \U$17813 ( \18190 , \18123 , \18188 );
or \U$17814 ( \18191 , \18176 , \18189 , \18190 );
xor \U$17815 ( \18192 , \17889 , \17893 );
xor \U$17816 ( \18193 , \18192 , \17898 );
xor \U$17817 ( \18194 , \17953 , \17957 );
xor \U$17818 ( \18195 , \18194 , \17962 );
and \U$17819 ( \18196 , \18193 , \18195 );
xor \U$17820 ( \18197 , \17970 , \17974 );
xor \U$17821 ( \18198 , \18197 , \17979 );
and \U$17822 ( \18199 , \18195 , \18198 );
and \U$17823 ( \18200 , \18193 , \18198 );
or \U$17824 ( \18201 , \18196 , \18199 , \18200 );
xor \U$17825 ( \18202 , \17905 , \17909 );
xor \U$17826 ( \18203 , \18202 , \17914 );
xor \U$17827 ( \18204 , \17922 , \17926 );
xor \U$17828 ( \18205 , \18204 , \2225 );
and \U$17829 ( \18206 , \18203 , \18205 );
and \U$17830 ( \18207 , \18201 , \18206 );
xor \U$17831 ( \18208 , \17789 , \17793 );
xor \U$17832 ( \18209 , \18208 , \17798 );
and \U$17833 ( \18210 , \18206 , \18209 );
and \U$17834 ( \18211 , \18201 , \18209 );
or \U$17835 ( \18212 , \18207 , \18210 , \18211 );
and \U$17836 ( \18213 , \18191 , \18212 );
xor \U$17837 ( \18214 , \17949 , \17965 );
xor \U$17838 ( \18215 , \18214 , \17982 );
xor \U$17839 ( \18216 , \18003 , \18005 );
xor \U$17840 ( \18217 , \18216 , \18008 );
and \U$17841 ( \18218 , \18215 , \18217 );
xor \U$17842 ( \18219 , \17990 , \17992 );
xor \U$17843 ( \18220 , \18219 , \17995 );
and \U$17844 ( \18221 , \18217 , \18220 );
and \U$17845 ( \18222 , \18215 , \18220 );
or \U$17846 ( \18223 , \18218 , \18221 , \18222 );
and \U$17847 ( \18224 , \18212 , \18223 );
and \U$17848 ( \18225 , \18191 , \18223 );
or \U$17849 ( \18226 , \18213 , \18224 , \18225 );
xor \U$17850 ( \18227 , \17933 , \17985 );
xor \U$17851 ( \18228 , \18227 , \17998 );
xor \U$17852 ( \18229 , \18011 , \18013 );
xor \U$17853 ( \18230 , \18229 , \18016 );
and \U$17854 ( \18231 , \18228 , \18230 );
xor \U$17855 ( \18232 , \18022 , \18024 );
xor \U$17856 ( \18233 , \18232 , \18027 );
and \U$17857 ( \18234 , \18230 , \18233 );
and \U$17858 ( \18235 , \18228 , \18233 );
or \U$17859 ( \18236 , \18231 , \18234 , \18235 );
and \U$17860 ( \18237 , \18226 , \18236 );
xor \U$17861 ( \18238 , \18035 , \18037 );
xor \U$17862 ( \18239 , \18238 , \18040 );
and \U$17863 ( \18240 , \18236 , \18239 );
and \U$17864 ( \18241 , \18226 , \18239 );
or \U$17865 ( \18242 , \18237 , \18240 , \18241 );
xor \U$17866 ( \18243 , \18033 , \18043 );
xor \U$17867 ( \18244 , \18243 , \18046 );
and \U$17868 ( \18245 , \18242 , \18244 );
xor \U$17869 ( \18246 , \18051 , \18053 );
xor \U$17870 ( \18247 , \18246 , \18056 );
and \U$17871 ( \18248 , \18244 , \18247 );
and \U$17872 ( \18249 , \18242 , \18247 );
or \U$17873 ( \18250 , \18245 , \18248 , \18249 );
xor \U$17874 ( \18251 , \18049 , \18059 );
xor \U$17875 ( \18252 , \18251 , \18062 );
and \U$17876 ( \18253 , \18250 , \18252 );
xor \U$17877 ( \18254 , \17850 , \17860 );
xor \U$17878 ( \18255 , \18254 , \17863 );
and \U$17879 ( \18256 , \18252 , \18255 );
and \U$17880 ( \18257 , \18250 , \18255 );
or \U$17881 ( \18258 , \18253 , \18256 , \18257 );
and \U$17882 ( \18259 , \18071 , \18258 );
xor \U$17883 ( \18260 , \18071 , \18258 );
xor \U$17884 ( \18261 , \18250 , \18252 );
xor \U$17885 ( \18262 , \18261 , \18255 );
and \U$17886 ( \18263 , \2902 , \10876 );
and \U$17887 ( \18264 , \2728 , \10873 );
nor \U$17888 ( \18265 , \18263 , \18264 );
xnor \U$17889 ( \18266 , \18265 , \9821 );
and \U$17890 ( \18267 , \3207 , \10063 );
and \U$17891 ( \18268 , \3069 , \10061 );
nor \U$17892 ( \18269 , \18267 , \18268 );
xnor \U$17893 ( \18270 , \18269 , \9824 );
and \U$17894 ( \18271 , \18266 , \18270 );
and \U$17895 ( \18272 , \18270 , \2516 );
and \U$17896 ( \18273 , \18266 , \2516 );
or \U$17897 ( \18274 , \18271 , \18272 , \18273 );
and \U$17898 ( \18275 , \3743 , \9495 );
and \U$17899 ( \18276 , \3326 , \9493 );
nor \U$17900 ( \18277 , \18275 , \18276 );
xnor \U$17901 ( \18278 , \18277 , \9185 );
and \U$17902 ( \18279 , \4073 , \8958 );
and \U$17903 ( \18280 , \3951 , \8956 );
nor \U$17904 ( \18281 , \18279 , \18280 );
xnor \U$17905 ( \18282 , \18281 , \8587 );
and \U$17906 ( \18283 , \18278 , \18282 );
and \U$17907 ( \18284 , \4334 , \8396 );
and \U$17908 ( \18285 , \4078 , \8394 );
nor \U$17909 ( \18286 , \18284 , \18285 );
xnor \U$17910 ( \18287 , \18286 , \8078 );
and \U$17911 ( \18288 , \18282 , \18287 );
and \U$17912 ( \18289 , \18278 , \18287 );
or \U$17913 ( \18290 , \18283 , \18288 , \18289 );
and \U$17914 ( \18291 , \18274 , \18290 );
and \U$17915 ( \18292 , \4833 , \7829 );
and \U$17916 ( \18293 , \4531 , \7827 );
nor \U$17917 ( \18294 , \18292 , \18293 );
xnor \U$17918 ( \18295 , \18294 , \7580 );
and \U$17919 ( \18296 , \5310 , \7300 );
and \U$17920 ( \18297 , \4841 , \7298 );
nor \U$17921 ( \18298 , \18296 , \18297 );
xnor \U$17922 ( \18299 , \18298 , \7040 );
and \U$17923 ( \18300 , \18295 , \18299 );
and \U$17924 ( \18301 , \5579 , \6806 );
and \U$17925 ( \18302 , \5315 , \6804 );
nor \U$17926 ( \18303 , \18301 , \18302 );
xnor \U$17927 ( \18304 , \18303 , \6491 );
and \U$17928 ( \18305 , \18299 , \18304 );
and \U$17929 ( \18306 , \18295 , \18304 );
or \U$17930 ( \18307 , \18300 , \18305 , \18306 );
and \U$17931 ( \18308 , \18290 , \18307 );
and \U$17932 ( \18309 , \18274 , \18307 );
or \U$17933 ( \18310 , \18291 , \18308 , \18309 );
and \U$17934 ( \18311 , \6210 , \6297 );
and \U$17935 ( \18312 , \5838 , \6295 );
nor \U$17936 ( \18313 , \18311 , \18312 );
xnor \U$17937 ( \18314 , \18313 , \5957 );
and \U$17938 ( \18315 , \6562 , \5708 );
and \U$17939 ( \18316 , \6219 , \5706 );
nor \U$17940 ( \18317 , \18315 , \18316 );
xnor \U$17941 ( \18318 , \18317 , \5467 );
and \U$17942 ( \18319 , \18314 , \18318 );
and \U$17943 ( \18320 , \7067 , \5242 );
and \U$17944 ( \18321 , \6764 , \5240 );
nor \U$17945 ( \18322 , \18320 , \18321 );
xnor \U$17946 ( \18323 , \18322 , \5054 );
and \U$17947 ( \18324 , \18318 , \18323 );
and \U$17948 ( \18325 , \18314 , \18323 );
or \U$17949 ( \18326 , \18319 , \18324 , \18325 );
and \U$17950 ( \18327 , \7765 , \4868 );
and \U$17951 ( \18328 , \7239 , \4866 );
nor \U$17952 ( \18329 , \18327 , \18328 );
xnor \U$17953 ( \18330 , \18329 , \4636 );
and \U$17954 ( \18331 , \8435 , \4417 );
and \U$17955 ( \18332 , \8189 , \4415 );
nor \U$17956 ( \18333 , \18331 , \18332 );
xnor \U$17957 ( \18334 , \18333 , \4274 );
and \U$17958 ( \18335 , \18330 , \18334 );
and \U$17959 ( \18336 , \8759 , \4094 );
and \U$17960 ( \18337 , \8440 , \4092 );
nor \U$17961 ( \18338 , \18336 , \18337 );
xnor \U$17962 ( \18339 , \18338 , \3848 );
and \U$17963 ( \18340 , \18334 , \18339 );
and \U$17964 ( \18341 , \18330 , \18339 );
or \U$17965 ( \18342 , \18335 , \18340 , \18341 );
and \U$17966 ( \18343 , \18326 , \18342 );
and \U$17967 ( \18344 , \9612 , \3699 );
and \U$17968 ( \18345 , \9043 , \3697 );
nor \U$17969 ( \18346 , \18344 , \18345 );
xnor \U$17970 ( \18347 , \18346 , \3512 );
and \U$17971 ( \18348 , \10223 , \3386 );
and \U$17972 ( \18349 , \9620 , \3384 );
nor \U$17973 ( \18350 , \18348 , \18349 );
xnor \U$17974 ( \18351 , \18350 , \3181 );
and \U$17975 ( \18352 , \18347 , \18351 );
and \U$17976 ( \18353 , \10409 , \2980 );
and \U$17977 ( \18354 , \10228 , \2978 );
nor \U$17978 ( \18355 , \18353 , \18354 );
xnor \U$17979 ( \18356 , \18355 , \2831 );
and \U$17980 ( \18357 , \18351 , \18356 );
and \U$17981 ( \18358 , \18347 , \18356 );
or \U$17982 ( \18359 , \18352 , \18357 , \18358 );
and \U$17983 ( \18360 , \18342 , \18359 );
and \U$17984 ( \18361 , \18326 , \18359 );
or \U$17985 ( \18362 , \18343 , \18360 , \18361 );
and \U$17986 ( \18363 , \18310 , \18362 );
xor \U$17987 ( \18364 , \18127 , \18131 );
xor \U$17988 ( \18365 , \18364 , \18136 );
xor \U$17989 ( \18366 , \18143 , \18147 );
xor \U$17990 ( \18367 , \18366 , \18152 );
and \U$17991 ( \18368 , \18365 , \18367 );
xor \U$17992 ( \18369 , \18160 , \18164 );
xor \U$17993 ( \18370 , \18369 , \18169 );
and \U$17994 ( \18371 , \18367 , \18370 );
and \U$17995 ( \18372 , \18365 , \18370 );
or \U$17996 ( \18373 , \18368 , \18371 , \18372 );
and \U$17997 ( \18374 , \18362 , \18373 );
and \U$17998 ( \18375 , \18310 , \18373 );
or \U$17999 ( \18376 , \18363 , \18374 , \18375 );
xor \U$18000 ( \18377 , \18087 , \18103 );
xor \U$18001 ( \18378 , \18377 , \18120 );
xor \U$18002 ( \18379 , \18139 , \18155 );
xor \U$18003 ( \18380 , \18379 , \18172 );
and \U$18004 ( \18381 , \18378 , \18380 );
xor \U$18005 ( \18382 , \18180 , \18182 );
xor \U$18006 ( \18383 , \18382 , \18185 );
and \U$18007 ( \18384 , \18380 , \18383 );
and \U$18008 ( \18385 , \18378 , \18383 );
or \U$18009 ( \18386 , \18381 , \18384 , \18385 );
and \U$18010 ( \18387 , \18376 , \18386 );
xor \U$18011 ( \18388 , \18075 , \18079 );
xor \U$18012 ( \18389 , \18388 , \18084 );
xor \U$18013 ( \18390 , \18091 , \18095 );
xor \U$18014 ( \18391 , \18390 , \18100 );
and \U$18015 ( \18392 , \18389 , \18391 );
xor \U$18016 ( \18393 , \18108 , \18112 );
xor \U$18017 ( \18394 , \18393 , \18117 );
and \U$18018 ( \18395 , \18391 , \18394 );
and \U$18019 ( \18396 , \18389 , \18394 );
or \U$18020 ( \18397 , \18392 , \18395 , \18396 );
xor \U$18021 ( \18398 , \18193 , \18195 );
xor \U$18022 ( \18399 , \18398 , \18198 );
and \U$18023 ( \18400 , \18397 , \18399 );
xor \U$18024 ( \18401 , \18203 , \18205 );
and \U$18025 ( \18402 , \18399 , \18401 );
and \U$18026 ( \18403 , \18397 , \18401 );
or \U$18027 ( \18404 , \18400 , \18402 , \18403 );
and \U$18028 ( \18405 , \18386 , \18404 );
and \U$18029 ( \18406 , \18376 , \18404 );
or \U$18030 ( \18407 , \18387 , \18405 , \18406 );
xor \U$18031 ( \18408 , \17901 , \17917 );
xor \U$18032 ( \18409 , \18408 , \17930 );
xor \U$18033 ( \18410 , \18201 , \18206 );
xor \U$18034 ( \18411 , \18410 , \18209 );
and \U$18035 ( \18412 , \18409 , \18411 );
xor \U$18036 ( \18413 , \18215 , \18217 );
xor \U$18037 ( \18414 , \18413 , \18220 );
and \U$18038 ( \18415 , \18411 , \18414 );
and \U$18039 ( \18416 , \18409 , \18414 );
or \U$18040 ( \18417 , \18412 , \18415 , \18416 );
and \U$18041 ( \18418 , \18407 , \18417 );
xor \U$18042 ( \18419 , \18228 , \18230 );
xor \U$18043 ( \18420 , \18419 , \18233 );
and \U$18044 ( \18421 , \18417 , \18420 );
and \U$18045 ( \18422 , \18407 , \18420 );
or \U$18046 ( \18423 , \18418 , \18421 , \18422 );
xor \U$18047 ( \18424 , \18001 , \18019 );
xor \U$18048 ( \18425 , \18424 , \18030 );
and \U$18049 ( \18426 , \18423 , \18425 );
xor \U$18050 ( \18427 , \18226 , \18236 );
xor \U$18051 ( \18428 , \18427 , \18239 );
and \U$18052 ( \18429 , \18425 , \18428 );
and \U$18053 ( \18430 , \18423 , \18428 );
or \U$18054 ( \18431 , \18426 , \18429 , \18430 );
xor \U$18055 ( \18432 , \18242 , \18244 );
xor \U$18056 ( \18433 , \18432 , \18247 );
and \U$18057 ( \18434 , \18431 , \18433 );
and \U$18058 ( \18435 , \18262 , \18434 );
xor \U$18059 ( \18436 , \18262 , \18434 );
xor \U$18060 ( \18437 , \18431 , \18433 );
and \U$18061 ( \18438 , \5315 , \7300 );
and \U$18062 ( \18439 , \5310 , \7298 );
nor \U$18063 ( \18440 , \18438 , \18439 );
xnor \U$18064 ( \18441 , \18440 , \7040 );
and \U$18065 ( \18442 , \5838 , \6806 );
and \U$18066 ( \18443 , \5579 , \6804 );
nor \U$18067 ( \18444 , \18442 , \18443 );
xnor \U$18068 ( \18445 , \18444 , \6491 );
and \U$18069 ( \18446 , \18441 , \18445 );
and \U$18070 ( \18447 , \6219 , \6297 );
and \U$18071 ( \18448 , \6210 , \6295 );
nor \U$18072 ( \18449 , \18447 , \18448 );
xnor \U$18073 ( \18450 , \18449 , \5957 );
and \U$18074 ( \18451 , \18445 , \18450 );
and \U$18075 ( \18452 , \18441 , \18450 );
or \U$18076 ( \18453 , \18446 , \18451 , \18452 );
and \U$18077 ( \18454 , \3069 , \10876 );
and \U$18078 ( \18455 , \2902 , \10873 );
nor \U$18079 ( \18456 , \18454 , \18455 );
xnor \U$18080 ( \18457 , \18456 , \9821 );
and \U$18081 ( \18458 , \3326 , \10063 );
and \U$18082 ( \18459 , \3207 , \10061 );
nor \U$18083 ( \18460 , \18458 , \18459 );
xnor \U$18084 ( \18461 , \18460 , \9824 );
and \U$18085 ( \18462 , \18457 , \18461 );
and \U$18086 ( \18463 , \3951 , \9495 );
and \U$18087 ( \18464 , \3743 , \9493 );
nor \U$18088 ( \18465 , \18463 , \18464 );
xnor \U$18089 ( \18466 , \18465 , \9185 );
and \U$18090 ( \18467 , \18461 , \18466 );
and \U$18091 ( \18468 , \18457 , \18466 );
or \U$18092 ( \18469 , \18462 , \18467 , \18468 );
and \U$18093 ( \18470 , \18453 , \18469 );
and \U$18094 ( \18471 , \4078 , \8958 );
and \U$18095 ( \18472 , \4073 , \8956 );
nor \U$18096 ( \18473 , \18471 , \18472 );
xnor \U$18097 ( \18474 , \18473 , \8587 );
and \U$18098 ( \18475 , \4531 , \8396 );
and \U$18099 ( \18476 , \4334 , \8394 );
nor \U$18100 ( \18477 , \18475 , \18476 );
xnor \U$18101 ( \18478 , \18477 , \8078 );
and \U$18102 ( \18479 , \18474 , \18478 );
and \U$18103 ( \18480 , \4841 , \7829 );
and \U$18104 ( \18481 , \4833 , \7827 );
nor \U$18105 ( \18482 , \18480 , \18481 );
xnor \U$18106 ( \18483 , \18482 , \7580 );
and \U$18107 ( \18484 , \18478 , \18483 );
and \U$18108 ( \18485 , \18474 , \18483 );
or \U$18109 ( \18486 , \18479 , \18484 , \18485 );
and \U$18110 ( \18487 , \18469 , \18486 );
and \U$18111 ( \18488 , \18453 , \18486 );
or \U$18112 ( \18489 , \18470 , \18487 , \18488 );
and \U$18113 ( \18490 , \8440 , \4417 );
and \U$18114 ( \18491 , \8435 , \4415 );
nor \U$18115 ( \18492 , \18490 , \18491 );
xnor \U$18116 ( \18493 , \18492 , \4274 );
and \U$18117 ( \18494 , \9043 , \4094 );
and \U$18118 ( \18495 , \8759 , \4092 );
nor \U$18119 ( \18496 , \18494 , \18495 );
xnor \U$18120 ( \18497 , \18496 , \3848 );
and \U$18121 ( \18498 , \18493 , \18497 );
and \U$18122 ( \18499 , \9620 , \3699 );
and \U$18123 ( \18500 , \9612 , \3697 );
nor \U$18124 ( \18501 , \18499 , \18500 );
xnor \U$18125 ( \18502 , \18501 , \3512 );
and \U$18126 ( \18503 , \18497 , \18502 );
and \U$18127 ( \18504 , \18493 , \18502 );
or \U$18128 ( \18505 , \18498 , \18503 , \18504 );
and \U$18129 ( \18506 , \6764 , \5708 );
and \U$18130 ( \18507 , \6562 , \5706 );
nor \U$18131 ( \18508 , \18506 , \18507 );
xnor \U$18132 ( \18509 , \18508 , \5467 );
and \U$18133 ( \18510 , \7239 , \5242 );
and \U$18134 ( \18511 , \7067 , \5240 );
nor \U$18135 ( \18512 , \18510 , \18511 );
xnor \U$18136 ( \18513 , \18512 , \5054 );
and \U$18137 ( \18514 , \18509 , \18513 );
and \U$18138 ( \18515 , \8189 , \4868 );
and \U$18139 ( \18516 , \7765 , \4866 );
nor \U$18140 ( \18517 , \18515 , \18516 );
xnor \U$18141 ( \18518 , \18517 , \4636 );
and \U$18142 ( \18519 , \18513 , \18518 );
and \U$18143 ( \18520 , \18509 , \18518 );
or \U$18144 ( \18521 , \18514 , \18519 , \18520 );
and \U$18145 ( \18522 , \18505 , \18521 );
and \U$18146 ( \18523 , \10228 , \3386 );
and \U$18147 ( \18524 , \10223 , \3384 );
nor \U$18148 ( \18525 , \18523 , \18524 );
xnor \U$18149 ( \18526 , \18525 , \3181 );
and \U$18150 ( \18527 , \11029 , \2980 );
and \U$18151 ( \18528 , \10409 , \2978 );
nor \U$18152 ( \18529 , \18527 , \18528 );
xnor \U$18153 ( \18530 , \18529 , \2831 );
and \U$18154 ( \18531 , \18526 , \18530 );
and \U$18155 ( \18532 , \18521 , \18531 );
and \U$18156 ( \18533 , \18505 , \18531 );
or \U$18157 ( \18534 , \18522 , \18532 , \18533 );
and \U$18158 ( \18535 , \18489 , \18534 );
nand \U$18159 ( \18536 , \11029 , \2656 );
xnor \U$18160 ( \18537 , \18536 , \2516 );
xor \U$18161 ( \18538 , \18330 , \18334 );
xor \U$18162 ( \18539 , \18538 , \18339 );
and \U$18163 ( \18540 , \18537 , \18539 );
xor \U$18164 ( \18541 , \18347 , \18351 );
xor \U$18165 ( \18542 , \18541 , \18356 );
and \U$18166 ( \18543 , \18539 , \18542 );
and \U$18167 ( \18544 , \18537 , \18542 );
or \U$18168 ( \18545 , \18540 , \18543 , \18544 );
and \U$18169 ( \18546 , \18534 , \18545 );
and \U$18170 ( \18547 , \18489 , \18545 );
or \U$18171 ( \18548 , \18535 , \18546 , \18547 );
xor \U$18172 ( \18549 , \18278 , \18282 );
xor \U$18173 ( \18550 , \18549 , \18287 );
xor \U$18174 ( \18551 , \18314 , \18318 );
xor \U$18175 ( \18552 , \18551 , \18323 );
and \U$18176 ( \18553 , \18550 , \18552 );
xor \U$18177 ( \18554 , \18295 , \18299 );
xor \U$18178 ( \18555 , \18554 , \18304 );
and \U$18179 ( \18556 , \18552 , \18555 );
and \U$18180 ( \18557 , \18550 , \18555 );
or \U$18181 ( \18558 , \18553 , \18556 , \18557 );
xor \U$18182 ( \18559 , \18365 , \18367 );
xor \U$18183 ( \18560 , \18559 , \18370 );
and \U$18184 ( \18561 , \18558 , \18560 );
xor \U$18185 ( \18562 , \18389 , \18391 );
xor \U$18186 ( \18563 , \18562 , \18394 );
and \U$18187 ( \18564 , \18560 , \18563 );
and \U$18188 ( \18565 , \18558 , \18563 );
or \U$18189 ( \18566 , \18561 , \18564 , \18565 );
and \U$18190 ( \18567 , \18548 , \18566 );
xor \U$18191 ( \18568 , \18274 , \18290 );
xor \U$18192 ( \18569 , \18568 , \18307 );
xor \U$18193 ( \18570 , \18326 , \18342 );
xor \U$18194 ( \18571 , \18570 , \18359 );
and \U$18195 ( \18572 , \18569 , \18571 );
and \U$18196 ( \18573 , \18566 , \18572 );
and \U$18197 ( \18574 , \18548 , \18572 );
or \U$18198 ( \18575 , \18567 , \18573 , \18574 );
xor \U$18199 ( \18576 , \18310 , \18362 );
xor \U$18200 ( \18577 , \18576 , \18373 );
xor \U$18201 ( \18578 , \18378 , \18380 );
xor \U$18202 ( \18579 , \18578 , \18383 );
and \U$18203 ( \18580 , \18577 , \18579 );
xor \U$18204 ( \18581 , \18397 , \18399 );
xor \U$18205 ( \18582 , \18581 , \18401 );
and \U$18206 ( \18583 , \18579 , \18582 );
and \U$18207 ( \18584 , \18577 , \18582 );
or \U$18208 ( \18585 , \18580 , \18583 , \18584 );
and \U$18209 ( \18586 , \18575 , \18585 );
xor \U$18210 ( \18587 , \18123 , \18175 );
xor \U$18211 ( \18588 , \18587 , \18188 );
and \U$18212 ( \18589 , \18585 , \18588 );
and \U$18213 ( \18590 , \18575 , \18588 );
or \U$18214 ( \18591 , \18586 , \18589 , \18590 );
xor \U$18215 ( \18592 , \18376 , \18386 );
xor \U$18216 ( \18593 , \18592 , \18404 );
xor \U$18217 ( \18594 , \18409 , \18411 );
xor \U$18218 ( \18595 , \18594 , \18414 );
and \U$18219 ( \18596 , \18593 , \18595 );
and \U$18220 ( \18597 , \18591 , \18596 );
xor \U$18221 ( \18598 , \18191 , \18212 );
xor \U$18222 ( \18599 , \18598 , \18223 );
and \U$18223 ( \18600 , \18596 , \18599 );
and \U$18224 ( \18601 , \18591 , \18599 );
or \U$18225 ( \18602 , \18597 , \18600 , \18601 );
xor \U$18226 ( \18603 , \18423 , \18425 );
xor \U$18227 ( \18604 , \18603 , \18428 );
and \U$18228 ( \18605 , \18602 , \18604 );
and \U$18229 ( \18606 , \18437 , \18605 );
xor \U$18230 ( \18607 , \18437 , \18605 );
xor \U$18231 ( \18608 , \18602 , \18604 );
xor \U$18232 ( \18609 , \18591 , \18596 );
xor \U$18233 ( \18610 , \18609 , \18599 );
xor \U$18234 ( \18611 , \18407 , \18417 );
xor \U$18235 ( \18612 , \18611 , \18420 );
and \U$18236 ( \18613 , \18610 , \18612 );
and \U$18237 ( \18614 , \18608 , \18613 );
xor \U$18238 ( \18615 , \18608 , \18613 );
xor \U$18239 ( \18616 , \18610 , \18612 );
and \U$18240 ( \18617 , \8435 , \4868 );
and \U$18241 ( \18618 , \8189 , \4866 );
nor \U$18242 ( \18619 , \18617 , \18618 );
xnor \U$18243 ( \18620 , \18619 , \4636 );
and \U$18244 ( \18621 , \8759 , \4417 );
and \U$18245 ( \18622 , \8440 , \4415 );
nor \U$18246 ( \18623 , \18621 , \18622 );
xnor \U$18247 ( \18624 , \18623 , \4274 );
and \U$18248 ( \18625 , \18620 , \18624 );
and \U$18249 ( \18626 , \9612 , \4094 );
and \U$18250 ( \18627 , \9043 , \4092 );
nor \U$18251 ( \18628 , \18626 , \18627 );
xnor \U$18252 ( \18629 , \18628 , \3848 );
and \U$18253 ( \18630 , \18624 , \18629 );
and \U$18254 ( \18631 , \18620 , \18629 );
or \U$18255 ( \18632 , \18625 , \18630 , \18631 );
and \U$18256 ( \18633 , \10223 , \3699 );
and \U$18257 ( \18634 , \9620 , \3697 );
nor \U$18258 ( \18635 , \18633 , \18634 );
xnor \U$18259 ( \18636 , \18635 , \3512 );
and \U$18260 ( \18637 , \10409 , \3386 );
and \U$18261 ( \18638 , \10228 , \3384 );
nor \U$18262 ( \18639 , \18637 , \18638 );
xnor \U$18263 ( \18640 , \18639 , \3181 );
and \U$18264 ( \18641 , \18636 , \18640 );
nand \U$18265 ( \18642 , \11029 , \2978 );
xnor \U$18266 ( \18643 , \18642 , \2831 );
and \U$18267 ( \18644 , \18640 , \18643 );
and \U$18268 ( \18645 , \18636 , \18643 );
or \U$18269 ( \18646 , \18641 , \18644 , \18645 );
and \U$18270 ( \18647 , \18632 , \18646 );
and \U$18271 ( \18648 , \6562 , \6297 );
and \U$18272 ( \18649 , \6219 , \6295 );
nor \U$18273 ( \18650 , \18648 , \18649 );
xnor \U$18274 ( \18651 , \18650 , \5957 );
and \U$18275 ( \18652 , \7067 , \5708 );
and \U$18276 ( \18653 , \6764 , \5706 );
nor \U$18277 ( \18654 , \18652 , \18653 );
xnor \U$18278 ( \18655 , \18654 , \5467 );
and \U$18279 ( \18656 , \18651 , \18655 );
and \U$18280 ( \18657 , \7765 , \5242 );
and \U$18281 ( \18658 , \7239 , \5240 );
nor \U$18282 ( \18659 , \18657 , \18658 );
xnor \U$18283 ( \18660 , \18659 , \5054 );
and \U$18284 ( \18661 , \18655 , \18660 );
and \U$18285 ( \18662 , \18651 , \18660 );
or \U$18286 ( \18663 , \18656 , \18661 , \18662 );
and \U$18287 ( \18664 , \18646 , \18663 );
and \U$18288 ( \18665 , \18632 , \18663 );
or \U$18289 ( \18666 , \18647 , \18664 , \18665 );
and \U$18290 ( \18667 , \5310 , \7829 );
and \U$18291 ( \18668 , \4841 , \7827 );
nor \U$18292 ( \18669 , \18667 , \18668 );
xnor \U$18293 ( \18670 , \18669 , \7580 );
and \U$18294 ( \18671 , \5579 , \7300 );
and \U$18295 ( \18672 , \5315 , \7298 );
nor \U$18296 ( \18673 , \18671 , \18672 );
xnor \U$18297 ( \18674 , \18673 , \7040 );
and \U$18298 ( \18675 , \18670 , \18674 );
and \U$18299 ( \18676 , \6210 , \6806 );
and \U$18300 ( \18677 , \5838 , \6804 );
nor \U$18301 ( \18678 , \18676 , \18677 );
xnor \U$18302 ( \18679 , \18678 , \6491 );
and \U$18303 ( \18680 , \18674 , \18679 );
and \U$18304 ( \18681 , \18670 , \18679 );
or \U$18305 ( \18682 , \18675 , \18680 , \18681 );
and \U$18306 ( \18683 , \3207 , \10876 );
and \U$18307 ( \18684 , \3069 , \10873 );
nor \U$18308 ( \18685 , \18683 , \18684 );
xnor \U$18309 ( \18686 , \18685 , \9821 );
and \U$18310 ( \18687 , \3743 , \10063 );
and \U$18311 ( \18688 , \3326 , \10061 );
nor \U$18312 ( \18689 , \18687 , \18688 );
xnor \U$18313 ( \18690 , \18689 , \9824 );
and \U$18314 ( \18691 , \18686 , \18690 );
and \U$18315 ( \18692 , \18690 , \2831 );
and \U$18316 ( \18693 , \18686 , \2831 );
or \U$18317 ( \18694 , \18691 , \18692 , \18693 );
and \U$18318 ( \18695 , \18682 , \18694 );
and \U$18319 ( \18696 , \4073 , \9495 );
and \U$18320 ( \18697 , \3951 , \9493 );
nor \U$18321 ( \18698 , \18696 , \18697 );
xnor \U$18322 ( \18699 , \18698 , \9185 );
and \U$18323 ( \18700 , \4334 , \8958 );
and \U$18324 ( \18701 , \4078 , \8956 );
nor \U$18325 ( \18702 , \18700 , \18701 );
xnor \U$18326 ( \18703 , \18702 , \8587 );
and \U$18327 ( \18704 , \18699 , \18703 );
and \U$18328 ( \18705 , \4833 , \8396 );
and \U$18329 ( \18706 , \4531 , \8394 );
nor \U$18330 ( \18707 , \18705 , \18706 );
xnor \U$18331 ( \18708 , \18707 , \8078 );
and \U$18332 ( \18709 , \18703 , \18708 );
and \U$18333 ( \18710 , \18699 , \18708 );
or \U$18334 ( \18711 , \18704 , \18709 , \18710 );
and \U$18335 ( \18712 , \18694 , \18711 );
and \U$18336 ( \18713 , \18682 , \18711 );
or \U$18337 ( \18714 , \18695 , \18712 , \18713 );
and \U$18338 ( \18715 , \18666 , \18714 );
xor \U$18339 ( \18716 , \18493 , \18497 );
xor \U$18340 ( \18717 , \18716 , \18502 );
xor \U$18341 ( \18718 , \18509 , \18513 );
xor \U$18342 ( \18719 , \18718 , \18518 );
and \U$18343 ( \18720 , \18717 , \18719 );
xor \U$18344 ( \18721 , \18526 , \18530 );
and \U$18345 ( \18722 , \18719 , \18721 );
and \U$18346 ( \18723 , \18717 , \18721 );
or \U$18347 ( \18724 , \18720 , \18722 , \18723 );
and \U$18348 ( \18725 , \18714 , \18724 );
and \U$18349 ( \18726 , \18666 , \18724 );
or \U$18350 ( \18727 , \18715 , \18725 , \18726 );
xor \U$18351 ( \18728 , \18441 , \18445 );
xor \U$18352 ( \18729 , \18728 , \18450 );
xor \U$18353 ( \18730 , \18457 , \18461 );
xor \U$18354 ( \18731 , \18730 , \18466 );
and \U$18355 ( \18732 , \18729 , \18731 );
xor \U$18356 ( \18733 , \18474 , \18478 );
xor \U$18357 ( \18734 , \18733 , \18483 );
and \U$18358 ( \18735 , \18731 , \18734 );
and \U$18359 ( \18736 , \18729 , \18734 );
or \U$18360 ( \18737 , \18732 , \18735 , \18736 );
xor \U$18361 ( \18738 , \18266 , \18270 );
xor \U$18362 ( \18739 , \18738 , \2516 );
and \U$18363 ( \18740 , \18737 , \18739 );
xor \U$18364 ( \18741 , \18550 , \18552 );
xor \U$18365 ( \18742 , \18741 , \18555 );
and \U$18366 ( \18743 , \18739 , \18742 );
and \U$18367 ( \18744 , \18737 , \18742 );
or \U$18368 ( \18745 , \18740 , \18743 , \18744 );
and \U$18369 ( \18746 , \18727 , \18745 );
xor \U$18370 ( \18747 , \18453 , \18469 );
xor \U$18371 ( \18748 , \18747 , \18486 );
xor \U$18372 ( \18749 , \18505 , \18521 );
xor \U$18373 ( \18750 , \18749 , \18531 );
and \U$18374 ( \18751 , \18748 , \18750 );
xor \U$18375 ( \18752 , \18537 , \18539 );
xor \U$18376 ( \18753 , \18752 , \18542 );
and \U$18377 ( \18754 , \18750 , \18753 );
and \U$18378 ( \18755 , \18748 , \18753 );
or \U$18379 ( \18756 , \18751 , \18754 , \18755 );
and \U$18380 ( \18757 , \18745 , \18756 );
and \U$18381 ( \18758 , \18727 , \18756 );
or \U$18382 ( \18759 , \18746 , \18757 , \18758 );
xor \U$18383 ( \18760 , \18489 , \18534 );
xor \U$18384 ( \18761 , \18760 , \18545 );
xor \U$18385 ( \18762 , \18558 , \18560 );
xor \U$18386 ( \18763 , \18762 , \18563 );
and \U$18387 ( \18764 , \18761 , \18763 );
xor \U$18388 ( \18765 , \18569 , \18571 );
and \U$18389 ( \18766 , \18763 , \18765 );
and \U$18390 ( \18767 , \18761 , \18765 );
or \U$18391 ( \18768 , \18764 , \18766 , \18767 );
and \U$18392 ( \18769 , \18759 , \18768 );
xor \U$18393 ( \18770 , \18577 , \18579 );
xor \U$18394 ( \18771 , \18770 , \18582 );
and \U$18395 ( \18772 , \18768 , \18771 );
and \U$18396 ( \18773 , \18759 , \18771 );
or \U$18397 ( \18774 , \18769 , \18772 , \18773 );
xor \U$18398 ( \18775 , \18575 , \18585 );
xor \U$18399 ( \18776 , \18775 , \18588 );
and \U$18400 ( \18777 , \18774 , \18776 );
xor \U$18401 ( \18778 , \18593 , \18595 );
and \U$18402 ( \18779 , \18776 , \18778 );
and \U$18403 ( \18780 , \18774 , \18778 );
or \U$18404 ( \18781 , \18777 , \18779 , \18780 );
and \U$18405 ( \18782 , \18616 , \18781 );
xor \U$18406 ( \18783 , \18616 , \18781 );
xor \U$18407 ( \18784 , \18774 , \18776 );
xor \U$18408 ( \18785 , \18784 , \18778 );
and \U$18409 ( \18786 , \4531 , \8958 );
and \U$18410 ( \18787 , \4334 , \8956 );
nor \U$18411 ( \18788 , \18786 , \18787 );
xnor \U$18412 ( \18789 , \18788 , \8587 );
and \U$18413 ( \18790 , \4841 , \8396 );
and \U$18414 ( \18791 , \4833 , \8394 );
nor \U$18415 ( \18792 , \18790 , \18791 );
xnor \U$18416 ( \18793 , \18792 , \8078 );
and \U$18417 ( \18794 , \18789 , \18793 );
and \U$18418 ( \18795 , \5315 , \7829 );
and \U$18419 ( \18796 , \5310 , \7827 );
nor \U$18420 ( \18797 , \18795 , \18796 );
xnor \U$18421 ( \18798 , \18797 , \7580 );
and \U$18422 ( \18799 , \18793 , \18798 );
and \U$18423 ( \18800 , \18789 , \18798 );
or \U$18424 ( \18801 , \18794 , \18799 , \18800 );
and \U$18425 ( \18802 , \3326 , \10876 );
and \U$18426 ( \18803 , \3207 , \10873 );
nor \U$18427 ( \18804 , \18802 , \18803 );
xnor \U$18428 ( \18805 , \18804 , \9821 );
and \U$18429 ( \18806 , \3951 , \10063 );
and \U$18430 ( \18807 , \3743 , \10061 );
nor \U$18431 ( \18808 , \18806 , \18807 );
xnor \U$18432 ( \18809 , \18808 , \9824 );
and \U$18433 ( \18810 , \18805 , \18809 );
and \U$18434 ( \18811 , \4078 , \9495 );
and \U$18435 ( \18812 , \4073 , \9493 );
nor \U$18436 ( \18813 , \18811 , \18812 );
xnor \U$18437 ( \18814 , \18813 , \9185 );
and \U$18438 ( \18815 , \18809 , \18814 );
and \U$18439 ( \18816 , \18805 , \18814 );
or \U$18440 ( \18817 , \18810 , \18815 , \18816 );
and \U$18441 ( \18818 , \18801 , \18817 );
and \U$18442 ( \18819 , \5838 , \7300 );
and \U$18443 ( \18820 , \5579 , \7298 );
nor \U$18444 ( \18821 , \18819 , \18820 );
xnor \U$18445 ( \18822 , \18821 , \7040 );
and \U$18446 ( \18823 , \6219 , \6806 );
and \U$18447 ( \18824 , \6210 , \6804 );
nor \U$18448 ( \18825 , \18823 , \18824 );
xnor \U$18449 ( \18826 , \18825 , \6491 );
and \U$18450 ( \18827 , \18822 , \18826 );
and \U$18451 ( \18828 , \6764 , \6297 );
and \U$18452 ( \18829 , \6562 , \6295 );
nor \U$18453 ( \18830 , \18828 , \18829 );
xnor \U$18454 ( \18831 , \18830 , \5957 );
and \U$18455 ( \18832 , \18826 , \18831 );
and \U$18456 ( \18833 , \18822 , \18831 );
or \U$18457 ( \18834 , \18827 , \18832 , \18833 );
and \U$18458 ( \18835 , \18817 , \18834 );
and \U$18459 ( \18836 , \18801 , \18834 );
or \U$18460 ( \18837 , \18818 , \18835 , \18836 );
xor \U$18461 ( \18838 , \18620 , \18624 );
xor \U$18462 ( \18839 , \18838 , \18629 );
xor \U$18463 ( \18840 , \18670 , \18674 );
xor \U$18464 ( \18841 , \18840 , \18679 );
and \U$18465 ( \18842 , \18839 , \18841 );
xor \U$18466 ( \18843 , \18651 , \18655 );
xor \U$18467 ( \18844 , \18843 , \18660 );
and \U$18468 ( \18845 , \18841 , \18844 );
and \U$18469 ( \18846 , \18839 , \18844 );
or \U$18470 ( \18847 , \18842 , \18845 , \18846 );
and \U$18471 ( \18848 , \18837 , \18847 );
and \U$18472 ( \18849 , \7239 , \5708 );
and \U$18473 ( \18850 , \7067 , \5706 );
nor \U$18474 ( \18851 , \18849 , \18850 );
xnor \U$18475 ( \18852 , \18851 , \5467 );
and \U$18476 ( \18853 , \8189 , \5242 );
and \U$18477 ( \18854 , \7765 , \5240 );
nor \U$18478 ( \18855 , \18853 , \18854 );
xnor \U$18479 ( \18856 , \18855 , \5054 );
and \U$18480 ( \18857 , \18852 , \18856 );
and \U$18481 ( \18858 , \8440 , \4868 );
and \U$18482 ( \18859 , \8435 , \4866 );
nor \U$18483 ( \18860 , \18858 , \18859 );
xnor \U$18484 ( \18861 , \18860 , \4636 );
and \U$18485 ( \18862 , \18856 , \18861 );
and \U$18486 ( \18863 , \18852 , \18861 );
or \U$18487 ( \18864 , \18857 , \18862 , \18863 );
and \U$18488 ( \18865 , \9043 , \4417 );
and \U$18489 ( \18866 , \8759 , \4415 );
nor \U$18490 ( \18867 , \18865 , \18866 );
xnor \U$18491 ( \18868 , \18867 , \4274 );
and \U$18492 ( \18869 , \9620 , \4094 );
and \U$18493 ( \18870 , \9612 , \4092 );
nor \U$18494 ( \18871 , \18869 , \18870 );
xnor \U$18495 ( \18872 , \18871 , \3848 );
and \U$18496 ( \18873 , \18868 , \18872 );
and \U$18497 ( \18874 , \10228 , \3699 );
and \U$18498 ( \18875 , \10223 , \3697 );
nor \U$18499 ( \18876 , \18874 , \18875 );
xnor \U$18500 ( \18877 , \18876 , \3512 );
and \U$18501 ( \18878 , \18872 , \18877 );
and \U$18502 ( \18879 , \18868 , \18877 );
or \U$18503 ( \18880 , \18873 , \18878 , \18879 );
and \U$18504 ( \18881 , \18864 , \18880 );
xor \U$18505 ( \18882 , \18636 , \18640 );
xor \U$18506 ( \18883 , \18882 , \18643 );
and \U$18507 ( \18884 , \18880 , \18883 );
and \U$18508 ( \18885 , \18864 , \18883 );
or \U$18509 ( \18886 , \18881 , \18884 , \18885 );
and \U$18510 ( \18887 , \18847 , \18886 );
and \U$18511 ( \18888 , \18837 , \18886 );
or \U$18512 ( \18889 , \18848 , \18887 , \18888 );
xor \U$18513 ( \18890 , \18632 , \18646 );
xor \U$18514 ( \18891 , \18890 , \18663 );
xor \U$18515 ( \18892 , \18729 , \18731 );
xor \U$18516 ( \18893 , \18892 , \18734 );
and \U$18517 ( \18894 , \18891 , \18893 );
xor \U$18518 ( \18895 , \18717 , \18719 );
xor \U$18519 ( \18896 , \18895 , \18721 );
and \U$18520 ( \18897 , \18893 , \18896 );
and \U$18521 ( \18898 , \18891 , \18896 );
or \U$18522 ( \18899 , \18894 , \18897 , \18898 );
and \U$18523 ( \18900 , \18889 , \18899 );
xor \U$18524 ( \18901 , \18748 , \18750 );
xor \U$18525 ( \18902 , \18901 , \18753 );
and \U$18526 ( \18903 , \18899 , \18902 );
and \U$18527 ( \18904 , \18889 , \18902 );
or \U$18528 ( \18905 , \18900 , \18903 , \18904 );
xor \U$18529 ( \18906 , \18727 , \18745 );
xor \U$18530 ( \18907 , \18906 , \18756 );
and \U$18531 ( \18908 , \18905 , \18907 );
xor \U$18532 ( \18909 , \18761 , \18763 );
xor \U$18533 ( \18910 , \18909 , \18765 );
and \U$18534 ( \18911 , \18907 , \18910 );
and \U$18535 ( \18912 , \18905 , \18910 );
or \U$18536 ( \18913 , \18908 , \18911 , \18912 );
xor \U$18537 ( \18914 , \18548 , \18566 );
xor \U$18538 ( \18915 , \18914 , \18572 );
and \U$18539 ( \18916 , \18913 , \18915 );
xor \U$18540 ( \18917 , \18759 , \18768 );
xor \U$18541 ( \18918 , \18917 , \18771 );
and \U$18542 ( \18919 , \18915 , \18918 );
and \U$18543 ( \18920 , \18913 , \18918 );
or \U$18544 ( \18921 , \18916 , \18919 , \18920 );
and \U$18545 ( \18922 , \18785 , \18921 );
xor \U$18546 ( \18923 , \18785 , \18921 );
xor \U$18547 ( \18924 , \18913 , \18915 );
xor \U$18548 ( \18925 , \18924 , \18918 );
and \U$18549 ( \18926 , \4334 , \9495 );
and \U$18550 ( \18927 , \4078 , \9493 );
nor \U$18551 ( \18928 , \18926 , \18927 );
xnor \U$18552 ( \18929 , \18928 , \9185 );
and \U$18553 ( \18930 , \4833 , \8958 );
and \U$18554 ( \18931 , \4531 , \8956 );
nor \U$18555 ( \18932 , \18930 , \18931 );
xnor \U$18556 ( \18933 , \18932 , \8587 );
and \U$18557 ( \18934 , \18929 , \18933 );
and \U$18558 ( \18935 , \5310 , \8396 );
and \U$18559 ( \18936 , \4841 , \8394 );
nor \U$18560 ( \18937 , \18935 , \18936 );
xnor \U$18561 ( \18938 , \18937 , \8078 );
and \U$18562 ( \18939 , \18933 , \18938 );
and \U$18563 ( \18940 , \18929 , \18938 );
or \U$18564 ( \18941 , \18934 , \18939 , \18940 );
and \U$18565 ( \18942 , \5579 , \7829 );
and \U$18566 ( \18943 , \5315 , \7827 );
nor \U$18567 ( \18944 , \18942 , \18943 );
xnor \U$18568 ( \18945 , \18944 , \7580 );
and \U$18569 ( \18946 , \6210 , \7300 );
and \U$18570 ( \18947 , \5838 , \7298 );
nor \U$18571 ( \18948 , \18946 , \18947 );
xnor \U$18572 ( \18949 , \18948 , \7040 );
and \U$18573 ( \18950 , \18945 , \18949 );
and \U$18574 ( \18951 , \6562 , \6806 );
and \U$18575 ( \18952 , \6219 , \6804 );
nor \U$18576 ( \18953 , \18951 , \18952 );
xnor \U$18577 ( \18954 , \18953 , \6491 );
and \U$18578 ( \18955 , \18949 , \18954 );
and \U$18579 ( \18956 , \18945 , \18954 );
or \U$18580 ( \18957 , \18950 , \18955 , \18956 );
and \U$18581 ( \18958 , \18941 , \18957 );
and \U$18582 ( \18959 , \3743 , \10876 );
and \U$18583 ( \18960 , \3326 , \10873 );
nor \U$18584 ( \18961 , \18959 , \18960 );
xnor \U$18585 ( \18962 , \18961 , \9821 );
and \U$18586 ( \18963 , \4073 , \10063 );
and \U$18587 ( \18964 , \3951 , \10061 );
nor \U$18588 ( \18965 , \18963 , \18964 );
xnor \U$18589 ( \18966 , \18965 , \9824 );
and \U$18590 ( \18967 , \18962 , \18966 );
and \U$18591 ( \18968 , \18966 , \3181 );
and \U$18592 ( \18969 , \18962 , \3181 );
or \U$18593 ( \18970 , \18967 , \18968 , \18969 );
and \U$18594 ( \18971 , \18957 , \18970 );
and \U$18595 ( \18972 , \18941 , \18970 );
or \U$18596 ( \18973 , \18958 , \18971 , \18972 );
and \U$18597 ( \18974 , \8759 , \4868 );
and \U$18598 ( \18975 , \8440 , \4866 );
nor \U$18599 ( \18976 , \18974 , \18975 );
xnor \U$18600 ( \18977 , \18976 , \4636 );
and \U$18601 ( \18978 , \9612 , \4417 );
and \U$18602 ( \18979 , \9043 , \4415 );
nor \U$18603 ( \18980 , \18978 , \18979 );
xnor \U$18604 ( \18981 , \18980 , \4274 );
and \U$18605 ( \18982 , \18977 , \18981 );
and \U$18606 ( \18983 , \10223 , \4094 );
and \U$18607 ( \18984 , \9620 , \4092 );
nor \U$18608 ( \18985 , \18983 , \18984 );
xnor \U$18609 ( \18986 , \18985 , \3848 );
and \U$18610 ( \18987 , \18981 , \18986 );
and \U$18611 ( \18988 , \18977 , \18986 );
or \U$18612 ( \18989 , \18982 , \18987 , \18988 );
and \U$18613 ( \18990 , \7067 , \6297 );
and \U$18614 ( \18991 , \6764 , \6295 );
nor \U$18615 ( \18992 , \18990 , \18991 );
xnor \U$18616 ( \18993 , \18992 , \5957 );
and \U$18617 ( \18994 , \7765 , \5708 );
and \U$18618 ( \18995 , \7239 , \5706 );
nor \U$18619 ( \18996 , \18994 , \18995 );
xnor \U$18620 ( \18997 , \18996 , \5467 );
and \U$18621 ( \18998 , \18993 , \18997 );
and \U$18622 ( \18999 , \8435 , \5242 );
and \U$18623 ( \19000 , \8189 , \5240 );
nor \U$18624 ( \19001 , \18999 , \19000 );
xnor \U$18625 ( \19002 , \19001 , \5054 );
and \U$18626 ( \19003 , \18997 , \19002 );
and \U$18627 ( \19004 , \18993 , \19002 );
or \U$18628 ( \19005 , \18998 , \19003 , \19004 );
and \U$18629 ( \19006 , \18989 , \19005 );
and \U$18630 ( \19007 , \11029 , \3386 );
and \U$18631 ( \19008 , \10409 , \3384 );
nor \U$18632 ( \19009 , \19007 , \19008 );
xnor \U$18633 ( \19010 , \19009 , \3181 );
and \U$18634 ( \19011 , \19005 , \19010 );
and \U$18635 ( \19012 , \18989 , \19010 );
or \U$18636 ( \19013 , \19006 , \19011 , \19012 );
and \U$18637 ( \19014 , \18973 , \19013 );
xor \U$18638 ( \19015 , \18852 , \18856 );
xor \U$18639 ( \19016 , \19015 , \18861 );
xor \U$18640 ( \19017 , \18868 , \18872 );
xor \U$18641 ( \19018 , \19017 , \18877 );
and \U$18642 ( \19019 , \19016 , \19018 );
xor \U$18643 ( \19020 , \18822 , \18826 );
xor \U$18644 ( \19021 , \19020 , \18831 );
and \U$18645 ( \19022 , \19018 , \19021 );
and \U$18646 ( \19023 , \19016 , \19021 );
or \U$18647 ( \19024 , \19019 , \19022 , \19023 );
and \U$18648 ( \19025 , \19013 , \19024 );
and \U$18649 ( \19026 , \18973 , \19024 );
or \U$18650 ( \19027 , \19014 , \19025 , \19026 );
xor \U$18651 ( \19028 , \18686 , \18690 );
xor \U$18652 ( \19029 , \19028 , \2831 );
xor \U$18653 ( \19030 , \18699 , \18703 );
xor \U$18654 ( \19031 , \19030 , \18708 );
and \U$18655 ( \19032 , \19029 , \19031 );
xor \U$18656 ( \19033 , \18839 , \18841 );
xor \U$18657 ( \19034 , \19033 , \18844 );
and \U$18658 ( \19035 , \19031 , \19034 );
and \U$18659 ( \19036 , \19029 , \19034 );
or \U$18660 ( \19037 , \19032 , \19035 , \19036 );
and \U$18661 ( \19038 , \19027 , \19037 );
xor \U$18662 ( \19039 , \18801 , \18817 );
xor \U$18663 ( \19040 , \19039 , \18834 );
xor \U$18664 ( \19041 , \18864 , \18880 );
xor \U$18665 ( \19042 , \19041 , \18883 );
and \U$18666 ( \19043 , \19040 , \19042 );
and \U$18667 ( \19044 , \19037 , \19043 );
and \U$18668 ( \19045 , \19027 , \19043 );
or \U$18669 ( \19046 , \19038 , \19044 , \19045 );
xor \U$18670 ( \19047 , \18682 , \18694 );
xor \U$18671 ( \19048 , \19047 , \18711 );
xor \U$18672 ( \19049 , \18837 , \18847 );
xor \U$18673 ( \19050 , \19049 , \18886 );
and \U$18674 ( \19051 , \19048 , \19050 );
xor \U$18675 ( \19052 , \18891 , \18893 );
xor \U$18676 ( \19053 , \19052 , \18896 );
and \U$18677 ( \19054 , \19050 , \19053 );
and \U$18678 ( \19055 , \19048 , \19053 );
or \U$18679 ( \19056 , \19051 , \19054 , \19055 );
and \U$18680 ( \19057 , \19046 , \19056 );
xor \U$18681 ( \19058 , \18737 , \18739 );
xor \U$18682 ( \19059 , \19058 , \18742 );
and \U$18683 ( \19060 , \19056 , \19059 );
and \U$18684 ( \19061 , \19046 , \19059 );
or \U$18685 ( \19062 , \19057 , \19060 , \19061 );
xor \U$18686 ( \19063 , \18666 , \18714 );
xor \U$18687 ( \19064 , \19063 , \18724 );
xor \U$18688 ( \19065 , \18889 , \18899 );
xor \U$18689 ( \19066 , \19065 , \18902 );
and \U$18690 ( \19067 , \19064 , \19066 );
and \U$18691 ( \19068 , \19062 , \19067 );
xor \U$18692 ( \19069 , \18905 , \18907 );
xor \U$18693 ( \19070 , \19069 , \18910 );
and \U$18694 ( \19071 , \19067 , \19070 );
and \U$18695 ( \19072 , \19062 , \19070 );
or \U$18696 ( \19073 , \19068 , \19071 , \19072 );
and \U$18697 ( \19074 , \18925 , \19073 );
xor \U$18698 ( \19075 , \18925 , \19073 );
xor \U$18699 ( \19076 , \19062 , \19067 );
xor \U$18700 ( \19077 , \19076 , \19070 );
and \U$18701 ( \19078 , \6219 , \7300 );
and \U$18702 ( \19079 , \6210 , \7298 );
nor \U$18703 ( \19080 , \19078 , \19079 );
xnor \U$18704 ( \19081 , \19080 , \7040 );
and \U$18705 ( \19082 , \6764 , \6806 );
and \U$18706 ( \19083 , \6562 , \6804 );
nor \U$18707 ( \19084 , \19082 , \19083 );
xnor \U$18708 ( \19085 , \19084 , \6491 );
and \U$18709 ( \19086 , \19081 , \19085 );
and \U$18710 ( \19087 , \7239 , \6297 );
and \U$18711 ( \19088 , \7067 , \6295 );
nor \U$18712 ( \19089 , \19087 , \19088 );
xnor \U$18713 ( \19090 , \19089 , \5957 );
and \U$18714 ( \19091 , \19085 , \19090 );
and \U$18715 ( \19092 , \19081 , \19090 );
or \U$18716 ( \19093 , \19086 , \19091 , \19092 );
and \U$18717 ( \19094 , \4841 , \8958 );
and \U$18718 ( \19095 , \4833 , \8956 );
nor \U$18719 ( \19096 , \19094 , \19095 );
xnor \U$18720 ( \19097 , \19096 , \8587 );
and \U$18721 ( \19098 , \5315 , \8396 );
and \U$18722 ( \19099 , \5310 , \8394 );
nor \U$18723 ( \19100 , \19098 , \19099 );
xnor \U$18724 ( \19101 , \19100 , \8078 );
and \U$18725 ( \19102 , \19097 , \19101 );
and \U$18726 ( \19103 , \5838 , \7829 );
and \U$18727 ( \19104 , \5579 , \7827 );
nor \U$18728 ( \19105 , \19103 , \19104 );
xnor \U$18729 ( \19106 , \19105 , \7580 );
and \U$18730 ( \19107 , \19101 , \19106 );
and \U$18731 ( \19108 , \19097 , \19106 );
or \U$18732 ( \19109 , \19102 , \19107 , \19108 );
and \U$18733 ( \19110 , \19093 , \19109 );
and \U$18734 ( \19111 , \3951 , \10876 );
and \U$18735 ( \19112 , \3743 , \10873 );
nor \U$18736 ( \19113 , \19111 , \19112 );
xnor \U$18737 ( \19114 , \19113 , \9821 );
and \U$18738 ( \19115 , \4078 , \10063 );
and \U$18739 ( \19116 , \4073 , \10061 );
nor \U$18740 ( \19117 , \19115 , \19116 );
xnor \U$18741 ( \19118 , \19117 , \9824 );
and \U$18742 ( \19119 , \19114 , \19118 );
and \U$18743 ( \19120 , \4531 , \9495 );
and \U$18744 ( \19121 , \4334 , \9493 );
nor \U$18745 ( \19122 , \19120 , \19121 );
xnor \U$18746 ( \19123 , \19122 , \9185 );
and \U$18747 ( \19124 , \19118 , \19123 );
and \U$18748 ( \19125 , \19114 , \19123 );
or \U$18749 ( \19126 , \19119 , \19124 , \19125 );
and \U$18750 ( \19127 , \19109 , \19126 );
and \U$18751 ( \19128 , \19093 , \19126 );
or \U$18752 ( \19129 , \19110 , \19127 , \19128 );
and \U$18753 ( \19130 , \9620 , \4417 );
and \U$18754 ( \19131 , \9612 , \4415 );
nor \U$18755 ( \19132 , \19130 , \19131 );
xnor \U$18756 ( \19133 , \19132 , \4274 );
and \U$18757 ( \19134 , \10228 , \4094 );
and \U$18758 ( \19135 , \10223 , \4092 );
nor \U$18759 ( \19136 , \19134 , \19135 );
xnor \U$18760 ( \19137 , \19136 , \3848 );
and \U$18761 ( \19138 , \19133 , \19137 );
and \U$18762 ( \19139 , \11029 , \3699 );
and \U$18763 ( \19140 , \10409 , \3697 );
nor \U$18764 ( \19141 , \19139 , \19140 );
xnor \U$18765 ( \19142 , \19141 , \3512 );
and \U$18766 ( \19143 , \19137 , \19142 );
and \U$18767 ( \19144 , \19133 , \19142 );
or \U$18768 ( \19145 , \19138 , \19143 , \19144 );
and \U$18769 ( \19146 , \8189 , \5708 );
and \U$18770 ( \19147 , \7765 , \5706 );
nor \U$18771 ( \19148 , \19146 , \19147 );
xnor \U$18772 ( \19149 , \19148 , \5467 );
and \U$18773 ( \19150 , \8440 , \5242 );
and \U$18774 ( \19151 , \8435 , \5240 );
nor \U$18775 ( \19152 , \19150 , \19151 );
xnor \U$18776 ( \19153 , \19152 , \5054 );
and \U$18777 ( \19154 , \19149 , \19153 );
and \U$18778 ( \19155 , \9043 , \4868 );
and \U$18779 ( \19156 , \8759 , \4866 );
nor \U$18780 ( \19157 , \19155 , \19156 );
xnor \U$18781 ( \19158 , \19157 , \4636 );
and \U$18782 ( \19159 , \19153 , \19158 );
and \U$18783 ( \19160 , \19149 , \19158 );
or \U$18784 ( \19161 , \19154 , \19159 , \19160 );
and \U$18785 ( \19162 , \19145 , \19161 );
and \U$18786 ( \19163 , \10409 , \3699 );
and \U$18787 ( \19164 , \10228 , \3697 );
nor \U$18788 ( \19165 , \19163 , \19164 );
xnor \U$18789 ( \19166 , \19165 , \3512 );
and \U$18790 ( \19167 , \19161 , \19166 );
and \U$18791 ( \19168 , \19145 , \19166 );
or \U$18792 ( \19169 , \19162 , \19167 , \19168 );
and \U$18793 ( \19170 , \19129 , \19169 );
nand \U$18794 ( \19171 , \11029 , \3384 );
xnor \U$18795 ( \19172 , \19171 , \3181 );
xor \U$18796 ( \19173 , \18977 , \18981 );
xor \U$18797 ( \19174 , \19173 , \18986 );
and \U$18798 ( \19175 , \19172 , \19174 );
xor \U$18799 ( \19176 , \18993 , \18997 );
xor \U$18800 ( \19177 , \19176 , \19002 );
and \U$18801 ( \19178 , \19174 , \19177 );
and \U$18802 ( \19179 , \19172 , \19177 );
or \U$18803 ( \19180 , \19175 , \19178 , \19179 );
and \U$18804 ( \19181 , \19169 , \19180 );
and \U$18805 ( \19182 , \19129 , \19180 );
or \U$18806 ( \19183 , \19170 , \19181 , \19182 );
xor \U$18807 ( \19184 , \18929 , \18933 );
xor \U$18808 ( \19185 , \19184 , \18938 );
xor \U$18809 ( \19186 , \18945 , \18949 );
xor \U$18810 ( \19187 , \19186 , \18954 );
and \U$18811 ( \19188 , \19185 , \19187 );
xor \U$18812 ( \19189 , \18962 , \18966 );
xor \U$18813 ( \19190 , \19189 , \3181 );
and \U$18814 ( \19191 , \19187 , \19190 );
and \U$18815 ( \19192 , \19185 , \19190 );
or \U$18816 ( \19193 , \19188 , \19191 , \19192 );
xor \U$18817 ( \19194 , \18789 , \18793 );
xor \U$18818 ( \19195 , \19194 , \18798 );
and \U$18819 ( \19196 , \19193 , \19195 );
xor \U$18820 ( \19197 , \18805 , \18809 );
xor \U$18821 ( \19198 , \19197 , \18814 );
and \U$18822 ( \19199 , \19195 , \19198 );
and \U$18823 ( \19200 , \19193 , \19198 );
or \U$18824 ( \19201 , \19196 , \19199 , \19200 );
and \U$18825 ( \19202 , \19183 , \19201 );
xor \U$18826 ( \19203 , \18941 , \18957 );
xor \U$18827 ( \19204 , \19203 , \18970 );
xor \U$18828 ( \19205 , \18989 , \19005 );
xor \U$18829 ( \19206 , \19205 , \19010 );
and \U$18830 ( \19207 , \19204 , \19206 );
xor \U$18831 ( \19208 , \19016 , \19018 );
xor \U$18832 ( \19209 , \19208 , \19021 );
and \U$18833 ( \19210 , \19206 , \19209 );
and \U$18834 ( \19211 , \19204 , \19209 );
or \U$18835 ( \19212 , \19207 , \19210 , \19211 );
and \U$18836 ( \19213 , \19201 , \19212 );
and \U$18837 ( \19214 , \19183 , \19212 );
or \U$18838 ( \19215 , \19202 , \19213 , \19214 );
xor \U$18839 ( \19216 , \18973 , \19013 );
xor \U$18840 ( \19217 , \19216 , \19024 );
xor \U$18841 ( \19218 , \19029 , \19031 );
xor \U$18842 ( \19219 , \19218 , \19034 );
and \U$18843 ( \19220 , \19217 , \19219 );
xor \U$18844 ( \19221 , \19040 , \19042 );
and \U$18845 ( \19222 , \19219 , \19221 );
and \U$18846 ( \19223 , \19217 , \19221 );
or \U$18847 ( \19224 , \19220 , \19222 , \19223 );
and \U$18848 ( \19225 , \19215 , \19224 );
xor \U$18849 ( \19226 , \19048 , \19050 );
xor \U$18850 ( \19227 , \19226 , \19053 );
and \U$18851 ( \19228 , \19224 , \19227 );
and \U$18852 ( \19229 , \19215 , \19227 );
or \U$18853 ( \19230 , \19225 , \19228 , \19229 );
xor \U$18854 ( \19231 , \19046 , \19056 );
xor \U$18855 ( \19232 , \19231 , \19059 );
and \U$18856 ( \19233 , \19230 , \19232 );
xor \U$18857 ( \19234 , \19064 , \19066 );
and \U$18858 ( \19235 , \19232 , \19234 );
and \U$18859 ( \19236 , \19230 , \19234 );
or \U$18860 ( \19237 , \19233 , \19235 , \19236 );
and \U$18861 ( \19238 , \19077 , \19237 );
xor \U$18862 ( \19239 , \19077 , \19237 );
xor \U$18863 ( \19240 , \19230 , \19232 );
xor \U$18864 ( \19241 , \19240 , \19234 );
and \U$18865 ( \19242 , \6210 , \7829 );
and \U$18866 ( \19243 , \5838 , \7827 );
nor \U$18867 ( \19244 , \19242 , \19243 );
xnor \U$18868 ( \19245 , \19244 , \7580 );
and \U$18869 ( \19246 , \6562 , \7300 );
and \U$18870 ( \19247 , \6219 , \7298 );
nor \U$18871 ( \19248 , \19246 , \19247 );
xnor \U$18872 ( \19249 , \19248 , \7040 );
and \U$18873 ( \19250 , \19245 , \19249 );
and \U$18874 ( \19251 , \7067 , \6806 );
and \U$18875 ( \19252 , \6764 , \6804 );
nor \U$18876 ( \19253 , \19251 , \19252 );
xnor \U$18877 ( \19254 , \19253 , \6491 );
and \U$18878 ( \19255 , \19249 , \19254 );
and \U$18879 ( \19256 , \19245 , \19254 );
or \U$18880 ( \19257 , \19250 , \19255 , \19256 );
and \U$18881 ( \19258 , \4833 , \9495 );
and \U$18882 ( \19259 , \4531 , \9493 );
nor \U$18883 ( \19260 , \19258 , \19259 );
xnor \U$18884 ( \19261 , \19260 , \9185 );
and \U$18885 ( \19262 , \5310 , \8958 );
and \U$18886 ( \19263 , \4841 , \8956 );
nor \U$18887 ( \19264 , \19262 , \19263 );
xnor \U$18888 ( \19265 , \19264 , \8587 );
and \U$18889 ( \19266 , \19261 , \19265 );
and \U$18890 ( \19267 , \5579 , \8396 );
and \U$18891 ( \19268 , \5315 , \8394 );
nor \U$18892 ( \19269 , \19267 , \19268 );
xnor \U$18893 ( \19270 , \19269 , \8078 );
and \U$18894 ( \19271 , \19265 , \19270 );
and \U$18895 ( \19272 , \19261 , \19270 );
or \U$18896 ( \19273 , \19266 , \19271 , \19272 );
and \U$18897 ( \19274 , \19257 , \19273 );
and \U$18898 ( \19275 , \4073 , \10876 );
and \U$18899 ( \19276 , \3951 , \10873 );
nor \U$18900 ( \19277 , \19275 , \19276 );
xnor \U$18901 ( \19278 , \19277 , \9821 );
and \U$18902 ( \19279 , \4334 , \10063 );
and \U$18903 ( \19280 , \4078 , \10061 );
nor \U$18904 ( \19281 , \19279 , \19280 );
xnor \U$18905 ( \19282 , \19281 , \9824 );
and \U$18906 ( \19283 , \19278 , \19282 );
and \U$18907 ( \19284 , \19282 , \3512 );
and \U$18908 ( \19285 , \19278 , \3512 );
or \U$18909 ( \19286 , \19283 , \19284 , \19285 );
and \U$18910 ( \19287 , \19273 , \19286 );
and \U$18911 ( \19288 , \19257 , \19286 );
or \U$18912 ( \19289 , \19274 , \19287 , \19288 );
and \U$18913 ( \19290 , \7765 , \6297 );
and \U$18914 ( \19291 , \7239 , \6295 );
nor \U$18915 ( \19292 , \19290 , \19291 );
xnor \U$18916 ( \19293 , \19292 , \5957 );
and \U$18917 ( \19294 , \8435 , \5708 );
and \U$18918 ( \19295 , \8189 , \5706 );
nor \U$18919 ( \19296 , \19294 , \19295 );
xnor \U$18920 ( \19297 , \19296 , \5467 );
and \U$18921 ( \19298 , \19293 , \19297 );
and \U$18922 ( \19299 , \8759 , \5242 );
and \U$18923 ( \19300 , \8440 , \5240 );
nor \U$18924 ( \19301 , \19299 , \19300 );
xnor \U$18925 ( \19302 , \19301 , \5054 );
and \U$18926 ( \19303 , \19297 , \19302 );
and \U$18927 ( \19304 , \19293 , \19302 );
or \U$18928 ( \19305 , \19298 , \19303 , \19304 );
and \U$18929 ( \19306 , \9612 , \4868 );
and \U$18930 ( \19307 , \9043 , \4866 );
nor \U$18931 ( \19308 , \19306 , \19307 );
xnor \U$18932 ( \19309 , \19308 , \4636 );
and \U$18933 ( \19310 , \10223 , \4417 );
and \U$18934 ( \19311 , \9620 , \4415 );
nor \U$18935 ( \19312 , \19310 , \19311 );
xnor \U$18936 ( \19313 , \19312 , \4274 );
and \U$18937 ( \19314 , \19309 , \19313 );
and \U$18938 ( \19315 , \10409 , \4094 );
and \U$18939 ( \19316 , \10228 , \4092 );
nor \U$18940 ( \19317 , \19315 , \19316 );
xnor \U$18941 ( \19318 , \19317 , \3848 );
and \U$18942 ( \19319 , \19313 , \19318 );
and \U$18943 ( \19320 , \19309 , \19318 );
or \U$18944 ( \19321 , \19314 , \19319 , \19320 );
and \U$18945 ( \19322 , \19305 , \19321 );
xor \U$18946 ( \19323 , \19133 , \19137 );
xor \U$18947 ( \19324 , \19323 , \19142 );
and \U$18948 ( \19325 , \19321 , \19324 );
and \U$18949 ( \19326 , \19305 , \19324 );
or \U$18950 ( \19327 , \19322 , \19325 , \19326 );
and \U$18951 ( \19328 , \19289 , \19327 );
xor \U$18952 ( \19329 , \19081 , \19085 );
xor \U$18953 ( \19330 , \19329 , \19090 );
xor \U$18954 ( \19331 , \19097 , \19101 );
xor \U$18955 ( \19332 , \19331 , \19106 );
and \U$18956 ( \19333 , \19330 , \19332 );
xor \U$18957 ( \19334 , \19149 , \19153 );
xor \U$18958 ( \19335 , \19334 , \19158 );
and \U$18959 ( \19336 , \19332 , \19335 );
and \U$18960 ( \19337 , \19330 , \19335 );
or \U$18961 ( \19338 , \19333 , \19336 , \19337 );
and \U$18962 ( \19339 , \19327 , \19338 );
and \U$18963 ( \19340 , \19289 , \19338 );
or \U$18964 ( \19341 , \19328 , \19339 , \19340 );
xor \U$18965 ( \19342 , \19145 , \19161 );
xor \U$18966 ( \19343 , \19342 , \19166 );
xor \U$18967 ( \19344 , \19185 , \19187 );
xor \U$18968 ( \19345 , \19344 , \19190 );
and \U$18969 ( \19346 , \19343 , \19345 );
xor \U$18970 ( \19347 , \19172 , \19174 );
xor \U$18971 ( \19348 , \19347 , \19177 );
and \U$18972 ( \19349 , \19345 , \19348 );
and \U$18973 ( \19350 , \19343 , \19348 );
or \U$18974 ( \19351 , \19346 , \19349 , \19350 );
and \U$18975 ( \19352 , \19341 , \19351 );
xor \U$18976 ( \19353 , \19204 , \19206 );
xor \U$18977 ( \19354 , \19353 , \19209 );
and \U$18978 ( \19355 , \19351 , \19354 );
and \U$18979 ( \19356 , \19341 , \19354 );
or \U$18980 ( \19357 , \19352 , \19355 , \19356 );
xor \U$18981 ( \19358 , \19129 , \19169 );
xor \U$18982 ( \19359 , \19358 , \19180 );
xor \U$18983 ( \19360 , \19193 , \19195 );
xor \U$18984 ( \19361 , \19360 , \19198 );
and \U$18985 ( \19362 , \19359 , \19361 );
and \U$18986 ( \19363 , \19357 , \19362 );
xor \U$18987 ( \19364 , \19217 , \19219 );
xor \U$18988 ( \19365 , \19364 , \19221 );
and \U$18989 ( \19366 , \19362 , \19365 );
and \U$18990 ( \19367 , \19357 , \19365 );
or \U$18991 ( \19368 , \19363 , \19366 , \19367 );
xor \U$18992 ( \19369 , \19027 , \19037 );
xor \U$18993 ( \19370 , \19369 , \19043 );
and \U$18994 ( \19371 , \19368 , \19370 );
xor \U$18995 ( \19372 , \19215 , \19224 );
xor \U$18996 ( \19373 , \19372 , \19227 );
and \U$18997 ( \19374 , \19370 , \19373 );
and \U$18998 ( \19375 , \19368 , \19373 );
or \U$18999 ( \19376 , \19371 , \19374 , \19375 );
and \U$19000 ( \19377 , \19241 , \19376 );
xor \U$19001 ( \19378 , \19241 , \19376 );
xor \U$19002 ( \19379 , \19368 , \19370 );
xor \U$19003 ( \19380 , \19379 , \19373 );
and \U$19004 ( \19381 , \4078 , \10876 );
and \U$19005 ( \19382 , \4073 , \10873 );
nor \U$19006 ( \19383 , \19381 , \19382 );
xnor \U$19007 ( \19384 , \19383 , \9821 );
and \U$19008 ( \19385 , \4531 , \10063 );
and \U$19009 ( \19386 , \4334 , \10061 );
nor \U$19010 ( \19387 , \19385 , \19386 );
xnor \U$19011 ( \19388 , \19387 , \9824 );
and \U$19012 ( \19389 , \19384 , \19388 );
and \U$19013 ( \19390 , \4841 , \9495 );
and \U$19014 ( \19391 , \4833 , \9493 );
nor \U$19015 ( \19392 , \19390 , \19391 );
xnor \U$19016 ( \19393 , \19392 , \9185 );
and \U$19017 ( \19394 , \19388 , \19393 );
and \U$19018 ( \19395 , \19384 , \19393 );
or \U$19019 ( \19396 , \19389 , \19394 , \19395 );
and \U$19020 ( \19397 , \6764 , \7300 );
and \U$19021 ( \19398 , \6562 , \7298 );
nor \U$19022 ( \19399 , \19397 , \19398 );
xnor \U$19023 ( \19400 , \19399 , \7040 );
and \U$19024 ( \19401 , \7239 , \6806 );
and \U$19025 ( \19402 , \7067 , \6804 );
nor \U$19026 ( \19403 , \19401 , \19402 );
xnor \U$19027 ( \19404 , \19403 , \6491 );
and \U$19028 ( \19405 , \19400 , \19404 );
and \U$19029 ( \19406 , \8189 , \6297 );
and \U$19030 ( \19407 , \7765 , \6295 );
nor \U$19031 ( \19408 , \19406 , \19407 );
xnor \U$19032 ( \19409 , \19408 , \5957 );
and \U$19033 ( \19410 , \19404 , \19409 );
and \U$19034 ( \19411 , \19400 , \19409 );
or \U$19035 ( \19412 , \19405 , \19410 , \19411 );
and \U$19036 ( \19413 , \19396 , \19412 );
and \U$19037 ( \19414 , \5315 , \8958 );
and \U$19038 ( \19415 , \5310 , \8956 );
nor \U$19039 ( \19416 , \19414 , \19415 );
xnor \U$19040 ( \19417 , \19416 , \8587 );
and \U$19041 ( \19418 , \5838 , \8396 );
and \U$19042 ( \19419 , \5579 , \8394 );
nor \U$19043 ( \19420 , \19418 , \19419 );
xnor \U$19044 ( \19421 , \19420 , \8078 );
and \U$19045 ( \19422 , \19417 , \19421 );
and \U$19046 ( \19423 , \6219 , \7829 );
and \U$19047 ( \19424 , \6210 , \7827 );
nor \U$19048 ( \19425 , \19423 , \19424 );
xnor \U$19049 ( \19426 , \19425 , \7580 );
and \U$19050 ( \19427 , \19421 , \19426 );
and \U$19051 ( \19428 , \19417 , \19426 );
or \U$19052 ( \19429 , \19422 , \19427 , \19428 );
and \U$19053 ( \19430 , \19412 , \19429 );
and \U$19054 ( \19431 , \19396 , \19429 );
or \U$19055 ( \19432 , \19413 , \19430 , \19431 );
xor \U$19056 ( \19433 , \19245 , \19249 );
xor \U$19057 ( \19434 , \19433 , \19254 );
xor \U$19058 ( \19435 , \19261 , \19265 );
xor \U$19059 ( \19436 , \19435 , \19270 );
and \U$19060 ( \19437 , \19434 , \19436 );
xor \U$19061 ( \19438 , \19293 , \19297 );
xor \U$19062 ( \19439 , \19438 , \19302 );
and \U$19063 ( \19440 , \19436 , \19439 );
and \U$19064 ( \19441 , \19434 , \19439 );
or \U$19065 ( \19442 , \19437 , \19440 , \19441 );
and \U$19066 ( \19443 , \19432 , \19442 );
and \U$19067 ( \19444 , \8440 , \5708 );
and \U$19068 ( \19445 , \8435 , \5706 );
nor \U$19069 ( \19446 , \19444 , \19445 );
xnor \U$19070 ( \19447 , \19446 , \5467 );
and \U$19071 ( \19448 , \9043 , \5242 );
and \U$19072 ( \19449 , \8759 , \5240 );
nor \U$19073 ( \19450 , \19448 , \19449 );
xnor \U$19074 ( \19451 , \19450 , \5054 );
and \U$19075 ( \19452 , \19447 , \19451 );
and \U$19076 ( \19453 , \9620 , \4868 );
and \U$19077 ( \19454 , \9612 , \4866 );
nor \U$19078 ( \19455 , \19453 , \19454 );
xnor \U$19079 ( \19456 , \19455 , \4636 );
and \U$19080 ( \19457 , \19451 , \19456 );
and \U$19081 ( \19458 , \19447 , \19456 );
or \U$19082 ( \19459 , \19452 , \19457 , \19458 );
nand \U$19083 ( \19460 , \11029 , \3697 );
xnor \U$19084 ( \19461 , \19460 , \3512 );
and \U$19085 ( \19462 , \19459 , \19461 );
xor \U$19086 ( \19463 , \19309 , \19313 );
xor \U$19087 ( \19464 , \19463 , \19318 );
and \U$19088 ( \19465 , \19461 , \19464 );
and \U$19089 ( \19466 , \19459 , \19464 );
or \U$19090 ( \19467 , \19462 , \19465 , \19466 );
and \U$19091 ( \19468 , \19442 , \19467 );
and \U$19092 ( \19469 , \19432 , \19467 );
or \U$19093 ( \19470 , \19443 , \19468 , \19469 );
xor \U$19094 ( \19471 , \19114 , \19118 );
xor \U$19095 ( \19472 , \19471 , \19123 );
xor \U$19096 ( \19473 , \19305 , \19321 );
xor \U$19097 ( \19474 , \19473 , \19324 );
and \U$19098 ( \19475 , \19472 , \19474 );
xor \U$19099 ( \19476 , \19330 , \19332 );
xor \U$19100 ( \19477 , \19476 , \19335 );
and \U$19101 ( \19478 , \19474 , \19477 );
and \U$19102 ( \19479 , \19472 , \19477 );
or \U$19103 ( \19480 , \19475 , \19478 , \19479 );
and \U$19104 ( \19481 , \19470 , \19480 );
xor \U$19105 ( \19482 , \19093 , \19109 );
xor \U$19106 ( \19483 , \19482 , \19126 );
and \U$19107 ( \19484 , \19480 , \19483 );
and \U$19108 ( \19485 , \19470 , \19483 );
or \U$19109 ( \19486 , \19481 , \19484 , \19485 );
xor \U$19110 ( \19487 , \19341 , \19351 );
xor \U$19111 ( \19488 , \19487 , \19354 );
and \U$19112 ( \19489 , \19486 , \19488 );
xor \U$19113 ( \19490 , \19359 , \19361 );
and \U$19114 ( \19491 , \19488 , \19490 );
and \U$19115 ( \19492 , \19486 , \19490 );
or \U$19116 ( \19493 , \19489 , \19491 , \19492 );
xor \U$19117 ( \19494 , \19183 , \19201 );
xor \U$19118 ( \19495 , \19494 , \19212 );
and \U$19119 ( \19496 , \19493 , \19495 );
xor \U$19120 ( \19497 , \19357 , \19362 );
xor \U$19121 ( \19498 , \19497 , \19365 );
and \U$19122 ( \19499 , \19495 , \19498 );
and \U$19123 ( \19500 , \19493 , \19498 );
or \U$19124 ( \19501 , \19496 , \19499 , \19500 );
and \U$19125 ( \19502 , \19380 , \19501 );
xor \U$19126 ( \19503 , \19380 , \19501 );
xor \U$19127 ( \19504 , \19493 , \19495 );
xor \U$19128 ( \19505 , \19504 , \19498 );
and \U$19129 ( \19506 , \8435 , \6297 );
and \U$19130 ( \19507 , \8189 , \6295 );
nor \U$19131 ( \19508 , \19506 , \19507 );
xnor \U$19132 ( \19509 , \19508 , \5957 );
and \U$19133 ( \19510 , \8759 , \5708 );
and \U$19134 ( \19511 , \8440 , \5706 );
nor \U$19135 ( \19512 , \19510 , \19511 );
xnor \U$19136 ( \19513 , \19512 , \5467 );
and \U$19137 ( \19514 , \19509 , \19513 );
and \U$19138 ( \19515 , \9612 , \5242 );
and \U$19139 ( \19516 , \9043 , \5240 );
nor \U$19140 ( \19517 , \19515 , \19516 );
xnor \U$19141 ( \19518 , \19517 , \5054 );
and \U$19142 ( \19519 , \19513 , \19518 );
and \U$19143 ( \19520 , \19509 , \19518 );
or \U$19144 ( \19521 , \19514 , \19519 , \19520 );
and \U$19145 ( \19522 , \10223 , \4868 );
and \U$19146 ( \19523 , \9620 , \4866 );
nor \U$19147 ( \19524 , \19522 , \19523 );
xnor \U$19148 ( \19525 , \19524 , \4636 );
and \U$19149 ( \19526 , \10409 , \4417 );
and \U$19150 ( \19527 , \10228 , \4415 );
nor \U$19151 ( \19528 , \19526 , \19527 );
xnor \U$19152 ( \19529 , \19528 , \4274 );
and \U$19153 ( \19530 , \19525 , \19529 );
nand \U$19154 ( \19531 , \11029 , \4092 );
xnor \U$19155 ( \19532 , \19531 , \3848 );
and \U$19156 ( \19533 , \19529 , \19532 );
and \U$19157 ( \19534 , \19525 , \19532 );
or \U$19158 ( \19535 , \19530 , \19533 , \19534 );
and \U$19159 ( \19536 , \19521 , \19535 );
and \U$19160 ( \19537 , \10228 , \4417 );
and \U$19161 ( \19538 , \10223 , \4415 );
nor \U$19162 ( \19539 , \19537 , \19538 );
xnor \U$19163 ( \19540 , \19539 , \4274 );
and \U$19164 ( \19541 , \19535 , \19540 );
and \U$19165 ( \19542 , \19521 , \19540 );
or \U$19166 ( \19543 , \19536 , \19541 , \19542 );
and \U$19167 ( \19544 , \6562 , \7829 );
and \U$19168 ( \19545 , \6219 , \7827 );
nor \U$19169 ( \19546 , \19544 , \19545 );
xnor \U$19170 ( \19547 , \19546 , \7580 );
and \U$19171 ( \19548 , \7067 , \7300 );
and \U$19172 ( \19549 , \6764 , \7298 );
nor \U$19173 ( \19550 , \19548 , \19549 );
xnor \U$19174 ( \19551 , \19550 , \7040 );
and \U$19175 ( \19552 , \19547 , \19551 );
and \U$19176 ( \19553 , \7765 , \6806 );
and \U$19177 ( \19554 , \7239 , \6804 );
nor \U$19178 ( \19555 , \19553 , \19554 );
xnor \U$19179 ( \19556 , \19555 , \6491 );
and \U$19180 ( \19557 , \19551 , \19556 );
and \U$19181 ( \19558 , \19547 , \19556 );
or \U$19182 ( \19559 , \19552 , \19557 , \19558 );
and \U$19183 ( \19560 , \4334 , \10876 );
and \U$19184 ( \19561 , \4078 , \10873 );
nor \U$19185 ( \19562 , \19560 , \19561 );
xnor \U$19186 ( \19563 , \19562 , \9821 );
and \U$19187 ( \19564 , \4833 , \10063 );
and \U$19188 ( \19565 , \4531 , \10061 );
nor \U$19189 ( \19566 , \19564 , \19565 );
xnor \U$19190 ( \19567 , \19566 , \9824 );
and \U$19191 ( \19568 , \19563 , \19567 );
and \U$19192 ( \19569 , \19567 , \3848 );
and \U$19193 ( \19570 , \19563 , \3848 );
or \U$19194 ( \19571 , \19568 , \19569 , \19570 );
and \U$19195 ( \19572 , \19559 , \19571 );
and \U$19196 ( \19573 , \5310 , \9495 );
and \U$19197 ( \19574 , \4841 , \9493 );
nor \U$19198 ( \19575 , \19573 , \19574 );
xnor \U$19199 ( \19576 , \19575 , \9185 );
and \U$19200 ( \19577 , \5579 , \8958 );
and \U$19201 ( \19578 , \5315 , \8956 );
nor \U$19202 ( \19579 , \19577 , \19578 );
xnor \U$19203 ( \19580 , \19579 , \8587 );
and \U$19204 ( \19581 , \19576 , \19580 );
and \U$19205 ( \19582 , \6210 , \8396 );
and \U$19206 ( \19583 , \5838 , \8394 );
nor \U$19207 ( \19584 , \19582 , \19583 );
xnor \U$19208 ( \19585 , \19584 , \8078 );
and \U$19209 ( \19586 , \19580 , \19585 );
and \U$19210 ( \19587 , \19576 , \19585 );
or \U$19211 ( \19588 , \19581 , \19586 , \19587 );
and \U$19212 ( \19589 , \19571 , \19588 );
and \U$19213 ( \19590 , \19559 , \19588 );
or \U$19214 ( \19591 , \19572 , \19589 , \19590 );
and \U$19215 ( \19592 , \19543 , \19591 );
and \U$19216 ( \19593 , \11029 , \4094 );
and \U$19217 ( \19594 , \10409 , \4092 );
nor \U$19218 ( \19595 , \19593 , \19594 );
xnor \U$19219 ( \19596 , \19595 , \3848 );
xor \U$19220 ( \19597 , \19447 , \19451 );
xor \U$19221 ( \19598 , \19597 , \19456 );
and \U$19222 ( \19599 , \19596 , \19598 );
xor \U$19223 ( \19600 , \19400 , \19404 );
xor \U$19224 ( \19601 , \19600 , \19409 );
and \U$19225 ( \19602 , \19598 , \19601 );
and \U$19226 ( \19603 , \19596 , \19601 );
or \U$19227 ( \19604 , \19599 , \19602 , \19603 );
and \U$19228 ( \19605 , \19591 , \19604 );
and \U$19229 ( \19606 , \19543 , \19604 );
or \U$19230 ( \19607 , \19592 , \19605 , \19606 );
xor \U$19231 ( \19608 , \19278 , \19282 );
xor \U$19232 ( \19609 , \19608 , \3512 );
xor \U$19233 ( \19610 , \19434 , \19436 );
xor \U$19234 ( \19611 , \19610 , \19439 );
and \U$19235 ( \19612 , \19609 , \19611 );
xor \U$19236 ( \19613 , \19459 , \19461 );
xor \U$19237 ( \19614 , \19613 , \19464 );
and \U$19238 ( \19615 , \19611 , \19614 );
and \U$19239 ( \19616 , \19609 , \19614 );
or \U$19240 ( \19617 , \19612 , \19615 , \19616 );
and \U$19241 ( \19618 , \19607 , \19617 );
xor \U$19242 ( \19619 , \19257 , \19273 );
xor \U$19243 ( \19620 , \19619 , \19286 );
and \U$19244 ( \19621 , \19617 , \19620 );
and \U$19245 ( \19622 , \19607 , \19620 );
or \U$19246 ( \19623 , \19618 , \19621 , \19622 );
xor \U$19247 ( \19624 , \19432 , \19442 );
xor \U$19248 ( \19625 , \19624 , \19467 );
xor \U$19249 ( \19626 , \19472 , \19474 );
xor \U$19250 ( \19627 , \19626 , \19477 );
and \U$19251 ( \19628 , \19625 , \19627 );
and \U$19252 ( \19629 , \19623 , \19628 );
xor \U$19253 ( \19630 , \19343 , \19345 );
xor \U$19254 ( \19631 , \19630 , \19348 );
and \U$19255 ( \19632 , \19628 , \19631 );
and \U$19256 ( \19633 , \19623 , \19631 );
or \U$19257 ( \19634 , \19629 , \19632 , \19633 );
xor \U$19258 ( \19635 , \19289 , \19327 );
xor \U$19259 ( \19636 , \19635 , \19338 );
xor \U$19260 ( \19637 , \19470 , \19480 );
xor \U$19261 ( \19638 , \19637 , \19483 );
and \U$19262 ( \19639 , \19636 , \19638 );
and \U$19263 ( \19640 , \19634 , \19639 );
xor \U$19264 ( \19641 , \19486 , \19488 );
xor \U$19265 ( \19642 , \19641 , \19490 );
and \U$19266 ( \19643 , \19639 , \19642 );
and \U$19267 ( \19644 , \19634 , \19642 );
or \U$19268 ( \19645 , \19640 , \19643 , \19644 );
and \U$19269 ( \19646 , \19505 , \19645 );
xor \U$19270 ( \19647 , \19505 , \19645 );
xor \U$19271 ( \19648 , \19634 , \19639 );
xor \U$19272 ( \19649 , \19648 , \19642 );
and \U$19273 ( \19650 , \5838 , \8958 );
and \U$19274 ( \19651 , \5579 , \8956 );
nor \U$19275 ( \19652 , \19650 , \19651 );
xnor \U$19276 ( \19653 , \19652 , \8587 );
and \U$19277 ( \19654 , \6219 , \8396 );
and \U$19278 ( \19655 , \6210 , \8394 );
nor \U$19279 ( \19656 , \19654 , \19655 );
xnor \U$19280 ( \19657 , \19656 , \8078 );
and \U$19281 ( \19658 , \19653 , \19657 );
and \U$19282 ( \19659 , \6764 , \7829 );
and \U$19283 ( \19660 , \6562 , \7827 );
nor \U$19284 ( \19661 , \19659 , \19660 );
xnor \U$19285 ( \19662 , \19661 , \7580 );
and \U$19286 ( \19663 , \19657 , \19662 );
and \U$19287 ( \19664 , \19653 , \19662 );
or \U$19288 ( \19665 , \19658 , \19663 , \19664 );
and \U$19289 ( \19666 , \4531 , \10876 );
and \U$19290 ( \19667 , \4334 , \10873 );
nor \U$19291 ( \19668 , \19666 , \19667 );
xnor \U$19292 ( \19669 , \19668 , \9821 );
and \U$19293 ( \19670 , \4841 , \10063 );
and \U$19294 ( \19671 , \4833 , \10061 );
nor \U$19295 ( \19672 , \19670 , \19671 );
xnor \U$19296 ( \19673 , \19672 , \9824 );
and \U$19297 ( \19674 , \19669 , \19673 );
and \U$19298 ( \19675 , \5315 , \9495 );
and \U$19299 ( \19676 , \5310 , \9493 );
nor \U$19300 ( \19677 , \19675 , \19676 );
xnor \U$19301 ( \19678 , \19677 , \9185 );
and \U$19302 ( \19679 , \19673 , \19678 );
and \U$19303 ( \19680 , \19669 , \19678 );
or \U$19304 ( \19681 , \19674 , \19679 , \19680 );
and \U$19305 ( \19682 , \19665 , \19681 );
and \U$19306 ( \19683 , \7239 , \7300 );
and \U$19307 ( \19684 , \7067 , \7298 );
nor \U$19308 ( \19685 , \19683 , \19684 );
xnor \U$19309 ( \19686 , \19685 , \7040 );
and \U$19310 ( \19687 , \8189 , \6806 );
and \U$19311 ( \19688 , \7765 , \6804 );
nor \U$19312 ( \19689 , \19687 , \19688 );
xnor \U$19313 ( \19690 , \19689 , \6491 );
and \U$19314 ( \19691 , \19686 , \19690 );
and \U$19315 ( \19692 , \8440 , \6297 );
and \U$19316 ( \19693 , \8435 , \6295 );
nor \U$19317 ( \19694 , \19692 , \19693 );
xnor \U$19318 ( \19695 , \19694 , \5957 );
and \U$19319 ( \19696 , \19690 , \19695 );
and \U$19320 ( \19697 , \19686 , \19695 );
or \U$19321 ( \19698 , \19691 , \19696 , \19697 );
and \U$19322 ( \19699 , \19681 , \19698 );
and \U$19323 ( \19700 , \19665 , \19698 );
or \U$19324 ( \19701 , \19682 , \19699 , \19700 );
xor \U$19325 ( \19702 , \19547 , \19551 );
xor \U$19326 ( \19703 , \19702 , \19556 );
xor \U$19327 ( \19704 , \19563 , \19567 );
xor \U$19328 ( \19705 , \19704 , \3848 );
and \U$19329 ( \19706 , \19703 , \19705 );
xor \U$19330 ( \19707 , \19576 , \19580 );
xor \U$19331 ( \19708 , \19707 , \19585 );
and \U$19332 ( \19709 , \19705 , \19708 );
and \U$19333 ( \19710 , \19703 , \19708 );
or \U$19334 ( \19711 , \19706 , \19709 , \19710 );
and \U$19335 ( \19712 , \19701 , \19711 );
and \U$19336 ( \19713 , \9043 , \5708 );
and \U$19337 ( \19714 , \8759 , \5706 );
nor \U$19338 ( \19715 , \19713 , \19714 );
xnor \U$19339 ( \19716 , \19715 , \5467 );
and \U$19340 ( \19717 , \9620 , \5242 );
and \U$19341 ( \19718 , \9612 , \5240 );
nor \U$19342 ( \19719 , \19717 , \19718 );
xnor \U$19343 ( \19720 , \19719 , \5054 );
and \U$19344 ( \19721 , \19716 , \19720 );
and \U$19345 ( \19722 , \10228 , \4868 );
and \U$19346 ( \19723 , \10223 , \4866 );
nor \U$19347 ( \19724 , \19722 , \19723 );
xnor \U$19348 ( \19725 , \19724 , \4636 );
and \U$19349 ( \19726 , \19720 , \19725 );
and \U$19350 ( \19727 , \19716 , \19725 );
or \U$19351 ( \19728 , \19721 , \19726 , \19727 );
xor \U$19352 ( \19729 , \19509 , \19513 );
xor \U$19353 ( \19730 , \19729 , \19518 );
and \U$19354 ( \19731 , \19728 , \19730 );
xor \U$19355 ( \19732 , \19525 , \19529 );
xor \U$19356 ( \19733 , \19732 , \19532 );
and \U$19357 ( \19734 , \19730 , \19733 );
and \U$19358 ( \19735 , \19728 , \19733 );
or \U$19359 ( \19736 , \19731 , \19734 , \19735 );
and \U$19360 ( \19737 , \19711 , \19736 );
and \U$19361 ( \19738 , \19701 , \19736 );
or \U$19362 ( \19739 , \19712 , \19737 , \19738 );
xor \U$19363 ( \19740 , \19384 , \19388 );
xor \U$19364 ( \19741 , \19740 , \19393 );
xor \U$19365 ( \19742 , \19417 , \19421 );
xor \U$19366 ( \19743 , \19742 , \19426 );
and \U$19367 ( \19744 , \19741 , \19743 );
xor \U$19368 ( \19745 , \19596 , \19598 );
xor \U$19369 ( \19746 , \19745 , \19601 );
and \U$19370 ( \19747 , \19743 , \19746 );
and \U$19371 ( \19748 , \19741 , \19746 );
or \U$19372 ( \19749 , \19744 , \19747 , \19748 );
and \U$19373 ( \19750 , \19739 , \19749 );
xor \U$19374 ( \19751 , \19396 , \19412 );
xor \U$19375 ( \19752 , \19751 , \19429 );
and \U$19376 ( \19753 , \19749 , \19752 );
and \U$19377 ( \19754 , \19739 , \19752 );
or \U$19378 ( \19755 , \19750 , \19753 , \19754 );
xor \U$19379 ( \19756 , \19607 , \19617 );
xor \U$19380 ( \19757 , \19756 , \19620 );
and \U$19381 ( \19758 , \19755 , \19757 );
xor \U$19382 ( \19759 , \19625 , \19627 );
and \U$19383 ( \19760 , \19757 , \19759 );
and \U$19384 ( \19761 , \19755 , \19759 );
or \U$19385 ( \19762 , \19758 , \19760 , \19761 );
xor \U$19386 ( \19763 , \19623 , \19628 );
xor \U$19387 ( \19764 , \19763 , \19631 );
and \U$19388 ( \19765 , \19762 , \19764 );
xor \U$19389 ( \19766 , \19636 , \19638 );
and \U$19390 ( \19767 , \19764 , \19766 );
and \U$19391 ( \19768 , \19762 , \19766 );
or \U$19392 ( \19769 , \19765 , \19767 , \19768 );
and \U$19393 ( \19770 , \19649 , \19769 );
xor \U$19394 ( \19771 , \19649 , \19769 );
xor \U$19395 ( \19772 , \19762 , \19764 );
xor \U$19396 ( \19773 , \19772 , \19766 );
and \U$19397 ( \19774 , \5579 , \9495 );
and \U$19398 ( \19775 , \5315 , \9493 );
nor \U$19399 ( \19776 , \19774 , \19775 );
xnor \U$19400 ( \19777 , \19776 , \9185 );
and \U$19401 ( \19778 , \6210 , \8958 );
and \U$19402 ( \19779 , \5838 , \8956 );
nor \U$19403 ( \19780 , \19778 , \19779 );
xnor \U$19404 ( \19781 , \19780 , \8587 );
and \U$19405 ( \19782 , \19777 , \19781 );
and \U$19406 ( \19783 , \6562 , \8396 );
and \U$19407 ( \19784 , \6219 , \8394 );
nor \U$19408 ( \19785 , \19783 , \19784 );
xnor \U$19409 ( \19786 , \19785 , \8078 );
and \U$19410 ( \19787 , \19781 , \19786 );
and \U$19411 ( \19788 , \19777 , \19786 );
or \U$19412 ( \19789 , \19782 , \19787 , \19788 );
and \U$19413 ( \19790 , \4833 , \10876 );
and \U$19414 ( \19791 , \4531 , \10873 );
nor \U$19415 ( \19792 , \19790 , \19791 );
xnor \U$19416 ( \19793 , \19792 , \9821 );
and \U$19417 ( \19794 , \5310 , \10063 );
and \U$19418 ( \19795 , \4841 , \10061 );
nor \U$19419 ( \19796 , \19794 , \19795 );
xnor \U$19420 ( \19797 , \19796 , \9824 );
and \U$19421 ( \19798 , \19793 , \19797 );
and \U$19422 ( \19799 , \19797 , \4274 );
and \U$19423 ( \19800 , \19793 , \4274 );
or \U$19424 ( \19801 , \19798 , \19799 , \19800 );
and \U$19425 ( \19802 , \19789 , \19801 );
and \U$19426 ( \19803 , \7067 , \7829 );
and \U$19427 ( \19804 , \6764 , \7827 );
nor \U$19428 ( \19805 , \19803 , \19804 );
xnor \U$19429 ( \19806 , \19805 , \7580 );
and \U$19430 ( \19807 , \7765 , \7300 );
and \U$19431 ( \19808 , \7239 , \7298 );
nor \U$19432 ( \19809 , \19807 , \19808 );
xnor \U$19433 ( \19810 , \19809 , \7040 );
and \U$19434 ( \19811 , \19806 , \19810 );
and \U$19435 ( \19812 , \8435 , \6806 );
and \U$19436 ( \19813 , \8189 , \6804 );
nor \U$19437 ( \19814 , \19812 , \19813 );
xnor \U$19438 ( \19815 , \19814 , \6491 );
and \U$19439 ( \19816 , \19810 , \19815 );
and \U$19440 ( \19817 , \19806 , \19815 );
or \U$19441 ( \19818 , \19811 , \19816 , \19817 );
and \U$19442 ( \19819 , \19801 , \19818 );
and \U$19443 ( \19820 , \19789 , \19818 );
or \U$19444 ( \19821 , \19802 , \19819 , \19820 );
and \U$19445 ( \19822 , \8759 , \6297 );
and \U$19446 ( \19823 , \8440 , \6295 );
nor \U$19447 ( \19824 , \19822 , \19823 );
xnor \U$19448 ( \19825 , \19824 , \5957 );
and \U$19449 ( \19826 , \9612 , \5708 );
and \U$19450 ( \19827 , \9043 , \5706 );
nor \U$19451 ( \19828 , \19826 , \19827 );
xnor \U$19452 ( \19829 , \19828 , \5467 );
and \U$19453 ( \19830 , \19825 , \19829 );
and \U$19454 ( \19831 , \10223 , \5242 );
and \U$19455 ( \19832 , \9620 , \5240 );
nor \U$19456 ( \19833 , \19831 , \19832 );
xnor \U$19457 ( \19834 , \19833 , \5054 );
and \U$19458 ( \19835 , \19829 , \19834 );
and \U$19459 ( \19836 , \19825 , \19834 );
or \U$19460 ( \19837 , \19830 , \19835 , \19836 );
and \U$19461 ( \19838 , \10409 , \4868 );
and \U$19462 ( \19839 , \10228 , \4866 );
nor \U$19463 ( \19840 , \19838 , \19839 );
xnor \U$19464 ( \19841 , \19840 , \4636 );
nand \U$19465 ( \19842 , \11029 , \4415 );
xnor \U$19466 ( \19843 , \19842 , \4274 );
and \U$19467 ( \19844 , \19841 , \19843 );
and \U$19468 ( \19845 , \19837 , \19844 );
and \U$19469 ( \19846 , \11029 , \4417 );
and \U$19470 ( \19847 , \10409 , \4415 );
nor \U$19471 ( \19848 , \19846 , \19847 );
xnor \U$19472 ( \19849 , \19848 , \4274 );
and \U$19473 ( \19850 , \19844 , \19849 );
and \U$19474 ( \19851 , \19837 , \19849 );
or \U$19475 ( \19852 , \19845 , \19850 , \19851 );
and \U$19476 ( \19853 , \19821 , \19852 );
xor \U$19477 ( \19854 , \19653 , \19657 );
xor \U$19478 ( \19855 , \19854 , \19662 );
xor \U$19479 ( \19856 , \19716 , \19720 );
xor \U$19480 ( \19857 , \19856 , \19725 );
and \U$19481 ( \19858 , \19855 , \19857 );
xor \U$19482 ( \19859 , \19686 , \19690 );
xor \U$19483 ( \19860 , \19859 , \19695 );
and \U$19484 ( \19861 , \19857 , \19860 );
and \U$19485 ( \19862 , \19855 , \19860 );
or \U$19486 ( \19863 , \19858 , \19861 , \19862 );
and \U$19487 ( \19864 , \19852 , \19863 );
and \U$19488 ( \19865 , \19821 , \19863 );
or \U$19489 ( \19866 , \19853 , \19864 , \19865 );
xor \U$19490 ( \19867 , \19665 , \19681 );
xor \U$19491 ( \19868 , \19867 , \19698 );
xor \U$19492 ( \19869 , \19703 , \19705 );
xor \U$19493 ( \19870 , \19869 , \19708 );
and \U$19494 ( \19871 , \19868 , \19870 );
xor \U$19495 ( \19872 , \19728 , \19730 );
xor \U$19496 ( \19873 , \19872 , \19733 );
and \U$19497 ( \19874 , \19870 , \19873 );
and \U$19498 ( \19875 , \19868 , \19873 );
or \U$19499 ( \19876 , \19871 , \19874 , \19875 );
and \U$19500 ( \19877 , \19866 , \19876 );
xor \U$19501 ( \19878 , \19521 , \19535 );
xor \U$19502 ( \19879 , \19878 , \19540 );
and \U$19503 ( \19880 , \19876 , \19879 );
and \U$19504 ( \19881 , \19866 , \19879 );
or \U$19505 ( \19882 , \19877 , \19880 , \19881 );
xor \U$19506 ( \19883 , \19559 , \19571 );
xor \U$19507 ( \19884 , \19883 , \19588 );
xor \U$19508 ( \19885 , \19701 , \19711 );
xor \U$19509 ( \19886 , \19885 , \19736 );
and \U$19510 ( \19887 , \19884 , \19886 );
xor \U$19511 ( \19888 , \19741 , \19743 );
xor \U$19512 ( \19889 , \19888 , \19746 );
and \U$19513 ( \19890 , \19886 , \19889 );
and \U$19514 ( \19891 , \19884 , \19889 );
or \U$19515 ( \19892 , \19887 , \19890 , \19891 );
and \U$19516 ( \19893 , \19882 , \19892 );
xor \U$19517 ( \19894 , \19609 , \19611 );
xor \U$19518 ( \19895 , \19894 , \19614 );
and \U$19519 ( \19896 , \19892 , \19895 );
and \U$19520 ( \19897 , \19882 , \19895 );
or \U$19521 ( \19898 , \19893 , \19896 , \19897 );
xor \U$19522 ( \19899 , \19543 , \19591 );
xor \U$19523 ( \19900 , \19899 , \19604 );
xor \U$19524 ( \19901 , \19739 , \19749 );
xor \U$19525 ( \19902 , \19901 , \19752 );
and \U$19526 ( \19903 , \19900 , \19902 );
and \U$19527 ( \19904 , \19898 , \19903 );
xor \U$19528 ( \19905 , \19755 , \19757 );
xor \U$19529 ( \19906 , \19905 , \19759 );
and \U$19530 ( \19907 , \19903 , \19906 );
and \U$19531 ( \19908 , \19898 , \19906 );
or \U$19532 ( \19909 , \19904 , \19907 , \19908 );
and \U$19533 ( \19910 , \19773 , \19909 );
xor \U$19534 ( \19911 , \19773 , \19909 );
xor \U$19535 ( \19912 , \19898 , \19903 );
xor \U$19536 ( \19913 , \19912 , \19906 );
and \U$19537 ( \19914 , \6219 , \8958 );
and \U$19538 ( \19915 , \6210 , \8956 );
nor \U$19539 ( \19916 , \19914 , \19915 );
xnor \U$19540 ( \19917 , \19916 , \8587 );
and \U$19541 ( \19918 , \6764 , \8396 );
and \U$19542 ( \19919 , \6562 , \8394 );
nor \U$19543 ( \19920 , \19918 , \19919 );
xnor \U$19544 ( \19921 , \19920 , \8078 );
and \U$19545 ( \19922 , \19917 , \19921 );
and \U$19546 ( \19923 , \7239 , \7829 );
and \U$19547 ( \19924 , \7067 , \7827 );
nor \U$19548 ( \19925 , \19923 , \19924 );
xnor \U$19549 ( \19926 , \19925 , \7580 );
and \U$19550 ( \19927 , \19921 , \19926 );
and \U$19551 ( \19928 , \19917 , \19926 );
or \U$19552 ( \19929 , \19922 , \19927 , \19928 );
and \U$19553 ( \19930 , \8189 , \7300 );
and \U$19554 ( \19931 , \7765 , \7298 );
nor \U$19555 ( \19932 , \19930 , \19931 );
xnor \U$19556 ( \19933 , \19932 , \7040 );
and \U$19557 ( \19934 , \8440 , \6806 );
and \U$19558 ( \19935 , \8435 , \6804 );
nor \U$19559 ( \19936 , \19934 , \19935 );
xnor \U$19560 ( \19937 , \19936 , \6491 );
and \U$19561 ( \19938 , \19933 , \19937 );
and \U$19562 ( \19939 , \9043 , \6297 );
and \U$19563 ( \19940 , \8759 , \6295 );
nor \U$19564 ( \19941 , \19939 , \19940 );
xnor \U$19565 ( \19942 , \19941 , \5957 );
and \U$19566 ( \19943 , \19937 , \19942 );
and \U$19567 ( \19944 , \19933 , \19942 );
or \U$19568 ( \19945 , \19938 , \19943 , \19944 );
and \U$19569 ( \19946 , \19929 , \19945 );
and \U$19570 ( \19947 , \4841 , \10876 );
and \U$19571 ( \19948 , \4833 , \10873 );
nor \U$19572 ( \19949 , \19947 , \19948 );
xnor \U$19573 ( \19950 , \19949 , \9821 );
and \U$19574 ( \19951 , \5315 , \10063 );
and \U$19575 ( \19952 , \5310 , \10061 );
nor \U$19576 ( \19953 , \19951 , \19952 );
xnor \U$19577 ( \19954 , \19953 , \9824 );
and \U$19578 ( \19955 , \19950 , \19954 );
and \U$19579 ( \19956 , \5838 , \9495 );
and \U$19580 ( \19957 , \5579 , \9493 );
nor \U$19581 ( \19958 , \19956 , \19957 );
xnor \U$19582 ( \19959 , \19958 , \9185 );
and \U$19583 ( \19960 , \19954 , \19959 );
and \U$19584 ( \19961 , \19950 , \19959 );
or \U$19585 ( \19962 , \19955 , \19960 , \19961 );
and \U$19586 ( \19963 , \19945 , \19962 );
and \U$19587 ( \19964 , \19929 , \19962 );
or \U$19588 ( \19965 , \19946 , \19963 , \19964 );
xor \U$19589 ( \19966 , \19777 , \19781 );
xor \U$19590 ( \19967 , \19966 , \19786 );
xor \U$19591 ( \19968 , \19793 , \19797 );
xor \U$19592 ( \19969 , \19968 , \4274 );
and \U$19593 ( \19970 , \19967 , \19969 );
xor \U$19594 ( \19971 , \19806 , \19810 );
xor \U$19595 ( \19972 , \19971 , \19815 );
and \U$19596 ( \19973 , \19969 , \19972 );
and \U$19597 ( \19974 , \19967 , \19972 );
or \U$19598 ( \19975 , \19970 , \19973 , \19974 );
and \U$19599 ( \19976 , \19965 , \19975 );
and \U$19600 ( \19977 , \9620 , \5708 );
and \U$19601 ( \19978 , \9612 , \5706 );
nor \U$19602 ( \19979 , \19977 , \19978 );
xnor \U$19603 ( \19980 , \19979 , \5467 );
and \U$19604 ( \19981 , \10228 , \5242 );
and \U$19605 ( \19982 , \10223 , \5240 );
nor \U$19606 ( \19983 , \19981 , \19982 );
xnor \U$19607 ( \19984 , \19983 , \5054 );
and \U$19608 ( \19985 , \19980 , \19984 );
and \U$19609 ( \19986 , \11029 , \4868 );
and \U$19610 ( \19987 , \10409 , \4866 );
nor \U$19611 ( \19988 , \19986 , \19987 );
xnor \U$19612 ( \19989 , \19988 , \4636 );
and \U$19613 ( \19990 , \19984 , \19989 );
and \U$19614 ( \19991 , \19980 , \19989 );
or \U$19615 ( \19992 , \19985 , \19990 , \19991 );
xor \U$19616 ( \19993 , \19825 , \19829 );
xor \U$19617 ( \19994 , \19993 , \19834 );
and \U$19618 ( \19995 , \19992 , \19994 );
xor \U$19619 ( \19996 , \19841 , \19843 );
and \U$19620 ( \19997 , \19994 , \19996 );
and \U$19621 ( \19998 , \19992 , \19996 );
or \U$19622 ( \19999 , \19995 , \19997 , \19998 );
and \U$19623 ( \20000 , \19975 , \19999 );
and \U$19624 ( \20001 , \19965 , \19999 );
or \U$19625 ( \20002 , \19976 , \20000 , \20001 );
xor \U$19626 ( \20003 , \19669 , \19673 );
xor \U$19627 ( \20004 , \20003 , \19678 );
xor \U$19628 ( \20005 , \19837 , \19844 );
xor \U$19629 ( \20006 , \20005 , \19849 );
and \U$19630 ( \20007 , \20004 , \20006 );
xor \U$19631 ( \20008 , \19855 , \19857 );
xor \U$19632 ( \20009 , \20008 , \19860 );
and \U$19633 ( \20010 , \20006 , \20009 );
and \U$19634 ( \20011 , \20004 , \20009 );
or \U$19635 ( \20012 , \20007 , \20010 , \20011 );
and \U$19636 ( \20013 , \20002 , \20012 );
xor \U$19637 ( \20014 , \19868 , \19870 );
xor \U$19638 ( \20015 , \20014 , \19873 );
and \U$19639 ( \20016 , \20012 , \20015 );
and \U$19640 ( \20017 , \20002 , \20015 );
or \U$19641 ( \20018 , \20013 , \20016 , \20017 );
xor \U$19642 ( \20019 , \19866 , \19876 );
xor \U$19643 ( \20020 , \20019 , \19879 );
and \U$19644 ( \20021 , \20018 , \20020 );
xor \U$19645 ( \20022 , \19884 , \19886 );
xor \U$19646 ( \20023 , \20022 , \19889 );
and \U$19647 ( \20024 , \20020 , \20023 );
and \U$19648 ( \20025 , \20018 , \20023 );
or \U$19649 ( \20026 , \20021 , \20024 , \20025 );
xor \U$19650 ( \20027 , \19882 , \19892 );
xor \U$19651 ( \20028 , \20027 , \19895 );
and \U$19652 ( \20029 , \20026 , \20028 );
xor \U$19653 ( \20030 , \19900 , \19902 );
and \U$19654 ( \20031 , \20028 , \20030 );
and \U$19655 ( \20032 , \20026 , \20030 );
or \U$19656 ( \20033 , \20029 , \20031 , \20032 );
and \U$19657 ( \20034 , \19913 , \20033 );
xor \U$19658 ( \20035 , \19913 , \20033 );
xor \U$19659 ( \20036 , \20026 , \20028 );
xor \U$19660 ( \20037 , \20036 , \20030 );
and \U$19661 ( \20038 , \6210 , \9495 );
and \U$19662 ( \20039 , \5838 , \9493 );
nor \U$19663 ( \20040 , \20038 , \20039 );
xnor \U$19664 ( \20041 , \20040 , \9185 );
and \U$19665 ( \20042 , \6562 , \8958 );
and \U$19666 ( \20043 , \6219 , \8956 );
nor \U$19667 ( \20044 , \20042 , \20043 );
xnor \U$19668 ( \20045 , \20044 , \8587 );
and \U$19669 ( \20046 , \20041 , \20045 );
and \U$19670 ( \20047 , \7067 , \8396 );
and \U$19671 ( \20048 , \6764 , \8394 );
nor \U$19672 ( \20049 , \20047 , \20048 );
xnor \U$19673 ( \20050 , \20049 , \8078 );
and \U$19674 ( \20051 , \20045 , \20050 );
and \U$19675 ( \20052 , \20041 , \20050 );
or \U$19676 ( \20053 , \20046 , \20051 , \20052 );
and \U$19677 ( \20054 , \7765 , \7829 );
and \U$19678 ( \20055 , \7239 , \7827 );
nor \U$19679 ( \20056 , \20054 , \20055 );
xnor \U$19680 ( \20057 , \20056 , \7580 );
and \U$19681 ( \20058 , \8435 , \7300 );
and \U$19682 ( \20059 , \8189 , \7298 );
nor \U$19683 ( \20060 , \20058 , \20059 );
xnor \U$19684 ( \20061 , \20060 , \7040 );
and \U$19685 ( \20062 , \20057 , \20061 );
and \U$19686 ( \20063 , \8759 , \6806 );
and \U$19687 ( \20064 , \8440 , \6804 );
nor \U$19688 ( \20065 , \20063 , \20064 );
xnor \U$19689 ( \20066 , \20065 , \6491 );
and \U$19690 ( \20067 , \20061 , \20066 );
and \U$19691 ( \20068 , \20057 , \20066 );
or \U$19692 ( \20069 , \20062 , \20067 , \20068 );
and \U$19693 ( \20070 , \20053 , \20069 );
and \U$19694 ( \20071 , \5310 , \10876 );
and \U$19695 ( \20072 , \4841 , \10873 );
nor \U$19696 ( \20073 , \20071 , \20072 );
xnor \U$19697 ( \20074 , \20073 , \9821 );
and \U$19698 ( \20075 , \5579 , \10063 );
and \U$19699 ( \20076 , \5315 , \10061 );
nor \U$19700 ( \20077 , \20075 , \20076 );
xnor \U$19701 ( \20078 , \20077 , \9824 );
and \U$19702 ( \20079 , \20074 , \20078 );
and \U$19703 ( \20080 , \20078 , \4636 );
and \U$19704 ( \20081 , \20074 , \4636 );
or \U$19705 ( \20082 , \20079 , \20080 , \20081 );
and \U$19706 ( \20083 , \20069 , \20082 );
and \U$19707 ( \20084 , \20053 , \20082 );
or \U$19708 ( \20085 , \20070 , \20083 , \20084 );
and \U$19709 ( \20086 , \9612 , \6297 );
and \U$19710 ( \20087 , \9043 , \6295 );
nor \U$19711 ( \20088 , \20086 , \20087 );
xnor \U$19712 ( \20089 , \20088 , \5957 );
and \U$19713 ( \20090 , \10223 , \5708 );
and \U$19714 ( \20091 , \9620 , \5706 );
nor \U$19715 ( \20092 , \20090 , \20091 );
xnor \U$19716 ( \20093 , \20092 , \5467 );
and \U$19717 ( \20094 , \20089 , \20093 );
and \U$19718 ( \20095 , \10409 , \5242 );
and \U$19719 ( \20096 , \10228 , \5240 );
nor \U$19720 ( \20097 , \20095 , \20096 );
xnor \U$19721 ( \20098 , \20097 , \5054 );
and \U$19722 ( \20099 , \20093 , \20098 );
and \U$19723 ( \20100 , \20089 , \20098 );
or \U$19724 ( \20101 , \20094 , \20099 , \20100 );
xor \U$19725 ( \20102 , \19933 , \19937 );
xor \U$19726 ( \20103 , \20102 , \19942 );
and \U$19727 ( \20104 , \20101 , \20103 );
xor \U$19728 ( \20105 , \19980 , \19984 );
xor \U$19729 ( \20106 , \20105 , \19989 );
and \U$19730 ( \20107 , \20103 , \20106 );
and \U$19731 ( \20108 , \20101 , \20106 );
or \U$19732 ( \20109 , \20104 , \20107 , \20108 );
and \U$19733 ( \20110 , \20085 , \20109 );
xor \U$19734 ( \20111 , \19917 , \19921 );
xor \U$19735 ( \20112 , \20111 , \19926 );
xor \U$19736 ( \20113 , \19950 , \19954 );
xor \U$19737 ( \20114 , \20113 , \19959 );
and \U$19738 ( \20115 , \20112 , \20114 );
and \U$19739 ( \20116 , \20109 , \20115 );
and \U$19740 ( \20117 , \20085 , \20115 );
or \U$19741 ( \20118 , \20110 , \20116 , \20117 );
xor \U$19742 ( \20119 , \19929 , \19945 );
xor \U$19743 ( \20120 , \20119 , \19962 );
xor \U$19744 ( \20121 , \19967 , \19969 );
xor \U$19745 ( \20122 , \20121 , \19972 );
and \U$19746 ( \20123 , \20120 , \20122 );
xor \U$19747 ( \20124 , \19992 , \19994 );
xor \U$19748 ( \20125 , \20124 , \19996 );
and \U$19749 ( \20126 , \20122 , \20125 );
and \U$19750 ( \20127 , \20120 , \20125 );
or \U$19751 ( \20128 , \20123 , \20126 , \20127 );
and \U$19752 ( \20129 , \20118 , \20128 );
xor \U$19753 ( \20130 , \19789 , \19801 );
xor \U$19754 ( \20131 , \20130 , \19818 );
and \U$19755 ( \20132 , \20128 , \20131 );
and \U$19756 ( \20133 , \20118 , \20131 );
or \U$19757 ( \20134 , \20129 , \20132 , \20133 );
xor \U$19758 ( \20135 , \19965 , \19975 );
xor \U$19759 ( \20136 , \20135 , \19999 );
xor \U$19760 ( \20137 , \20004 , \20006 );
xor \U$19761 ( \20138 , \20137 , \20009 );
and \U$19762 ( \20139 , \20136 , \20138 );
and \U$19763 ( \20140 , \20134 , \20139 );
xor \U$19764 ( \20141 , \19821 , \19852 );
xor \U$19765 ( \20142 , \20141 , \19863 );
and \U$19766 ( \20143 , \20139 , \20142 );
and \U$19767 ( \20144 , \20134 , \20142 );
or \U$19768 ( \20145 , \20140 , \20143 , \20144 );
xor \U$19769 ( \20146 , \20018 , \20020 );
xor \U$19770 ( \20147 , \20146 , \20023 );
and \U$19771 ( \20148 , \20145 , \20147 );
and \U$19772 ( \20149 , \20037 , \20148 );
xor \U$19773 ( \20150 , \20037 , \20148 );
xor \U$19774 ( \20151 , \20145 , \20147 );
xor \U$19775 ( \20152 , \20134 , \20139 );
xor \U$19776 ( \20153 , \20152 , \20142 );
xor \U$19777 ( \20154 , \20002 , \20012 );
xor \U$19778 ( \20155 , \20154 , \20015 );
and \U$19779 ( \20156 , \20153 , \20155 );
and \U$19780 ( \20157 , \20151 , \20156 );
xor \U$19781 ( \20158 , \20151 , \20156 );
xor \U$19782 ( \20159 , \20153 , \20155 );
and \U$19783 ( \20160 , \5315 , \10876 );
and \U$19784 ( \20161 , \5310 , \10873 );
nor \U$19785 ( \20162 , \20160 , \20161 );
xnor \U$19786 ( \20163 , \20162 , \9821 );
and \U$19787 ( \20164 , \5838 , \10063 );
and \U$19788 ( \20165 , \5579 , \10061 );
nor \U$19789 ( \20166 , \20164 , \20165 );
xnor \U$19790 ( \20167 , \20166 , \9824 );
and \U$19791 ( \20168 , \20163 , \20167 );
and \U$19792 ( \20169 , \6219 , \9495 );
and \U$19793 ( \20170 , \6210 , \9493 );
nor \U$19794 ( \20171 , \20169 , \20170 );
xnor \U$19795 ( \20172 , \20171 , \9185 );
and \U$19796 ( \20173 , \20167 , \20172 );
and \U$19797 ( \20174 , \20163 , \20172 );
or \U$19798 ( \20175 , \20168 , \20173 , \20174 );
and \U$19799 ( \20176 , \8440 , \7300 );
and \U$19800 ( \20177 , \8435 , \7298 );
nor \U$19801 ( \20178 , \20176 , \20177 );
xnor \U$19802 ( \20179 , \20178 , \7040 );
and \U$19803 ( \20180 , \9043 , \6806 );
and \U$19804 ( \20181 , \8759 , \6804 );
nor \U$19805 ( \20182 , \20180 , \20181 );
xnor \U$19806 ( \20183 , \20182 , \6491 );
and \U$19807 ( \20184 , \20179 , \20183 );
and \U$19808 ( \20185 , \9620 , \6297 );
and \U$19809 ( \20186 , \9612 , \6295 );
nor \U$19810 ( \20187 , \20185 , \20186 );
xnor \U$19811 ( \20188 , \20187 , \5957 );
and \U$19812 ( \20189 , \20183 , \20188 );
and \U$19813 ( \20190 , \20179 , \20188 );
or \U$19814 ( \20191 , \20184 , \20189 , \20190 );
and \U$19815 ( \20192 , \20175 , \20191 );
and \U$19816 ( \20193 , \6764 , \8958 );
and \U$19817 ( \20194 , \6562 , \8956 );
nor \U$19818 ( \20195 , \20193 , \20194 );
xnor \U$19819 ( \20196 , \20195 , \8587 );
and \U$19820 ( \20197 , \7239 , \8396 );
and \U$19821 ( \20198 , \7067 , \8394 );
nor \U$19822 ( \20199 , \20197 , \20198 );
xnor \U$19823 ( \20200 , \20199 , \8078 );
and \U$19824 ( \20201 , \20196 , \20200 );
and \U$19825 ( \20202 , \8189 , \7829 );
and \U$19826 ( \20203 , \7765 , \7827 );
nor \U$19827 ( \20204 , \20202 , \20203 );
xnor \U$19828 ( \20205 , \20204 , \7580 );
and \U$19829 ( \20206 , \20200 , \20205 );
and \U$19830 ( \20207 , \20196 , \20205 );
or \U$19831 ( \20208 , \20201 , \20206 , \20207 );
and \U$19832 ( \20209 , \20191 , \20208 );
and \U$19833 ( \20210 , \20175 , \20208 );
or \U$19834 ( \20211 , \20192 , \20209 , \20210 );
nand \U$19835 ( \20212 , \11029 , \4866 );
xnor \U$19836 ( \20213 , \20212 , \4636 );
xor \U$19837 ( \20214 , \20057 , \20061 );
xor \U$19838 ( \20215 , \20214 , \20066 );
and \U$19839 ( \20216 , \20213 , \20215 );
xor \U$19840 ( \20217 , \20089 , \20093 );
xor \U$19841 ( \20218 , \20217 , \20098 );
and \U$19842 ( \20219 , \20215 , \20218 );
and \U$19843 ( \20220 , \20213 , \20218 );
or \U$19844 ( \20221 , \20216 , \20219 , \20220 );
and \U$19845 ( \20222 , \20211 , \20221 );
xor \U$19846 ( \20223 , \20041 , \20045 );
xor \U$19847 ( \20224 , \20223 , \20050 );
xor \U$19848 ( \20225 , \20074 , \20078 );
xor \U$19849 ( \20226 , \20225 , \4636 );
and \U$19850 ( \20227 , \20224 , \20226 );
and \U$19851 ( \20228 , \20221 , \20227 );
and \U$19852 ( \20229 , \20211 , \20227 );
or \U$19853 ( \20230 , \20222 , \20228 , \20229 );
xor \U$19854 ( \20231 , \20053 , \20069 );
xor \U$19855 ( \20232 , \20231 , \20082 );
xor \U$19856 ( \20233 , \20101 , \20103 );
xor \U$19857 ( \20234 , \20233 , \20106 );
and \U$19858 ( \20235 , \20232 , \20234 );
xor \U$19859 ( \20236 , \20112 , \20114 );
and \U$19860 ( \20237 , \20234 , \20236 );
and \U$19861 ( \20238 , \20232 , \20236 );
or \U$19862 ( \20239 , \20235 , \20237 , \20238 );
and \U$19863 ( \20240 , \20230 , \20239 );
xor \U$19864 ( \20241 , \20120 , \20122 );
xor \U$19865 ( \20242 , \20241 , \20125 );
and \U$19866 ( \20243 , \20239 , \20242 );
and \U$19867 ( \20244 , \20230 , \20242 );
or \U$19868 ( \20245 , \20240 , \20243 , \20244 );
xor \U$19869 ( \20246 , \20118 , \20128 );
xor \U$19870 ( \20247 , \20246 , \20131 );
and \U$19871 ( \20248 , \20245 , \20247 );
xor \U$19872 ( \20249 , \20136 , \20138 );
and \U$19873 ( \20250 , \20247 , \20249 );
and \U$19874 ( \20251 , \20245 , \20249 );
or \U$19875 ( \20252 , \20248 , \20250 , \20251 );
and \U$19876 ( \20253 , \20159 , \20252 );
xor \U$19877 ( \20254 , \20159 , \20252 );
xor \U$19878 ( \20255 , \20245 , \20247 );
xor \U$19879 ( \20256 , \20255 , \20249 );
and \U$19880 ( \20257 , \10223 , \6297 );
and \U$19881 ( \20258 , \9620 , \6295 );
nor \U$19882 ( \20259 , \20257 , \20258 );
xnor \U$19883 ( \20260 , \20259 , \5957 );
and \U$19884 ( \20261 , \10409 , \5708 );
and \U$19885 ( \20262 , \10228 , \5706 );
nor \U$19886 ( \20263 , \20261 , \20262 );
xnor \U$19887 ( \20264 , \20263 , \5467 );
and \U$19888 ( \20265 , \20260 , \20264 );
nand \U$19889 ( \20266 , \11029 , \5240 );
xnor \U$19890 ( \20267 , \20266 , \5054 );
and \U$19891 ( \20268 , \20264 , \20267 );
and \U$19892 ( \20269 , \20260 , \20267 );
or \U$19893 ( \20270 , \20265 , \20268 , \20269 );
and \U$19894 ( \20271 , \10228 , \5708 );
and \U$19895 ( \20272 , \10223 , \5706 );
nor \U$19896 ( \20273 , \20271 , \20272 );
xnor \U$19897 ( \20274 , \20273 , \5467 );
and \U$19898 ( \20275 , \20270 , \20274 );
and \U$19899 ( \20276 , \11029 , \5242 );
and \U$19900 ( \20277 , \10409 , \5240 );
nor \U$19901 ( \20278 , \20276 , \20277 );
xnor \U$19902 ( \20279 , \20278 , \5054 );
and \U$19903 ( \20280 , \20274 , \20279 );
and \U$19904 ( \20281 , \20270 , \20279 );
or \U$19905 ( \20282 , \20275 , \20280 , \20281 );
and \U$19906 ( \20283 , \5579 , \10876 );
and \U$19907 ( \20284 , \5315 , \10873 );
nor \U$19908 ( \20285 , \20283 , \20284 );
xnor \U$19909 ( \20286 , \20285 , \9821 );
and \U$19910 ( \20287 , \6210 , \10063 );
and \U$19911 ( \20288 , \5838 , \10061 );
nor \U$19912 ( \20289 , \20287 , \20288 );
xnor \U$19913 ( \20290 , \20289 , \9824 );
and \U$19914 ( \20291 , \20286 , \20290 );
and \U$19915 ( \20292 , \20290 , \5054 );
and \U$19916 ( \20293 , \20286 , \5054 );
or \U$19917 ( \20294 , \20291 , \20292 , \20293 );
and \U$19918 ( \20295 , \6562 , \9495 );
and \U$19919 ( \20296 , \6219 , \9493 );
nor \U$19920 ( \20297 , \20295 , \20296 );
xnor \U$19921 ( \20298 , \20297 , \9185 );
and \U$19922 ( \20299 , \7067 , \8958 );
and \U$19923 ( \20300 , \6764 , \8956 );
nor \U$19924 ( \20301 , \20299 , \20300 );
xnor \U$19925 ( \20302 , \20301 , \8587 );
and \U$19926 ( \20303 , \20298 , \20302 );
and \U$19927 ( \20304 , \7765 , \8396 );
and \U$19928 ( \20305 , \7239 , \8394 );
nor \U$19929 ( \20306 , \20304 , \20305 );
xnor \U$19930 ( \20307 , \20306 , \8078 );
and \U$19931 ( \20308 , \20302 , \20307 );
and \U$19932 ( \20309 , \20298 , \20307 );
or \U$19933 ( \20310 , \20303 , \20308 , \20309 );
and \U$19934 ( \20311 , \20294 , \20310 );
and \U$19935 ( \20312 , \8435 , \7829 );
and \U$19936 ( \20313 , \8189 , \7827 );
nor \U$19937 ( \20314 , \20312 , \20313 );
xnor \U$19938 ( \20315 , \20314 , \7580 );
and \U$19939 ( \20316 , \8759 , \7300 );
and \U$19940 ( \20317 , \8440 , \7298 );
nor \U$19941 ( \20318 , \20316 , \20317 );
xnor \U$19942 ( \20319 , \20318 , \7040 );
and \U$19943 ( \20320 , \20315 , \20319 );
and \U$19944 ( \20321 , \9612 , \6806 );
and \U$19945 ( \20322 , \9043 , \6804 );
nor \U$19946 ( \20323 , \20321 , \20322 );
xnor \U$19947 ( \20324 , \20323 , \6491 );
and \U$19948 ( \20325 , \20319 , \20324 );
and \U$19949 ( \20326 , \20315 , \20324 );
or \U$19950 ( \20327 , \20320 , \20325 , \20326 );
and \U$19951 ( \20328 , \20310 , \20327 );
and \U$19952 ( \20329 , \20294 , \20327 );
or \U$19953 ( \20330 , \20311 , \20328 , \20329 );
and \U$19954 ( \20331 , \20282 , \20330 );
xor \U$19955 ( \20332 , \20163 , \20167 );
xor \U$19956 ( \20333 , \20332 , \20172 );
xor \U$19957 ( \20334 , \20179 , \20183 );
xor \U$19958 ( \20335 , \20334 , \20188 );
and \U$19959 ( \20336 , \20333 , \20335 );
xor \U$19960 ( \20337 , \20196 , \20200 );
xor \U$19961 ( \20338 , \20337 , \20205 );
and \U$19962 ( \20339 , \20335 , \20338 );
and \U$19963 ( \20340 , \20333 , \20338 );
or \U$19964 ( \20341 , \20336 , \20339 , \20340 );
and \U$19965 ( \20342 , \20330 , \20341 );
and \U$19966 ( \20343 , \20282 , \20341 );
or \U$19967 ( \20344 , \20331 , \20342 , \20343 );
xor \U$19968 ( \20345 , \20175 , \20191 );
xor \U$19969 ( \20346 , \20345 , \20208 );
xor \U$19970 ( \20347 , \20213 , \20215 );
xor \U$19971 ( \20348 , \20347 , \20218 );
and \U$19972 ( \20349 , \20346 , \20348 );
xor \U$19973 ( \20350 , \20224 , \20226 );
and \U$19974 ( \20351 , \20348 , \20350 );
and \U$19975 ( \20352 , \20346 , \20350 );
or \U$19976 ( \20353 , \20349 , \20351 , \20352 );
and \U$19977 ( \20354 , \20344 , \20353 );
xor \U$19978 ( \20355 , \20232 , \20234 );
xor \U$19979 ( \20356 , \20355 , \20236 );
and \U$19980 ( \20357 , \20353 , \20356 );
and \U$19981 ( \20358 , \20344 , \20356 );
or \U$19982 ( \20359 , \20354 , \20357 , \20358 );
xor \U$19983 ( \20360 , \20085 , \20109 );
xor \U$19984 ( \20361 , \20360 , \20115 );
and \U$19985 ( \20362 , \20359 , \20361 );
xor \U$19986 ( \20363 , \20230 , \20239 );
xor \U$19987 ( \20364 , \20363 , \20242 );
and \U$19988 ( \20365 , \20361 , \20364 );
and \U$19989 ( \20366 , \20359 , \20364 );
or \U$19990 ( \20367 , \20362 , \20365 , \20366 );
and \U$19991 ( \20368 , \20256 , \20367 );
xor \U$19992 ( \20369 , \20256 , \20367 );
xor \U$19993 ( \20370 , \20359 , \20361 );
xor \U$19994 ( \20371 , \20370 , \20364 );
and \U$19995 ( \20372 , \9043 , \7300 );
and \U$19996 ( \20373 , \8759 , \7298 );
nor \U$19997 ( \20374 , \20372 , \20373 );
xnor \U$19998 ( \20375 , \20374 , \7040 );
and \U$19999 ( \20376 , \9620 , \6806 );
and \U$20000 ( \20377 , \9612 , \6804 );
nor \U$20001 ( \20378 , \20376 , \20377 );
xnor \U$20002 ( \20379 , \20378 , \6491 );
and \U$20003 ( \20380 , \20375 , \20379 );
and \U$20004 ( \20381 , \10228 , \6297 );
and \U$20005 ( \20382 , \10223 , \6295 );
nor \U$20006 ( \20383 , \20381 , \20382 );
xnor \U$20007 ( \20384 , \20383 , \5957 );
and \U$20008 ( \20385 , \20379 , \20384 );
and \U$20009 ( \20386 , \20375 , \20384 );
or \U$20010 ( \20387 , \20380 , \20385 , \20386 );
and \U$20011 ( \20388 , \5838 , \10876 );
and \U$20012 ( \20389 , \5579 , \10873 );
nor \U$20013 ( \20390 , \20388 , \20389 );
xnor \U$20014 ( \20391 , \20390 , \9821 );
and \U$20015 ( \20392 , \6219 , \10063 );
and \U$20016 ( \20393 , \6210 , \10061 );
nor \U$20017 ( \20394 , \20392 , \20393 );
xnor \U$20018 ( \20395 , \20394 , \9824 );
and \U$20019 ( \20396 , \20391 , \20395 );
and \U$20020 ( \20397 , \6764 , \9495 );
and \U$20021 ( \20398 , \6562 , \9493 );
nor \U$20022 ( \20399 , \20397 , \20398 );
xnor \U$20023 ( \20400 , \20399 , \9185 );
and \U$20024 ( \20401 , \20395 , \20400 );
and \U$20025 ( \20402 , \20391 , \20400 );
or \U$20026 ( \20403 , \20396 , \20401 , \20402 );
and \U$20027 ( \20404 , \20387 , \20403 );
and \U$20028 ( \20405 , \7239 , \8958 );
and \U$20029 ( \20406 , \7067 , \8956 );
nor \U$20030 ( \20407 , \20405 , \20406 );
xnor \U$20031 ( \20408 , \20407 , \8587 );
and \U$20032 ( \20409 , \8189 , \8396 );
and \U$20033 ( \20410 , \7765 , \8394 );
nor \U$20034 ( \20411 , \20409 , \20410 );
xnor \U$20035 ( \20412 , \20411 , \8078 );
and \U$20036 ( \20413 , \20408 , \20412 );
and \U$20037 ( \20414 , \8440 , \7829 );
and \U$20038 ( \20415 , \8435 , \7827 );
nor \U$20039 ( \20416 , \20414 , \20415 );
xnor \U$20040 ( \20417 , \20416 , \7580 );
and \U$20041 ( \20418 , \20412 , \20417 );
and \U$20042 ( \20419 , \20408 , \20417 );
or \U$20043 ( \20420 , \20413 , \20418 , \20419 );
and \U$20044 ( \20421 , \20403 , \20420 );
and \U$20045 ( \20422 , \20387 , \20420 );
or \U$20046 ( \20423 , \20404 , \20421 , \20422 );
xor \U$20047 ( \20424 , \20298 , \20302 );
xor \U$20048 ( \20425 , \20424 , \20307 );
xor \U$20049 ( \20426 , \20260 , \20264 );
xor \U$20050 ( \20427 , \20426 , \20267 );
and \U$20051 ( \20428 , \20425 , \20427 );
xor \U$20052 ( \20429 , \20315 , \20319 );
xor \U$20053 ( \20430 , \20429 , \20324 );
and \U$20054 ( \20431 , \20427 , \20430 );
and \U$20055 ( \20432 , \20425 , \20430 );
or \U$20056 ( \20433 , \20428 , \20431 , \20432 );
and \U$20057 ( \20434 , \20423 , \20433 );
xor \U$20058 ( \20435 , \20333 , \20335 );
xor \U$20059 ( \20436 , \20435 , \20338 );
and \U$20060 ( \20437 , \20433 , \20436 );
and \U$20061 ( \20438 , \20423 , \20436 );
or \U$20062 ( \20439 , \20434 , \20437 , \20438 );
xor \U$20063 ( \20440 , \20282 , \20330 );
xor \U$20064 ( \20441 , \20440 , \20341 );
and \U$20065 ( \20442 , \20439 , \20441 );
xor \U$20066 ( \20443 , \20346 , \20348 );
xor \U$20067 ( \20444 , \20443 , \20350 );
and \U$20068 ( \20445 , \20441 , \20444 );
and \U$20069 ( \20446 , \20439 , \20444 );
or \U$20070 ( \20447 , \20442 , \20445 , \20446 );
xor \U$20071 ( \20448 , \20211 , \20221 );
xor \U$20072 ( \20449 , \20448 , \20227 );
and \U$20073 ( \20450 , \20447 , \20449 );
xor \U$20074 ( \20451 , \20344 , \20353 );
xor \U$20075 ( \20452 , \20451 , \20356 );
and \U$20076 ( \20453 , \20449 , \20452 );
and \U$20077 ( \20454 , \20447 , \20452 );
or \U$20078 ( \20455 , \20450 , \20453 , \20454 );
and \U$20079 ( \20456 , \20371 , \20455 );
xor \U$20080 ( \20457 , \20371 , \20455 );
xor \U$20081 ( \20458 , \20447 , \20449 );
xor \U$20082 ( \20459 , \20458 , \20452 );
and \U$20083 ( \20460 , \6210 , \10876 );
and \U$20084 ( \20461 , \5838 , \10873 );
nor \U$20085 ( \20462 , \20460 , \20461 );
xnor \U$20086 ( \20463 , \20462 , \9821 );
and \U$20087 ( \20464 , \6562 , \10063 );
and \U$20088 ( \20465 , \6219 , \10061 );
nor \U$20089 ( \20466 , \20464 , \20465 );
xnor \U$20090 ( \20467 , \20466 , \9824 );
and \U$20091 ( \20468 , \20463 , \20467 );
and \U$20092 ( \20469 , \20467 , \5467 );
and \U$20093 ( \20470 , \20463 , \5467 );
or \U$20094 ( \20471 , \20468 , \20469 , \20470 );
and \U$20095 ( \20472 , \8759 , \7829 );
and \U$20096 ( \20473 , \8440 , \7827 );
nor \U$20097 ( \20474 , \20472 , \20473 );
xnor \U$20098 ( \20475 , \20474 , \7580 );
and \U$20099 ( \20476 , \9612 , \7300 );
and \U$20100 ( \20477 , \9043 , \7298 );
nor \U$20101 ( \20478 , \20476 , \20477 );
xnor \U$20102 ( \20479 , \20478 , \7040 );
and \U$20103 ( \20480 , \20475 , \20479 );
and \U$20104 ( \20481 , \10223 , \6806 );
and \U$20105 ( \20482 , \9620 , \6804 );
nor \U$20106 ( \20483 , \20481 , \20482 );
xnor \U$20107 ( \20484 , \20483 , \6491 );
and \U$20108 ( \20485 , \20479 , \20484 );
and \U$20109 ( \20486 , \20475 , \20484 );
or \U$20110 ( \20487 , \20480 , \20485 , \20486 );
and \U$20111 ( \20488 , \20471 , \20487 );
and \U$20112 ( \20489 , \7067 , \9495 );
and \U$20113 ( \20490 , \6764 , \9493 );
nor \U$20114 ( \20491 , \20489 , \20490 );
xnor \U$20115 ( \20492 , \20491 , \9185 );
and \U$20116 ( \20493 , \7765 , \8958 );
and \U$20117 ( \20494 , \7239 , \8956 );
nor \U$20118 ( \20495 , \20493 , \20494 );
xnor \U$20119 ( \20496 , \20495 , \8587 );
and \U$20120 ( \20497 , \20492 , \20496 );
and \U$20121 ( \20498 , \8435 , \8396 );
and \U$20122 ( \20499 , \8189 , \8394 );
nor \U$20123 ( \20500 , \20498 , \20499 );
xnor \U$20124 ( \20501 , \20500 , \8078 );
and \U$20125 ( \20502 , \20496 , \20501 );
and \U$20126 ( \20503 , \20492 , \20501 );
or \U$20127 ( \20504 , \20497 , \20502 , \20503 );
and \U$20128 ( \20505 , \20487 , \20504 );
and \U$20129 ( \20506 , \20471 , \20504 );
or \U$20130 ( \20507 , \20488 , \20505 , \20506 );
and \U$20131 ( \20508 , \11029 , \5708 );
and \U$20132 ( \20509 , \10409 , \5706 );
nor \U$20133 ( \20510 , \20508 , \20509 );
xnor \U$20134 ( \20511 , \20510 , \5467 );
xor \U$20135 ( \20512 , \20375 , \20379 );
xor \U$20136 ( \20513 , \20512 , \20384 );
and \U$20137 ( \20514 , \20511 , \20513 );
xor \U$20138 ( \20515 , \20408 , \20412 );
xor \U$20139 ( \20516 , \20515 , \20417 );
and \U$20140 ( \20517 , \20513 , \20516 );
and \U$20141 ( \20518 , \20511 , \20516 );
or \U$20142 ( \20519 , \20514 , \20517 , \20518 );
and \U$20143 ( \20520 , \20507 , \20519 );
xor \U$20144 ( \20521 , \20286 , \20290 );
xor \U$20145 ( \20522 , \20521 , \5054 );
and \U$20146 ( \20523 , \20519 , \20522 );
and \U$20147 ( \20524 , \20507 , \20522 );
or \U$20148 ( \20525 , \20520 , \20523 , \20524 );
xor \U$20149 ( \20526 , \20387 , \20403 );
xor \U$20150 ( \20527 , \20526 , \20420 );
xor \U$20151 ( \20528 , \20425 , \20427 );
xor \U$20152 ( \20529 , \20528 , \20430 );
and \U$20153 ( \20530 , \20527 , \20529 );
and \U$20154 ( \20531 , \20525 , \20530 );
xor \U$20155 ( \20532 , \20270 , \20274 );
xor \U$20156 ( \20533 , \20532 , \20279 );
and \U$20157 ( \20534 , \20530 , \20533 );
and \U$20158 ( \20535 , \20525 , \20533 );
or \U$20159 ( \20536 , \20531 , \20534 , \20535 );
xor \U$20160 ( \20537 , \20294 , \20310 );
xor \U$20161 ( \20538 , \20537 , \20327 );
xor \U$20162 ( \20539 , \20423 , \20433 );
xor \U$20163 ( \20540 , \20539 , \20436 );
and \U$20164 ( \20541 , \20538 , \20540 );
and \U$20165 ( \20542 , \20536 , \20541 );
xor \U$20166 ( \20543 , \20439 , \20441 );
xor \U$20167 ( \20544 , \20543 , \20444 );
and \U$20168 ( \20545 , \20541 , \20544 );
and \U$20169 ( \20546 , \20536 , \20544 );
or \U$20170 ( \20547 , \20542 , \20545 , \20546 );
and \U$20171 ( \20548 , \20459 , \20547 );
xor \U$20172 ( \20549 , \20459 , \20547 );
xor \U$20173 ( \20550 , \20536 , \20541 );
xor \U$20174 ( \20551 , \20550 , \20544 );
and \U$20175 ( \20552 , \8189 , \8958 );
and \U$20176 ( \20553 , \7765 , \8956 );
nor \U$20177 ( \20554 , \20552 , \20553 );
xnor \U$20178 ( \20555 , \20554 , \8587 );
and \U$20179 ( \20556 , \8440 , \8396 );
and \U$20180 ( \20557 , \8435 , \8394 );
nor \U$20181 ( \20558 , \20556 , \20557 );
xnor \U$20182 ( \20559 , \20558 , \8078 );
and \U$20183 ( \20560 , \20555 , \20559 );
and \U$20184 ( \20561 , \9043 , \7829 );
and \U$20185 ( \20562 , \8759 , \7827 );
nor \U$20186 ( \20563 , \20561 , \20562 );
xnor \U$20187 ( \20564 , \20563 , \7580 );
and \U$20188 ( \20565 , \20559 , \20564 );
and \U$20189 ( \20566 , \20555 , \20564 );
or \U$20190 ( \20567 , \20560 , \20565 , \20566 );
and \U$20191 ( \20568 , \6219 , \10876 );
and \U$20192 ( \20569 , \6210 , \10873 );
nor \U$20193 ( \20570 , \20568 , \20569 );
xnor \U$20194 ( \20571 , \20570 , \9821 );
and \U$20195 ( \20572 , \6764 , \10063 );
and \U$20196 ( \20573 , \6562 , \10061 );
nor \U$20197 ( \20574 , \20572 , \20573 );
xnor \U$20198 ( \20575 , \20574 , \9824 );
and \U$20199 ( \20576 , \20571 , \20575 );
and \U$20200 ( \20577 , \7239 , \9495 );
and \U$20201 ( \20578 , \7067 , \9493 );
nor \U$20202 ( \20579 , \20577 , \20578 );
xnor \U$20203 ( \20580 , \20579 , \9185 );
and \U$20204 ( \20581 , \20575 , \20580 );
and \U$20205 ( \20582 , \20571 , \20580 );
or \U$20206 ( \20583 , \20576 , \20581 , \20582 );
and \U$20207 ( \20584 , \20567 , \20583 );
and \U$20208 ( \20585 , \9620 , \7300 );
and \U$20209 ( \20586 , \9612 , \7298 );
nor \U$20210 ( \20587 , \20585 , \20586 );
xnor \U$20211 ( \20588 , \20587 , \7040 );
and \U$20212 ( \20589 , \10228 , \6806 );
and \U$20213 ( \20590 , \10223 , \6804 );
nor \U$20214 ( \20591 , \20589 , \20590 );
xnor \U$20215 ( \20592 , \20591 , \6491 );
and \U$20216 ( \20593 , \20588 , \20592 );
and \U$20217 ( \20594 , \11029 , \6297 );
and \U$20218 ( \20595 , \10409 , \6295 );
nor \U$20219 ( \20596 , \20594 , \20595 );
xnor \U$20220 ( \20597 , \20596 , \5957 );
and \U$20221 ( \20598 , \20592 , \20597 );
and \U$20222 ( \20599 , \20588 , \20597 );
or \U$20223 ( \20600 , \20593 , \20598 , \20599 );
and \U$20224 ( \20601 , \20583 , \20600 );
and \U$20225 ( \20602 , \20567 , \20600 );
or \U$20226 ( \20603 , \20584 , \20601 , \20602 );
and \U$20227 ( \20604 , \10409 , \6297 );
and \U$20228 ( \20605 , \10228 , \6295 );
nor \U$20229 ( \20606 , \20604 , \20605 );
xnor \U$20230 ( \20607 , \20606 , \5957 );
nand \U$20231 ( \20608 , \11029 , \5706 );
xnor \U$20232 ( \20609 , \20608 , \5467 );
and \U$20233 ( \20610 , \20607 , \20609 );
xor \U$20234 ( \20611 , \20475 , \20479 );
xor \U$20235 ( \20612 , \20611 , \20484 );
and \U$20236 ( \20613 , \20609 , \20612 );
and \U$20237 ( \20614 , \20607 , \20612 );
or \U$20238 ( \20615 , \20610 , \20613 , \20614 );
and \U$20239 ( \20616 , \20603 , \20615 );
xor \U$20240 ( \20617 , \20391 , \20395 );
xor \U$20241 ( \20618 , \20617 , \20400 );
and \U$20242 ( \20619 , \20615 , \20618 );
and \U$20243 ( \20620 , \20603 , \20618 );
or \U$20244 ( \20621 , \20616 , \20619 , \20620 );
xor \U$20245 ( \20622 , \20507 , \20519 );
xor \U$20246 ( \20623 , \20622 , \20522 );
and \U$20247 ( \20624 , \20621 , \20623 );
xor \U$20248 ( \20625 , \20527 , \20529 );
and \U$20249 ( \20626 , \20623 , \20625 );
and \U$20250 ( \20627 , \20621 , \20625 );
or \U$20251 ( \20628 , \20624 , \20626 , \20627 );
xor \U$20252 ( \20629 , \20525 , \20530 );
xor \U$20253 ( \20630 , \20629 , \20533 );
and \U$20254 ( \20631 , \20628 , \20630 );
xor \U$20255 ( \20632 , \20538 , \20540 );
and \U$20256 ( \20633 , \20630 , \20632 );
and \U$20257 ( \20634 , \20628 , \20632 );
or \U$20258 ( \20635 , \20631 , \20633 , \20634 );
and \U$20259 ( \20636 , \20551 , \20635 );
xor \U$20260 ( \20637 , \20551 , \20635 );
xor \U$20261 ( \20638 , \20628 , \20630 );
xor \U$20262 ( \20639 , \20638 , \20632 );
and \U$20263 ( \20640 , \7765 , \9495 );
and \U$20264 ( \20641 , \7239 , \9493 );
nor \U$20265 ( \20642 , \20640 , \20641 );
xnor \U$20266 ( \20643 , \20642 , \9185 );
and \U$20267 ( \20644 , \8435 , \8958 );
and \U$20268 ( \20645 , \8189 , \8956 );
nor \U$20269 ( \20646 , \20644 , \20645 );
xnor \U$20270 ( \20647 , \20646 , \8587 );
and \U$20271 ( \20648 , \20643 , \20647 );
and \U$20272 ( \20649 , \8759 , \8396 );
and \U$20273 ( \20650 , \8440 , \8394 );
nor \U$20274 ( \20651 , \20649 , \20650 );
xnor \U$20275 ( \20652 , \20651 , \8078 );
and \U$20276 ( \20653 , \20647 , \20652 );
and \U$20277 ( \20654 , \20643 , \20652 );
or \U$20278 ( \20655 , \20648 , \20653 , \20654 );
and \U$20279 ( \20656 , \6562 , \10876 );
and \U$20280 ( \20657 , \6219 , \10873 );
nor \U$20281 ( \20658 , \20656 , \20657 );
xnor \U$20282 ( \20659 , \20658 , \9821 );
and \U$20283 ( \20660 , \7067 , \10063 );
and \U$20284 ( \20661 , \6764 , \10061 );
nor \U$20285 ( \20662 , \20660 , \20661 );
xnor \U$20286 ( \20663 , \20662 , \9824 );
and \U$20287 ( \20664 , \20659 , \20663 );
and \U$20288 ( \20665 , \20663 , \5957 );
and \U$20289 ( \20666 , \20659 , \5957 );
or \U$20290 ( \20667 , \20664 , \20665 , \20666 );
and \U$20291 ( \20668 , \20655 , \20667 );
and \U$20292 ( \20669 , \9612 , \7829 );
and \U$20293 ( \20670 , \9043 , \7827 );
nor \U$20294 ( \20671 , \20669 , \20670 );
xnor \U$20295 ( \20672 , \20671 , \7580 );
and \U$20296 ( \20673 , \10223 , \7300 );
and \U$20297 ( \20674 , \9620 , \7298 );
nor \U$20298 ( \20675 , \20673 , \20674 );
xnor \U$20299 ( \20676 , \20675 , \7040 );
and \U$20300 ( \20677 , \20672 , \20676 );
and \U$20301 ( \20678 , \10409 , \6806 );
and \U$20302 ( \20679 , \10228 , \6804 );
nor \U$20303 ( \20680 , \20678 , \20679 );
xnor \U$20304 ( \20681 , \20680 , \6491 );
and \U$20305 ( \20682 , \20676 , \20681 );
and \U$20306 ( \20683 , \20672 , \20681 );
or \U$20307 ( \20684 , \20677 , \20682 , \20683 );
and \U$20308 ( \20685 , \20667 , \20684 );
and \U$20309 ( \20686 , \20655 , \20684 );
or \U$20310 ( \20687 , \20668 , \20685 , \20686 );
xor \U$20311 ( \20688 , \20555 , \20559 );
xor \U$20312 ( \20689 , \20688 , \20564 );
xor \U$20313 ( \20690 , \20571 , \20575 );
xor \U$20314 ( \20691 , \20690 , \20580 );
and \U$20315 ( \20692 , \20689 , \20691 );
xor \U$20316 ( \20693 , \20588 , \20592 );
xor \U$20317 ( \20694 , \20693 , \20597 );
and \U$20318 ( \20695 , \20691 , \20694 );
and \U$20319 ( \20696 , \20689 , \20694 );
or \U$20320 ( \20697 , \20692 , \20695 , \20696 );
and \U$20321 ( \20698 , \20687 , \20697 );
xor \U$20322 ( \20699 , \20492 , \20496 );
xor \U$20323 ( \20700 , \20699 , \20501 );
and \U$20324 ( \20701 , \20697 , \20700 );
and \U$20325 ( \20702 , \20687 , \20700 );
or \U$20326 ( \20703 , \20698 , \20701 , \20702 );
xor \U$20327 ( \20704 , \20463 , \20467 );
xor \U$20328 ( \20705 , \20704 , \5467 );
xor \U$20329 ( \20706 , \20567 , \20583 );
xor \U$20330 ( \20707 , \20706 , \20600 );
and \U$20331 ( \20708 , \20705 , \20707 );
xor \U$20332 ( \20709 , \20607 , \20609 );
xor \U$20333 ( \20710 , \20709 , \20612 );
and \U$20334 ( \20711 , \20707 , \20710 );
and \U$20335 ( \20712 , \20705 , \20710 );
or \U$20336 ( \20713 , \20708 , \20711 , \20712 );
and \U$20337 ( \20714 , \20703 , \20713 );
xor \U$20338 ( \20715 , \20511 , \20513 );
xor \U$20339 ( \20716 , \20715 , \20516 );
and \U$20340 ( \20717 , \20713 , \20716 );
and \U$20341 ( \20718 , \20703 , \20716 );
or \U$20342 ( \20719 , \20714 , \20717 , \20718 );
xor \U$20343 ( \20720 , \20471 , \20487 );
xor \U$20344 ( \20721 , \20720 , \20504 );
xor \U$20345 ( \20722 , \20603 , \20615 );
xor \U$20346 ( \20723 , \20722 , \20618 );
and \U$20347 ( \20724 , \20721 , \20723 );
and \U$20348 ( \20725 , \20719 , \20724 );
xor \U$20349 ( \20726 , \20621 , \20623 );
xor \U$20350 ( \20727 , \20726 , \20625 );
and \U$20351 ( \20728 , \20724 , \20727 );
and \U$20352 ( \20729 , \20719 , \20727 );
or \U$20353 ( \20730 , \20725 , \20728 , \20729 );
and \U$20354 ( \20731 , \20639 , \20730 );
xor \U$20355 ( \20732 , \20639 , \20730 );
xor \U$20356 ( \20733 , \20719 , \20724 );
xor \U$20357 ( \20734 , \20733 , \20727 );
and \U$20358 ( \20735 , \6764 , \10876 );
and \U$20359 ( \20736 , \6562 , \10873 );
nor \U$20360 ( \20737 , \20735 , \20736 );
xnor \U$20361 ( \20738 , \20737 , \9821 );
and \U$20362 ( \20739 , \7239 , \10063 );
and \U$20363 ( \20740 , \7067 , \10061 );
nor \U$20364 ( \20741 , \20739 , \20740 );
xnor \U$20365 ( \20742 , \20741 , \9824 );
and \U$20366 ( \20743 , \20738 , \20742 );
and \U$20367 ( \20744 , \8189 , \9495 );
and \U$20368 ( \20745 , \7765 , \9493 );
nor \U$20369 ( \20746 , \20744 , \20745 );
xnor \U$20370 ( \20747 , \20746 , \9185 );
and \U$20371 ( \20748 , \20742 , \20747 );
and \U$20372 ( \20749 , \20738 , \20747 );
or \U$20373 ( \20750 , \20743 , \20748 , \20749 );
and \U$20374 ( \20751 , \8440 , \8958 );
and \U$20375 ( \20752 , \8435 , \8956 );
nor \U$20376 ( \20753 , \20751 , \20752 );
xnor \U$20377 ( \20754 , \20753 , \8587 );
and \U$20378 ( \20755 , \9043 , \8396 );
and \U$20379 ( \20756 , \8759 , \8394 );
nor \U$20380 ( \20757 , \20755 , \20756 );
xnor \U$20381 ( \20758 , \20757 , \8078 );
and \U$20382 ( \20759 , \20754 , \20758 );
and \U$20383 ( \20760 , \9620 , \7829 );
and \U$20384 ( \20761 , \9612 , \7827 );
nor \U$20385 ( \20762 , \20760 , \20761 );
xnor \U$20386 ( \20763 , \20762 , \7580 );
and \U$20387 ( \20764 , \20758 , \20763 );
and \U$20388 ( \20765 , \20754 , \20763 );
or \U$20389 ( \20766 , \20759 , \20764 , \20765 );
and \U$20390 ( \20767 , \20750 , \20766 );
and \U$20391 ( \20768 , \10228 , \7300 );
and \U$20392 ( \20769 , \10223 , \7298 );
nor \U$20393 ( \20770 , \20768 , \20769 );
xnor \U$20394 ( \20771 , \20770 , \7040 );
and \U$20395 ( \20772 , \11029 , \6806 );
and \U$20396 ( \20773 , \10409 , \6804 );
nor \U$20397 ( \20774 , \20772 , \20773 );
xnor \U$20398 ( \20775 , \20774 , \6491 );
and \U$20399 ( \20776 , \20771 , \20775 );
and \U$20400 ( \20777 , \20766 , \20776 );
and \U$20401 ( \20778 , \20750 , \20776 );
or \U$20402 ( \20779 , \20767 , \20777 , \20778 );
nand \U$20403 ( \20780 , \11029 , \6295 );
xnor \U$20404 ( \20781 , \20780 , \5957 );
xor \U$20405 ( \20782 , \20643 , \20647 );
xor \U$20406 ( \20783 , \20782 , \20652 );
and \U$20407 ( \20784 , \20781 , \20783 );
xor \U$20408 ( \20785 , \20672 , \20676 );
xor \U$20409 ( \20786 , \20785 , \20681 );
and \U$20410 ( \20787 , \20783 , \20786 );
and \U$20411 ( \20788 , \20781 , \20786 );
or \U$20412 ( \20789 , \20784 , \20787 , \20788 );
and \U$20413 ( \20790 , \20779 , \20789 );
xor \U$20414 ( \20791 , \20689 , \20691 );
xor \U$20415 ( \20792 , \20791 , \20694 );
and \U$20416 ( \20793 , \20789 , \20792 );
and \U$20417 ( \20794 , \20779 , \20792 );
or \U$20418 ( \20795 , \20790 , \20793 , \20794 );
xor \U$20419 ( \20796 , \20687 , \20697 );
xor \U$20420 ( \20797 , \20796 , \20700 );
and \U$20421 ( \20798 , \20795 , \20797 );
xor \U$20422 ( \20799 , \20705 , \20707 );
xor \U$20423 ( \20800 , \20799 , \20710 );
and \U$20424 ( \20801 , \20797 , \20800 );
and \U$20425 ( \20802 , \20795 , \20800 );
or \U$20426 ( \20803 , \20798 , \20801 , \20802 );
xor \U$20427 ( \20804 , \20703 , \20713 );
xor \U$20428 ( \20805 , \20804 , \20716 );
and \U$20429 ( \20806 , \20803 , \20805 );
xor \U$20430 ( \20807 , \20721 , \20723 );
and \U$20431 ( \20808 , \20805 , \20807 );
and \U$20432 ( \20809 , \20803 , \20807 );
or \U$20433 ( \20810 , \20806 , \20808 , \20809 );
and \U$20434 ( \20811 , \20734 , \20810 );
xor \U$20435 ( \20812 , \20734 , \20810 );
xor \U$20436 ( \20813 , \20803 , \20805 );
xor \U$20437 ( \20814 , \20813 , \20807 );
and \U$20438 ( \20815 , \10223 , \7829 );
and \U$20439 ( \20816 , \9620 , \7827 );
nor \U$20440 ( \20817 , \20815 , \20816 );
xnor \U$20441 ( \20818 , \20817 , \7580 );
and \U$20442 ( \20819 , \10409 , \7300 );
and \U$20443 ( \20820 , \10228 , \7298 );
nor \U$20444 ( \20821 , \20819 , \20820 );
xnor \U$20445 ( \20822 , \20821 , \7040 );
and \U$20446 ( \20823 , \20818 , \20822 );
nand \U$20447 ( \20824 , \11029 , \6804 );
xnor \U$20448 ( \20825 , \20824 , \6491 );
and \U$20449 ( \20826 , \20822 , \20825 );
and \U$20450 ( \20827 , \20818 , \20825 );
or \U$20451 ( \20828 , \20823 , \20826 , \20827 );
and \U$20452 ( \20829 , \7067 , \10876 );
and \U$20453 ( \20830 , \6764 , \10873 );
nor \U$20454 ( \20831 , \20829 , \20830 );
xnor \U$20455 ( \20832 , \20831 , \9821 );
and \U$20456 ( \20833 , \7765 , \10063 );
and \U$20457 ( \20834 , \7239 , \10061 );
nor \U$20458 ( \20835 , \20833 , \20834 );
xnor \U$20459 ( \20836 , \20835 , \9824 );
and \U$20460 ( \20837 , \20832 , \20836 );
and \U$20461 ( \20838 , \20836 , \6491 );
and \U$20462 ( \20839 , \20832 , \6491 );
or \U$20463 ( \20840 , \20837 , \20838 , \20839 );
and \U$20464 ( \20841 , \20828 , \20840 );
and \U$20465 ( \20842 , \8435 , \9495 );
and \U$20466 ( \20843 , \8189 , \9493 );
nor \U$20467 ( \20844 , \20842 , \20843 );
xnor \U$20468 ( \20845 , \20844 , \9185 );
and \U$20469 ( \20846 , \8759 , \8958 );
and \U$20470 ( \20847 , \8440 , \8956 );
nor \U$20471 ( \20848 , \20846 , \20847 );
xnor \U$20472 ( \20849 , \20848 , \8587 );
and \U$20473 ( \20850 , \20845 , \20849 );
and \U$20474 ( \20851 , \9612 , \8396 );
and \U$20475 ( \20852 , \9043 , \8394 );
nor \U$20476 ( \20853 , \20851 , \20852 );
xnor \U$20477 ( \20854 , \20853 , \8078 );
and \U$20478 ( \20855 , \20849 , \20854 );
and \U$20479 ( \20856 , \20845 , \20854 );
or \U$20480 ( \20857 , \20850 , \20855 , \20856 );
and \U$20481 ( \20858 , \20840 , \20857 );
and \U$20482 ( \20859 , \20828 , \20857 );
or \U$20483 ( \20860 , \20841 , \20858 , \20859 );
xor \U$20484 ( \20861 , \20738 , \20742 );
xor \U$20485 ( \20862 , \20861 , \20747 );
xor \U$20486 ( \20863 , \20754 , \20758 );
xor \U$20487 ( \20864 , \20863 , \20763 );
and \U$20488 ( \20865 , \20862 , \20864 );
xor \U$20489 ( \20866 , \20771 , \20775 );
and \U$20490 ( \20867 , \20864 , \20866 );
and \U$20491 ( \20868 , \20862 , \20866 );
or \U$20492 ( \20869 , \20865 , \20867 , \20868 );
and \U$20493 ( \20870 , \20860 , \20869 );
xor \U$20494 ( \20871 , \20659 , \20663 );
xor \U$20495 ( \20872 , \20871 , \5957 );
and \U$20496 ( \20873 , \20869 , \20872 );
and \U$20497 ( \20874 , \20860 , \20872 );
or \U$20498 ( \20875 , \20870 , \20873 , \20874 );
xor \U$20499 ( \20876 , \20750 , \20766 );
xor \U$20500 ( \20877 , \20876 , \20776 );
xor \U$20501 ( \20878 , \20781 , \20783 );
xor \U$20502 ( \20879 , \20878 , \20786 );
and \U$20503 ( \20880 , \20877 , \20879 );
and \U$20504 ( \20881 , \20875 , \20880 );
xor \U$20505 ( \20882 , \20655 , \20667 );
xor \U$20506 ( \20883 , \20882 , \20684 );
and \U$20507 ( \20884 , \20880 , \20883 );
and \U$20508 ( \20885 , \20875 , \20883 );
or \U$20509 ( \20886 , \20881 , \20884 , \20885 );
xor \U$20510 ( \20887 , \20795 , \20797 );
xor \U$20511 ( \20888 , \20887 , \20800 );
and \U$20512 ( \20889 , \20886 , \20888 );
and \U$20513 ( \20890 , \20814 , \20889 );
xor \U$20514 ( \20891 , \20814 , \20889 );
xor \U$20515 ( \20892 , \20886 , \20888 );
xor \U$20516 ( \20893 , \20875 , \20880 );
xor \U$20517 ( \20894 , \20893 , \20883 );
xor \U$20518 ( \20895 , \20779 , \20789 );
xor \U$20519 ( \20896 , \20895 , \20792 );
and \U$20520 ( \20897 , \20894 , \20896 );
and \U$20521 ( \20898 , \20892 , \20897 );
xor \U$20522 ( \20899 , \20892 , \20897 );
xor \U$20523 ( \20900 , \20894 , \20896 );
and \U$20524 ( \20901 , \7239 , \10876 );
and \U$20525 ( \20902 , \7067 , \10873 );
nor \U$20526 ( \20903 , \20901 , \20902 );
xnor \U$20527 ( \20904 , \20903 , \9821 );
and \U$20528 ( \20905 , \8189 , \10063 );
and \U$20529 ( \20906 , \7765 , \10061 );
nor \U$20530 ( \20907 , \20905 , \20906 );
xnor \U$20531 ( \20908 , \20907 , \9824 );
and \U$20532 ( \20909 , \20904 , \20908 );
and \U$20533 ( \20910 , \8440 , \9495 );
and \U$20534 ( \20911 , \8435 , \9493 );
nor \U$20535 ( \20912 , \20910 , \20911 );
xnor \U$20536 ( \20913 , \20912 , \9185 );
and \U$20537 ( \20914 , \20908 , \20913 );
and \U$20538 ( \20915 , \20904 , \20913 );
or \U$20539 ( \20916 , \20909 , \20914 , \20915 );
and \U$20540 ( \20917 , \9043 , \8958 );
and \U$20541 ( \20918 , \8759 , \8956 );
nor \U$20542 ( \20919 , \20917 , \20918 );
xnor \U$20543 ( \20920 , \20919 , \8587 );
and \U$20544 ( \20921 , \9620 , \8396 );
and \U$20545 ( \20922 , \9612 , \8394 );
nor \U$20546 ( \20923 , \20921 , \20922 );
xnor \U$20547 ( \20924 , \20923 , \8078 );
and \U$20548 ( \20925 , \20920 , \20924 );
and \U$20549 ( \20926 , \10228 , \7829 );
and \U$20550 ( \20927 , \10223 , \7827 );
nor \U$20551 ( \20928 , \20926 , \20927 );
xnor \U$20552 ( \20929 , \20928 , \7580 );
and \U$20553 ( \20930 , \20924 , \20929 );
and \U$20554 ( \20931 , \20920 , \20929 );
or \U$20555 ( \20932 , \20925 , \20930 , \20931 );
and \U$20556 ( \20933 , \20916 , \20932 );
xor \U$20557 ( \20934 , \20818 , \20822 );
xor \U$20558 ( \20935 , \20934 , \20825 );
and \U$20559 ( \20936 , \20932 , \20935 );
and \U$20560 ( \20937 , \20916 , \20935 );
or \U$20561 ( \20938 , \20933 , \20936 , \20937 );
xor \U$20562 ( \20939 , \20832 , \20836 );
xor \U$20563 ( \20940 , \20939 , \6491 );
xor \U$20564 ( \20941 , \20845 , \20849 );
xor \U$20565 ( \20942 , \20941 , \20854 );
and \U$20566 ( \20943 , \20940 , \20942 );
and \U$20567 ( \20944 , \20938 , \20943 );
xor \U$20568 ( \20945 , \20862 , \20864 );
xor \U$20569 ( \20946 , \20945 , \20866 );
and \U$20570 ( \20947 , \20943 , \20946 );
and \U$20571 ( \20948 , \20938 , \20946 );
or \U$20572 ( \20949 , \20944 , \20947 , \20948 );
xor \U$20573 ( \20950 , \20860 , \20869 );
xor \U$20574 ( \20951 , \20950 , \20872 );
and \U$20575 ( \20952 , \20949 , \20951 );
xor \U$20576 ( \20953 , \20877 , \20879 );
and \U$20577 ( \20954 , \20951 , \20953 );
and \U$20578 ( \20955 , \20949 , \20953 );
or \U$20579 ( \20956 , \20952 , \20954 , \20955 );
and \U$20580 ( \20957 , \20900 , \20956 );
xor \U$20581 ( \20958 , \20900 , \20956 );
xor \U$20582 ( \20959 , \20949 , \20951 );
xor \U$20583 ( \20960 , \20959 , \20953 );
and \U$20584 ( \20961 , \7765 , \10876 );
and \U$20585 ( \20962 , \7239 , \10873 );
nor \U$20586 ( \20963 , \20961 , \20962 );
xnor \U$20587 ( \20964 , \20963 , \9821 );
and \U$20588 ( \20965 , \8435 , \10063 );
and \U$20589 ( \20966 , \8189 , \10061 );
nor \U$20590 ( \20967 , \20965 , \20966 );
xnor \U$20591 ( \20968 , \20967 , \9824 );
and \U$20592 ( \20969 , \20964 , \20968 );
and \U$20593 ( \20970 , \20968 , \7040 );
and \U$20594 ( \20971 , \20964 , \7040 );
or \U$20595 ( \20972 , \20969 , \20970 , \20971 );
and \U$20596 ( \20973 , \8759 , \9495 );
and \U$20597 ( \20974 , \8440 , \9493 );
nor \U$20598 ( \20975 , \20973 , \20974 );
xnor \U$20599 ( \20976 , \20975 , \9185 );
and \U$20600 ( \20977 , \9612 , \8958 );
and \U$20601 ( \20978 , \9043 , \8956 );
nor \U$20602 ( \20979 , \20977 , \20978 );
xnor \U$20603 ( \20980 , \20979 , \8587 );
and \U$20604 ( \20981 , \20976 , \20980 );
and \U$20605 ( \20982 , \10223 , \8396 );
and \U$20606 ( \20983 , \9620 , \8394 );
nor \U$20607 ( \20984 , \20982 , \20983 );
xnor \U$20608 ( \20985 , \20984 , \8078 );
and \U$20609 ( \20986 , \20980 , \20985 );
and \U$20610 ( \20987 , \20976 , \20985 );
or \U$20611 ( \20988 , \20981 , \20986 , \20987 );
and \U$20612 ( \20989 , \20972 , \20988 );
and \U$20613 ( \20990 , \11029 , \7300 );
and \U$20614 ( \20991 , \10409 , \7298 );
nor \U$20615 ( \20992 , \20990 , \20991 );
xnor \U$20616 ( \20993 , \20992 , \7040 );
and \U$20617 ( \20994 , \20988 , \20993 );
and \U$20618 ( \20995 , \20972 , \20993 );
or \U$20619 ( \20996 , \20989 , \20994 , \20995 );
xor \U$20620 ( \20997 , \20916 , \20932 );
xor \U$20621 ( \20998 , \20997 , \20935 );
and \U$20622 ( \20999 , \20996 , \20998 );
xor \U$20623 ( \21000 , \20940 , \20942 );
and \U$20624 ( \21001 , \20998 , \21000 );
and \U$20625 ( \21002 , \20996 , \21000 );
or \U$20626 ( \21003 , \20999 , \21001 , \21002 );
xor \U$20627 ( \21004 , \20828 , \20840 );
xor \U$20628 ( \21005 , \21004 , \20857 );
and \U$20629 ( \21006 , \21003 , \21005 );
xor \U$20630 ( \21007 , \20938 , \20943 );
xor \U$20631 ( \21008 , \21007 , \20946 );
and \U$20632 ( \21009 , \21005 , \21008 );
and \U$20633 ( \21010 , \21003 , \21008 );
or \U$20634 ( \21011 , \21006 , \21009 , \21010 );
and \U$20635 ( \21012 , \20960 , \21011 );
xor \U$20636 ( \21013 , \20960 , \21011 );
xor \U$20637 ( \21014 , \21003 , \21005 );
xor \U$20638 ( \21015 , \21014 , \21008 );
and \U$20639 ( \21016 , \9620 , \8958 );
and \U$20640 ( \21017 , \9612 , \8956 );
nor \U$20641 ( \21018 , \21016 , \21017 );
xnor \U$20642 ( \21019 , \21018 , \8587 );
and \U$20643 ( \21020 , \10228 , \8396 );
and \U$20644 ( \21021 , \10223 , \8394 );
nor \U$20645 ( \21022 , \21020 , \21021 );
xnor \U$20646 ( \21023 , \21022 , \8078 );
and \U$20647 ( \21024 , \21019 , \21023 );
and \U$20648 ( \21025 , \11029 , \7829 );
and \U$20649 ( \21026 , \10409 , \7827 );
nor \U$20650 ( \21027 , \21025 , \21026 );
xnor \U$20651 ( \21028 , \21027 , \7580 );
and \U$20652 ( \21029 , \21023 , \21028 );
and \U$20653 ( \21030 , \21019 , \21028 );
or \U$20654 ( \21031 , \21024 , \21029 , \21030 );
and \U$20655 ( \21032 , \8189 , \10876 );
and \U$20656 ( \21033 , \7765 , \10873 );
nor \U$20657 ( \21034 , \21032 , \21033 );
xnor \U$20658 ( \21035 , \21034 , \9821 );
and \U$20659 ( \21036 , \8440 , \10063 );
and \U$20660 ( \21037 , \8435 , \10061 );
nor \U$20661 ( \21038 , \21036 , \21037 );
xnor \U$20662 ( \21039 , \21038 , \9824 );
and \U$20663 ( \21040 , \21035 , \21039 );
and \U$20664 ( \21041 , \9043 , \9495 );
and \U$20665 ( \21042 , \8759 , \9493 );
nor \U$20666 ( \21043 , \21041 , \21042 );
xnor \U$20667 ( \21044 , \21043 , \9185 );
and \U$20668 ( \21045 , \21039 , \21044 );
and \U$20669 ( \21046 , \21035 , \21044 );
or \U$20670 ( \21047 , \21040 , \21045 , \21046 );
and \U$20671 ( \21048 , \21031 , \21047 );
and \U$20672 ( \21049 , \10409 , \7829 );
and \U$20673 ( \21050 , \10228 , \7827 );
nor \U$20674 ( \21051 , \21049 , \21050 );
xnor \U$20675 ( \21052 , \21051 , \7580 );
and \U$20676 ( \21053 , \21047 , \21052 );
and \U$20677 ( \21054 , \21031 , \21052 );
or \U$20678 ( \21055 , \21048 , \21053 , \21054 );
nand \U$20679 ( \21056 , \11029 , \7298 );
xnor \U$20680 ( \21057 , \21056 , \7040 );
xor \U$20681 ( \21058 , \20964 , \20968 );
xor \U$20682 ( \21059 , \21058 , \7040 );
and \U$20683 ( \21060 , \21057 , \21059 );
xor \U$20684 ( \21061 , \20976 , \20980 );
xor \U$20685 ( \21062 , \21061 , \20985 );
and \U$20686 ( \21063 , \21059 , \21062 );
and \U$20687 ( \21064 , \21057 , \21062 );
or \U$20688 ( \21065 , \21060 , \21063 , \21064 );
and \U$20689 ( \21066 , \21055 , \21065 );
xor \U$20690 ( \21067 , \20920 , \20924 );
xor \U$20691 ( \21068 , \21067 , \20929 );
and \U$20692 ( \21069 , \21065 , \21068 );
and \U$20693 ( \21070 , \21055 , \21068 );
or \U$20694 ( \21071 , \21066 , \21069 , \21070 );
xor \U$20695 ( \21072 , \20904 , \20908 );
xor \U$20696 ( \21073 , \21072 , \20913 );
xor \U$20697 ( \21074 , \20972 , \20988 );
xor \U$20698 ( \21075 , \21074 , \20993 );
and \U$20699 ( \21076 , \21073 , \21075 );
and \U$20700 ( \21077 , \21071 , \21076 );
xor \U$20701 ( \21078 , \20996 , \20998 );
xor \U$20702 ( \21079 , \21078 , \21000 );
and \U$20703 ( \21080 , \21076 , \21079 );
and \U$20704 ( \21081 , \21071 , \21079 );
or \U$20705 ( \21082 , \21077 , \21080 , \21081 );
and \U$20706 ( \21083 , \21015 , \21082 );
xor \U$20707 ( \21084 , \21015 , \21082 );
xor \U$20708 ( \21085 , \21071 , \21076 );
xor \U$20709 ( \21086 , \21085 , \21079 );
and \U$20710 ( \21087 , \9612 , \9495 );
and \U$20711 ( \21088 , \9043 , \9493 );
nor \U$20712 ( \21089 , \21087 , \21088 );
xnor \U$20713 ( \21090 , \21089 , \9185 );
and \U$20714 ( \21091 , \10223 , \8958 );
and \U$20715 ( \21092 , \9620 , \8956 );
nor \U$20716 ( \21093 , \21091 , \21092 );
xnor \U$20717 ( \21094 , \21093 , \8587 );
and \U$20718 ( \21095 , \21090 , \21094 );
and \U$20719 ( \21096 , \10409 , \8396 );
and \U$20720 ( \21097 , \10228 , \8394 );
nor \U$20721 ( \21098 , \21096 , \21097 );
xnor \U$20722 ( \21099 , \21098 , \8078 );
and \U$20723 ( \21100 , \21094 , \21099 );
and \U$20724 ( \21101 , \21090 , \21099 );
or \U$20725 ( \21102 , \21095 , \21100 , \21101 );
and \U$20726 ( \21103 , \8435 , \10876 );
and \U$20727 ( \21104 , \8189 , \10873 );
nor \U$20728 ( \21105 , \21103 , \21104 );
xnor \U$20729 ( \21106 , \21105 , \9821 );
and \U$20730 ( \21107 , \8759 , \10063 );
and \U$20731 ( \21108 , \8440 , \10061 );
nor \U$20732 ( \21109 , \21107 , \21108 );
xnor \U$20733 ( \21110 , \21109 , \9824 );
and \U$20734 ( \21111 , \21106 , \21110 );
and \U$20735 ( \21112 , \21110 , \7580 );
and \U$20736 ( \21113 , \21106 , \7580 );
or \U$20737 ( \21114 , \21111 , \21112 , \21113 );
and \U$20738 ( \21115 , \21102 , \21114 );
xor \U$20739 ( \21116 , \21019 , \21023 );
xor \U$20740 ( \21117 , \21116 , \21028 );
and \U$20741 ( \21118 , \21114 , \21117 );
and \U$20742 ( \21119 , \21102 , \21117 );
or \U$20743 ( \21120 , \21115 , \21118 , \21119 );
xor \U$20744 ( \21121 , \21031 , \21047 );
xor \U$20745 ( \21122 , \21121 , \21052 );
and \U$20746 ( \21123 , \21120 , \21122 );
xor \U$20747 ( \21124 , \21057 , \21059 );
xor \U$20748 ( \21125 , \21124 , \21062 );
and \U$20749 ( \21126 , \21122 , \21125 );
and \U$20750 ( \21127 , \21120 , \21125 );
or \U$20751 ( \21128 , \21123 , \21126 , \21127 );
xor \U$20752 ( \21129 , \21055 , \21065 );
xor \U$20753 ( \21130 , \21129 , \21068 );
and \U$20754 ( \21131 , \21128 , \21130 );
xor \U$20755 ( \21132 , \21073 , \21075 );
and \U$20756 ( \21133 , \21130 , \21132 );
and \U$20757 ( \21134 , \21128 , \21132 );
or \U$20758 ( \21135 , \21131 , \21133 , \21134 );
and \U$20759 ( \21136 , \21086 , \21135 );
xor \U$20760 ( \21137 , \21086 , \21135 );
xor \U$20761 ( \21138 , \21128 , \21130 );
xor \U$20762 ( \21139 , \21138 , \21132 );
and \U$20763 ( \21140 , \8440 , \10876 );
and \U$20764 ( \21141 , \8435 , \10873 );
nor \U$20765 ( \21142 , \21140 , \21141 );
xnor \U$20766 ( \21143 , \21142 , \9821 );
and \U$20767 ( \21144 , \9043 , \10063 );
and \U$20768 ( \21145 , \8759 , \10061 );
nor \U$20769 ( \21146 , \21144 , \21145 );
xnor \U$20770 ( \21147 , \21146 , \9824 );
and \U$20771 ( \21148 , \21143 , \21147 );
and \U$20772 ( \21149 , \9620 , \9495 );
and \U$20773 ( \21150 , \9612 , \9493 );
nor \U$20774 ( \21151 , \21149 , \21150 );
xnor \U$20775 ( \21152 , \21151 , \9185 );
and \U$20776 ( \21153 , \21147 , \21152 );
and \U$20777 ( \21154 , \21143 , \21152 );
or \U$20778 ( \21155 , \21148 , \21153 , \21154 );
nand \U$20779 ( \21156 , \11029 , \7827 );
xnor \U$20780 ( \21157 , \21156 , \7580 );
and \U$20781 ( \21158 , \21155 , \21157 );
xor \U$20782 ( \21159 , \21090 , \21094 );
xor \U$20783 ( \21160 , \21159 , \21099 );
and \U$20784 ( \21161 , \21157 , \21160 );
and \U$20785 ( \21162 , \21155 , \21160 );
or \U$20786 ( \21163 , \21158 , \21161 , \21162 );
xor \U$20787 ( \21164 , \21035 , \21039 );
xor \U$20788 ( \21165 , \21164 , \21044 );
and \U$20789 ( \21166 , \21163 , \21165 );
xor \U$20790 ( \21167 , \21102 , \21114 );
xor \U$20791 ( \21168 , \21167 , \21117 );
and \U$20792 ( \21169 , \21165 , \21168 );
and \U$20793 ( \21170 , \21163 , \21168 );
or \U$20794 ( \21171 , \21166 , \21169 , \21170 );
xor \U$20795 ( \21172 , \21120 , \21122 );
xor \U$20796 ( \21173 , \21172 , \21125 );
and \U$20797 ( \21174 , \21171 , \21173 );
and \U$20798 ( \21175 , \21139 , \21174 );
xor \U$20799 ( \21176 , \21139 , \21174 );
xor \U$20800 ( \21177 , \21171 , \21173 );
and \U$20801 ( \21178 , \10223 , \9495 );
and \U$20802 ( \21179 , \9620 , \9493 );
nor \U$20803 ( \21180 , \21178 , \21179 );
xnor \U$20804 ( \21181 , \21180 , \9185 );
and \U$20805 ( \21182 , \10409 , \8958 );
and \U$20806 ( \21183 , \10228 , \8956 );
nor \U$20807 ( \21184 , \21182 , \21183 );
xnor \U$20808 ( \21185 , \21184 , \8587 );
and \U$20809 ( \21186 , \21181 , \21185 );
nand \U$20810 ( \21187 , \11029 , \8394 );
xnor \U$20811 ( \21188 , \21187 , \8078 );
and \U$20812 ( \21189 , \21185 , \21188 );
and \U$20813 ( \21190 , \21181 , \21188 );
or \U$20814 ( \21191 , \21186 , \21189 , \21190 );
and \U$20815 ( \21192 , \8759 , \10876 );
and \U$20816 ( \21193 , \8440 , \10873 );
nor \U$20817 ( \21194 , \21192 , \21193 );
xnor \U$20818 ( \21195 , \21194 , \9821 );
and \U$20819 ( \21196 , \9612 , \10063 );
and \U$20820 ( \21197 , \9043 , \10061 );
nor \U$20821 ( \21198 , \21196 , \21197 );
xnor \U$20822 ( \21199 , \21198 , \9824 );
and \U$20823 ( \21200 , \21195 , \21199 );
and \U$20824 ( \21201 , \21199 , \8078 );
and \U$20825 ( \21202 , \21195 , \8078 );
or \U$20826 ( \21203 , \21200 , \21201 , \21202 );
and \U$20827 ( \21204 , \21191 , \21203 );
and \U$20828 ( \21205 , \10228 , \8958 );
and \U$20829 ( \21206 , \10223 , \8956 );
nor \U$20830 ( \21207 , \21205 , \21206 );
xnor \U$20831 ( \21208 , \21207 , \8587 );
and \U$20832 ( \21209 , \21203 , \21208 );
and \U$20833 ( \21210 , \21191 , \21208 );
or \U$20834 ( \21211 , \21204 , \21209 , \21210 );
and \U$20835 ( \21212 , \11029 , \8396 );
and \U$20836 ( \21213 , \10409 , \8394 );
nor \U$20837 ( \21214 , \21212 , \21213 );
xnor \U$20838 ( \21215 , \21214 , \8078 );
xor \U$20839 ( \21216 , \21143 , \21147 );
xor \U$20840 ( \21217 , \21216 , \21152 );
and \U$20841 ( \21218 , \21215 , \21217 );
and \U$20842 ( \21219 , \21211 , \21218 );
xor \U$20843 ( \21220 , \21106 , \21110 );
xor \U$20844 ( \21221 , \21220 , \7580 );
and \U$20845 ( \21222 , \21218 , \21221 );
and \U$20846 ( \21223 , \21211 , \21221 );
or \U$20847 ( \21224 , \21219 , \21222 , \21223 );
xor \U$20848 ( \21225 , \21163 , \21165 );
xor \U$20849 ( \21226 , \21225 , \21168 );
and \U$20850 ( \21227 , \21224 , \21226 );
and \U$20851 ( \21228 , \21177 , \21227 );
xor \U$20852 ( \21229 , \21177 , \21227 );
xor \U$20853 ( \21230 , \21224 , \21226 );
xor \U$20854 ( \21231 , \21155 , \21157 );
xor \U$20855 ( \21232 , \21231 , \21160 );
xor \U$20856 ( \21233 , \21211 , \21218 );
xor \U$20857 ( \21234 , \21233 , \21221 );
and \U$20858 ( \21235 , \21232 , \21234 );
and \U$20859 ( \21236 , \21230 , \21235 );
xor \U$20860 ( \21237 , \21230 , \21235 );
xor \U$20861 ( \21238 , \21232 , \21234 );
and \U$20862 ( \21239 , \9043 , \10876 );
and \U$20863 ( \21240 , \8759 , \10873 );
nor \U$20864 ( \21241 , \21239 , \21240 );
xnor \U$20865 ( \21242 , \21241 , \9821 );
and \U$20866 ( \21243 , \9620 , \10063 );
and \U$20867 ( \21244 , \9612 , \10061 );
nor \U$20868 ( \21245 , \21243 , \21244 );
xnor \U$20869 ( \21246 , \21245 , \9824 );
and \U$20870 ( \21247 , \21242 , \21246 );
and \U$20871 ( \21248 , \10228 , \9495 );
and \U$20872 ( \21249 , \10223 , \9493 );
nor \U$20873 ( \21250 , \21248 , \21249 );
xnor \U$20874 ( \21251 , \21250 , \9185 );
and \U$20875 ( \21252 , \21246 , \21251 );
and \U$20876 ( \21253 , \21242 , \21251 );
or \U$20877 ( \21254 , \21247 , \21252 , \21253 );
xor \U$20878 ( \21255 , \21181 , \21185 );
xor \U$20879 ( \21256 , \21255 , \21188 );
and \U$20880 ( \21257 , \21254 , \21256 );
xor \U$20881 ( \21258 , \21195 , \21199 );
xor \U$20882 ( \21259 , \21258 , \8078 );
and \U$20883 ( \21260 , \21256 , \21259 );
and \U$20884 ( \21261 , \21254 , \21259 );
or \U$20885 ( \21262 , \21257 , \21260 , \21261 );
xor \U$20886 ( \21263 , \21191 , \21203 );
xor \U$20887 ( \21264 , \21263 , \21208 );
and \U$20888 ( \21265 , \21262 , \21264 );
xor \U$20889 ( \21266 , \21215 , \21217 );
and \U$20890 ( \21267 , \21264 , \21266 );
and \U$20891 ( \21268 , \21262 , \21266 );
or \U$20892 ( \21269 , \21265 , \21267 , \21268 );
and \U$20893 ( \21270 , \21238 , \21269 );
xor \U$20894 ( \21271 , \21238 , \21269 );
xor \U$20895 ( \21272 , \21262 , \21264 );
xor \U$20896 ( \21273 , \21272 , \21266 );
and \U$20897 ( \21274 , \9612 , \10876 );
and \U$20898 ( \21275 , \9043 , \10873 );
nor \U$20899 ( \21276 , \21274 , \21275 );
xnor \U$20900 ( \21277 , \21276 , \9821 );
and \U$20901 ( \21278 , \10223 , \10063 );
and \U$20902 ( \21279 , \9620 , \10061 );
nor \U$20903 ( \21280 , \21278 , \21279 );
xnor \U$20904 ( \21281 , \21280 , \9824 );
and \U$20905 ( \21282 , \21277 , \21281 );
and \U$20906 ( \21283 , \21281 , \8587 );
and \U$20907 ( \21284 , \21277 , \8587 );
or \U$20908 ( \21285 , \21282 , \21283 , \21284 );
and \U$20909 ( \21286 , \10409 , \9495 );
and \U$20910 ( \21287 , \10228 , \9493 );
nor \U$20911 ( \21288 , \21286 , \21287 );
xnor \U$20912 ( \21289 , \21288 , \9185 );
nand \U$20913 ( \21290 , \11029 , \8956 );
xnor \U$20914 ( \21291 , \21290 , \8587 );
and \U$20915 ( \21292 , \21289 , \21291 );
and \U$20916 ( \21293 , \21285 , \21292 );
and \U$20917 ( \21294 , \11029 , \8958 );
and \U$20918 ( \21295 , \10409 , \8956 );
nor \U$20919 ( \21296 , \21294 , \21295 );
xnor \U$20920 ( \21297 , \21296 , \8587 );
and \U$20921 ( \21298 , \21292 , \21297 );
and \U$20922 ( \21299 , \21285 , \21297 );
or \U$20923 ( \21300 , \21293 , \21298 , \21299 );
xor \U$20924 ( \21301 , \21254 , \21256 );
xor \U$20925 ( \21302 , \21301 , \21259 );
and \U$20926 ( \21303 , \21300 , \21302 );
and \U$20927 ( \21304 , \21273 , \21303 );
xor \U$20928 ( \21305 , \21273 , \21303 );
xor \U$20929 ( \21306 , \21300 , \21302 );
xor \U$20930 ( \21307 , \21242 , \21246 );
xor \U$20931 ( \21308 , \21307 , \21251 );
xor \U$20932 ( \21309 , \21285 , \21292 );
xor \U$20933 ( \21310 , \21309 , \21297 );
and \U$20934 ( \21311 , \21308 , \21310 );
and \U$20935 ( \21312 , \21306 , \21311 );
xor \U$20936 ( \21313 , \21306 , \21311 );
xor \U$20937 ( \21314 , \21308 , \21310 );
and \U$20938 ( \21315 , \9620 , \10876 );
and \U$20939 ( \21316 , \9612 , \10873 );
nor \U$20940 ( \21317 , \21315 , \21316 );
xnor \U$20941 ( \21318 , \21317 , \9821 );
and \U$20942 ( \21319 , \10228 , \10063 );
and \U$20943 ( \21320 , \10223 , \10061 );
nor \U$20944 ( \21321 , \21319 , \21320 );
xnor \U$20945 ( \21322 , \21321 , \9824 );
and \U$20946 ( \21323 , \21318 , \21322 );
and \U$20947 ( \21324 , \11029 , \9495 );
and \U$20948 ( \21325 , \10409 , \9493 );
nor \U$20949 ( \21326 , \21324 , \21325 );
xnor \U$20950 ( \21327 , \21326 , \9185 );
and \U$20951 ( \21328 , \21322 , \21327 );
and \U$20952 ( \21329 , \21318 , \21327 );
or \U$20953 ( \21330 , \21323 , \21328 , \21329 );
xor \U$20954 ( \21331 , \21277 , \21281 );
xor \U$20955 ( \21332 , \21331 , \8587 );
and \U$20956 ( \21333 , \21330 , \21332 );
xor \U$20957 ( \21334 , \21289 , \21291 );
and \U$20958 ( \21335 , \21332 , \21334 );
and \U$20959 ( \21336 , \21330 , \21334 );
or \U$20960 ( \21337 , \21333 , \21335 , \21336 );
and \U$20961 ( \21338 , \21314 , \21337 );
xor \U$20962 ( \21339 , \21314 , \21337 );
xor \U$20963 ( \21340 , \21330 , \21332 );
xor \U$20964 ( \21341 , \21340 , \21334 );
and \U$20965 ( \21342 , \10223 , \10876 );
and \U$20966 ( \21343 , \9620 , \10873 );
nor \U$20967 ( \21344 , \21342 , \21343 );
xnor \U$20968 ( \21345 , \21344 , \9821 );
and \U$20969 ( \21346 , \10409 , \10063 );
and \U$20970 ( \21347 , \10228 , \10061 );
nor \U$20971 ( \21348 , \21346 , \21347 );
xnor \U$20972 ( \21349 , \21348 , \9824 );
and \U$20973 ( \21350 , \21345 , \21349 );
and \U$20974 ( \21351 , \21349 , \9185 );
and \U$20975 ( \21352 , \21345 , \9185 );
or \U$20976 ( \21353 , \21350 , \21351 , \21352 );
xor \U$20977 ( \21354 , \21318 , \21322 );
xor \U$20978 ( \21355 , \21354 , \21327 );
and \U$20979 ( \21356 , \21353 , \21355 );
and \U$20980 ( \21357 , \21341 , \21356 );
xor \U$20981 ( \21358 , \21341 , \21356 );
xor \U$20982 ( \21359 , \21353 , \21355 );
nand \U$20983 ( \21360 , \11029 , \9493 );
xnor \U$20984 ( \21361 , \21360 , \9185 );
xor \U$20985 ( \21362 , \21345 , \21349 );
xor \U$20986 ( \21363 , \21362 , \9185 );
and \U$20987 ( \21364 , \21361 , \21363 );
and \U$20988 ( \21365 , \21359 , \21364 );
xor \U$20989 ( \21366 , \21359 , \21364 );
xor \U$20990 ( \21367 , \21361 , \21363 );
and \U$20991 ( \21368 , \10228 , \10876 );
and \U$20992 ( \21369 , \10223 , \10873 );
nor \U$20993 ( \21370 , \21368 , \21369 );
xnor \U$20994 ( \21371 , \21370 , \9821 );
and \U$20995 ( \21372 , \11029 , \10063 );
and \U$20996 ( \21373 , \10409 , \10061 );
nor \U$20997 ( \21374 , \21372 , \21373 );
xnor \U$20998 ( \21375 , \21374 , \9824 );
and \U$20999 ( \21376 , \21371 , \21375 );
and \U$21000 ( \21377 , \21367 , \21376 );
xor \U$21001 ( \21378 , \21367 , \21376 );
xor \U$21002 ( \21379 , \21371 , \21375 );
and \U$21003 ( \21380 , \10409 , \10876 );
and \U$21004 ( \21381 , \10228 , \10873 );
nor \U$21005 ( \21382 , \21380 , \21381 );
xnor \U$21006 ( \21383 , \21382 , \9821 );
and \U$21007 ( \21384 , \21383 , \9824 );
and \U$21008 ( \21385 , \21379 , \21384 );
xor \U$21009 ( \21386 , \21379 , \21384 );
nand \U$21010 ( \21387 , \11029 , \10061 );
xnor \U$21011 ( \21388 , \21387 , \9824 );
xor \U$21012 ( \21389 , \21383 , \9824 );
and \U$21013 ( \21390 , \21388 , \21389 );
xor \U$21014 ( \21391 , \21388 , \21389 );
and \U$21015 ( \21392 , \11029 , \10876 );
and \U$21016 ( \21393 , \10409 , \10873 );
nor \U$21017 ( \21394 , \21392 , \21393 );
xnor \U$21018 ( \21395 , \21394 , \9821 );
nand \U$21019 ( \21396 , \11029 , \10873 );
xnor \U$21020 ( \21397 , \21396 , \9821 );
and \U$21021 ( \21398 , \21397 , \9821 );
and \U$21022 ( \21399 , \21395 , \21398 );
and \U$21023 ( \21400 , \21391 , \21399 );
or \U$21024 ( \21401 , \21390 , \21400 );
and \U$21025 ( \21402 , \21386 , \21401 );
or \U$21026 ( \21403 , \21385 , \21402 );
and \U$21027 ( \21404 , \21378 , \21403 );
or \U$21028 ( \21405 , \21377 , \21404 );
and \U$21029 ( \21406 , \21366 , \21405 );
or \U$21030 ( \21407 , \21365 , \21406 );
and \U$21031 ( \21408 , \21358 , \21407 );
or \U$21032 ( \21409 , \21357 , \21408 );
and \U$21033 ( \21410 , \21339 , \21409 );
or \U$21034 ( \21411 , \21338 , \21410 );
and \U$21035 ( \21412 , \21313 , \21411 );
or \U$21036 ( \21413 , \21312 , \21412 );
and \U$21037 ( \21414 , \21305 , \21413 );
or \U$21038 ( \21415 , \21304 , \21414 );
and \U$21039 ( \21416 , \21271 , \21415 );
or \U$21040 ( \21417 , \21270 , \21416 );
and \U$21041 ( \21418 , \21237 , \21417 );
or \U$21042 ( \21419 , \21236 , \21418 );
and \U$21043 ( \21420 , \21229 , \21419 );
or \U$21044 ( \21421 , \21228 , \21420 );
and \U$21045 ( \21422 , \21176 , \21421 );
or \U$21046 ( \21423 , \21175 , \21422 );
and \U$21047 ( \21424 , \21137 , \21423 );
or \U$21048 ( \21425 , \21136 , \21424 );
and \U$21049 ( \21426 , \21084 , \21425 );
or \U$21050 ( \21427 , \21083 , \21426 );
and \U$21051 ( \21428 , \21013 , \21427 );
or \U$21052 ( \21429 , \21012 , \21428 );
and \U$21053 ( \21430 , \20958 , \21429 );
or \U$21054 ( \21431 , \20957 , \21430 );
and \U$21055 ( \21432 , \20899 , \21431 );
or \U$21056 ( \21433 , \20898 , \21432 );
and \U$21057 ( \21434 , \20891 , \21433 );
or \U$21058 ( \21435 , \20890 , \21434 );
and \U$21059 ( \21436 , \20812 , \21435 );
or \U$21060 ( \21437 , \20811 , \21436 );
and \U$21061 ( \21438 , \20732 , \21437 );
or \U$21062 ( \21439 , \20731 , \21438 );
and \U$21063 ( \21440 , \20637 , \21439 );
or \U$21064 ( \21441 , \20636 , \21440 );
and \U$21065 ( \21442 , \20549 , \21441 );
or \U$21066 ( \21443 , \20548 , \21442 );
and \U$21067 ( \21444 , \20457 , \21443 );
or \U$21068 ( \21445 , \20456 , \21444 );
and \U$21069 ( \21446 , \20369 , \21445 );
or \U$21070 ( \21447 , \20368 , \21446 );
and \U$21071 ( \21448 , \20254 , \21447 );
or \U$21072 ( \21449 , \20253 , \21448 );
and \U$21073 ( \21450 , \20158 , \21449 );
or \U$21074 ( \21451 , \20157 , \21450 );
and \U$21075 ( \21452 , \20150 , \21451 );
or \U$21076 ( \21453 , \20149 , \21452 );
and \U$21077 ( \21454 , \20035 , \21453 );
or \U$21078 ( \21455 , \20034 , \21454 );
and \U$21079 ( \21456 , \19911 , \21455 );
or \U$21080 ( \21457 , \19910 , \21456 );
and \U$21081 ( \21458 , \19771 , \21457 );
or \U$21082 ( \21459 , \19770 , \21458 );
and \U$21083 ( \21460 , \19647 , \21459 );
or \U$21084 ( \21461 , \19646 , \21460 );
and \U$21085 ( \21462 , \19503 , \21461 );
or \U$21086 ( \21463 , \19502 , \21462 );
and \U$21087 ( \21464 , \19378 , \21463 );
or \U$21088 ( \21465 , \19377 , \21464 );
and \U$21089 ( \21466 , \19239 , \21465 );
or \U$21090 ( \21467 , \19238 , \21466 );
and \U$21091 ( \21468 , \19075 , \21467 );
or \U$21092 ( \21469 , \19074 , \21468 );
and \U$21093 ( \21470 , \18923 , \21469 );
or \U$21094 ( \21471 , \18922 , \21470 );
and \U$21095 ( \21472 , \18783 , \21471 );
or \U$21096 ( \21473 , \18782 , \21472 );
and \U$21097 ( \21474 , \18615 , \21473 );
or \U$21098 ( \21475 , \18614 , \21474 );
and \U$21099 ( \21476 , \18607 , \21475 );
or \U$21100 ( \21477 , \18606 , \21476 );
and \U$21101 ( \21478 , \18436 , \21477 );
or \U$21102 ( \21479 , \18435 , \21478 );
and \U$21103 ( \21480 , \18260 , \21479 );
or \U$21104 ( \21481 , \18259 , \21480 );
and \U$21105 ( \21482 , \18070 , \21481 );
or \U$21106 ( \21483 , \18069 , \21482 );
and \U$21107 ( \21484 , \17883 , \21483 );
or \U$21108 ( \21485 , \17882 , \21484 );
and \U$21109 ( \21486 , \17698 , \21485 );
or \U$21110 ( \21487 , \17697 , \21486 );
and \U$21111 ( \21488 , \17490 , \21487 );
or \U$21112 ( \21489 , \17489 , \21488 );
and \U$21113 ( \21490 , \17294 , \21489 );
or \U$21114 ( \21491 , \17293 , \21490 );
and \U$21115 ( \21492 , \17097 , \21491 );
or \U$21116 ( \21493 , \17096 , \21492 );
and \U$21117 ( \21494 , \16884 , \21493 );
or \U$21118 ( \21495 , \16883 , \21494 );
and \U$21119 ( \21496 , \16673 , \21495 );
or \U$21120 ( \21497 , \16672 , \21496 );
and \U$21121 ( \21498 , \16442 , \21497 );
or \U$21122 ( \21499 , \16441 , \21498 );
and \U$21123 ( \21500 , \16212 , \21499 );
or \U$21124 ( \21501 , \16211 , \21500 );
and \U$21125 ( \21502 , \15993 , \21501 );
or \U$21126 ( \21503 , \15992 , \21502 );
and \U$21127 ( \21504 , \15768 , \21503 );
or \U$21128 ( \21505 , \15767 , \21504 );
and \U$21129 ( \21506 , \15518 , \21505 );
or \U$21130 ( \21507 , \15517 , \21506 );
and \U$21131 ( \21508 , \15288 , \21507 );
or \U$21132 ( \21509 , \15287 , \21508 );
and \U$21133 ( \21510 , \15042 , \21509 );
or \U$21134 ( \21511 , \15041 , \21510 );
and \U$21135 ( \21512 , \15034 , \21511 );
or \U$21136 ( \21513 , \15033 , \21512 );
and \U$21137 ( \21514 , \14773 , \21513 );
or \U$21138 ( \21515 , \14772 , \21514 );
and \U$21139 ( \21516 , \14511 , \21515 );
or \U$21140 ( \21517 , \14510 , \21516 );
and \U$21141 ( \21518 , \14241 , \21517 );
or \U$21142 ( \21519 , \14240 , \21518 );
and \U$21143 ( \21520 , \13964 , \21519 );
or \U$21144 ( \21521 , \13963 , \21520 );
and \U$21145 ( \21522 , \13688 , \21521 );
or \U$21146 ( \21523 , \13687 , \21522 );
and \U$21147 ( \21524 , \13417 , \21523 );
or \U$21148 ( \21525 , \13416 , \21524 );
and \U$21149 ( \21526 , \13114 , \21525 );
or \U$21150 ( \21527 , \13113 , \21526 );
and \U$21151 ( \21528 , \12835 , \21527 );
or \U$21152 ( \21529 , \12834 , \21528 );
and \U$21153 ( \21530 , \12550 , \21529 );
or \U$21154 ( \21531 , \12549 , \21530 );
and \U$21155 ( \21532 , \12234 , \21531 );
or \U$21156 ( \21533 , \12233 , \21532 );
and \U$21157 ( \21534 , \11934 , \21533 );
or \U$21158 ( \21535 , \11933 , \21534 );
and \U$21159 ( \21536 , \11618 , \21535 );
or \U$21160 ( \21537 , \11617 , \21536 );
and \U$21161 ( \21538 , \11300 , \21537 );
or \U$21162 ( \21539 , \11299 , \21538 );
and \U$21163 ( \21540 , \10989 , \21539 );
or \U$21164 ( \21541 , \10988 , \21540 );
and \U$21165 ( \21542 , \10676 , \21541 );
or \U$21166 ( \21543 , \10675 , \21542 );
and \U$21167 ( \21544 , \10360 , \21543 );
or \U$21168 ( \21545 , \10359 , \21544 );
and \U$21169 ( \21546 , \10042 , \21545 );
or \U$21170 ( \21547 , \10041 , \21546 );
and \U$21171 ( \21548 , \9733 , \21547 );
or \U$21172 ( \21549 , \9732 , \21548 );
and \U$21173 ( \21550 , \9437 , \21549 );
or \U$21174 ( \21551 , \9436 , \21550 );
and \U$21175 ( \21552 , \9136 , \21551 );
or \U$21176 ( \21553 , \9135 , \21552 );
and \U$21177 ( \21554 , \8848 , \21553 );
or \U$21178 ( \21555 , \8847 , \21554 );
and \U$21179 ( \21556 , \8565 , \21555 );
or \U$21180 ( \21557 , \8564 , \21556 );
and \U$21181 ( \21558 , \8270 , \21557 );
or \U$21182 ( \21559 , \8269 , \21558 );
and \U$21183 ( \21560 , \8004 , \21559 );
or \U$21184 ( \21561 , \8003 , \21560 );
and \U$21185 ( \21562 , \7738 , \21561 );
or \U$21186 ( \21563 , \7737 , \21562 );
and \U$21187 ( \21564 , \7477 , \21563 );
or \U$21188 ( \21565 , \7476 , \21564 );
and \U$21189 ( \21566 , \7212 , \21565 );
or \U$21190 ( \21567 , \7211 , \21566 );
and \U$21191 ( \21568 , \6949 , \21567 );
or \U$21192 ( \21569 , \6948 , \21568 );
and \U$21193 ( \21570 , \6692 , \21569 );
or \U$21194 ( \21571 , \6691 , \21570 );
and \U$21195 ( \21572 , \6436 , \21571 );
or \U$21196 ( \21573 , \6435 , \21572 );
and \U$21197 ( \21574 , \6183 , \21573 );
or \U$21198 ( \21575 , \6182 , \21574 );
and \U$21199 ( \21576 , \5935 , \21575 );
or \U$21200 ( \21577 , \5934 , \21576 );
and \U$21201 ( \21578 , \5703 , \21577 );
or \U$21202 ( \21579 , \5702 , \21578 );
and \U$21203 ( \21580 , \5460 , \21579 );
or \U$21204 ( \21581 , \5459 , \21580 );
and \U$21205 ( \21582 , \5031 , \21581 );
or \U$21206 ( \21583 , \5030 , \21582 );
and \U$21207 ( \21584 , \4821 , \21583 );
or \U$21208 ( \21585 , \4820 , \21584 );
and \U$21209 ( \21586 , \4614 , \21585 );
or \U$21210 ( \21587 , \4613 , \21586 );
and \U$21211 ( \21588 , \4412 , \21587 );
or \U$21212 ( \21589 , \4411 , \21588 );
and \U$21213 ( \21590 , \4216 , \21589 );
or \U$21214 ( \21591 , \4215 , \21590 );
and \U$21215 ( \21592 , \4019 , \21591 );
or \U$21216 ( \21593 , \4018 , \21592 );
and \U$21217 ( \21594 , \3842 , \21593 );
or \U$21218 ( \21595 , \3841 , \21594 );
and \U$21219 ( \21596 , \3661 , \21595 );
or \U$21220 ( \21597 , \3660 , \21596 );
and \U$21221 ( \21598 , \3490 , \21597 );
or \U$21222 ( \21599 , \3489 , \21598 );
and \U$21223 ( \21600 , \3315 , \21599 );
or \U$21224 ( \21601 , \3314 , \21600 );
and \U$21225 ( \21602 , \3142 , \21601 );
or \U$21226 ( \21603 , \3141 , \21602 );
and \U$21227 ( \21604 , \2975 , \21603 );
or \U$21228 ( \21605 , \2974 , \21604 );
and \U$21229 ( \21606 , \2809 , \21605 );
or \U$21230 ( \21607 , \2808 , \21606 );
and \U$21231 ( \21608 , \2636 , \21607 );
or \U$21232 ( \21609 , \2635 , \21608 );
and \U$21233 ( \21610 , \2356 , \21609 );
or \U$21234 ( \21611 , \2355 , \21610 );
and \U$21235 ( \21612 , \2219 , \21611 );
or \U$21236 ( \21613 , \2218 , \21612 );
and \U$21237 ( \21614 , \2086 , \21613 );
or \U$21238 ( \21615 , \2085 , \21614 );
and \U$21239 ( \21616 , \1965 , \21615 );
or \U$21240 ( \21617 , \1964 , \21616 );
and \U$21241 ( \21618 , \1842 , \21617 );
or \U$21242 ( \21619 , \1841 , \21618 );
and \U$21243 ( \21620 , \1726 , \21619 );
or \U$21244 ( \21621 , \1725 , \21620 );
and \U$21245 ( \21622 , \1611 , \21621 );
or \U$21246 ( \21623 , \1610 , \21622 );
and \U$21247 ( \21624 , \1497 , \21623 );
or \U$21248 ( \21625 , \1496 , \21624 );
and \U$21249 ( \21626 , \1383 , \21625 );
or \U$21250 ( \21627 , \1382 , \21626 );
and \U$21251 ( \21628 , \1201 , \21627 );
or \U$21252 ( \21629 , \1200 , \21628 );
and \U$21253 ( \21630 , \1122 , \21629 );
or \U$21254 ( \21631 , \1121 , \21630 );
and \U$21255 ( \21632 , \1039 , \21631 );
or \U$21256 ( \21633 , \1038 , \21632 );
and \U$21257 ( \21634 , \958 , \21633 );
or \U$21258 ( \21635 , \957 , \21634 );
and \U$21259 ( \21636 , \883 , \21635 );
or \U$21260 ( \21637 , \882 , \21636 );
and \U$21261 ( \21638 , \809 , \21637 );
or \U$21262 ( \21639 , \808 , \21638 );
and \U$21263 ( \21640 , \689 , \21639 );
or \U$21264 ( \21641 , \688 , \21640 );
and \U$21265 ( \21642 , \636 , \21641 );
or \U$21266 ( \21643 , \635 , \21642 );
and \U$21267 ( \21644 , \586 , \21643 );
or \U$21268 ( \21645 , \585 , \21644 );
and \U$21269 ( \21646 , \534 , \21645 );
or \U$21270 ( \21647 , \533 , \21646 );
and \U$21271 ( \21648 , \464 , \21647 );
or \U$21272 ( \21649 , \463 , \21648 );
xor \U$21273 ( \21650 , \417 , \21649 );
buf gaed4_GF_PartitionCandidate( \21651_nGaed4 , \21650 );
buf \U$21274 ( \21652 , \21651_nGaed4 );
buf \U$21275 ( \21653 , RIc229590_129);
buf \U$21276 ( \21654 , RIc2275b0_1);
buf \U$21277 ( \21655 , RIc227538_2);
xor \U$21278 ( \21656 , \21654 , \21655 );
buf \U$21279 ( \21657 , RIc2274c0_3);
xor \U$21280 ( \21658 , \21655 , \21657 );
not \U$21281 ( \21659 , \21658 );
and \U$21282 ( \21660 , \21656 , \21659 );
and \U$21283 ( \21661 , \21653 , \21660 );
not \U$21284 ( \21662 , \21661 );
and \U$21285 ( \21663 , \21655 , \21657 );
not \U$21286 ( \21664 , \21663 );
and \U$21287 ( \21665 , \21654 , \21664 );
xnor \U$21288 ( \21666 , \21662 , \21665 );
buf \U$21289 ( \21667 , RIc229608_130);
and \U$21290 ( \21668 , \21667 , \21654 );
or \U$21291 ( \21669 , \21666 , \21668 );
not \U$21292 ( \21670 , \21665 );
xor \U$21293 ( \21671 , \21669 , \21670 );
and \U$21294 ( \21672 , \21653 , \21654 );
xor \U$21295 ( \21673 , \21671 , \21672 );
buf \U$21296 ( \21674 , RIc227448_4);
buf \U$21297 ( \21675 , RIc2273d0_5);
and \U$21298 ( \21676 , \21674 , \21675 );
not \U$21299 ( \21677 , \21676 );
and \U$21300 ( \21678 , \21657 , \21677 );
not \U$21301 ( \21679 , \21678 );
and \U$21302 ( \21680 , \21667 , \21660 );
and \U$21303 ( \21681 , \21653 , \21658 );
nor \U$21304 ( \21682 , \21680 , \21681 );
xnor \U$21305 ( \21683 , \21682 , \21665 );
and \U$21306 ( \21684 , \21679 , \21683 );
buf \U$21307 ( \21685 , RIc229680_131);
and \U$21308 ( \21686 , \21685 , \21654 );
and \U$21309 ( \21687 , \21683 , \21686 );
and \U$21310 ( \21688 , \21679 , \21686 );
or \U$21311 ( \21689 , \21684 , \21687 , \21688 );
xnor \U$21312 ( \21690 , \21666 , \21668 );
and \U$21313 ( \21691 , \21689 , \21690 );
xor \U$21314 ( \21692 , \21673 , \21691 );
xor \U$21315 ( \21693 , \21689 , \21690 );
xor \U$21316 ( \21694 , \21657 , \21674 );
xor \U$21317 ( \21695 , \21674 , \21675 );
not \U$21318 ( \21696 , \21695 );
and \U$21319 ( \21697 , \21694 , \21696 );
and \U$21320 ( \21698 , \21653 , \21697 );
not \U$21321 ( \21699 , \21698 );
xnor \U$21322 ( \21700 , \21699 , \21678 );
and \U$21323 ( \21701 , \21685 , \21660 );
and \U$21324 ( \21702 , \21667 , \21658 );
nor \U$21325 ( \21703 , \21701 , \21702 );
xnor \U$21326 ( \21704 , \21703 , \21665 );
and \U$21327 ( \21705 , \21700 , \21704 );
buf \U$21328 ( \21706 , RIc2296f8_132);
and \U$21329 ( \21707 , \21706 , \21654 );
and \U$21330 ( \21708 , \21704 , \21707 );
and \U$21331 ( \21709 , \21700 , \21707 );
or \U$21332 ( \21710 , \21705 , \21708 , \21709 );
buf \U$21333 ( \21711 , RIc227358_6);
buf \U$21334 ( \21712 , RIc2272e0_7);
and \U$21335 ( \21713 , \21711 , \21712 );
not \U$21336 ( \21714 , \21713 );
and \U$21337 ( \21715 , \21675 , \21714 );
not \U$21338 ( \21716 , \21715 );
and \U$21339 ( \21717 , \21667 , \21697 );
and \U$21340 ( \21718 , \21653 , \21695 );
nor \U$21341 ( \21719 , \21717 , \21718 );
xnor \U$21342 ( \21720 , \21719 , \21678 );
and \U$21343 ( \21721 , \21716 , \21720 );
and \U$21344 ( \21722 , \21706 , \21660 );
and \U$21345 ( \21723 , \21685 , \21658 );
nor \U$21346 ( \21724 , \21722 , \21723 );
xnor \U$21347 ( \21725 , \21724 , \21665 );
and \U$21348 ( \21726 , \21720 , \21725 );
and \U$21349 ( \21727 , \21716 , \21725 );
or \U$21350 ( \21728 , \21721 , \21726 , \21727 );
xor \U$21351 ( \21729 , \21700 , \21704 );
xor \U$21352 ( \21730 , \21729 , \21707 );
or \U$21353 ( \21731 , \21728 , \21730 );
and \U$21354 ( \21732 , \21710 , \21731 );
xor \U$21355 ( \21733 , \21679 , \21683 );
xor \U$21356 ( \21734 , \21733 , \21686 );
and \U$21357 ( \21735 , \21731 , \21734 );
and \U$21358 ( \21736 , \21710 , \21734 );
or \U$21359 ( \21737 , \21732 , \21735 , \21736 );
and \U$21360 ( \21738 , \21693 , \21737 );
xor \U$21361 ( \21739 , \21693 , \21737 );
xor \U$21362 ( \21740 , \21710 , \21731 );
xor \U$21363 ( \21741 , \21740 , \21734 );
xor \U$21364 ( \21742 , \21675 , \21711 );
xor \U$21365 ( \21743 , \21711 , \21712 );
not \U$21366 ( \21744 , \21743 );
and \U$21367 ( \21745 , \21742 , \21744 );
and \U$21368 ( \21746 , \21653 , \21745 );
not \U$21369 ( \21747 , \21746 );
xnor \U$21370 ( \21748 , \21747 , \21715 );
and \U$21371 ( \21749 , \21685 , \21697 );
and \U$21372 ( \21750 , \21667 , \21695 );
nor \U$21373 ( \21751 , \21749 , \21750 );
xnor \U$21374 ( \21752 , \21751 , \21678 );
and \U$21375 ( \21753 , \21748 , \21752 );
buf \U$21376 ( \21754 , RIc229770_133);
and \U$21377 ( \21755 , \21754 , \21660 );
and \U$21378 ( \21756 , \21706 , \21658 );
nor \U$21379 ( \21757 , \21755 , \21756 );
xnor \U$21380 ( \21758 , \21757 , \21665 );
and \U$21381 ( \21759 , \21752 , \21758 );
and \U$21382 ( \21760 , \21748 , \21758 );
or \U$21383 ( \21761 , \21753 , \21759 , \21760 );
buf \U$21384 ( \21762 , RIc2297e8_134);
and \U$21385 ( \21763 , \21762 , \21654 );
buf \U$21386 ( \21764 , \21763 );
and \U$21387 ( \21765 , \21761 , \21764 );
and \U$21388 ( \21766 , \21754 , \21654 );
and \U$21389 ( \21767 , \21764 , \21766 );
and \U$21390 ( \21768 , \21761 , \21766 );
or \U$21391 ( \21769 , \21765 , \21767 , \21768 );
buf \U$21392 ( \21770 , RIc227268_8);
buf \U$21393 ( \21771 , RIc2271f0_9);
and \U$21394 ( \21772 , \21770 , \21771 );
not \U$21395 ( \21773 , \21772 );
and \U$21396 ( \21774 , \21712 , \21773 );
not \U$21397 ( \21775 , \21774 );
and \U$21398 ( \21776 , \21667 , \21745 );
and \U$21399 ( \21777 , \21653 , \21743 );
nor \U$21400 ( \21778 , \21776 , \21777 );
xnor \U$21401 ( \21779 , \21778 , \21715 );
and \U$21402 ( \21780 , \21775 , \21779 );
and \U$21403 ( \21781 , \21706 , \21697 );
and \U$21404 ( \21782 , \21685 , \21695 );
nor \U$21405 ( \21783 , \21781 , \21782 );
xnor \U$21406 ( \21784 , \21783 , \21678 );
and \U$21407 ( \21785 , \21779 , \21784 );
and \U$21408 ( \21786 , \21775 , \21784 );
or \U$21409 ( \21787 , \21780 , \21785 , \21786 );
xor \U$21410 ( \21788 , \21748 , \21752 );
xor \U$21411 ( \21789 , \21788 , \21758 );
and \U$21412 ( \21790 , \21787 , \21789 );
not \U$21413 ( \21791 , \21763 );
and \U$21414 ( \21792 , \21789 , \21791 );
and \U$21415 ( \21793 , \21787 , \21791 );
or \U$21416 ( \21794 , \21790 , \21792 , \21793 );
xor \U$21417 ( \21795 , \21716 , \21720 );
xor \U$21418 ( \21796 , \21795 , \21725 );
and \U$21419 ( \21797 , \21794 , \21796 );
xor \U$21420 ( \21798 , \21761 , \21764 );
xor \U$21421 ( \21799 , \21798 , \21766 );
and \U$21422 ( \21800 , \21796 , \21799 );
and \U$21423 ( \21801 , \21794 , \21799 );
or \U$21424 ( \21802 , \21797 , \21800 , \21801 );
and \U$21425 ( \21803 , \21769 , \21802 );
xnor \U$21426 ( \21804 , \21728 , \21730 );
and \U$21427 ( \21805 , \21802 , \21804 );
and \U$21428 ( \21806 , \21769 , \21804 );
or \U$21429 ( \21807 , \21803 , \21805 , \21806 );
and \U$21430 ( \21808 , \21741 , \21807 );
xor \U$21431 ( \21809 , \21741 , \21807 );
xor \U$21432 ( \21810 , \21769 , \21802 );
xor \U$21433 ( \21811 , \21810 , \21804 );
xor \U$21434 ( \21812 , \21712 , \21770 );
xor \U$21435 ( \21813 , \21770 , \21771 );
not \U$21436 ( \21814 , \21813 );
and \U$21437 ( \21815 , \21812 , \21814 );
and \U$21438 ( \21816 , \21653 , \21815 );
not \U$21439 ( \21817 , \21816 );
xnor \U$21440 ( \21818 , \21817 , \21774 );
and \U$21441 ( \21819 , \21685 , \21745 );
and \U$21442 ( \21820 , \21667 , \21743 );
nor \U$21443 ( \21821 , \21819 , \21820 );
xnor \U$21444 ( \21822 , \21821 , \21715 );
and \U$21445 ( \21823 , \21818 , \21822 );
and \U$21446 ( \21824 , \21754 , \21697 );
and \U$21447 ( \21825 , \21706 , \21695 );
nor \U$21448 ( \21826 , \21824 , \21825 );
xnor \U$21449 ( \21827 , \21826 , \21678 );
and \U$21450 ( \21828 , \21822 , \21827 );
and \U$21451 ( \21829 , \21818 , \21827 );
or \U$21452 ( \21830 , \21823 , \21828 , \21829 );
buf \U$21453 ( \21831 , RIc229860_135);
and \U$21454 ( \21832 , \21831 , \21660 );
and \U$21455 ( \21833 , \21762 , \21658 );
nor \U$21456 ( \21834 , \21832 , \21833 );
xnor \U$21457 ( \21835 , \21834 , \21665 );
buf \U$21458 ( \21836 , RIc2298d8_136);
and \U$21459 ( \21837 , \21836 , \21654 );
or \U$21460 ( \21838 , \21835 , \21837 );
and \U$21461 ( \21839 , \21830 , \21838 );
and \U$21462 ( \21840 , \21762 , \21660 );
and \U$21463 ( \21841 , \21754 , \21658 );
nor \U$21464 ( \21842 , \21840 , \21841 );
xnor \U$21465 ( \21843 , \21842 , \21665 );
and \U$21466 ( \21844 , \21838 , \21843 );
and \U$21467 ( \21845 , \21830 , \21843 );
or \U$21468 ( \21846 , \21839 , \21844 , \21845 );
and \U$21469 ( \21847 , \21831 , \21654 );
xor \U$21470 ( \21848 , \21775 , \21779 );
xor \U$21471 ( \21849 , \21848 , \21784 );
and \U$21472 ( \21850 , \21847 , \21849 );
and \U$21473 ( \21851 , \21846 , \21850 );
xor \U$21474 ( \21852 , \21787 , \21789 );
xor \U$21475 ( \21853 , \21852 , \21791 );
and \U$21476 ( \21854 , \21850 , \21853 );
and \U$21477 ( \21855 , \21846 , \21853 );
or \U$21478 ( \21856 , \21851 , \21854 , \21855 );
xor \U$21479 ( \21857 , \21794 , \21796 );
xor \U$21480 ( \21858 , \21857 , \21799 );
and \U$21481 ( \21859 , \21856 , \21858 );
and \U$21482 ( \21860 , \21811 , \21859 );
xor \U$21483 ( \21861 , \21811 , \21859 );
xor \U$21484 ( \21862 , \21856 , \21858 );
buf \U$21485 ( \21863 , RIc227178_10);
buf \U$21486 ( \21864 , RIc227100_11);
and \U$21487 ( \21865 , \21863 , \21864 );
not \U$21488 ( \21866 , \21865 );
and \U$21489 ( \21867 , \21771 , \21866 );
not \U$21490 ( \21868 , \21867 );
and \U$21491 ( \21869 , \21667 , \21815 );
and \U$21492 ( \21870 , \21653 , \21813 );
nor \U$21493 ( \21871 , \21869 , \21870 );
xnor \U$21494 ( \21872 , \21871 , \21774 );
and \U$21495 ( \21873 , \21868 , \21872 );
and \U$21496 ( \21874 , \21706 , \21745 );
and \U$21497 ( \21875 , \21685 , \21743 );
nor \U$21498 ( \21876 , \21874 , \21875 );
xnor \U$21499 ( \21877 , \21876 , \21715 );
and \U$21500 ( \21878 , \21872 , \21877 );
and \U$21501 ( \21879 , \21868 , \21877 );
or \U$21502 ( \21880 , \21873 , \21878 , \21879 );
and \U$21503 ( \21881 , \21762 , \21697 );
and \U$21504 ( \21882 , \21754 , \21695 );
nor \U$21505 ( \21883 , \21881 , \21882 );
xnor \U$21506 ( \21884 , \21883 , \21678 );
and \U$21507 ( \21885 , \21836 , \21660 );
and \U$21508 ( \21886 , \21831 , \21658 );
nor \U$21509 ( \21887 , \21885 , \21886 );
xnor \U$21510 ( \21888 , \21887 , \21665 );
and \U$21511 ( \21889 , \21884 , \21888 );
buf \U$21512 ( \21890 , RIc229950_137);
and \U$21513 ( \21891 , \21890 , \21654 );
and \U$21514 ( \21892 , \21888 , \21891 );
and \U$21515 ( \21893 , \21884 , \21891 );
or \U$21516 ( \21894 , \21889 , \21892 , \21893 );
and \U$21517 ( \21895 , \21880 , \21894 );
xnor \U$21518 ( \21896 , \21835 , \21837 );
and \U$21519 ( \21897 , \21894 , \21896 );
and \U$21520 ( \21898 , \21880 , \21896 );
or \U$21521 ( \21899 , \21895 , \21897 , \21898 );
xor \U$21522 ( \21900 , \21830 , \21838 );
xor \U$21523 ( \21901 , \21900 , \21843 );
and \U$21524 ( \21902 , \21899 , \21901 );
xor \U$21525 ( \21903 , \21847 , \21849 );
and \U$21526 ( \21904 , \21901 , \21903 );
and \U$21527 ( \21905 , \21899 , \21903 );
or \U$21528 ( \21906 , \21902 , \21904 , \21905 );
xor \U$21529 ( \21907 , \21846 , \21850 );
xor \U$21530 ( \21908 , \21907 , \21853 );
and \U$21531 ( \21909 , \21906 , \21908 );
and \U$21532 ( \21910 , \21862 , \21909 );
xor \U$21533 ( \21911 , \21862 , \21909 );
xor \U$21534 ( \21912 , \21906 , \21908 );
xor \U$21535 ( \21913 , \21771 , \21863 );
xor \U$21536 ( \21914 , \21863 , \21864 );
not \U$21537 ( \21915 , \21914 );
and \U$21538 ( \21916 , \21913 , \21915 );
and \U$21539 ( \21917 , \21653 , \21916 );
not \U$21540 ( \21918 , \21917 );
xnor \U$21541 ( \21919 , \21918 , \21867 );
and \U$21542 ( \21920 , \21685 , \21815 );
and \U$21543 ( \21921 , \21667 , \21813 );
nor \U$21544 ( \21922 , \21920 , \21921 );
xnor \U$21545 ( \21923 , \21922 , \21774 );
and \U$21546 ( \21924 , \21919 , \21923 );
and \U$21547 ( \21925 , \21754 , \21745 );
and \U$21548 ( \21926 , \21706 , \21743 );
nor \U$21549 ( \21927 , \21925 , \21926 );
xnor \U$21550 ( \21928 , \21927 , \21715 );
and \U$21551 ( \21929 , \21923 , \21928 );
and \U$21552 ( \21930 , \21919 , \21928 );
or \U$21553 ( \21931 , \21924 , \21929 , \21930 );
and \U$21554 ( \21932 , \21831 , \21697 );
and \U$21555 ( \21933 , \21762 , \21695 );
nor \U$21556 ( \21934 , \21932 , \21933 );
xnor \U$21557 ( \21935 , \21934 , \21678 );
and \U$21558 ( \21936 , \21890 , \21660 );
and \U$21559 ( \21937 , \21836 , \21658 );
nor \U$21560 ( \21938 , \21936 , \21937 );
xnor \U$21561 ( \21939 , \21938 , \21665 );
and \U$21562 ( \21940 , \21935 , \21939 );
buf \U$21563 ( \21941 , RIc2299c8_138);
and \U$21564 ( \21942 , \21941 , \21654 );
and \U$21565 ( \21943 , \21939 , \21942 );
and \U$21566 ( \21944 , \21935 , \21942 );
or \U$21567 ( \21945 , \21940 , \21943 , \21944 );
and \U$21568 ( \21946 , \21931 , \21945 );
xor \U$21569 ( \21947 , \21884 , \21888 );
xor \U$21570 ( \21948 , \21947 , \21891 );
and \U$21571 ( \21949 , \21945 , \21948 );
and \U$21572 ( \21950 , \21931 , \21948 );
or \U$21573 ( \21951 , \21946 , \21949 , \21950 );
xor \U$21574 ( \21952 , \21818 , \21822 );
xor \U$21575 ( \21953 , \21952 , \21827 );
and \U$21576 ( \21954 , \21951 , \21953 );
xor \U$21577 ( \21955 , \21880 , \21894 );
xor \U$21578 ( \21956 , \21955 , \21896 );
and \U$21579 ( \21957 , \21953 , \21956 );
and \U$21580 ( \21958 , \21951 , \21956 );
or \U$21581 ( \21959 , \21954 , \21957 , \21958 );
xor \U$21582 ( \21960 , \21899 , \21901 );
xor \U$21583 ( \21961 , \21960 , \21903 );
and \U$21584 ( \21962 , \21959 , \21961 );
and \U$21585 ( \21963 , \21912 , \21962 );
xor \U$21586 ( \21964 , \21912 , \21962 );
xor \U$21587 ( \21965 , \21959 , \21961 );
and \U$21588 ( \21966 , \21762 , \21745 );
and \U$21589 ( \21967 , \21754 , \21743 );
nor \U$21590 ( \21968 , \21966 , \21967 );
xnor \U$21591 ( \21969 , \21968 , \21715 );
and \U$21592 ( \21970 , \21836 , \21697 );
and \U$21593 ( \21971 , \21831 , \21695 );
nor \U$21594 ( \21972 , \21970 , \21971 );
xnor \U$21595 ( \21973 , \21972 , \21678 );
and \U$21596 ( \21974 , \21969 , \21973 );
and \U$21597 ( \21975 , \21941 , \21660 );
and \U$21598 ( \21976 , \21890 , \21658 );
nor \U$21599 ( \21977 , \21975 , \21976 );
xnor \U$21600 ( \21978 , \21977 , \21665 );
and \U$21601 ( \21979 , \21973 , \21978 );
and \U$21602 ( \21980 , \21969 , \21978 );
or \U$21603 ( \21981 , \21974 , \21979 , \21980 );
buf \U$21604 ( \21982 , RIc227088_12);
buf \U$21605 ( \21983 , RIc227010_13);
and \U$21606 ( \21984 , \21982 , \21983 );
not \U$21607 ( \21985 , \21984 );
and \U$21608 ( \21986 , \21864 , \21985 );
not \U$21609 ( \21987 , \21986 );
and \U$21610 ( \21988 , \21667 , \21916 );
and \U$21611 ( \21989 , \21653 , \21914 );
nor \U$21612 ( \21990 , \21988 , \21989 );
xnor \U$21613 ( \21991 , \21990 , \21867 );
and \U$21614 ( \21992 , \21987 , \21991 );
and \U$21615 ( \21993 , \21706 , \21815 );
and \U$21616 ( \21994 , \21685 , \21813 );
nor \U$21617 ( \21995 , \21993 , \21994 );
xnor \U$21618 ( \21996 , \21995 , \21774 );
and \U$21619 ( \21997 , \21991 , \21996 );
and \U$21620 ( \21998 , \21987 , \21996 );
or \U$21621 ( \21999 , \21992 , \21997 , \21998 );
or \U$21622 ( \22000 , \21981 , \21999 );
xor \U$21623 ( \22001 , \21868 , \21872 );
xor \U$21624 ( \22002 , \22001 , \21877 );
and \U$21625 ( \22003 , \22000 , \22002 );
xor \U$21626 ( \22004 , \21931 , \21945 );
xor \U$21627 ( \22005 , \22004 , \21948 );
and \U$21628 ( \22006 , \22002 , \22005 );
and \U$21629 ( \22007 , \22000 , \22005 );
or \U$21630 ( \22008 , \22003 , \22006 , \22007 );
and \U$21631 ( \22009 , \21831 , \21745 );
and \U$21632 ( \22010 , \21762 , \21743 );
nor \U$21633 ( \22011 , \22009 , \22010 );
xnor \U$21634 ( \22012 , \22011 , \21715 );
and \U$21635 ( \22013 , \21890 , \21697 );
and \U$21636 ( \22014 , \21836 , \21695 );
nor \U$21637 ( \22015 , \22013 , \22014 );
xnor \U$21638 ( \22016 , \22015 , \21678 );
and \U$21639 ( \22017 , \22012 , \22016 );
buf \U$21640 ( \22018 , RIc229a40_139);
and \U$21641 ( \22019 , \22018 , \21660 );
and \U$21642 ( \22020 , \21941 , \21658 );
nor \U$21643 ( \22021 , \22019 , \22020 );
xnor \U$21644 ( \22022 , \22021 , \21665 );
and \U$21645 ( \22023 , \22016 , \22022 );
and \U$21646 ( \22024 , \22012 , \22022 );
or \U$21647 ( \22025 , \22017 , \22023 , \22024 );
xor \U$21648 ( \22026 , \21864 , \21982 );
xor \U$21649 ( \22027 , \21982 , \21983 );
not \U$21650 ( \22028 , \22027 );
and \U$21651 ( \22029 , \22026 , \22028 );
and \U$21652 ( \22030 , \21653 , \22029 );
not \U$21653 ( \22031 , \22030 );
xnor \U$21654 ( \22032 , \22031 , \21986 );
and \U$21655 ( \22033 , \21685 , \21916 );
and \U$21656 ( \22034 , \21667 , \21914 );
nor \U$21657 ( \22035 , \22033 , \22034 );
xnor \U$21658 ( \22036 , \22035 , \21867 );
and \U$21659 ( \22037 , \22032 , \22036 );
and \U$21660 ( \22038 , \21754 , \21815 );
and \U$21661 ( \22039 , \21706 , \21813 );
nor \U$21662 ( \22040 , \22038 , \22039 );
xnor \U$21663 ( \22041 , \22040 , \21774 );
and \U$21664 ( \22042 , \22036 , \22041 );
and \U$21665 ( \22043 , \22032 , \22041 );
or \U$21666 ( \22044 , \22037 , \22042 , \22043 );
and \U$21667 ( \22045 , \22025 , \22044 );
buf \U$21668 ( \22046 , RIc229ab8_140);
and \U$21669 ( \22047 , \22046 , \21654 );
buf \U$21670 ( \22048 , \22047 );
and \U$21671 ( \22049 , \22044 , \22048 );
and \U$21672 ( \22050 , \22025 , \22048 );
or \U$21673 ( \22051 , \22045 , \22049 , \22050 );
and \U$21674 ( \22052 , \22018 , \21654 );
xor \U$21675 ( \22053 , \21969 , \21973 );
xor \U$21676 ( \22054 , \22053 , \21978 );
and \U$21677 ( \22055 , \22052 , \22054 );
xor \U$21678 ( \22056 , \21987 , \21991 );
xor \U$21679 ( \22057 , \22056 , \21996 );
and \U$21680 ( \22058 , \22054 , \22057 );
and \U$21681 ( \22059 , \22052 , \22057 );
or \U$21682 ( \22060 , \22055 , \22058 , \22059 );
and \U$21683 ( \22061 , \22051 , \22060 );
xor \U$21684 ( \22062 , \21935 , \21939 );
xor \U$21685 ( \22063 , \22062 , \21942 );
and \U$21686 ( \22064 , \22060 , \22063 );
and \U$21687 ( \22065 , \22051 , \22063 );
or \U$21688 ( \22066 , \22061 , \22064 , \22065 );
xor \U$21689 ( \22067 , \21919 , \21923 );
xor \U$21690 ( \22068 , \22067 , \21928 );
xnor \U$21691 ( \22069 , \21981 , \21999 );
and \U$21692 ( \22070 , \22068 , \22069 );
and \U$21693 ( \22071 , \22066 , \22070 );
xor \U$21694 ( \22072 , \22000 , \22002 );
xor \U$21695 ( \22073 , \22072 , \22005 );
and \U$21696 ( \22074 , \22070 , \22073 );
and \U$21697 ( \22075 , \22066 , \22073 );
or \U$21698 ( \22076 , \22071 , \22074 , \22075 );
and \U$21699 ( \22077 , \22008 , \22076 );
xor \U$21700 ( \22078 , \21951 , \21953 );
xor \U$21701 ( \22079 , \22078 , \21956 );
and \U$21702 ( \22080 , \22076 , \22079 );
and \U$21703 ( \22081 , \22008 , \22079 );
or \U$21704 ( \22082 , \22077 , \22080 , \22081 );
and \U$21705 ( \22083 , \21965 , \22082 );
xor \U$21706 ( \22084 , \21965 , \22082 );
xor \U$21707 ( \22085 , \22008 , \22076 );
xor \U$21708 ( \22086 , \22085 , \22079 );
buf \U$21709 ( \22087 , RIc226f98_14);
buf \U$21710 ( \22088 , RIc226f20_15);
and \U$21711 ( \22089 , \22087 , \22088 );
not \U$21712 ( \22090 , \22089 );
and \U$21713 ( \22091 , \21983 , \22090 );
not \U$21714 ( \22092 , \22091 );
and \U$21715 ( \22093 , \21667 , \22029 );
and \U$21716 ( \22094 , \21653 , \22027 );
nor \U$21717 ( \22095 , \22093 , \22094 );
xnor \U$21718 ( \22096 , \22095 , \21986 );
and \U$21719 ( \22097 , \22092 , \22096 );
and \U$21720 ( \22098 , \21706 , \21916 );
and \U$21721 ( \22099 , \21685 , \21914 );
nor \U$21722 ( \22100 , \22098 , \22099 );
xnor \U$21723 ( \22101 , \22100 , \21867 );
and \U$21724 ( \22102 , \22096 , \22101 );
and \U$21725 ( \22103 , \22092 , \22101 );
or \U$21726 ( \22104 , \22097 , \22102 , \22103 );
and \U$21727 ( \22105 , \21762 , \21815 );
and \U$21728 ( \22106 , \21754 , \21813 );
nor \U$21729 ( \22107 , \22105 , \22106 );
xnor \U$21730 ( \22108 , \22107 , \21774 );
and \U$21731 ( \22109 , \21836 , \21745 );
and \U$21732 ( \22110 , \21831 , \21743 );
nor \U$21733 ( \22111 , \22109 , \22110 );
xnor \U$21734 ( \22112 , \22111 , \21715 );
and \U$21735 ( \22113 , \22108 , \22112 );
and \U$21736 ( \22114 , \21941 , \21697 );
and \U$21737 ( \22115 , \21890 , \21695 );
nor \U$21738 ( \22116 , \22114 , \22115 );
xnor \U$21739 ( \22117 , \22116 , \21678 );
and \U$21740 ( \22118 , \22112 , \22117 );
and \U$21741 ( \22119 , \22108 , \22117 );
or \U$21742 ( \22120 , \22113 , \22118 , \22119 );
and \U$21743 ( \22121 , \22104 , \22120 );
and \U$21744 ( \22122 , \22046 , \21660 );
and \U$21745 ( \22123 , \22018 , \21658 );
nor \U$21746 ( \22124 , \22122 , \22123 );
xnor \U$21747 ( \22125 , \22124 , \21665 );
buf \U$21748 ( \22126 , RIc229b30_141);
and \U$21749 ( \22127 , \22126 , \21654 );
and \U$21750 ( \22128 , \22125 , \22127 );
and \U$21751 ( \22129 , \22120 , \22128 );
and \U$21752 ( \22130 , \22104 , \22128 );
or \U$21753 ( \22131 , \22121 , \22129 , \22130 );
xor \U$21754 ( \22132 , \22012 , \22016 );
xor \U$21755 ( \22133 , \22132 , \22022 );
xor \U$21756 ( \22134 , \22032 , \22036 );
xor \U$21757 ( \22135 , \22134 , \22041 );
and \U$21758 ( \22136 , \22133 , \22135 );
not \U$21759 ( \22137 , \22047 );
and \U$21760 ( \22138 , \22135 , \22137 );
and \U$21761 ( \22139 , \22133 , \22137 );
or \U$21762 ( \22140 , \22136 , \22138 , \22139 );
and \U$21763 ( \22141 , \22131 , \22140 );
xor \U$21764 ( \22142 , \22052 , \22054 );
xor \U$21765 ( \22143 , \22142 , \22057 );
and \U$21766 ( \22144 , \22140 , \22143 );
and \U$21767 ( \22145 , \22131 , \22143 );
or \U$21768 ( \22146 , \22141 , \22144 , \22145 );
xor \U$21769 ( \22147 , \22051 , \22060 );
xor \U$21770 ( \22148 , \22147 , \22063 );
and \U$21771 ( \22149 , \22146 , \22148 );
xor \U$21772 ( \22150 , \22068 , \22069 );
and \U$21773 ( \22151 , \22148 , \22150 );
and \U$21774 ( \22152 , \22146 , \22150 );
or \U$21775 ( \22153 , \22149 , \22151 , \22152 );
xor \U$21776 ( \22154 , \22066 , \22070 );
xor \U$21777 ( \22155 , \22154 , \22073 );
and \U$21778 ( \22156 , \22153 , \22155 );
and \U$21779 ( \22157 , \22086 , \22156 );
xor \U$21780 ( \22158 , \22086 , \22156 );
xor \U$21781 ( \22159 , \22153 , \22155 );
xor \U$21782 ( \22160 , \21983 , \22087 );
xor \U$21783 ( \22161 , \22087 , \22088 );
not \U$21784 ( \22162 , \22161 );
and \U$21785 ( \22163 , \22160 , \22162 );
and \U$21786 ( \22164 , \21653 , \22163 );
not \U$21787 ( \22165 , \22164 );
xnor \U$21788 ( \22166 , \22165 , \22091 );
and \U$21789 ( \22167 , \21685 , \22029 );
and \U$21790 ( \22168 , \21667 , \22027 );
nor \U$21791 ( \22169 , \22167 , \22168 );
xnor \U$21792 ( \22170 , \22169 , \21986 );
and \U$21793 ( \22171 , \22166 , \22170 );
and \U$21794 ( \22172 , \21754 , \21916 );
and \U$21795 ( \22173 , \21706 , \21914 );
nor \U$21796 ( \22174 , \22172 , \22173 );
xnor \U$21797 ( \22175 , \22174 , \21867 );
and \U$21798 ( \22176 , \22170 , \22175 );
and \U$21799 ( \22177 , \22166 , \22175 );
or \U$21800 ( \22178 , \22171 , \22176 , \22177 );
and \U$21801 ( \22179 , \21831 , \21815 );
and \U$21802 ( \22180 , \21762 , \21813 );
nor \U$21803 ( \22181 , \22179 , \22180 );
xnor \U$21804 ( \22182 , \22181 , \21774 );
and \U$21805 ( \22183 , \21890 , \21745 );
and \U$21806 ( \22184 , \21836 , \21743 );
nor \U$21807 ( \22185 , \22183 , \22184 );
xnor \U$21808 ( \22186 , \22185 , \21715 );
and \U$21809 ( \22187 , \22182 , \22186 );
and \U$21810 ( \22188 , \22018 , \21697 );
and \U$21811 ( \22189 , \21941 , \21695 );
nor \U$21812 ( \22190 , \22188 , \22189 );
xnor \U$21813 ( \22191 , \22190 , \21678 );
and \U$21814 ( \22192 , \22186 , \22191 );
and \U$21815 ( \22193 , \22182 , \22191 );
or \U$21816 ( \22194 , \22187 , \22192 , \22193 );
and \U$21817 ( \22195 , \22178 , \22194 );
and \U$21818 ( \22196 , \22126 , \21660 );
and \U$21819 ( \22197 , \22046 , \21658 );
nor \U$21820 ( \22198 , \22196 , \22197 );
xnor \U$21821 ( \22199 , \22198 , \21665 );
buf \U$21822 ( \22200 , RIc229ba8_142);
and \U$21823 ( \22201 , \22200 , \21654 );
or \U$21824 ( \22202 , \22199 , \22201 );
and \U$21825 ( \22203 , \22194 , \22202 );
and \U$21826 ( \22204 , \22178 , \22202 );
or \U$21827 ( \22205 , \22195 , \22203 , \22204 );
xor \U$21828 ( \22206 , \22092 , \22096 );
xor \U$21829 ( \22207 , \22206 , \22101 );
xor \U$21830 ( \22208 , \22108 , \22112 );
xor \U$21831 ( \22209 , \22208 , \22117 );
and \U$21832 ( \22210 , \22207 , \22209 );
xor \U$21833 ( \22211 , \22125 , \22127 );
and \U$21834 ( \22212 , \22209 , \22211 );
and \U$21835 ( \22213 , \22207 , \22211 );
or \U$21836 ( \22214 , \22210 , \22212 , \22213 );
and \U$21837 ( \22215 , \22205 , \22214 );
xor \U$21838 ( \22216 , \22133 , \22135 );
xor \U$21839 ( \22217 , \22216 , \22137 );
and \U$21840 ( \22218 , \22214 , \22217 );
and \U$21841 ( \22219 , \22205 , \22217 );
or \U$21842 ( \22220 , \22215 , \22218 , \22219 );
xor \U$21843 ( \22221 , \22025 , \22044 );
xor \U$21844 ( \22222 , \22221 , \22048 );
and \U$21845 ( \22223 , \22220 , \22222 );
xor \U$21846 ( \22224 , \22131 , \22140 );
xor \U$21847 ( \22225 , \22224 , \22143 );
and \U$21848 ( \22226 , \22222 , \22225 );
and \U$21849 ( \22227 , \22220 , \22225 );
or \U$21850 ( \22228 , \22223 , \22226 , \22227 );
xor \U$21851 ( \22229 , \22146 , \22148 );
xor \U$21852 ( \22230 , \22229 , \22150 );
and \U$21853 ( \22231 , \22228 , \22230 );
and \U$21854 ( \22232 , \22159 , \22231 );
xor \U$21855 ( \22233 , \22159 , \22231 );
xor \U$21856 ( \22234 , \22228 , \22230 );
buf \U$21857 ( \22235 , RIc226ea8_16);
buf \U$21858 ( \22236 , RIc226e30_17);
and \U$21859 ( \22237 , \22235 , \22236 );
not \U$21860 ( \22238 , \22237 );
and \U$21861 ( \22239 , \22088 , \22238 );
not \U$21862 ( \22240 , \22239 );
and \U$21863 ( \22241 , \21667 , \22163 );
and \U$21864 ( \22242 , \21653 , \22161 );
nor \U$21865 ( \22243 , \22241 , \22242 );
xnor \U$21866 ( \22244 , \22243 , \22091 );
and \U$21867 ( \22245 , \22240 , \22244 );
and \U$21868 ( \22246 , \21706 , \22029 );
and \U$21869 ( \22247 , \21685 , \22027 );
nor \U$21870 ( \22248 , \22246 , \22247 );
xnor \U$21871 ( \22249 , \22248 , \21986 );
and \U$21872 ( \22250 , \22244 , \22249 );
and \U$21873 ( \22251 , \22240 , \22249 );
or \U$21874 ( \22252 , \22245 , \22250 , \22251 );
and \U$21875 ( \22253 , \22046 , \21697 );
and \U$21876 ( \22254 , \22018 , \21695 );
nor \U$21877 ( \22255 , \22253 , \22254 );
xnor \U$21878 ( \22256 , \22255 , \21678 );
and \U$21879 ( \22257 , \22200 , \21660 );
and \U$21880 ( \22258 , \22126 , \21658 );
nor \U$21881 ( \22259 , \22257 , \22258 );
xnor \U$21882 ( \22260 , \22259 , \21665 );
and \U$21883 ( \22261 , \22256 , \22260 );
buf \U$21884 ( \22262 , RIc229c20_143);
and \U$21885 ( \22263 , \22262 , \21654 );
and \U$21886 ( \22264 , \22260 , \22263 );
and \U$21887 ( \22265 , \22256 , \22263 );
or \U$21888 ( \22266 , \22261 , \22264 , \22265 );
and \U$21889 ( \22267 , \22252 , \22266 );
and \U$21890 ( \22268 , \21762 , \21916 );
and \U$21891 ( \22269 , \21754 , \21914 );
nor \U$21892 ( \22270 , \22268 , \22269 );
xnor \U$21893 ( \22271 , \22270 , \21867 );
and \U$21894 ( \22272 , \21836 , \21815 );
and \U$21895 ( \22273 , \21831 , \21813 );
nor \U$21896 ( \22274 , \22272 , \22273 );
xnor \U$21897 ( \22275 , \22274 , \21774 );
and \U$21898 ( \22276 , \22271 , \22275 );
and \U$21899 ( \22277 , \21941 , \21745 );
and \U$21900 ( \22278 , \21890 , \21743 );
nor \U$21901 ( \22279 , \22277 , \22278 );
xnor \U$21902 ( \22280 , \22279 , \21715 );
and \U$21903 ( \22281 , \22275 , \22280 );
and \U$21904 ( \22282 , \22271 , \22280 );
or \U$21905 ( \22283 , \22276 , \22281 , \22282 );
and \U$21906 ( \22284 , \22266 , \22283 );
and \U$21907 ( \22285 , \22252 , \22283 );
or \U$21908 ( \22286 , \22267 , \22284 , \22285 );
xor \U$21909 ( \22287 , \22166 , \22170 );
xor \U$21910 ( \22288 , \22287 , \22175 );
xor \U$21911 ( \22289 , \22182 , \22186 );
xor \U$21912 ( \22290 , \22289 , \22191 );
and \U$21913 ( \22291 , \22288 , \22290 );
xnor \U$21914 ( \22292 , \22199 , \22201 );
and \U$21915 ( \22293 , \22290 , \22292 );
and \U$21916 ( \22294 , \22288 , \22292 );
or \U$21917 ( \22295 , \22291 , \22293 , \22294 );
and \U$21918 ( \22296 , \22286 , \22295 );
xor \U$21919 ( \22297 , \22207 , \22209 );
xor \U$21920 ( \22298 , \22297 , \22211 );
and \U$21921 ( \22299 , \22295 , \22298 );
and \U$21922 ( \22300 , \22286 , \22298 );
or \U$21923 ( \22301 , \22296 , \22299 , \22300 );
xor \U$21924 ( \22302 , \22104 , \22120 );
xor \U$21925 ( \22303 , \22302 , \22128 );
and \U$21926 ( \22304 , \22301 , \22303 );
xor \U$21927 ( \22305 , \22205 , \22214 );
xor \U$21928 ( \22306 , \22305 , \22217 );
and \U$21929 ( \22307 , \22303 , \22306 );
and \U$21930 ( \22308 , \22301 , \22306 );
or \U$21931 ( \22309 , \22304 , \22307 , \22308 );
xor \U$21932 ( \22310 , \22220 , \22222 );
xor \U$21933 ( \22311 , \22310 , \22225 );
and \U$21934 ( \22312 , \22309 , \22311 );
and \U$21935 ( \22313 , \22234 , \22312 );
xor \U$21936 ( \22314 , \22234 , \22312 );
xor \U$21937 ( \22315 , \22309 , \22311 );
and \U$21938 ( \22316 , \22126 , \21697 );
and \U$21939 ( \22317 , \22046 , \21695 );
nor \U$21940 ( \22318 , \22316 , \22317 );
xnor \U$21941 ( \22319 , \22318 , \21678 );
and \U$21942 ( \22320 , \22262 , \21660 );
and \U$21943 ( \22321 , \22200 , \21658 );
nor \U$21944 ( \22322 , \22320 , \22321 );
xnor \U$21945 ( \22323 , \22322 , \21665 );
and \U$21946 ( \22324 , \22319 , \22323 );
buf \U$21947 ( \22325 , RIc229c98_144);
and \U$21948 ( \22326 , \22325 , \21654 );
and \U$21949 ( \22327 , \22323 , \22326 );
and \U$21950 ( \22328 , \22319 , \22326 );
or \U$21951 ( \22329 , \22324 , \22327 , \22328 );
xor \U$21952 ( \22330 , \22088 , \22235 );
xor \U$21953 ( \22331 , \22235 , \22236 );
not \U$21954 ( \22332 , \22331 );
and \U$21955 ( \22333 , \22330 , \22332 );
and \U$21956 ( \22334 , \21653 , \22333 );
not \U$21957 ( \22335 , \22334 );
xnor \U$21958 ( \22336 , \22335 , \22239 );
and \U$21959 ( \22337 , \21685 , \22163 );
and \U$21960 ( \22338 , \21667 , \22161 );
nor \U$21961 ( \22339 , \22337 , \22338 );
xnor \U$21962 ( \22340 , \22339 , \22091 );
and \U$21963 ( \22341 , \22336 , \22340 );
and \U$21964 ( \22342 , \21754 , \22029 );
and \U$21965 ( \22343 , \21706 , \22027 );
nor \U$21966 ( \22344 , \22342 , \22343 );
xnor \U$21967 ( \22345 , \22344 , \21986 );
and \U$21968 ( \22346 , \22340 , \22345 );
and \U$21969 ( \22347 , \22336 , \22345 );
or \U$21970 ( \22348 , \22341 , \22346 , \22347 );
and \U$21971 ( \22349 , \22329 , \22348 );
and \U$21972 ( \22350 , \21831 , \21916 );
and \U$21973 ( \22351 , \21762 , \21914 );
nor \U$21974 ( \22352 , \22350 , \22351 );
xnor \U$21975 ( \22353 , \22352 , \21867 );
and \U$21976 ( \22354 , \21890 , \21815 );
and \U$21977 ( \22355 , \21836 , \21813 );
nor \U$21978 ( \22356 , \22354 , \22355 );
xnor \U$21979 ( \22357 , \22356 , \21774 );
and \U$21980 ( \22358 , \22353 , \22357 );
and \U$21981 ( \22359 , \22018 , \21745 );
and \U$21982 ( \22360 , \21941 , \21743 );
nor \U$21983 ( \22361 , \22359 , \22360 );
xnor \U$21984 ( \22362 , \22361 , \21715 );
and \U$21985 ( \22363 , \22357 , \22362 );
and \U$21986 ( \22364 , \22353 , \22362 );
or \U$21987 ( \22365 , \22358 , \22363 , \22364 );
and \U$21988 ( \22366 , \22348 , \22365 );
and \U$21989 ( \22367 , \22329 , \22365 );
or \U$21990 ( \22368 , \22349 , \22366 , \22367 );
xor \U$21991 ( \22369 , \22240 , \22244 );
xor \U$21992 ( \22370 , \22369 , \22249 );
xor \U$21993 ( \22371 , \22256 , \22260 );
xor \U$21994 ( \22372 , \22371 , \22263 );
and \U$21995 ( \22373 , \22370 , \22372 );
xor \U$21996 ( \22374 , \22271 , \22275 );
xor \U$21997 ( \22375 , \22374 , \22280 );
and \U$21998 ( \22376 , \22372 , \22375 );
and \U$21999 ( \22377 , \22370 , \22375 );
or \U$22000 ( \22378 , \22373 , \22376 , \22377 );
and \U$22001 ( \22379 , \22368 , \22378 );
xor \U$22002 ( \22380 , \22288 , \22290 );
xor \U$22003 ( \22381 , \22380 , \22292 );
and \U$22004 ( \22382 , \22378 , \22381 );
and \U$22005 ( \22383 , \22368 , \22381 );
or \U$22006 ( \22384 , \22379 , \22382 , \22383 );
xor \U$22007 ( \22385 , \22178 , \22194 );
xor \U$22008 ( \22386 , \22385 , \22202 );
and \U$22009 ( \22387 , \22384 , \22386 );
xor \U$22010 ( \22388 , \22286 , \22295 );
xor \U$22011 ( \22389 , \22388 , \22298 );
and \U$22012 ( \22390 , \22386 , \22389 );
and \U$22013 ( \22391 , \22384 , \22389 );
or \U$22014 ( \22392 , \22387 , \22390 , \22391 );
xor \U$22015 ( \22393 , \22301 , \22303 );
xor \U$22016 ( \22394 , \22393 , \22306 );
and \U$22017 ( \22395 , \22392 , \22394 );
and \U$22018 ( \22396 , \22315 , \22395 );
xor \U$22019 ( \22397 , \22315 , \22395 );
xor \U$22020 ( \22398 , \22392 , \22394 );
and \U$22021 ( \22399 , \21762 , \22029 );
and \U$22022 ( \22400 , \21754 , \22027 );
nor \U$22023 ( \22401 , \22399 , \22400 );
xnor \U$22024 ( \22402 , \22401 , \21986 );
and \U$22025 ( \22403 , \21836 , \21916 );
and \U$22026 ( \22404 , \21831 , \21914 );
nor \U$22027 ( \22405 , \22403 , \22404 );
xnor \U$22028 ( \22406 , \22405 , \21867 );
and \U$22029 ( \22407 , \22402 , \22406 );
and \U$22030 ( \22408 , \21941 , \21815 );
and \U$22031 ( \22409 , \21890 , \21813 );
nor \U$22032 ( \22410 , \22408 , \22409 );
xnor \U$22033 ( \22411 , \22410 , \21774 );
and \U$22034 ( \22412 , \22406 , \22411 );
and \U$22035 ( \22413 , \22402 , \22411 );
or \U$22036 ( \22414 , \22407 , \22412 , \22413 );
buf \U$22037 ( \22415 , RIc226db8_18);
buf \U$22038 ( \22416 , RIc226d40_19);
and \U$22039 ( \22417 , \22415 , \22416 );
not \U$22040 ( \22418 , \22417 );
and \U$22041 ( \22419 , \22236 , \22418 );
not \U$22042 ( \22420 , \22419 );
and \U$22043 ( \22421 , \21667 , \22333 );
and \U$22044 ( \22422 , \21653 , \22331 );
nor \U$22045 ( \22423 , \22421 , \22422 );
xnor \U$22046 ( \22424 , \22423 , \22239 );
and \U$22047 ( \22425 , \22420 , \22424 );
and \U$22048 ( \22426 , \21706 , \22163 );
and \U$22049 ( \22427 , \21685 , \22161 );
nor \U$22050 ( \22428 , \22426 , \22427 );
xnor \U$22051 ( \22429 , \22428 , \22091 );
and \U$22052 ( \22430 , \22424 , \22429 );
and \U$22053 ( \22431 , \22420 , \22429 );
or \U$22054 ( \22432 , \22425 , \22430 , \22431 );
and \U$22055 ( \22433 , \22414 , \22432 );
and \U$22056 ( \22434 , \22046 , \21745 );
and \U$22057 ( \22435 , \22018 , \21743 );
nor \U$22058 ( \22436 , \22434 , \22435 );
xnor \U$22059 ( \22437 , \22436 , \21715 );
and \U$22060 ( \22438 , \22200 , \21697 );
and \U$22061 ( \22439 , \22126 , \21695 );
nor \U$22062 ( \22440 , \22438 , \22439 );
xnor \U$22063 ( \22441 , \22440 , \21678 );
and \U$22064 ( \22442 , \22437 , \22441 );
and \U$22065 ( \22443 , \22325 , \21660 );
and \U$22066 ( \22444 , \22262 , \21658 );
nor \U$22067 ( \22445 , \22443 , \22444 );
xnor \U$22068 ( \22446 , \22445 , \21665 );
and \U$22069 ( \22447 , \22441 , \22446 );
and \U$22070 ( \22448 , \22437 , \22446 );
or \U$22071 ( \22449 , \22442 , \22447 , \22448 );
and \U$22072 ( \22450 , \22432 , \22449 );
and \U$22073 ( \22451 , \22414 , \22449 );
or \U$22074 ( \22452 , \22433 , \22450 , \22451 );
xor \U$22075 ( \22453 , \22319 , \22323 );
xor \U$22076 ( \22454 , \22453 , \22326 );
xor \U$22077 ( \22455 , \22353 , \22357 );
xor \U$22078 ( \22456 , \22455 , \22362 );
or \U$22079 ( \22457 , \22454 , \22456 );
and \U$22080 ( \22458 , \22452 , \22457 );
xor \U$22081 ( \22459 , \22370 , \22372 );
xor \U$22082 ( \22460 , \22459 , \22375 );
and \U$22083 ( \22461 , \22457 , \22460 );
and \U$22084 ( \22462 , \22452 , \22460 );
or \U$22085 ( \22463 , \22458 , \22461 , \22462 );
xor \U$22086 ( \22464 , \22252 , \22266 );
xor \U$22087 ( \22465 , \22464 , \22283 );
and \U$22088 ( \22466 , \22463 , \22465 );
xor \U$22089 ( \22467 , \22368 , \22378 );
xor \U$22090 ( \22468 , \22467 , \22381 );
and \U$22091 ( \22469 , \22465 , \22468 );
and \U$22092 ( \22470 , \22463 , \22468 );
or \U$22093 ( \22471 , \22466 , \22469 , \22470 );
xor \U$22094 ( \22472 , \22384 , \22386 );
xor \U$22095 ( \22473 , \22472 , \22389 );
and \U$22096 ( \22474 , \22471 , \22473 );
and \U$22097 ( \22475 , \22398 , \22474 );
xor \U$22098 ( \22476 , \22398 , \22474 );
xor \U$22099 ( \22477 , \22471 , \22473 );
and \U$22100 ( \22478 , \21831 , \22029 );
and \U$22101 ( \22479 , \21762 , \22027 );
nor \U$22102 ( \22480 , \22478 , \22479 );
xnor \U$22103 ( \22481 , \22480 , \21986 );
and \U$22104 ( \22482 , \21890 , \21916 );
and \U$22105 ( \22483 , \21836 , \21914 );
nor \U$22106 ( \22484 , \22482 , \22483 );
xnor \U$22107 ( \22485 , \22484 , \21867 );
and \U$22108 ( \22486 , \22481 , \22485 );
and \U$22109 ( \22487 , \22018 , \21815 );
and \U$22110 ( \22488 , \21941 , \21813 );
nor \U$22111 ( \22489 , \22487 , \22488 );
xnor \U$22112 ( \22490 , \22489 , \21774 );
and \U$22113 ( \22491 , \22485 , \22490 );
and \U$22114 ( \22492 , \22481 , \22490 );
or \U$22115 ( \22493 , \22486 , \22491 , \22492 );
xor \U$22116 ( \22494 , \22236 , \22415 );
xor \U$22117 ( \22495 , \22415 , \22416 );
not \U$22118 ( \22496 , \22495 );
and \U$22119 ( \22497 , \22494 , \22496 );
and \U$22120 ( \22498 , \21653 , \22497 );
not \U$22121 ( \22499 , \22498 );
xnor \U$22122 ( \22500 , \22499 , \22419 );
and \U$22123 ( \22501 , \21685 , \22333 );
and \U$22124 ( \22502 , \21667 , \22331 );
nor \U$22125 ( \22503 , \22501 , \22502 );
xnor \U$22126 ( \22504 , \22503 , \22239 );
and \U$22127 ( \22505 , \22500 , \22504 );
and \U$22128 ( \22506 , \21754 , \22163 );
and \U$22129 ( \22507 , \21706 , \22161 );
nor \U$22130 ( \22508 , \22506 , \22507 );
xnor \U$22131 ( \22509 , \22508 , \22091 );
and \U$22132 ( \22510 , \22504 , \22509 );
and \U$22133 ( \22511 , \22500 , \22509 );
or \U$22134 ( \22512 , \22505 , \22510 , \22511 );
and \U$22135 ( \22513 , \22493 , \22512 );
and \U$22136 ( \22514 , \22126 , \21745 );
and \U$22137 ( \22515 , \22046 , \21743 );
nor \U$22138 ( \22516 , \22514 , \22515 );
xnor \U$22139 ( \22517 , \22516 , \21715 );
and \U$22140 ( \22518 , \22262 , \21697 );
and \U$22141 ( \22519 , \22200 , \21695 );
nor \U$22142 ( \22520 , \22518 , \22519 );
xnor \U$22143 ( \22521 , \22520 , \21678 );
and \U$22144 ( \22522 , \22517 , \22521 );
buf \U$22145 ( \22523 , RIc229d10_145);
and \U$22146 ( \22524 , \22523 , \21660 );
and \U$22147 ( \22525 , \22325 , \21658 );
nor \U$22148 ( \22526 , \22524 , \22525 );
xnor \U$22149 ( \22527 , \22526 , \21665 );
and \U$22150 ( \22528 , \22521 , \22527 );
and \U$22151 ( \22529 , \22517 , \22527 );
or \U$22152 ( \22530 , \22522 , \22528 , \22529 );
and \U$22153 ( \22531 , \22512 , \22530 );
and \U$22154 ( \22532 , \22493 , \22530 );
or \U$22155 ( \22533 , \22513 , \22531 , \22532 );
and \U$22156 ( \22534 , \22523 , \21654 );
xor \U$22157 ( \22535 , \22402 , \22406 );
xor \U$22158 ( \22536 , \22535 , \22411 );
and \U$22159 ( \22537 , \22534 , \22536 );
xor \U$22160 ( \22538 , \22437 , \22441 );
xor \U$22161 ( \22539 , \22538 , \22446 );
and \U$22162 ( \22540 , \22536 , \22539 );
and \U$22163 ( \22541 , \22534 , \22539 );
or \U$22164 ( \22542 , \22537 , \22540 , \22541 );
and \U$22165 ( \22543 , \22533 , \22542 );
xor \U$22166 ( \22544 , \22336 , \22340 );
xor \U$22167 ( \22545 , \22544 , \22345 );
and \U$22168 ( \22546 , \22542 , \22545 );
and \U$22169 ( \22547 , \22533 , \22545 );
or \U$22170 ( \22548 , \22543 , \22546 , \22547 );
xor \U$22171 ( \22549 , \22329 , \22348 );
xor \U$22172 ( \22550 , \22549 , \22365 );
and \U$22173 ( \22551 , \22548 , \22550 );
xor \U$22174 ( \22552 , \22452 , \22457 );
xor \U$22175 ( \22553 , \22552 , \22460 );
and \U$22176 ( \22554 , \22550 , \22553 );
and \U$22177 ( \22555 , \22548 , \22553 );
or \U$22178 ( \22556 , \22551 , \22554 , \22555 );
buf \U$22179 ( \22557 , RIc226cc8_20);
buf \U$22180 ( \22558 , RIc226c50_21);
and \U$22181 ( \22559 , \22557 , \22558 );
not \U$22182 ( \22560 , \22559 );
and \U$22183 ( \22561 , \22416 , \22560 );
not \U$22184 ( \22562 , \22561 );
and \U$22185 ( \22563 , \21667 , \22497 );
and \U$22186 ( \22564 , \21653 , \22495 );
nor \U$22187 ( \22565 , \22563 , \22564 );
xnor \U$22188 ( \22566 , \22565 , \22419 );
and \U$22189 ( \22567 , \22562 , \22566 );
and \U$22190 ( \22568 , \21706 , \22333 );
and \U$22191 ( \22569 , \21685 , \22331 );
nor \U$22192 ( \22570 , \22568 , \22569 );
xnor \U$22193 ( \22571 , \22570 , \22239 );
and \U$22194 ( \22572 , \22566 , \22571 );
and \U$22195 ( \22573 , \22562 , \22571 );
or \U$22196 ( \22574 , \22567 , \22572 , \22573 );
and \U$22197 ( \22575 , \21762 , \22163 );
and \U$22198 ( \22576 , \21754 , \22161 );
nor \U$22199 ( \22577 , \22575 , \22576 );
xnor \U$22200 ( \22578 , \22577 , \22091 );
and \U$22201 ( \22579 , \21836 , \22029 );
and \U$22202 ( \22580 , \21831 , \22027 );
nor \U$22203 ( \22581 , \22579 , \22580 );
xnor \U$22204 ( \22582 , \22581 , \21986 );
and \U$22205 ( \22583 , \22578 , \22582 );
and \U$22206 ( \22584 , \21941 , \21916 );
and \U$22207 ( \22585 , \21890 , \21914 );
nor \U$22208 ( \22586 , \22584 , \22585 );
xnor \U$22209 ( \22587 , \22586 , \21867 );
and \U$22210 ( \22588 , \22582 , \22587 );
and \U$22211 ( \22589 , \22578 , \22587 );
or \U$22212 ( \22590 , \22583 , \22588 , \22589 );
and \U$22213 ( \22591 , \22574 , \22590 );
and \U$22214 ( \22592 , \22046 , \21815 );
and \U$22215 ( \22593 , \22018 , \21813 );
nor \U$22216 ( \22594 , \22592 , \22593 );
xnor \U$22217 ( \22595 , \22594 , \21774 );
and \U$22218 ( \22596 , \22200 , \21745 );
and \U$22219 ( \22597 , \22126 , \21743 );
nor \U$22220 ( \22598 , \22596 , \22597 );
xnor \U$22221 ( \22599 , \22598 , \21715 );
and \U$22222 ( \22600 , \22595 , \22599 );
and \U$22223 ( \22601 , \22325 , \21697 );
and \U$22224 ( \22602 , \22262 , \21695 );
nor \U$22225 ( \22603 , \22601 , \22602 );
xnor \U$22226 ( \22604 , \22603 , \21678 );
and \U$22227 ( \22605 , \22599 , \22604 );
and \U$22228 ( \22606 , \22595 , \22604 );
or \U$22229 ( \22607 , \22600 , \22605 , \22606 );
and \U$22230 ( \22608 , \22590 , \22607 );
and \U$22231 ( \22609 , \22574 , \22607 );
or \U$22232 ( \22610 , \22591 , \22608 , \22609 );
buf \U$22233 ( \22611 , RIc229d88_146);
and \U$22234 ( \22612 , \22611 , \21654 );
xor \U$22235 ( \22613 , \22517 , \22521 );
xor \U$22236 ( \22614 , \22613 , \22527 );
or \U$22237 ( \22615 , \22612 , \22614 );
and \U$22238 ( \22616 , \22610 , \22615 );
xor \U$22239 ( \22617 , \22481 , \22485 );
xor \U$22240 ( \22618 , \22617 , \22490 );
xor \U$22241 ( \22619 , \22500 , \22504 );
xor \U$22242 ( \22620 , \22619 , \22509 );
and \U$22243 ( \22621 , \22618 , \22620 );
and \U$22244 ( \22622 , \22615 , \22621 );
and \U$22245 ( \22623 , \22610 , \22621 );
or \U$22246 ( \22624 , \22616 , \22622 , \22623 );
xor \U$22247 ( \22625 , \22420 , \22424 );
xor \U$22248 ( \22626 , \22625 , \22429 );
xor \U$22249 ( \22627 , \22493 , \22512 );
xor \U$22250 ( \22628 , \22627 , \22530 );
and \U$22251 ( \22629 , \22626 , \22628 );
xor \U$22252 ( \22630 , \22534 , \22536 );
xor \U$22253 ( \22631 , \22630 , \22539 );
and \U$22254 ( \22632 , \22628 , \22631 );
and \U$22255 ( \22633 , \22626 , \22631 );
or \U$22256 ( \22634 , \22629 , \22632 , \22633 );
and \U$22257 ( \22635 , \22624 , \22634 );
xnor \U$22258 ( \22636 , \22454 , \22456 );
and \U$22259 ( \22637 , \22634 , \22636 );
and \U$22260 ( \22638 , \22624 , \22636 );
or \U$22261 ( \22639 , \22635 , \22637 , \22638 );
xor \U$22262 ( \22640 , \22414 , \22432 );
xor \U$22263 ( \22641 , \22640 , \22449 );
xor \U$22264 ( \22642 , \22533 , \22542 );
xor \U$22265 ( \22643 , \22642 , \22545 );
and \U$22266 ( \22644 , \22641 , \22643 );
and \U$22267 ( \22645 , \22639 , \22644 );
xor \U$22268 ( \22646 , \22548 , \22550 );
xor \U$22269 ( \22647 , \22646 , \22553 );
and \U$22270 ( \22648 , \22644 , \22647 );
and \U$22271 ( \22649 , \22639 , \22647 );
or \U$22272 ( \22650 , \22645 , \22648 , \22649 );
and \U$22273 ( \22651 , \22556 , \22650 );
xor \U$22274 ( \22652 , \22463 , \22465 );
xor \U$22275 ( \22653 , \22652 , \22468 );
and \U$22276 ( \22654 , \22650 , \22653 );
and \U$22277 ( \22655 , \22556 , \22653 );
or \U$22278 ( \22656 , \22651 , \22654 , \22655 );
and \U$22279 ( \22657 , \22477 , \22656 );
xor \U$22280 ( \22658 , \22477 , \22656 );
xor \U$22281 ( \22659 , \22556 , \22650 );
xor \U$22282 ( \22660 , \22659 , \22653 );
and \U$22283 ( \22661 , \22126 , \21815 );
and \U$22284 ( \22662 , \22046 , \21813 );
nor \U$22285 ( \22663 , \22661 , \22662 );
xnor \U$22286 ( \22664 , \22663 , \21774 );
and \U$22287 ( \22665 , \22262 , \21745 );
and \U$22288 ( \22666 , \22200 , \21743 );
nor \U$22289 ( \22667 , \22665 , \22666 );
xnor \U$22290 ( \22668 , \22667 , \21715 );
and \U$22291 ( \22669 , \22664 , \22668 );
and \U$22292 ( \22670 , \22523 , \21697 );
and \U$22293 ( \22671 , \22325 , \21695 );
nor \U$22294 ( \22672 , \22670 , \22671 );
xnor \U$22295 ( \22673 , \22672 , \21678 );
and \U$22296 ( \22674 , \22668 , \22673 );
and \U$22297 ( \22675 , \22664 , \22673 );
or \U$22298 ( \22676 , \22669 , \22674 , \22675 );
and \U$22299 ( \22677 , \21831 , \22163 );
and \U$22300 ( \22678 , \21762 , \22161 );
nor \U$22301 ( \22679 , \22677 , \22678 );
xnor \U$22302 ( \22680 , \22679 , \22091 );
and \U$22303 ( \22681 , \21890 , \22029 );
and \U$22304 ( \22682 , \21836 , \22027 );
nor \U$22305 ( \22683 , \22681 , \22682 );
xnor \U$22306 ( \22684 , \22683 , \21986 );
and \U$22307 ( \22685 , \22680 , \22684 );
and \U$22308 ( \22686 , \22018 , \21916 );
and \U$22309 ( \22687 , \21941 , \21914 );
nor \U$22310 ( \22688 , \22686 , \22687 );
xnor \U$22311 ( \22689 , \22688 , \21867 );
and \U$22312 ( \22690 , \22684 , \22689 );
and \U$22313 ( \22691 , \22680 , \22689 );
or \U$22314 ( \22692 , \22685 , \22690 , \22691 );
and \U$22315 ( \22693 , \22676 , \22692 );
xor \U$22316 ( \22694 , \22416 , \22557 );
xor \U$22317 ( \22695 , \22557 , \22558 );
not \U$22318 ( \22696 , \22695 );
and \U$22319 ( \22697 , \22694 , \22696 );
and \U$22320 ( \22698 , \21653 , \22697 );
not \U$22321 ( \22699 , \22698 );
xnor \U$22322 ( \22700 , \22699 , \22561 );
and \U$22323 ( \22701 , \21685 , \22497 );
and \U$22324 ( \22702 , \21667 , \22495 );
nor \U$22325 ( \22703 , \22701 , \22702 );
xnor \U$22326 ( \22704 , \22703 , \22419 );
and \U$22327 ( \22705 , \22700 , \22704 );
and \U$22328 ( \22706 , \21754 , \22333 );
and \U$22329 ( \22707 , \21706 , \22331 );
nor \U$22330 ( \22708 , \22706 , \22707 );
xnor \U$22331 ( \22709 , \22708 , \22239 );
and \U$22332 ( \22710 , \22704 , \22709 );
and \U$22333 ( \22711 , \22700 , \22709 );
or \U$22334 ( \22712 , \22705 , \22710 , \22711 );
and \U$22335 ( \22713 , \22692 , \22712 );
and \U$22336 ( \22714 , \22676 , \22712 );
or \U$22337 ( \22715 , \22693 , \22713 , \22714 );
buf \U$22338 ( \22716 , RIc229e00_147);
and \U$22339 ( \22717 , \22716 , \21660 );
and \U$22340 ( \22718 , \22611 , \21658 );
nor \U$22341 ( \22719 , \22717 , \22718 );
xnor \U$22342 ( \22720 , \22719 , \21665 );
buf \U$22343 ( \22721 , RIc229e78_148);
and \U$22344 ( \22722 , \22721 , \21654 );
or \U$22345 ( \22723 , \22720 , \22722 );
and \U$22346 ( \22724 , \22611 , \21660 );
and \U$22347 ( \22725 , \22523 , \21658 );
nor \U$22348 ( \22726 , \22724 , \22725 );
xnor \U$22349 ( \22727 , \22726 , \21665 );
and \U$22350 ( \22728 , \22723 , \22727 );
and \U$22351 ( \22729 , \22716 , \21654 );
and \U$22352 ( \22730 , \22727 , \22729 );
and \U$22353 ( \22731 , \22723 , \22729 );
or \U$22354 ( \22732 , \22728 , \22730 , \22731 );
and \U$22355 ( \22733 , \22715 , \22732 );
xor \U$22356 ( \22734 , \22562 , \22566 );
xor \U$22357 ( \22735 , \22734 , \22571 );
xor \U$22358 ( \22736 , \22578 , \22582 );
xor \U$22359 ( \22737 , \22736 , \22587 );
and \U$22360 ( \22738 , \22735 , \22737 );
xor \U$22361 ( \22739 , \22595 , \22599 );
xor \U$22362 ( \22740 , \22739 , \22604 );
and \U$22363 ( \22741 , \22737 , \22740 );
and \U$22364 ( \22742 , \22735 , \22740 );
or \U$22365 ( \22743 , \22738 , \22741 , \22742 );
and \U$22366 ( \22744 , \22732 , \22743 );
and \U$22367 ( \22745 , \22715 , \22743 );
or \U$22368 ( \22746 , \22733 , \22744 , \22745 );
xor \U$22369 ( \22747 , \22574 , \22590 );
xor \U$22370 ( \22748 , \22747 , \22607 );
xnor \U$22371 ( \22749 , \22612 , \22614 );
and \U$22372 ( \22750 , \22748 , \22749 );
xor \U$22373 ( \22751 , \22618 , \22620 );
and \U$22374 ( \22752 , \22749 , \22751 );
and \U$22375 ( \22753 , \22748 , \22751 );
or \U$22376 ( \22754 , \22750 , \22752 , \22753 );
and \U$22377 ( \22755 , \22746 , \22754 );
xor \U$22378 ( \22756 , \22626 , \22628 );
xor \U$22379 ( \22757 , \22756 , \22631 );
and \U$22380 ( \22758 , \22754 , \22757 );
and \U$22381 ( \22759 , \22746 , \22757 );
or \U$22382 ( \22760 , \22755 , \22758 , \22759 );
xor \U$22383 ( \22761 , \22624 , \22634 );
xor \U$22384 ( \22762 , \22761 , \22636 );
and \U$22385 ( \22763 , \22760 , \22762 );
xor \U$22386 ( \22764 , \22641 , \22643 );
and \U$22387 ( \22765 , \22762 , \22764 );
and \U$22388 ( \22766 , \22760 , \22764 );
or \U$22389 ( \22767 , \22763 , \22765 , \22766 );
xor \U$22390 ( \22768 , \22639 , \22644 );
xor \U$22391 ( \22769 , \22768 , \22647 );
and \U$22392 ( \22770 , \22767 , \22769 );
and \U$22393 ( \22771 , \22660 , \22770 );
xor \U$22394 ( \22772 , \22660 , \22770 );
xor \U$22395 ( \22773 , \22767 , \22769 );
buf \U$22396 ( \22774 , RIc226bd8_22);
buf \U$22397 ( \22775 , RIc226b60_23);
and \U$22398 ( \22776 , \22774 , \22775 );
not \U$22399 ( \22777 , \22776 );
and \U$22400 ( \22778 , \22558 , \22777 );
not \U$22401 ( \22779 , \22778 );
and \U$22402 ( \22780 , \21667 , \22697 );
and \U$22403 ( \22781 , \21653 , \22695 );
nor \U$22404 ( \22782 , \22780 , \22781 );
xnor \U$22405 ( \22783 , \22782 , \22561 );
and \U$22406 ( \22784 , \22779 , \22783 );
and \U$22407 ( \22785 , \21706 , \22497 );
and \U$22408 ( \22786 , \21685 , \22495 );
nor \U$22409 ( \22787 , \22785 , \22786 );
xnor \U$22410 ( \22788 , \22787 , \22419 );
and \U$22411 ( \22789 , \22783 , \22788 );
and \U$22412 ( \22790 , \22779 , \22788 );
or \U$22413 ( \22791 , \22784 , \22789 , \22790 );
and \U$22414 ( \22792 , \22046 , \21916 );
and \U$22415 ( \22793 , \22018 , \21914 );
nor \U$22416 ( \22794 , \22792 , \22793 );
xnor \U$22417 ( \22795 , \22794 , \21867 );
and \U$22418 ( \22796 , \22200 , \21815 );
and \U$22419 ( \22797 , \22126 , \21813 );
nor \U$22420 ( \22798 , \22796 , \22797 );
xnor \U$22421 ( \22799 , \22798 , \21774 );
and \U$22422 ( \22800 , \22795 , \22799 );
and \U$22423 ( \22801 , \22325 , \21745 );
and \U$22424 ( \22802 , \22262 , \21743 );
nor \U$22425 ( \22803 , \22801 , \22802 );
xnor \U$22426 ( \22804 , \22803 , \21715 );
and \U$22427 ( \22805 , \22799 , \22804 );
and \U$22428 ( \22806 , \22795 , \22804 );
or \U$22429 ( \22807 , \22800 , \22805 , \22806 );
and \U$22430 ( \22808 , \22791 , \22807 );
and \U$22431 ( \22809 , \21762 , \22333 );
and \U$22432 ( \22810 , \21754 , \22331 );
nor \U$22433 ( \22811 , \22809 , \22810 );
xnor \U$22434 ( \22812 , \22811 , \22239 );
and \U$22435 ( \22813 , \21836 , \22163 );
and \U$22436 ( \22814 , \21831 , \22161 );
nor \U$22437 ( \22815 , \22813 , \22814 );
xnor \U$22438 ( \22816 , \22815 , \22091 );
and \U$22439 ( \22817 , \22812 , \22816 );
and \U$22440 ( \22818 , \21941 , \22029 );
and \U$22441 ( \22819 , \21890 , \22027 );
nor \U$22442 ( \22820 , \22818 , \22819 );
xnor \U$22443 ( \22821 , \22820 , \21986 );
and \U$22444 ( \22822 , \22816 , \22821 );
and \U$22445 ( \22823 , \22812 , \22821 );
or \U$22446 ( \22824 , \22817 , \22822 , \22823 );
and \U$22447 ( \22825 , \22807 , \22824 );
and \U$22448 ( \22826 , \22791 , \22824 );
or \U$22449 ( \22827 , \22808 , \22825 , \22826 );
and \U$22450 ( \22828 , \22611 , \21697 );
and \U$22451 ( \22829 , \22523 , \21695 );
nor \U$22452 ( \22830 , \22828 , \22829 );
xnor \U$22453 ( \22831 , \22830 , \21678 );
and \U$22454 ( \22832 , \22721 , \21660 );
and \U$22455 ( \22833 , \22716 , \21658 );
nor \U$22456 ( \22834 , \22832 , \22833 );
xnor \U$22457 ( \22835 , \22834 , \21665 );
and \U$22458 ( \22836 , \22831 , \22835 );
buf \U$22459 ( \22837 , RIc229ef0_149);
and \U$22460 ( \22838 , \22837 , \21654 );
and \U$22461 ( \22839 , \22835 , \22838 );
and \U$22462 ( \22840 , \22831 , \22838 );
or \U$22463 ( \22841 , \22836 , \22839 , \22840 );
xor \U$22464 ( \22842 , \22664 , \22668 );
xor \U$22465 ( \22843 , \22842 , \22673 );
and \U$22466 ( \22844 , \22841 , \22843 );
xnor \U$22467 ( \22845 , \22720 , \22722 );
and \U$22468 ( \22846 , \22843 , \22845 );
and \U$22469 ( \22847 , \22841 , \22845 );
or \U$22470 ( \22848 , \22844 , \22846 , \22847 );
and \U$22471 ( \22849 , \22827 , \22848 );
xor \U$22472 ( \22850 , \22680 , \22684 );
xor \U$22473 ( \22851 , \22850 , \22689 );
xor \U$22474 ( \22852 , \22700 , \22704 );
xor \U$22475 ( \22853 , \22852 , \22709 );
and \U$22476 ( \22854 , \22851 , \22853 );
and \U$22477 ( \22855 , \22848 , \22854 );
and \U$22478 ( \22856 , \22827 , \22854 );
or \U$22479 ( \22857 , \22849 , \22855 , \22856 );
xor \U$22480 ( \22858 , \22676 , \22692 );
xor \U$22481 ( \22859 , \22858 , \22712 );
xor \U$22482 ( \22860 , \22723 , \22727 );
xor \U$22483 ( \22861 , \22860 , \22729 );
and \U$22484 ( \22862 , \22859 , \22861 );
xor \U$22485 ( \22863 , \22735 , \22737 );
xor \U$22486 ( \22864 , \22863 , \22740 );
and \U$22487 ( \22865 , \22861 , \22864 );
and \U$22488 ( \22866 , \22859 , \22864 );
or \U$22489 ( \22867 , \22862 , \22865 , \22866 );
and \U$22490 ( \22868 , \22857 , \22867 );
xor \U$22491 ( \22869 , \22748 , \22749 );
xor \U$22492 ( \22870 , \22869 , \22751 );
and \U$22493 ( \22871 , \22867 , \22870 );
and \U$22494 ( \22872 , \22857 , \22870 );
or \U$22495 ( \22873 , \22868 , \22871 , \22872 );
xor \U$22496 ( \22874 , \22610 , \22615 );
xor \U$22497 ( \22875 , \22874 , \22621 );
and \U$22498 ( \22876 , \22873 , \22875 );
xor \U$22499 ( \22877 , \22746 , \22754 );
xor \U$22500 ( \22878 , \22877 , \22757 );
and \U$22501 ( \22879 , \22875 , \22878 );
and \U$22502 ( \22880 , \22873 , \22878 );
or \U$22503 ( \22881 , \22876 , \22879 , \22880 );
xor \U$22504 ( \22882 , \22760 , \22762 );
xor \U$22505 ( \22883 , \22882 , \22764 );
and \U$22506 ( \22884 , \22881 , \22883 );
and \U$22507 ( \22885 , \22773 , \22884 );
xor \U$22508 ( \22886 , \22773 , \22884 );
xor \U$22509 ( \22887 , \22881 , \22883 );
xor \U$22510 ( \22888 , \22558 , \22774 );
xor \U$22511 ( \22889 , \22774 , \22775 );
not \U$22512 ( \22890 , \22889 );
and \U$22513 ( \22891 , \22888 , \22890 );
and \U$22514 ( \22892 , \21653 , \22891 );
not \U$22515 ( \22893 , \22892 );
xnor \U$22516 ( \22894 , \22893 , \22778 );
and \U$22517 ( \22895 , \21685 , \22697 );
and \U$22518 ( \22896 , \21667 , \22695 );
nor \U$22519 ( \22897 , \22895 , \22896 );
xnor \U$22520 ( \22898 , \22897 , \22561 );
and \U$22521 ( \22899 , \22894 , \22898 );
and \U$22522 ( \22900 , \21754 , \22497 );
and \U$22523 ( \22901 , \21706 , \22495 );
nor \U$22524 ( \22902 , \22900 , \22901 );
xnor \U$22525 ( \22903 , \22902 , \22419 );
and \U$22526 ( \22904 , \22898 , \22903 );
and \U$22527 ( \22905 , \22894 , \22903 );
or \U$22528 ( \22906 , \22899 , \22904 , \22905 );
and \U$22529 ( \22907 , \22126 , \21916 );
and \U$22530 ( \22908 , \22046 , \21914 );
nor \U$22531 ( \22909 , \22907 , \22908 );
xnor \U$22532 ( \22910 , \22909 , \21867 );
and \U$22533 ( \22911 , \22262 , \21815 );
and \U$22534 ( \22912 , \22200 , \21813 );
nor \U$22535 ( \22913 , \22911 , \22912 );
xnor \U$22536 ( \22914 , \22913 , \21774 );
and \U$22537 ( \22915 , \22910 , \22914 );
and \U$22538 ( \22916 , \22523 , \21745 );
and \U$22539 ( \22917 , \22325 , \21743 );
nor \U$22540 ( \22918 , \22916 , \22917 );
xnor \U$22541 ( \22919 , \22918 , \21715 );
and \U$22542 ( \22920 , \22914 , \22919 );
and \U$22543 ( \22921 , \22910 , \22919 );
or \U$22544 ( \22922 , \22915 , \22920 , \22921 );
and \U$22545 ( \22923 , \22906 , \22922 );
and \U$22546 ( \22924 , \21831 , \22333 );
and \U$22547 ( \22925 , \21762 , \22331 );
nor \U$22548 ( \22926 , \22924 , \22925 );
xnor \U$22549 ( \22927 , \22926 , \22239 );
and \U$22550 ( \22928 , \21890 , \22163 );
and \U$22551 ( \22929 , \21836 , \22161 );
nor \U$22552 ( \22930 , \22928 , \22929 );
xnor \U$22553 ( \22931 , \22930 , \22091 );
and \U$22554 ( \22932 , \22927 , \22931 );
and \U$22555 ( \22933 , \22018 , \22029 );
and \U$22556 ( \22934 , \21941 , \22027 );
nor \U$22557 ( \22935 , \22933 , \22934 );
xnor \U$22558 ( \22936 , \22935 , \21986 );
and \U$22559 ( \22937 , \22931 , \22936 );
and \U$22560 ( \22938 , \22927 , \22936 );
or \U$22561 ( \22939 , \22932 , \22937 , \22938 );
and \U$22562 ( \22940 , \22922 , \22939 );
and \U$22563 ( \22941 , \22906 , \22939 );
or \U$22564 ( \22942 , \22923 , \22940 , \22941 );
and \U$22565 ( \22943 , \22716 , \21697 );
and \U$22566 ( \22944 , \22611 , \21695 );
nor \U$22567 ( \22945 , \22943 , \22944 );
xnor \U$22568 ( \22946 , \22945 , \21678 );
and \U$22569 ( \22947 , \22837 , \21660 );
and \U$22570 ( \22948 , \22721 , \21658 );
nor \U$22571 ( \22949 , \22947 , \22948 );
xnor \U$22572 ( \22950 , \22949 , \21665 );
and \U$22573 ( \22951 , \22946 , \22950 );
buf \U$22574 ( \22952 , RIc229f68_150);
and \U$22575 ( \22953 , \22952 , \21654 );
and \U$22576 ( \22954 , \22950 , \22953 );
and \U$22577 ( \22955 , \22946 , \22953 );
or \U$22578 ( \22956 , \22951 , \22954 , \22955 );
xor \U$22579 ( \22957 , \22831 , \22835 );
xor \U$22580 ( \22958 , \22957 , \22838 );
and \U$22581 ( \22959 , \22956 , \22958 );
xor \U$22582 ( \22960 , \22795 , \22799 );
xor \U$22583 ( \22961 , \22960 , \22804 );
and \U$22584 ( \22962 , \22958 , \22961 );
and \U$22585 ( \22963 , \22956 , \22961 );
or \U$22586 ( \22964 , \22959 , \22962 , \22963 );
and \U$22587 ( \22965 , \22942 , \22964 );
xor \U$22588 ( \22966 , \22779 , \22783 );
xor \U$22589 ( \22967 , \22966 , \22788 );
xor \U$22590 ( \22968 , \22812 , \22816 );
xor \U$22591 ( \22969 , \22968 , \22821 );
and \U$22592 ( \22970 , \22967 , \22969 );
and \U$22593 ( \22971 , \22964 , \22970 );
and \U$22594 ( \22972 , \22942 , \22970 );
or \U$22595 ( \22973 , \22965 , \22971 , \22972 );
xor \U$22596 ( \22974 , \22791 , \22807 );
xor \U$22597 ( \22975 , \22974 , \22824 );
xor \U$22598 ( \22976 , \22841 , \22843 );
xor \U$22599 ( \22977 , \22976 , \22845 );
and \U$22600 ( \22978 , \22975 , \22977 );
xor \U$22601 ( \22979 , \22851 , \22853 );
and \U$22602 ( \22980 , \22977 , \22979 );
and \U$22603 ( \22981 , \22975 , \22979 );
or \U$22604 ( \22982 , \22978 , \22980 , \22981 );
and \U$22605 ( \22983 , \22973 , \22982 );
xor \U$22606 ( \22984 , \22859 , \22861 );
xor \U$22607 ( \22985 , \22984 , \22864 );
and \U$22608 ( \22986 , \22982 , \22985 );
and \U$22609 ( \22987 , \22973 , \22985 );
or \U$22610 ( \22988 , \22983 , \22986 , \22987 );
xor \U$22611 ( \22989 , \22715 , \22732 );
xor \U$22612 ( \22990 , \22989 , \22743 );
and \U$22613 ( \22991 , \22988 , \22990 );
xor \U$22614 ( \22992 , \22857 , \22867 );
xor \U$22615 ( \22993 , \22992 , \22870 );
and \U$22616 ( \22994 , \22990 , \22993 );
and \U$22617 ( \22995 , \22988 , \22993 );
or \U$22618 ( \22996 , \22991 , \22994 , \22995 );
xor \U$22619 ( \22997 , \22873 , \22875 );
xor \U$22620 ( \22998 , \22997 , \22878 );
and \U$22621 ( \22999 , \22996 , \22998 );
and \U$22622 ( \23000 , \22887 , \22999 );
xor \U$22623 ( \23001 , \22887 , \22999 );
xor \U$22624 ( \23002 , \22996 , \22998 );
buf \U$22625 ( \23003 , RIc226ae8_24);
buf \U$22626 ( \23004 , RIc226a70_25);
and \U$22627 ( \23005 , \23003 , \23004 );
not \U$22628 ( \23006 , \23005 );
and \U$22629 ( \23007 , \22775 , \23006 );
not \U$22630 ( \23008 , \23007 );
and \U$22631 ( \23009 , \21667 , \22891 );
and \U$22632 ( \23010 , \21653 , \22889 );
nor \U$22633 ( \23011 , \23009 , \23010 );
xnor \U$22634 ( \23012 , \23011 , \22778 );
and \U$22635 ( \23013 , \23008 , \23012 );
and \U$22636 ( \23014 , \21706 , \22697 );
and \U$22637 ( \23015 , \21685 , \22695 );
nor \U$22638 ( \23016 , \23014 , \23015 );
xnor \U$22639 ( \23017 , \23016 , \22561 );
and \U$22640 ( \23018 , \23012 , \23017 );
and \U$22641 ( \23019 , \23008 , \23017 );
or \U$22642 ( \23020 , \23013 , \23018 , \23019 );
and \U$22643 ( \23021 , \21762 , \22497 );
and \U$22644 ( \23022 , \21754 , \22495 );
nor \U$22645 ( \23023 , \23021 , \23022 );
xnor \U$22646 ( \23024 , \23023 , \22419 );
and \U$22647 ( \23025 , \21836 , \22333 );
and \U$22648 ( \23026 , \21831 , \22331 );
nor \U$22649 ( \23027 , \23025 , \23026 );
xnor \U$22650 ( \23028 , \23027 , \22239 );
and \U$22651 ( \23029 , \23024 , \23028 );
and \U$22652 ( \23030 , \21941 , \22163 );
and \U$22653 ( \23031 , \21890 , \22161 );
nor \U$22654 ( \23032 , \23030 , \23031 );
xnor \U$22655 ( \23033 , \23032 , \22091 );
and \U$22656 ( \23034 , \23028 , \23033 );
and \U$22657 ( \23035 , \23024 , \23033 );
or \U$22658 ( \23036 , \23029 , \23034 , \23035 );
and \U$22659 ( \23037 , \23020 , \23036 );
and \U$22660 ( \23038 , \22046 , \22029 );
and \U$22661 ( \23039 , \22018 , \22027 );
nor \U$22662 ( \23040 , \23038 , \23039 );
xnor \U$22663 ( \23041 , \23040 , \21986 );
and \U$22664 ( \23042 , \22200 , \21916 );
and \U$22665 ( \23043 , \22126 , \21914 );
nor \U$22666 ( \23044 , \23042 , \23043 );
xnor \U$22667 ( \23045 , \23044 , \21867 );
and \U$22668 ( \23046 , \23041 , \23045 );
and \U$22669 ( \23047 , \22325 , \21815 );
and \U$22670 ( \23048 , \22262 , \21813 );
nor \U$22671 ( \23049 , \23047 , \23048 );
xnor \U$22672 ( \23050 , \23049 , \21774 );
and \U$22673 ( \23051 , \23045 , \23050 );
and \U$22674 ( \23052 , \23041 , \23050 );
or \U$22675 ( \23053 , \23046 , \23051 , \23052 );
and \U$22676 ( \23054 , \23036 , \23053 );
and \U$22677 ( \23055 , \23020 , \23053 );
or \U$22678 ( \23056 , \23037 , \23054 , \23055 );
xor \U$22679 ( \23057 , \22894 , \22898 );
xor \U$22680 ( \23058 , \23057 , \22903 );
xor \U$22681 ( \23059 , \22910 , \22914 );
xor \U$22682 ( \23060 , \23059 , \22919 );
and \U$22683 ( \23061 , \23058 , \23060 );
xor \U$22684 ( \23062 , \22927 , \22931 );
xor \U$22685 ( \23063 , \23062 , \22936 );
and \U$22686 ( \23064 , \23060 , \23063 );
and \U$22687 ( \23065 , \23058 , \23063 );
or \U$22688 ( \23066 , \23061 , \23064 , \23065 );
and \U$22689 ( \23067 , \23056 , \23066 );
and \U$22690 ( \23068 , \22611 , \21745 );
and \U$22691 ( \23069 , \22523 , \21743 );
nor \U$22692 ( \23070 , \23068 , \23069 );
xnor \U$22693 ( \23071 , \23070 , \21715 );
and \U$22694 ( \23072 , \22721 , \21697 );
and \U$22695 ( \23073 , \22716 , \21695 );
nor \U$22696 ( \23074 , \23072 , \23073 );
xnor \U$22697 ( \23075 , \23074 , \21678 );
and \U$22698 ( \23076 , \23071 , \23075 );
and \U$22699 ( \23077 , \22952 , \21660 );
and \U$22700 ( \23078 , \22837 , \21658 );
nor \U$22701 ( \23079 , \23077 , \23078 );
xnor \U$22702 ( \23080 , \23079 , \21665 );
and \U$22703 ( \23081 , \23075 , \23080 );
and \U$22704 ( \23082 , \23071 , \23080 );
or \U$22705 ( \23083 , \23076 , \23081 , \23082 );
xor \U$22706 ( \23084 , \22946 , \22950 );
xor \U$22707 ( \23085 , \23084 , \22953 );
or \U$22708 ( \23086 , \23083 , \23085 );
and \U$22709 ( \23087 , \23066 , \23086 );
and \U$22710 ( \23088 , \23056 , \23086 );
or \U$22711 ( \23089 , \23067 , \23087 , \23088 );
xor \U$22712 ( \23090 , \22906 , \22922 );
xor \U$22713 ( \23091 , \23090 , \22939 );
xor \U$22714 ( \23092 , \22956 , \22958 );
xor \U$22715 ( \23093 , \23092 , \22961 );
and \U$22716 ( \23094 , \23091 , \23093 );
xor \U$22717 ( \23095 , \22967 , \22969 );
and \U$22718 ( \23096 , \23093 , \23095 );
and \U$22719 ( \23097 , \23091 , \23095 );
or \U$22720 ( \23098 , \23094 , \23096 , \23097 );
and \U$22721 ( \23099 , \23089 , \23098 );
xor \U$22722 ( \23100 , \22975 , \22977 );
xor \U$22723 ( \23101 , \23100 , \22979 );
and \U$22724 ( \23102 , \23098 , \23101 );
and \U$22725 ( \23103 , \23089 , \23101 );
or \U$22726 ( \23104 , \23099 , \23102 , \23103 );
xor \U$22727 ( \23105 , \22827 , \22848 );
xor \U$22728 ( \23106 , \23105 , \22854 );
and \U$22729 ( \23107 , \23104 , \23106 );
xor \U$22730 ( \23108 , \22973 , \22982 );
xor \U$22731 ( \23109 , \23108 , \22985 );
and \U$22732 ( \23110 , \23106 , \23109 );
and \U$22733 ( \23111 , \23104 , \23109 );
or \U$22734 ( \23112 , \23107 , \23110 , \23111 );
xor \U$22735 ( \23113 , \22988 , \22990 );
xor \U$22736 ( \23114 , \23113 , \22993 );
and \U$22737 ( \23115 , \23112 , \23114 );
and \U$22738 ( \23116 , \23002 , \23115 );
xor \U$22739 ( \23117 , \23002 , \23115 );
xor \U$22740 ( \23118 , \23112 , \23114 );
and \U$22741 ( \23119 , \22716 , \21745 );
and \U$22742 ( \23120 , \22611 , \21743 );
nor \U$22743 ( \23121 , \23119 , \23120 );
xnor \U$22744 ( \23122 , \23121 , \21715 );
and \U$22745 ( \23123 , \22837 , \21697 );
and \U$22746 ( \23124 , \22721 , \21695 );
nor \U$22747 ( \23125 , \23123 , \23124 );
xnor \U$22748 ( \23126 , \23125 , \21678 );
and \U$22749 ( \23127 , \23122 , \23126 );
buf \U$22750 ( \23128 , RIc229fe0_151);
and \U$22751 ( \23129 , \23128 , \21660 );
and \U$22752 ( \23130 , \22952 , \21658 );
nor \U$22753 ( \23131 , \23129 , \23130 );
xnor \U$22754 ( \23132 , \23131 , \21665 );
and \U$22755 ( \23133 , \23126 , \23132 );
and \U$22756 ( \23134 , \23122 , \23132 );
or \U$22757 ( \23135 , \23127 , \23133 , \23134 );
buf \U$22758 ( \23136 , RIc22a058_152);
and \U$22759 ( \23137 , \23136 , \21654 );
buf \U$22760 ( \23138 , \23137 );
and \U$22761 ( \23139 , \23135 , \23138 );
and \U$22762 ( \23140 , \23128 , \21654 );
and \U$22763 ( \23141 , \23138 , \23140 );
and \U$22764 ( \23142 , \23135 , \23140 );
or \U$22765 ( \23143 , \23139 , \23141 , \23142 );
and \U$22766 ( \23144 , \21831 , \22497 );
and \U$22767 ( \23145 , \21762 , \22495 );
nor \U$22768 ( \23146 , \23144 , \23145 );
xnor \U$22769 ( \23147 , \23146 , \22419 );
and \U$22770 ( \23148 , \21890 , \22333 );
and \U$22771 ( \23149 , \21836 , \22331 );
nor \U$22772 ( \23150 , \23148 , \23149 );
xnor \U$22773 ( \23151 , \23150 , \22239 );
and \U$22774 ( \23152 , \23147 , \23151 );
and \U$22775 ( \23153 , \22018 , \22163 );
and \U$22776 ( \23154 , \21941 , \22161 );
nor \U$22777 ( \23155 , \23153 , \23154 );
xnor \U$22778 ( \23156 , \23155 , \22091 );
and \U$22779 ( \23157 , \23151 , \23156 );
and \U$22780 ( \23158 , \23147 , \23156 );
or \U$22781 ( \23159 , \23152 , \23157 , \23158 );
xor \U$22782 ( \23160 , \22775 , \23003 );
xor \U$22783 ( \23161 , \23003 , \23004 );
not \U$22784 ( \23162 , \23161 );
and \U$22785 ( \23163 , \23160 , \23162 );
and \U$22786 ( \23164 , \21653 , \23163 );
not \U$22787 ( \23165 , \23164 );
xnor \U$22788 ( \23166 , \23165 , \23007 );
and \U$22789 ( \23167 , \21685 , \22891 );
and \U$22790 ( \23168 , \21667 , \22889 );
nor \U$22791 ( \23169 , \23167 , \23168 );
xnor \U$22792 ( \23170 , \23169 , \22778 );
and \U$22793 ( \23171 , \23166 , \23170 );
and \U$22794 ( \23172 , \21754 , \22697 );
and \U$22795 ( \23173 , \21706 , \22695 );
nor \U$22796 ( \23174 , \23172 , \23173 );
xnor \U$22797 ( \23175 , \23174 , \22561 );
and \U$22798 ( \23176 , \23170 , \23175 );
and \U$22799 ( \23177 , \23166 , \23175 );
or \U$22800 ( \23178 , \23171 , \23176 , \23177 );
and \U$22801 ( \23179 , \23159 , \23178 );
and \U$22802 ( \23180 , \22126 , \22029 );
and \U$22803 ( \23181 , \22046 , \22027 );
nor \U$22804 ( \23182 , \23180 , \23181 );
xnor \U$22805 ( \23183 , \23182 , \21986 );
and \U$22806 ( \23184 , \22262 , \21916 );
and \U$22807 ( \23185 , \22200 , \21914 );
nor \U$22808 ( \23186 , \23184 , \23185 );
xnor \U$22809 ( \23187 , \23186 , \21867 );
and \U$22810 ( \23188 , \23183 , \23187 );
and \U$22811 ( \23189 , \22523 , \21815 );
and \U$22812 ( \23190 , \22325 , \21813 );
nor \U$22813 ( \23191 , \23189 , \23190 );
xnor \U$22814 ( \23192 , \23191 , \21774 );
and \U$22815 ( \23193 , \23187 , \23192 );
and \U$22816 ( \23194 , \23183 , \23192 );
or \U$22817 ( \23195 , \23188 , \23193 , \23194 );
and \U$22818 ( \23196 , \23178 , \23195 );
and \U$22819 ( \23197 , \23159 , \23195 );
or \U$22820 ( \23198 , \23179 , \23196 , \23197 );
and \U$22821 ( \23199 , \23143 , \23198 );
xor \U$22822 ( \23200 , \23024 , \23028 );
xor \U$22823 ( \23201 , \23200 , \23033 );
xor \U$22824 ( \23202 , \23071 , \23075 );
xor \U$22825 ( \23203 , \23202 , \23080 );
and \U$22826 ( \23204 , \23201 , \23203 );
xor \U$22827 ( \23205 , \23041 , \23045 );
xor \U$22828 ( \23206 , \23205 , \23050 );
and \U$22829 ( \23207 , \23203 , \23206 );
and \U$22830 ( \23208 , \23201 , \23206 );
or \U$22831 ( \23209 , \23204 , \23207 , \23208 );
and \U$22832 ( \23210 , \23198 , \23209 );
and \U$22833 ( \23211 , \23143 , \23209 );
or \U$22834 ( \23212 , \23199 , \23210 , \23211 );
xor \U$22835 ( \23213 , \23020 , \23036 );
xor \U$22836 ( \23214 , \23213 , \23053 );
xor \U$22837 ( \23215 , \23058 , \23060 );
xor \U$22838 ( \23216 , \23215 , \23063 );
and \U$22839 ( \23217 , \23214 , \23216 );
xnor \U$22840 ( \23218 , \23083 , \23085 );
and \U$22841 ( \23219 , \23216 , \23218 );
and \U$22842 ( \23220 , \23214 , \23218 );
or \U$22843 ( \23221 , \23217 , \23219 , \23220 );
and \U$22844 ( \23222 , \23212 , \23221 );
xor \U$22845 ( \23223 , \23091 , \23093 );
xor \U$22846 ( \23224 , \23223 , \23095 );
and \U$22847 ( \23225 , \23221 , \23224 );
and \U$22848 ( \23226 , \23212 , \23224 );
or \U$22849 ( \23227 , \23222 , \23225 , \23226 );
xor \U$22850 ( \23228 , \22942 , \22964 );
xor \U$22851 ( \23229 , \23228 , \22970 );
and \U$22852 ( \23230 , \23227 , \23229 );
xor \U$22853 ( \23231 , \23089 , \23098 );
xor \U$22854 ( \23232 , \23231 , \23101 );
and \U$22855 ( \23233 , \23229 , \23232 );
and \U$22856 ( \23234 , \23227 , \23232 );
or \U$22857 ( \23235 , \23230 , \23233 , \23234 );
xor \U$22858 ( \23236 , \23104 , \23106 );
xor \U$22859 ( \23237 , \23236 , \23109 );
and \U$22860 ( \23238 , \23235 , \23237 );
and \U$22861 ( \23239 , \23118 , \23238 );
xor \U$22862 ( \23240 , \23118 , \23238 );
xor \U$22863 ( \23241 , \23235 , \23237 );
and \U$22864 ( \23242 , \22046 , \22163 );
and \U$22865 ( \23243 , \22018 , \22161 );
nor \U$22866 ( \23244 , \23242 , \23243 );
xnor \U$22867 ( \23245 , \23244 , \22091 );
and \U$22868 ( \23246 , \22200 , \22029 );
and \U$22869 ( \23247 , \22126 , \22027 );
nor \U$22870 ( \23248 , \23246 , \23247 );
xnor \U$22871 ( \23249 , \23248 , \21986 );
and \U$22872 ( \23250 , \23245 , \23249 );
and \U$22873 ( \23251 , \22325 , \21916 );
and \U$22874 ( \23252 , \22262 , \21914 );
nor \U$22875 ( \23253 , \23251 , \23252 );
xnor \U$22876 ( \23254 , \23253 , \21867 );
and \U$22877 ( \23255 , \23249 , \23254 );
and \U$22878 ( \23256 , \23245 , \23254 );
or \U$22879 ( \23257 , \23250 , \23255 , \23256 );
and \U$22880 ( \23258 , \21762 , \22697 );
and \U$22881 ( \23259 , \21754 , \22695 );
nor \U$22882 ( \23260 , \23258 , \23259 );
xnor \U$22883 ( \23261 , \23260 , \22561 );
and \U$22884 ( \23262 , \21836 , \22497 );
and \U$22885 ( \23263 , \21831 , \22495 );
nor \U$22886 ( \23264 , \23262 , \23263 );
xnor \U$22887 ( \23265 , \23264 , \22419 );
and \U$22888 ( \23266 , \23261 , \23265 );
and \U$22889 ( \23267 , \21941 , \22333 );
and \U$22890 ( \23268 , \21890 , \22331 );
nor \U$22891 ( \23269 , \23267 , \23268 );
xnor \U$22892 ( \23270 , \23269 , \22239 );
and \U$22893 ( \23271 , \23265 , \23270 );
and \U$22894 ( \23272 , \23261 , \23270 );
or \U$22895 ( \23273 , \23266 , \23271 , \23272 );
and \U$22896 ( \23274 , \23257 , \23273 );
buf \U$22897 ( \23275 , RIc2269f8_26);
buf \U$22898 ( \23276 , RIc226980_27);
and \U$22899 ( \23277 , \23275 , \23276 );
not \U$22900 ( \23278 , \23277 );
and \U$22901 ( \23279 , \23004 , \23278 );
not \U$22902 ( \23280 , \23279 );
and \U$22903 ( \23281 , \21667 , \23163 );
and \U$22904 ( \23282 , \21653 , \23161 );
nor \U$22905 ( \23283 , \23281 , \23282 );
xnor \U$22906 ( \23284 , \23283 , \23007 );
and \U$22907 ( \23285 , \23280 , \23284 );
and \U$22908 ( \23286 , \21706 , \22891 );
and \U$22909 ( \23287 , \21685 , \22889 );
nor \U$22910 ( \23288 , \23286 , \23287 );
xnor \U$22911 ( \23289 , \23288 , \22778 );
and \U$22912 ( \23290 , \23284 , \23289 );
and \U$22913 ( \23291 , \23280 , \23289 );
or \U$22914 ( \23292 , \23285 , \23290 , \23291 );
and \U$22915 ( \23293 , \23273 , \23292 );
and \U$22916 ( \23294 , \23257 , \23292 );
or \U$22917 ( \23295 , \23274 , \23293 , \23294 );
xor \U$22918 ( \23296 , \23147 , \23151 );
xor \U$22919 ( \23297 , \23296 , \23156 );
xor \U$22920 ( \23298 , \23166 , \23170 );
xor \U$22921 ( \23299 , \23298 , \23175 );
and \U$22922 ( \23300 , \23297 , \23299 );
xor \U$22923 ( \23301 , \23183 , \23187 );
xor \U$22924 ( \23302 , \23301 , \23192 );
and \U$22925 ( \23303 , \23299 , \23302 );
and \U$22926 ( \23304 , \23297 , \23302 );
or \U$22927 ( \23305 , \23300 , \23303 , \23304 );
and \U$22928 ( \23306 , \23295 , \23305 );
and \U$22929 ( \23307 , \22611 , \21815 );
and \U$22930 ( \23308 , \22523 , \21813 );
nor \U$22931 ( \23309 , \23307 , \23308 );
xnor \U$22932 ( \23310 , \23309 , \21774 );
and \U$22933 ( \23311 , \22721 , \21745 );
and \U$22934 ( \23312 , \22716 , \21743 );
nor \U$22935 ( \23313 , \23311 , \23312 );
xnor \U$22936 ( \23314 , \23313 , \21715 );
and \U$22937 ( \23315 , \23310 , \23314 );
and \U$22938 ( \23316 , \22952 , \21697 );
and \U$22939 ( \23317 , \22837 , \21695 );
nor \U$22940 ( \23318 , \23316 , \23317 );
xnor \U$22941 ( \23319 , \23318 , \21678 );
and \U$22942 ( \23320 , \23314 , \23319 );
and \U$22943 ( \23321 , \23310 , \23319 );
or \U$22944 ( \23322 , \23315 , \23320 , \23321 );
xor \U$22945 ( \23323 , \23122 , \23126 );
xor \U$22946 ( \23324 , \23323 , \23132 );
and \U$22947 ( \23325 , \23322 , \23324 );
not \U$22948 ( \23326 , \23137 );
and \U$22949 ( \23327 , \23324 , \23326 );
and \U$22950 ( \23328 , \23322 , \23326 );
or \U$22951 ( \23329 , \23325 , \23327 , \23328 );
and \U$22952 ( \23330 , \23305 , \23329 );
and \U$22953 ( \23331 , \23295 , \23329 );
or \U$22954 ( \23332 , \23306 , \23330 , \23331 );
xor \U$22955 ( \23333 , \23008 , \23012 );
xor \U$22956 ( \23334 , \23333 , \23017 );
xor \U$22957 ( \23335 , \23135 , \23138 );
xor \U$22958 ( \23336 , \23335 , \23140 );
and \U$22959 ( \23337 , \23334 , \23336 );
xor \U$22960 ( \23338 , \23201 , \23203 );
xor \U$22961 ( \23339 , \23338 , \23206 );
and \U$22962 ( \23340 , \23336 , \23339 );
and \U$22963 ( \23341 , \23334 , \23339 );
or \U$22964 ( \23342 , \23337 , \23340 , \23341 );
and \U$22965 ( \23343 , \23332 , \23342 );
xor \U$22966 ( \23344 , \23214 , \23216 );
xor \U$22967 ( \23345 , \23344 , \23218 );
and \U$22968 ( \23346 , \23342 , \23345 );
and \U$22969 ( \23347 , \23332 , \23345 );
or \U$22970 ( \23348 , \23343 , \23346 , \23347 );
xor \U$22971 ( \23349 , \23056 , \23066 );
xor \U$22972 ( \23350 , \23349 , \23086 );
and \U$22973 ( \23351 , \23348 , \23350 );
xor \U$22974 ( \23352 , \23212 , \23221 );
xor \U$22975 ( \23353 , \23352 , \23224 );
and \U$22976 ( \23354 , \23350 , \23353 );
and \U$22977 ( \23355 , \23348 , \23353 );
or \U$22978 ( \23356 , \23351 , \23354 , \23355 );
xor \U$22979 ( \23357 , \23227 , \23229 );
xor \U$22980 ( \23358 , \23357 , \23232 );
and \U$22981 ( \23359 , \23356 , \23358 );
and \U$22982 ( \23360 , \23241 , \23359 );
xor \U$22983 ( \23361 , \23241 , \23359 );
xor \U$22984 ( \23362 , \23356 , \23358 );
and \U$22985 ( \23363 , \22716 , \21815 );
and \U$22986 ( \23364 , \22611 , \21813 );
nor \U$22987 ( \23365 , \23363 , \23364 );
xnor \U$22988 ( \23366 , \23365 , \21774 );
and \U$22989 ( \23367 , \22837 , \21745 );
and \U$22990 ( \23368 , \22721 , \21743 );
nor \U$22991 ( \23369 , \23367 , \23368 );
xnor \U$22992 ( \23370 , \23369 , \21715 );
and \U$22993 ( \23371 , \23366 , \23370 );
and \U$22994 ( \23372 , \23128 , \21697 );
and \U$22995 ( \23373 , \22952 , \21695 );
nor \U$22996 ( \23374 , \23372 , \23373 );
xnor \U$22997 ( \23375 , \23374 , \21678 );
and \U$22998 ( \23376 , \23370 , \23375 );
and \U$22999 ( \23377 , \23366 , \23375 );
or \U$23000 ( \23378 , \23371 , \23376 , \23377 );
buf \U$23001 ( \23379 , RIc22a0d0_153);
and \U$23002 ( \23380 , \23379 , \21660 );
and \U$23003 ( \23381 , \23136 , \21658 );
nor \U$23004 ( \23382 , \23380 , \23381 );
xnor \U$23005 ( \23383 , \23382 , \21665 );
buf \U$23006 ( \23384 , RIc22a148_154);
and \U$23007 ( \23385 , \23384 , \21654 );
or \U$23008 ( \23386 , \23383 , \23385 );
and \U$23009 ( \23387 , \23378 , \23386 );
and \U$23010 ( \23388 , \23136 , \21660 );
and \U$23011 ( \23389 , \23128 , \21658 );
nor \U$23012 ( \23390 , \23388 , \23389 );
xnor \U$23013 ( \23391 , \23390 , \21665 );
and \U$23014 ( \23392 , \23386 , \23391 );
and \U$23015 ( \23393 , \23378 , \23391 );
or \U$23016 ( \23394 , \23387 , \23392 , \23393 );
and \U$23017 ( \23395 , \22126 , \22163 );
and \U$23018 ( \23396 , \22046 , \22161 );
nor \U$23019 ( \23397 , \23395 , \23396 );
xnor \U$23020 ( \23398 , \23397 , \22091 );
and \U$23021 ( \23399 , \22262 , \22029 );
and \U$23022 ( \23400 , \22200 , \22027 );
nor \U$23023 ( \23401 , \23399 , \23400 );
xnor \U$23024 ( \23402 , \23401 , \21986 );
and \U$23025 ( \23403 , \23398 , \23402 );
and \U$23026 ( \23404 , \22523 , \21916 );
and \U$23027 ( \23405 , \22325 , \21914 );
nor \U$23028 ( \23406 , \23404 , \23405 );
xnor \U$23029 ( \23407 , \23406 , \21867 );
and \U$23030 ( \23408 , \23402 , \23407 );
and \U$23031 ( \23409 , \23398 , \23407 );
or \U$23032 ( \23410 , \23403 , \23408 , \23409 );
and \U$23033 ( \23411 , \21831 , \22697 );
and \U$23034 ( \23412 , \21762 , \22695 );
nor \U$23035 ( \23413 , \23411 , \23412 );
xnor \U$23036 ( \23414 , \23413 , \22561 );
and \U$23037 ( \23415 , \21890 , \22497 );
and \U$23038 ( \23416 , \21836 , \22495 );
nor \U$23039 ( \23417 , \23415 , \23416 );
xnor \U$23040 ( \23418 , \23417 , \22419 );
and \U$23041 ( \23419 , \23414 , \23418 );
and \U$23042 ( \23420 , \22018 , \22333 );
and \U$23043 ( \23421 , \21941 , \22331 );
nor \U$23044 ( \23422 , \23420 , \23421 );
xnor \U$23045 ( \23423 , \23422 , \22239 );
and \U$23046 ( \23424 , \23418 , \23423 );
and \U$23047 ( \23425 , \23414 , \23423 );
or \U$23048 ( \23426 , \23419 , \23424 , \23425 );
and \U$23049 ( \23427 , \23410 , \23426 );
xor \U$23050 ( \23428 , \23004 , \23275 );
xor \U$23051 ( \23429 , \23275 , \23276 );
not \U$23052 ( \23430 , \23429 );
and \U$23053 ( \23431 , \23428 , \23430 );
and \U$23054 ( \23432 , \21653 , \23431 );
not \U$23055 ( \23433 , \23432 );
xnor \U$23056 ( \23434 , \23433 , \23279 );
and \U$23057 ( \23435 , \21685 , \23163 );
and \U$23058 ( \23436 , \21667 , \23161 );
nor \U$23059 ( \23437 , \23435 , \23436 );
xnor \U$23060 ( \23438 , \23437 , \23007 );
and \U$23061 ( \23439 , \23434 , \23438 );
and \U$23062 ( \23440 , \21754 , \22891 );
and \U$23063 ( \23441 , \21706 , \22889 );
nor \U$23064 ( \23442 , \23440 , \23441 );
xnor \U$23065 ( \23443 , \23442 , \22778 );
and \U$23066 ( \23444 , \23438 , \23443 );
and \U$23067 ( \23445 , \23434 , \23443 );
or \U$23068 ( \23446 , \23439 , \23444 , \23445 );
and \U$23069 ( \23447 , \23426 , \23446 );
and \U$23070 ( \23448 , \23410 , \23446 );
or \U$23071 ( \23449 , \23427 , \23447 , \23448 );
and \U$23072 ( \23450 , \23394 , \23449 );
and \U$23073 ( \23451 , \23379 , \21654 );
xor \U$23074 ( \23452 , \23245 , \23249 );
xor \U$23075 ( \23453 , \23452 , \23254 );
and \U$23076 ( \23454 , \23451 , \23453 );
xor \U$23077 ( \23455 , \23310 , \23314 );
xor \U$23078 ( \23456 , \23455 , \23319 );
and \U$23079 ( \23457 , \23453 , \23456 );
and \U$23080 ( \23458 , \23451 , \23456 );
or \U$23081 ( \23459 , \23454 , \23457 , \23458 );
and \U$23082 ( \23460 , \23449 , \23459 );
and \U$23083 ( \23461 , \23394 , \23459 );
or \U$23084 ( \23462 , \23450 , \23460 , \23461 );
xor \U$23085 ( \23463 , \23257 , \23273 );
xor \U$23086 ( \23464 , \23463 , \23292 );
xor \U$23087 ( \23465 , \23297 , \23299 );
xor \U$23088 ( \23466 , \23465 , \23302 );
and \U$23089 ( \23467 , \23464 , \23466 );
xor \U$23090 ( \23468 , \23322 , \23324 );
xor \U$23091 ( \23469 , \23468 , \23326 );
and \U$23092 ( \23470 , \23466 , \23469 );
and \U$23093 ( \23471 , \23464 , \23469 );
or \U$23094 ( \23472 , \23467 , \23470 , \23471 );
and \U$23095 ( \23473 , \23462 , \23472 );
xor \U$23096 ( \23474 , \23159 , \23178 );
xor \U$23097 ( \23475 , \23474 , \23195 );
and \U$23098 ( \23476 , \23472 , \23475 );
and \U$23099 ( \23477 , \23462 , \23475 );
or \U$23100 ( \23478 , \23473 , \23476 , \23477 );
xor \U$23101 ( \23479 , \23295 , \23305 );
xor \U$23102 ( \23480 , \23479 , \23329 );
xor \U$23103 ( \23481 , \23334 , \23336 );
xor \U$23104 ( \23482 , \23481 , \23339 );
and \U$23105 ( \23483 , \23480 , \23482 );
and \U$23106 ( \23484 , \23478 , \23483 );
xor \U$23107 ( \23485 , \23143 , \23198 );
xor \U$23108 ( \23486 , \23485 , \23209 );
and \U$23109 ( \23487 , \23483 , \23486 );
and \U$23110 ( \23488 , \23478 , \23486 );
or \U$23111 ( \23489 , \23484 , \23487 , \23488 );
xor \U$23112 ( \23490 , \23348 , \23350 );
xor \U$23113 ( \23491 , \23490 , \23353 );
and \U$23114 ( \23492 , \23489 , \23491 );
and \U$23115 ( \23493 , \23362 , \23492 );
xor \U$23116 ( \23494 , \23362 , \23492 );
xor \U$23117 ( \23495 , \23489 , \23491 );
buf \U$23118 ( \23496 , RIc226908_28);
buf \U$23119 ( \23497 , RIc226890_29);
and \U$23120 ( \23498 , \23496 , \23497 );
not \U$23121 ( \23499 , \23498 );
and \U$23122 ( \23500 , \23276 , \23499 );
not \U$23123 ( \23501 , \23500 );
and \U$23124 ( \23502 , \21667 , \23431 );
and \U$23125 ( \23503 , \21653 , \23429 );
nor \U$23126 ( \23504 , \23502 , \23503 );
xnor \U$23127 ( \23505 , \23504 , \23279 );
and \U$23128 ( \23506 , \23501 , \23505 );
and \U$23129 ( \23507 , \21706 , \23163 );
and \U$23130 ( \23508 , \21685 , \23161 );
nor \U$23131 ( \23509 , \23507 , \23508 );
xnor \U$23132 ( \23510 , \23509 , \23007 );
and \U$23133 ( \23511 , \23505 , \23510 );
and \U$23134 ( \23512 , \23501 , \23510 );
or \U$23135 ( \23513 , \23506 , \23511 , \23512 );
and \U$23136 ( \23514 , \21762 , \22891 );
and \U$23137 ( \23515 , \21754 , \22889 );
nor \U$23138 ( \23516 , \23514 , \23515 );
xnor \U$23139 ( \23517 , \23516 , \22778 );
and \U$23140 ( \23518 , \21836 , \22697 );
and \U$23141 ( \23519 , \21831 , \22695 );
nor \U$23142 ( \23520 , \23518 , \23519 );
xnor \U$23143 ( \23521 , \23520 , \22561 );
and \U$23144 ( \23522 , \23517 , \23521 );
and \U$23145 ( \23523 , \21941 , \22497 );
and \U$23146 ( \23524 , \21890 , \22495 );
nor \U$23147 ( \23525 , \23523 , \23524 );
xnor \U$23148 ( \23526 , \23525 , \22419 );
and \U$23149 ( \23527 , \23521 , \23526 );
and \U$23150 ( \23528 , \23517 , \23526 );
or \U$23151 ( \23529 , \23522 , \23527 , \23528 );
and \U$23152 ( \23530 , \23513 , \23529 );
and \U$23153 ( \23531 , \22046 , \22333 );
and \U$23154 ( \23532 , \22018 , \22331 );
nor \U$23155 ( \23533 , \23531 , \23532 );
xnor \U$23156 ( \23534 , \23533 , \22239 );
and \U$23157 ( \23535 , \22200 , \22163 );
and \U$23158 ( \23536 , \22126 , \22161 );
nor \U$23159 ( \23537 , \23535 , \23536 );
xnor \U$23160 ( \23538 , \23537 , \22091 );
and \U$23161 ( \23539 , \23534 , \23538 );
and \U$23162 ( \23540 , \22325 , \22029 );
and \U$23163 ( \23541 , \22262 , \22027 );
nor \U$23164 ( \23542 , \23540 , \23541 );
xnor \U$23165 ( \23543 , \23542 , \21986 );
and \U$23166 ( \23544 , \23538 , \23543 );
and \U$23167 ( \23545 , \23534 , \23543 );
or \U$23168 ( \23546 , \23539 , \23544 , \23545 );
and \U$23169 ( \23547 , \23529 , \23546 );
and \U$23170 ( \23548 , \23513 , \23546 );
or \U$23171 ( \23549 , \23530 , \23547 , \23548 );
xor \U$23172 ( \23550 , \23398 , \23402 );
xor \U$23173 ( \23551 , \23550 , \23407 );
xor \U$23174 ( \23552 , \23414 , \23418 );
xor \U$23175 ( \23553 , \23552 , \23423 );
and \U$23176 ( \23554 , \23551 , \23553 );
xor \U$23177 ( \23555 , \23366 , \23370 );
xor \U$23178 ( \23556 , \23555 , \23375 );
and \U$23179 ( \23557 , \23553 , \23556 );
and \U$23180 ( \23558 , \23551 , \23556 );
or \U$23181 ( \23559 , \23554 , \23557 , \23558 );
and \U$23182 ( \23560 , \23549 , \23559 );
and \U$23183 ( \23561 , \23136 , \21697 );
and \U$23184 ( \23562 , \23128 , \21695 );
nor \U$23185 ( \23563 , \23561 , \23562 );
xnor \U$23186 ( \23564 , \23563 , \21678 );
and \U$23187 ( \23565 , \23384 , \21660 );
and \U$23188 ( \23566 , \23379 , \21658 );
nor \U$23189 ( \23567 , \23565 , \23566 );
xnor \U$23190 ( \23568 , \23567 , \21665 );
and \U$23191 ( \23569 , \23564 , \23568 );
buf \U$23192 ( \23570 , RIc22a1c0_155);
and \U$23193 ( \23571 , \23570 , \21654 );
and \U$23194 ( \23572 , \23568 , \23571 );
and \U$23195 ( \23573 , \23564 , \23571 );
or \U$23196 ( \23574 , \23569 , \23572 , \23573 );
and \U$23197 ( \23575 , \22611 , \21916 );
and \U$23198 ( \23576 , \22523 , \21914 );
nor \U$23199 ( \23577 , \23575 , \23576 );
xnor \U$23200 ( \23578 , \23577 , \21867 );
and \U$23201 ( \23579 , \22721 , \21815 );
and \U$23202 ( \23580 , \22716 , \21813 );
nor \U$23203 ( \23581 , \23579 , \23580 );
xnor \U$23204 ( \23582 , \23581 , \21774 );
and \U$23205 ( \23583 , \23578 , \23582 );
and \U$23206 ( \23584 , \22952 , \21745 );
and \U$23207 ( \23585 , \22837 , \21743 );
nor \U$23208 ( \23586 , \23584 , \23585 );
xnor \U$23209 ( \23587 , \23586 , \21715 );
and \U$23210 ( \23588 , \23582 , \23587 );
and \U$23211 ( \23589 , \23578 , \23587 );
or \U$23212 ( \23590 , \23583 , \23588 , \23589 );
and \U$23213 ( \23591 , \23574 , \23590 );
xnor \U$23214 ( \23592 , \23383 , \23385 );
and \U$23215 ( \23593 , \23590 , \23592 );
and \U$23216 ( \23594 , \23574 , \23592 );
or \U$23217 ( \23595 , \23591 , \23593 , \23594 );
and \U$23218 ( \23596 , \23559 , \23595 );
and \U$23219 ( \23597 , \23549 , \23595 );
or \U$23220 ( \23598 , \23560 , \23596 , \23597 );
xor \U$23221 ( \23599 , \23261 , \23265 );
xor \U$23222 ( \23600 , \23599 , \23270 );
xor \U$23223 ( \23601 , \23280 , \23284 );
xor \U$23224 ( \23602 , \23601 , \23289 );
and \U$23225 ( \23603 , \23600 , \23602 );
xor \U$23226 ( \23604 , \23451 , \23453 );
xor \U$23227 ( \23605 , \23604 , \23456 );
and \U$23228 ( \23606 , \23602 , \23605 );
and \U$23229 ( \23607 , \23600 , \23605 );
or \U$23230 ( \23608 , \23603 , \23606 , \23607 );
and \U$23231 ( \23609 , \23598 , \23608 );
xor \U$23232 ( \23610 , \23464 , \23466 );
xor \U$23233 ( \23611 , \23610 , \23469 );
and \U$23234 ( \23612 , \23608 , \23611 );
and \U$23235 ( \23613 , \23598 , \23611 );
or \U$23236 ( \23614 , \23609 , \23612 , \23613 );
xor \U$23237 ( \23615 , \23462 , \23472 );
xor \U$23238 ( \23616 , \23615 , \23475 );
and \U$23239 ( \23617 , \23614 , \23616 );
xor \U$23240 ( \23618 , \23480 , \23482 );
and \U$23241 ( \23619 , \23616 , \23618 );
and \U$23242 ( \23620 , \23614 , \23618 );
or \U$23243 ( \23621 , \23617 , \23619 , \23620 );
xor \U$23244 ( \23622 , \23478 , \23483 );
xor \U$23245 ( \23623 , \23622 , \23486 );
and \U$23246 ( \23624 , \23621 , \23623 );
xor \U$23247 ( \23625 , \23332 , \23342 );
xor \U$23248 ( \23626 , \23625 , \23345 );
and \U$23249 ( \23627 , \23623 , \23626 );
and \U$23250 ( \23628 , \23621 , \23626 );
or \U$23251 ( \23629 , \23624 , \23627 , \23628 );
and \U$23252 ( \23630 , \23495 , \23629 );
xor \U$23253 ( \23631 , \23495 , \23629 );
xor \U$23254 ( \23632 , \23621 , \23623 );
xor \U$23255 ( \23633 , \23632 , \23626 );
xor \U$23256 ( \23634 , \23276 , \23496 );
xor \U$23257 ( \23635 , \23496 , \23497 );
not \U$23258 ( \23636 , \23635 );
and \U$23259 ( \23637 , \23634 , \23636 );
and \U$23260 ( \23638 , \21653 , \23637 );
not \U$23261 ( \23639 , \23638 );
xnor \U$23262 ( \23640 , \23639 , \23500 );
and \U$23263 ( \23641 , \21685 , \23431 );
and \U$23264 ( \23642 , \21667 , \23429 );
nor \U$23265 ( \23643 , \23641 , \23642 );
xnor \U$23266 ( \23644 , \23643 , \23279 );
and \U$23267 ( \23645 , \23640 , \23644 );
and \U$23268 ( \23646 , \21754 , \23163 );
and \U$23269 ( \23647 , \21706 , \23161 );
nor \U$23270 ( \23648 , \23646 , \23647 );
xnor \U$23271 ( \23649 , \23648 , \23007 );
and \U$23272 ( \23650 , \23644 , \23649 );
and \U$23273 ( \23651 , \23640 , \23649 );
or \U$23274 ( \23652 , \23645 , \23650 , \23651 );
and \U$23275 ( \23653 , \21831 , \22891 );
and \U$23276 ( \23654 , \21762 , \22889 );
nor \U$23277 ( \23655 , \23653 , \23654 );
xnor \U$23278 ( \23656 , \23655 , \22778 );
and \U$23279 ( \23657 , \21890 , \22697 );
and \U$23280 ( \23658 , \21836 , \22695 );
nor \U$23281 ( \23659 , \23657 , \23658 );
xnor \U$23282 ( \23660 , \23659 , \22561 );
and \U$23283 ( \23661 , \23656 , \23660 );
and \U$23284 ( \23662 , \22018 , \22497 );
and \U$23285 ( \23663 , \21941 , \22495 );
nor \U$23286 ( \23664 , \23662 , \23663 );
xnor \U$23287 ( \23665 , \23664 , \22419 );
and \U$23288 ( \23666 , \23660 , \23665 );
and \U$23289 ( \23667 , \23656 , \23665 );
or \U$23290 ( \23668 , \23661 , \23666 , \23667 );
and \U$23291 ( \23669 , \23652 , \23668 );
and \U$23292 ( \23670 , \22126 , \22333 );
and \U$23293 ( \23671 , \22046 , \22331 );
nor \U$23294 ( \23672 , \23670 , \23671 );
xnor \U$23295 ( \23673 , \23672 , \22239 );
and \U$23296 ( \23674 , \22262 , \22163 );
and \U$23297 ( \23675 , \22200 , \22161 );
nor \U$23298 ( \23676 , \23674 , \23675 );
xnor \U$23299 ( \23677 , \23676 , \22091 );
and \U$23300 ( \23678 , \23673 , \23677 );
and \U$23301 ( \23679 , \22523 , \22029 );
and \U$23302 ( \23680 , \22325 , \22027 );
nor \U$23303 ( \23681 , \23679 , \23680 );
xnor \U$23304 ( \23682 , \23681 , \21986 );
and \U$23305 ( \23683 , \23677 , \23682 );
and \U$23306 ( \23684 , \23673 , \23682 );
or \U$23307 ( \23685 , \23678 , \23683 , \23684 );
and \U$23308 ( \23686 , \23668 , \23685 );
and \U$23309 ( \23687 , \23652 , \23685 );
or \U$23310 ( \23688 , \23669 , \23686 , \23687 );
and \U$23311 ( \23689 , \22716 , \21916 );
and \U$23312 ( \23690 , \22611 , \21914 );
nor \U$23313 ( \23691 , \23689 , \23690 );
xnor \U$23314 ( \23692 , \23691 , \21867 );
and \U$23315 ( \23693 , \22837 , \21815 );
and \U$23316 ( \23694 , \22721 , \21813 );
nor \U$23317 ( \23695 , \23693 , \23694 );
xnor \U$23318 ( \23696 , \23695 , \21774 );
and \U$23319 ( \23697 , \23692 , \23696 );
and \U$23320 ( \23698 , \23128 , \21745 );
and \U$23321 ( \23699 , \22952 , \21743 );
nor \U$23322 ( \23700 , \23698 , \23699 );
xnor \U$23323 ( \23701 , \23700 , \21715 );
and \U$23324 ( \23702 , \23696 , \23701 );
and \U$23325 ( \23703 , \23692 , \23701 );
or \U$23326 ( \23704 , \23697 , \23702 , \23703 );
and \U$23327 ( \23705 , \23379 , \21697 );
and \U$23328 ( \23706 , \23136 , \21695 );
nor \U$23329 ( \23707 , \23705 , \23706 );
xnor \U$23330 ( \23708 , \23707 , \21678 );
and \U$23331 ( \23709 , \23570 , \21660 );
and \U$23332 ( \23710 , \23384 , \21658 );
nor \U$23333 ( \23711 , \23709 , \23710 );
xnor \U$23334 ( \23712 , \23711 , \21665 );
and \U$23335 ( \23713 , \23708 , \23712 );
buf \U$23336 ( \23714 , RIc22a238_156);
and \U$23337 ( \23715 , \23714 , \21654 );
and \U$23338 ( \23716 , \23712 , \23715 );
and \U$23339 ( \23717 , \23708 , \23715 );
or \U$23340 ( \23718 , \23713 , \23716 , \23717 );
and \U$23341 ( \23719 , \23704 , \23718 );
xor \U$23342 ( \23720 , \23564 , \23568 );
xor \U$23343 ( \23721 , \23720 , \23571 );
and \U$23344 ( \23722 , \23718 , \23721 );
and \U$23345 ( \23723 , \23704 , \23721 );
or \U$23346 ( \23724 , \23719 , \23722 , \23723 );
and \U$23347 ( \23725 , \23688 , \23724 );
xor \U$23348 ( \23726 , \23517 , \23521 );
xor \U$23349 ( \23727 , \23726 , \23526 );
xor \U$23350 ( \23728 , \23578 , \23582 );
xor \U$23351 ( \23729 , \23728 , \23587 );
and \U$23352 ( \23730 , \23727 , \23729 );
xor \U$23353 ( \23731 , \23534 , \23538 );
xor \U$23354 ( \23732 , \23731 , \23543 );
and \U$23355 ( \23733 , \23729 , \23732 );
and \U$23356 ( \23734 , \23727 , \23732 );
or \U$23357 ( \23735 , \23730 , \23733 , \23734 );
and \U$23358 ( \23736 , \23724 , \23735 );
and \U$23359 ( \23737 , \23688 , \23735 );
or \U$23360 ( \23738 , \23725 , \23736 , \23737 );
xor \U$23361 ( \23739 , \23434 , \23438 );
xor \U$23362 ( \23740 , \23739 , \23443 );
xor \U$23363 ( \23741 , \23551 , \23553 );
xor \U$23364 ( \23742 , \23741 , \23556 );
and \U$23365 ( \23743 , \23740 , \23742 );
xor \U$23366 ( \23744 , \23574 , \23590 );
xor \U$23367 ( \23745 , \23744 , \23592 );
and \U$23368 ( \23746 , \23742 , \23745 );
and \U$23369 ( \23747 , \23740 , \23745 );
or \U$23370 ( \23748 , \23743 , \23746 , \23747 );
and \U$23371 ( \23749 , \23738 , \23748 );
xor \U$23372 ( \23750 , \23378 , \23386 );
xor \U$23373 ( \23751 , \23750 , \23391 );
and \U$23374 ( \23752 , \23748 , \23751 );
and \U$23375 ( \23753 , \23738 , \23751 );
or \U$23376 ( \23754 , \23749 , \23752 , \23753 );
xor \U$23377 ( \23755 , \23410 , \23426 );
xor \U$23378 ( \23756 , \23755 , \23446 );
xor \U$23379 ( \23757 , \23549 , \23559 );
xor \U$23380 ( \23758 , \23757 , \23595 );
and \U$23381 ( \23759 , \23756 , \23758 );
xor \U$23382 ( \23760 , \23600 , \23602 );
xor \U$23383 ( \23761 , \23760 , \23605 );
and \U$23384 ( \23762 , \23758 , \23761 );
and \U$23385 ( \23763 , \23756 , \23761 );
or \U$23386 ( \23764 , \23759 , \23762 , \23763 );
and \U$23387 ( \23765 , \23754 , \23764 );
xor \U$23388 ( \23766 , \23394 , \23449 );
xor \U$23389 ( \23767 , \23766 , \23459 );
and \U$23390 ( \23768 , \23764 , \23767 );
and \U$23391 ( \23769 , \23754 , \23767 );
or \U$23392 ( \23770 , \23765 , \23768 , \23769 );
and \U$23393 ( \23771 , \21762 , \23163 );
and \U$23394 ( \23772 , \21754 , \23161 );
nor \U$23395 ( \23773 , \23771 , \23772 );
xnor \U$23396 ( \23774 , \23773 , \23007 );
and \U$23397 ( \23775 , \21836 , \22891 );
and \U$23398 ( \23776 , \21831 , \22889 );
nor \U$23399 ( \23777 , \23775 , \23776 );
xnor \U$23400 ( \23778 , \23777 , \22778 );
and \U$23401 ( \23779 , \23774 , \23778 );
and \U$23402 ( \23780 , \21941 , \22697 );
and \U$23403 ( \23781 , \21890 , \22695 );
nor \U$23404 ( \23782 , \23780 , \23781 );
xnor \U$23405 ( \23783 , \23782 , \22561 );
and \U$23406 ( \23784 , \23778 , \23783 );
and \U$23407 ( \23785 , \23774 , \23783 );
or \U$23408 ( \23786 , \23779 , \23784 , \23785 );
buf \U$23409 ( \23787 , RIc226818_30);
buf \U$23410 ( \23788 , RIc2267a0_31);
and \U$23411 ( \23789 , \23787 , \23788 );
not \U$23412 ( \23790 , \23789 );
and \U$23413 ( \23791 , \23497 , \23790 );
not \U$23414 ( \23792 , \23791 );
and \U$23415 ( \23793 , \21667 , \23637 );
and \U$23416 ( \23794 , \21653 , \23635 );
nor \U$23417 ( \23795 , \23793 , \23794 );
xnor \U$23418 ( \23796 , \23795 , \23500 );
and \U$23419 ( \23797 , \23792 , \23796 );
and \U$23420 ( \23798 , \21706 , \23431 );
and \U$23421 ( \23799 , \21685 , \23429 );
nor \U$23422 ( \23800 , \23798 , \23799 );
xnor \U$23423 ( \23801 , \23800 , \23279 );
and \U$23424 ( \23802 , \23796 , \23801 );
and \U$23425 ( \23803 , \23792 , \23801 );
or \U$23426 ( \23804 , \23797 , \23802 , \23803 );
and \U$23427 ( \23805 , \23786 , \23804 );
and \U$23428 ( \23806 , \22046 , \22497 );
and \U$23429 ( \23807 , \22018 , \22495 );
nor \U$23430 ( \23808 , \23806 , \23807 );
xnor \U$23431 ( \23809 , \23808 , \22419 );
and \U$23432 ( \23810 , \22200 , \22333 );
and \U$23433 ( \23811 , \22126 , \22331 );
nor \U$23434 ( \23812 , \23810 , \23811 );
xnor \U$23435 ( \23813 , \23812 , \22239 );
and \U$23436 ( \23814 , \23809 , \23813 );
and \U$23437 ( \23815 , \22325 , \22163 );
and \U$23438 ( \23816 , \22262 , \22161 );
nor \U$23439 ( \23817 , \23815 , \23816 );
xnor \U$23440 ( \23818 , \23817 , \22091 );
and \U$23441 ( \23819 , \23813 , \23818 );
and \U$23442 ( \23820 , \23809 , \23818 );
or \U$23443 ( \23821 , \23814 , \23819 , \23820 );
and \U$23444 ( \23822 , \23804 , \23821 );
and \U$23445 ( \23823 , \23786 , \23821 );
or \U$23446 ( \23824 , \23805 , \23822 , \23823 );
xor \U$23447 ( \23825 , \23692 , \23696 );
xor \U$23448 ( \23826 , \23825 , \23701 );
xor \U$23449 ( \23827 , \23708 , \23712 );
xor \U$23450 ( \23828 , \23827 , \23715 );
and \U$23451 ( \23829 , \23826 , \23828 );
xor \U$23452 ( \23830 , \23673 , \23677 );
xor \U$23453 ( \23831 , \23830 , \23682 );
and \U$23454 ( \23832 , \23828 , \23831 );
and \U$23455 ( \23833 , \23826 , \23831 );
or \U$23456 ( \23834 , \23829 , \23832 , \23833 );
and \U$23457 ( \23835 , \23824 , \23834 );
and \U$23458 ( \23836 , \23136 , \21745 );
and \U$23459 ( \23837 , \23128 , \21743 );
nor \U$23460 ( \23838 , \23836 , \23837 );
xnor \U$23461 ( \23839 , \23838 , \21715 );
and \U$23462 ( \23840 , \23384 , \21697 );
and \U$23463 ( \23841 , \23379 , \21695 );
nor \U$23464 ( \23842 , \23840 , \23841 );
xnor \U$23465 ( \23843 , \23842 , \21678 );
and \U$23466 ( \23844 , \23839 , \23843 );
and \U$23467 ( \23845 , \23714 , \21660 );
and \U$23468 ( \23846 , \23570 , \21658 );
nor \U$23469 ( \23847 , \23845 , \23846 );
xnor \U$23470 ( \23848 , \23847 , \21665 );
and \U$23471 ( \23849 , \23843 , \23848 );
and \U$23472 ( \23850 , \23839 , \23848 );
or \U$23473 ( \23851 , \23844 , \23849 , \23850 );
and \U$23474 ( \23852 , \22611 , \22029 );
and \U$23475 ( \23853 , \22523 , \22027 );
nor \U$23476 ( \23854 , \23852 , \23853 );
xnor \U$23477 ( \23855 , \23854 , \21986 );
and \U$23478 ( \23856 , \22721 , \21916 );
and \U$23479 ( \23857 , \22716 , \21914 );
nor \U$23480 ( \23858 , \23856 , \23857 );
xnor \U$23481 ( \23859 , \23858 , \21867 );
and \U$23482 ( \23860 , \23855 , \23859 );
and \U$23483 ( \23861 , \22952 , \21815 );
and \U$23484 ( \23862 , \22837 , \21813 );
nor \U$23485 ( \23863 , \23861 , \23862 );
xnor \U$23486 ( \23864 , \23863 , \21774 );
and \U$23487 ( \23865 , \23859 , \23864 );
and \U$23488 ( \23866 , \23855 , \23864 );
or \U$23489 ( \23867 , \23860 , \23865 , \23866 );
or \U$23490 ( \23868 , \23851 , \23867 );
and \U$23491 ( \23869 , \23834 , \23868 );
and \U$23492 ( \23870 , \23824 , \23868 );
or \U$23493 ( \23871 , \23835 , \23869 , \23870 );
xor \U$23494 ( \23872 , \23501 , \23505 );
xor \U$23495 ( \23873 , \23872 , \23510 );
xor \U$23496 ( \23874 , \23704 , \23718 );
xor \U$23497 ( \23875 , \23874 , \23721 );
and \U$23498 ( \23876 , \23873 , \23875 );
xor \U$23499 ( \23877 , \23727 , \23729 );
xor \U$23500 ( \23878 , \23877 , \23732 );
and \U$23501 ( \23879 , \23875 , \23878 );
and \U$23502 ( \23880 , \23873 , \23878 );
or \U$23503 ( \23881 , \23876 , \23879 , \23880 );
and \U$23504 ( \23882 , \23871 , \23881 );
xor \U$23505 ( \23883 , \23513 , \23529 );
xor \U$23506 ( \23884 , \23883 , \23546 );
and \U$23507 ( \23885 , \23881 , \23884 );
and \U$23508 ( \23886 , \23871 , \23884 );
or \U$23509 ( \23887 , \23882 , \23885 , \23886 );
xor \U$23510 ( \23888 , \23738 , \23748 );
xor \U$23511 ( \23889 , \23888 , \23751 );
and \U$23512 ( \23890 , \23887 , \23889 );
xor \U$23513 ( \23891 , \23756 , \23758 );
xor \U$23514 ( \23892 , \23891 , \23761 );
and \U$23515 ( \23893 , \23889 , \23892 );
and \U$23516 ( \23894 , \23887 , \23892 );
or \U$23517 ( \23895 , \23890 , \23893 , \23894 );
xor \U$23518 ( \23896 , \23754 , \23764 );
xor \U$23519 ( \23897 , \23896 , \23767 );
and \U$23520 ( \23898 , \23895 , \23897 );
xor \U$23521 ( \23899 , \23598 , \23608 );
xor \U$23522 ( \23900 , \23899 , \23611 );
and \U$23523 ( \23901 , \23897 , \23900 );
and \U$23524 ( \23902 , \23895 , \23900 );
or \U$23525 ( \23903 , \23898 , \23901 , \23902 );
and \U$23526 ( \23904 , \23770 , \23903 );
xor \U$23527 ( \23905 , \23614 , \23616 );
xor \U$23528 ( \23906 , \23905 , \23618 );
and \U$23529 ( \23907 , \23903 , \23906 );
and \U$23530 ( \23908 , \23770 , \23906 );
or \U$23531 ( \23909 , \23904 , \23907 , \23908 );
and \U$23532 ( \23910 , \23633 , \23909 );
xor \U$23533 ( \23911 , \23633 , \23909 );
xor \U$23534 ( \23912 , \23770 , \23903 );
xor \U$23535 ( \23913 , \23912 , \23906 );
and \U$23536 ( \23914 , \21831 , \23163 );
and \U$23537 ( \23915 , \21762 , \23161 );
nor \U$23538 ( \23916 , \23914 , \23915 );
xnor \U$23539 ( \23917 , \23916 , \23007 );
and \U$23540 ( \23918 , \21890 , \22891 );
and \U$23541 ( \23919 , \21836 , \22889 );
nor \U$23542 ( \23920 , \23918 , \23919 );
xnor \U$23543 ( \23921 , \23920 , \22778 );
and \U$23544 ( \23922 , \23917 , \23921 );
and \U$23545 ( \23923 , \22018 , \22697 );
and \U$23546 ( \23924 , \21941 , \22695 );
nor \U$23547 ( \23925 , \23923 , \23924 );
xnor \U$23548 ( \23926 , \23925 , \22561 );
and \U$23549 ( \23927 , \23921 , \23926 );
and \U$23550 ( \23928 , \23917 , \23926 );
or \U$23551 ( \23929 , \23922 , \23927 , \23928 );
xor \U$23552 ( \23930 , \23497 , \23787 );
xor \U$23553 ( \23931 , \23787 , \23788 );
not \U$23554 ( \23932 , \23931 );
and \U$23555 ( \23933 , \23930 , \23932 );
and \U$23556 ( \23934 , \21653 , \23933 );
not \U$23557 ( \23935 , \23934 );
xnor \U$23558 ( \23936 , \23935 , \23791 );
and \U$23559 ( \23937 , \21685 , \23637 );
and \U$23560 ( \23938 , \21667 , \23635 );
nor \U$23561 ( \23939 , \23937 , \23938 );
xnor \U$23562 ( \23940 , \23939 , \23500 );
and \U$23563 ( \23941 , \23936 , \23940 );
and \U$23564 ( \23942 , \21754 , \23431 );
and \U$23565 ( \23943 , \21706 , \23429 );
nor \U$23566 ( \23944 , \23942 , \23943 );
xnor \U$23567 ( \23945 , \23944 , \23279 );
and \U$23568 ( \23946 , \23940 , \23945 );
and \U$23569 ( \23947 , \23936 , \23945 );
or \U$23570 ( \23948 , \23941 , \23946 , \23947 );
and \U$23571 ( \23949 , \23929 , \23948 );
and \U$23572 ( \23950 , \22126 , \22497 );
and \U$23573 ( \23951 , \22046 , \22495 );
nor \U$23574 ( \23952 , \23950 , \23951 );
xnor \U$23575 ( \23953 , \23952 , \22419 );
and \U$23576 ( \23954 , \22262 , \22333 );
and \U$23577 ( \23955 , \22200 , \22331 );
nor \U$23578 ( \23956 , \23954 , \23955 );
xnor \U$23579 ( \23957 , \23956 , \22239 );
and \U$23580 ( \23958 , \23953 , \23957 );
and \U$23581 ( \23959 , \22523 , \22163 );
and \U$23582 ( \23960 , \22325 , \22161 );
nor \U$23583 ( \23961 , \23959 , \23960 );
xnor \U$23584 ( \23962 , \23961 , \22091 );
and \U$23585 ( \23963 , \23957 , \23962 );
and \U$23586 ( \23964 , \23953 , \23962 );
or \U$23587 ( \23965 , \23958 , \23963 , \23964 );
and \U$23588 ( \23966 , \23948 , \23965 );
and \U$23589 ( \23967 , \23929 , \23965 );
or \U$23590 ( \23968 , \23949 , \23966 , \23967 );
and \U$23591 ( \23969 , \23379 , \21745 );
and \U$23592 ( \23970 , \23136 , \21743 );
nor \U$23593 ( \23971 , \23969 , \23970 );
xnor \U$23594 ( \23972 , \23971 , \21715 );
and \U$23595 ( \23973 , \23570 , \21697 );
and \U$23596 ( \23974 , \23384 , \21695 );
nor \U$23597 ( \23975 , \23973 , \23974 );
xnor \U$23598 ( \23976 , \23975 , \21678 );
and \U$23599 ( \23977 , \23972 , \23976 );
buf \U$23600 ( \23978 , RIc22a2b0_157);
and \U$23601 ( \23979 , \23978 , \21660 );
and \U$23602 ( \23980 , \23714 , \21658 );
nor \U$23603 ( \23981 , \23979 , \23980 );
xnor \U$23604 ( \23982 , \23981 , \21665 );
and \U$23605 ( \23983 , \23976 , \23982 );
and \U$23606 ( \23984 , \23972 , \23982 );
or \U$23607 ( \23985 , \23977 , \23983 , \23984 );
and \U$23608 ( \23986 , \22716 , \22029 );
and \U$23609 ( \23987 , \22611 , \22027 );
nor \U$23610 ( \23988 , \23986 , \23987 );
xnor \U$23611 ( \23989 , \23988 , \21986 );
and \U$23612 ( \23990 , \22837 , \21916 );
and \U$23613 ( \23991 , \22721 , \21914 );
nor \U$23614 ( \23992 , \23990 , \23991 );
xnor \U$23615 ( \23993 , \23992 , \21867 );
and \U$23616 ( \23994 , \23989 , \23993 );
and \U$23617 ( \23995 , \23128 , \21815 );
and \U$23618 ( \23996 , \22952 , \21813 );
nor \U$23619 ( \23997 , \23995 , \23996 );
xnor \U$23620 ( \23998 , \23997 , \21774 );
and \U$23621 ( \23999 , \23993 , \23998 );
and \U$23622 ( \24000 , \23989 , \23998 );
or \U$23623 ( \24001 , \23994 , \23999 , \24000 );
and \U$23624 ( \24002 , \23985 , \24001 );
buf \U$23625 ( \24003 , RIc22a328_158);
and \U$23626 ( \24004 , \24003 , \21654 );
buf \U$23627 ( \24005 , \24004 );
and \U$23628 ( \24006 , \24001 , \24005 );
and \U$23629 ( \24007 , \23985 , \24005 );
or \U$23630 ( \24008 , \24002 , \24006 , \24007 );
and \U$23631 ( \24009 , \23968 , \24008 );
and \U$23632 ( \24010 , \23978 , \21654 );
xor \U$23633 ( \24011 , \23839 , \23843 );
xor \U$23634 ( \24012 , \24011 , \23848 );
and \U$23635 ( \24013 , \24010 , \24012 );
xor \U$23636 ( \24014 , \23855 , \23859 );
xor \U$23637 ( \24015 , \24014 , \23864 );
and \U$23638 ( \24016 , \24012 , \24015 );
and \U$23639 ( \24017 , \24010 , \24015 );
or \U$23640 ( \24018 , \24013 , \24016 , \24017 );
and \U$23641 ( \24019 , \24008 , \24018 );
and \U$23642 ( \24020 , \23968 , \24018 );
or \U$23643 ( \24021 , \24009 , \24019 , \24020 );
xor \U$23644 ( \24022 , \23774 , \23778 );
xor \U$23645 ( \24023 , \24022 , \23783 );
xor \U$23646 ( \24024 , \23792 , \23796 );
xor \U$23647 ( \24025 , \24024 , \23801 );
and \U$23648 ( \24026 , \24023 , \24025 );
xor \U$23649 ( \24027 , \23809 , \23813 );
xor \U$23650 ( \24028 , \24027 , \23818 );
and \U$23651 ( \24029 , \24025 , \24028 );
and \U$23652 ( \24030 , \24023 , \24028 );
or \U$23653 ( \24031 , \24026 , \24029 , \24030 );
xor \U$23654 ( \24032 , \23640 , \23644 );
xor \U$23655 ( \24033 , \24032 , \23649 );
and \U$23656 ( \24034 , \24031 , \24033 );
xor \U$23657 ( \24035 , \23656 , \23660 );
xor \U$23658 ( \24036 , \24035 , \23665 );
and \U$23659 ( \24037 , \24033 , \24036 );
and \U$23660 ( \24038 , \24031 , \24036 );
or \U$23661 ( \24039 , \24034 , \24037 , \24038 );
and \U$23662 ( \24040 , \24021 , \24039 );
xor \U$23663 ( \24041 , \23786 , \23804 );
xor \U$23664 ( \24042 , \24041 , \23821 );
xor \U$23665 ( \24043 , \23826 , \23828 );
xor \U$23666 ( \24044 , \24043 , \23831 );
and \U$23667 ( \24045 , \24042 , \24044 );
xnor \U$23668 ( \24046 , \23851 , \23867 );
and \U$23669 ( \24047 , \24044 , \24046 );
and \U$23670 ( \24048 , \24042 , \24046 );
or \U$23671 ( \24049 , \24045 , \24047 , \24048 );
and \U$23672 ( \24050 , \24039 , \24049 );
and \U$23673 ( \24051 , \24021 , \24049 );
or \U$23674 ( \24052 , \24040 , \24050 , \24051 );
xor \U$23675 ( \24053 , \23652 , \23668 );
xor \U$23676 ( \24054 , \24053 , \23685 );
xor \U$23677 ( \24055 , \23824 , \23834 );
xor \U$23678 ( \24056 , \24055 , \23868 );
and \U$23679 ( \24057 , \24054 , \24056 );
xor \U$23680 ( \24058 , \23873 , \23875 );
xor \U$23681 ( \24059 , \24058 , \23878 );
and \U$23682 ( \24060 , \24056 , \24059 );
and \U$23683 ( \24061 , \24054 , \24059 );
or \U$23684 ( \24062 , \24057 , \24060 , \24061 );
and \U$23685 ( \24063 , \24052 , \24062 );
xor \U$23686 ( \24064 , \23740 , \23742 );
xor \U$23687 ( \24065 , \24064 , \23745 );
and \U$23688 ( \24066 , \24062 , \24065 );
and \U$23689 ( \24067 , \24052 , \24065 );
or \U$23690 ( \24068 , \24063 , \24066 , \24067 );
xor \U$23691 ( \24069 , \23688 , \23724 );
xor \U$23692 ( \24070 , \24069 , \23735 );
xor \U$23693 ( \24071 , \23871 , \23881 );
xor \U$23694 ( \24072 , \24071 , \23884 );
and \U$23695 ( \24073 , \24070 , \24072 );
and \U$23696 ( \24074 , \24068 , \24073 );
xor \U$23697 ( \24075 , \23887 , \23889 );
xor \U$23698 ( \24076 , \24075 , \23892 );
and \U$23699 ( \24077 , \24073 , \24076 );
and \U$23700 ( \24078 , \24068 , \24076 );
or \U$23701 ( \24079 , \24074 , \24077 , \24078 );
xor \U$23702 ( \24080 , \23895 , \23897 );
xor \U$23703 ( \24081 , \24080 , \23900 );
and \U$23704 ( \24082 , \24079 , \24081 );
and \U$23705 ( \24083 , \23913 , \24082 );
xor \U$23706 ( \24084 , \23913 , \24082 );
xor \U$23707 ( \24085 , \24079 , \24081 );
and \U$23708 ( \24086 , \22046 , \22697 );
and \U$23709 ( \24087 , \22018 , \22695 );
nor \U$23710 ( \24088 , \24086 , \24087 );
xnor \U$23711 ( \24089 , \24088 , \22561 );
and \U$23712 ( \24090 , \22200 , \22497 );
and \U$23713 ( \24091 , \22126 , \22495 );
nor \U$23714 ( \24092 , \24090 , \24091 );
xnor \U$23715 ( \24093 , \24092 , \22419 );
and \U$23716 ( \24094 , \24089 , \24093 );
and \U$23717 ( \24095 , \22325 , \22333 );
and \U$23718 ( \24096 , \22262 , \22331 );
nor \U$23719 ( \24097 , \24095 , \24096 );
xnor \U$23720 ( \24098 , \24097 , \22239 );
and \U$23721 ( \24099 , \24093 , \24098 );
and \U$23722 ( \24100 , \24089 , \24098 );
or \U$23723 ( \24101 , \24094 , \24099 , \24100 );
buf \U$23724 ( \24102 , RIc226728_32);
buf \U$23725 ( \24103 , RIc2266b0_33);
and \U$23726 ( \24104 , \24102 , \24103 );
not \U$23727 ( \24105 , \24104 );
and \U$23728 ( \24106 , \23788 , \24105 );
not \U$23729 ( \24107 , \24106 );
and \U$23730 ( \24108 , \21667 , \23933 );
and \U$23731 ( \24109 , \21653 , \23931 );
nor \U$23732 ( \24110 , \24108 , \24109 );
xnor \U$23733 ( \24111 , \24110 , \23791 );
and \U$23734 ( \24112 , \24107 , \24111 );
and \U$23735 ( \24113 , \21706 , \23637 );
and \U$23736 ( \24114 , \21685 , \23635 );
nor \U$23737 ( \24115 , \24113 , \24114 );
xnor \U$23738 ( \24116 , \24115 , \23500 );
and \U$23739 ( \24117 , \24111 , \24116 );
and \U$23740 ( \24118 , \24107 , \24116 );
or \U$23741 ( \24119 , \24112 , \24117 , \24118 );
and \U$23742 ( \24120 , \24101 , \24119 );
and \U$23743 ( \24121 , \21762 , \23431 );
and \U$23744 ( \24122 , \21754 , \23429 );
nor \U$23745 ( \24123 , \24121 , \24122 );
xnor \U$23746 ( \24124 , \24123 , \23279 );
and \U$23747 ( \24125 , \21836 , \23163 );
and \U$23748 ( \24126 , \21831 , \23161 );
nor \U$23749 ( \24127 , \24125 , \24126 );
xnor \U$23750 ( \24128 , \24127 , \23007 );
and \U$23751 ( \24129 , \24124 , \24128 );
and \U$23752 ( \24130 , \21941 , \22891 );
and \U$23753 ( \24131 , \21890 , \22889 );
nor \U$23754 ( \24132 , \24130 , \24131 );
xnor \U$23755 ( \24133 , \24132 , \22778 );
and \U$23756 ( \24134 , \24128 , \24133 );
and \U$23757 ( \24135 , \24124 , \24133 );
or \U$23758 ( \24136 , \24129 , \24134 , \24135 );
and \U$23759 ( \24137 , \24119 , \24136 );
and \U$23760 ( \24138 , \24101 , \24136 );
or \U$23761 ( \24139 , \24120 , \24137 , \24138 );
and \U$23762 ( \24140 , \23136 , \21815 );
and \U$23763 ( \24141 , \23128 , \21813 );
nor \U$23764 ( \24142 , \24140 , \24141 );
xnor \U$23765 ( \24143 , \24142 , \21774 );
and \U$23766 ( \24144 , \23384 , \21745 );
and \U$23767 ( \24145 , \23379 , \21743 );
nor \U$23768 ( \24146 , \24144 , \24145 );
xnor \U$23769 ( \24147 , \24146 , \21715 );
and \U$23770 ( \24148 , \24143 , \24147 );
and \U$23771 ( \24149 , \23714 , \21697 );
and \U$23772 ( \24150 , \23570 , \21695 );
nor \U$23773 ( \24151 , \24149 , \24150 );
xnor \U$23774 ( \24152 , \24151 , \21678 );
and \U$23775 ( \24153 , \24147 , \24152 );
and \U$23776 ( \24154 , \24143 , \24152 );
or \U$23777 ( \24155 , \24148 , \24153 , \24154 );
and \U$23778 ( \24156 , \22611 , \22163 );
and \U$23779 ( \24157 , \22523 , \22161 );
nor \U$23780 ( \24158 , \24156 , \24157 );
xnor \U$23781 ( \24159 , \24158 , \22091 );
and \U$23782 ( \24160 , \22721 , \22029 );
and \U$23783 ( \24161 , \22716 , \22027 );
nor \U$23784 ( \24162 , \24160 , \24161 );
xnor \U$23785 ( \24163 , \24162 , \21986 );
and \U$23786 ( \24164 , \24159 , \24163 );
and \U$23787 ( \24165 , \22952 , \21916 );
and \U$23788 ( \24166 , \22837 , \21914 );
nor \U$23789 ( \24167 , \24165 , \24166 );
xnor \U$23790 ( \24168 , \24167 , \21867 );
and \U$23791 ( \24169 , \24163 , \24168 );
and \U$23792 ( \24170 , \24159 , \24168 );
or \U$23793 ( \24171 , \24164 , \24169 , \24170 );
and \U$23794 ( \24172 , \24155 , \24171 );
and \U$23795 ( \24173 , \24003 , \21660 );
and \U$23796 ( \24174 , \23978 , \21658 );
nor \U$23797 ( \24175 , \24173 , \24174 );
xnor \U$23798 ( \24176 , \24175 , \21665 );
buf \U$23799 ( \24177 , RIc22a3a0_159);
and \U$23800 ( \24178 , \24177 , \21654 );
and \U$23801 ( \24179 , \24176 , \24178 );
and \U$23802 ( \24180 , \24171 , \24179 );
and \U$23803 ( \24181 , \24155 , \24179 );
or \U$23804 ( \24182 , \24172 , \24180 , \24181 );
and \U$23805 ( \24183 , \24139 , \24182 );
xor \U$23806 ( \24184 , \23972 , \23976 );
xor \U$23807 ( \24185 , \24184 , \23982 );
xor \U$23808 ( \24186 , \23989 , \23993 );
xor \U$23809 ( \24187 , \24186 , \23998 );
and \U$23810 ( \24188 , \24185 , \24187 );
not \U$23811 ( \24189 , \24004 );
and \U$23812 ( \24190 , \24187 , \24189 );
and \U$23813 ( \24191 , \24185 , \24189 );
or \U$23814 ( \24192 , \24188 , \24190 , \24191 );
and \U$23815 ( \24193 , \24182 , \24192 );
and \U$23816 ( \24194 , \24139 , \24192 );
or \U$23817 ( \24195 , \24183 , \24193 , \24194 );
xor \U$23818 ( \24196 , \23917 , \23921 );
xor \U$23819 ( \24197 , \24196 , \23926 );
xor \U$23820 ( \24198 , \23936 , \23940 );
xor \U$23821 ( \24199 , \24198 , \23945 );
and \U$23822 ( \24200 , \24197 , \24199 );
xor \U$23823 ( \24201 , \23953 , \23957 );
xor \U$23824 ( \24202 , \24201 , \23962 );
and \U$23825 ( \24203 , \24199 , \24202 );
and \U$23826 ( \24204 , \24197 , \24202 );
or \U$23827 ( \24205 , \24200 , \24203 , \24204 );
xor \U$23828 ( \24206 , \24023 , \24025 );
xor \U$23829 ( \24207 , \24206 , \24028 );
and \U$23830 ( \24208 , \24205 , \24207 );
xor \U$23831 ( \24209 , \24010 , \24012 );
xor \U$23832 ( \24210 , \24209 , \24015 );
and \U$23833 ( \24211 , \24207 , \24210 );
and \U$23834 ( \24212 , \24205 , \24210 );
or \U$23835 ( \24213 , \24208 , \24211 , \24212 );
and \U$23836 ( \24214 , \24195 , \24213 );
xor \U$23837 ( \24215 , \23929 , \23948 );
xor \U$23838 ( \24216 , \24215 , \23965 );
xor \U$23839 ( \24217 , \23985 , \24001 );
xor \U$23840 ( \24218 , \24217 , \24005 );
and \U$23841 ( \24219 , \24216 , \24218 );
and \U$23842 ( \24220 , \24213 , \24219 );
and \U$23843 ( \24221 , \24195 , \24219 );
or \U$23844 ( \24222 , \24214 , \24220 , \24221 );
xor \U$23845 ( \24223 , \23968 , \24008 );
xor \U$23846 ( \24224 , \24223 , \24018 );
xor \U$23847 ( \24225 , \24031 , \24033 );
xor \U$23848 ( \24226 , \24225 , \24036 );
and \U$23849 ( \24227 , \24224 , \24226 );
xor \U$23850 ( \24228 , \24042 , \24044 );
xor \U$23851 ( \24229 , \24228 , \24046 );
and \U$23852 ( \24230 , \24226 , \24229 );
and \U$23853 ( \24231 , \24224 , \24229 );
or \U$23854 ( \24232 , \24227 , \24230 , \24231 );
and \U$23855 ( \24233 , \24222 , \24232 );
xor \U$23856 ( \24234 , \24054 , \24056 );
xor \U$23857 ( \24235 , \24234 , \24059 );
and \U$23858 ( \24236 , \24232 , \24235 );
and \U$23859 ( \24237 , \24222 , \24235 );
or \U$23860 ( \24238 , \24233 , \24236 , \24237 );
xor \U$23861 ( \24239 , \24052 , \24062 );
xor \U$23862 ( \24240 , \24239 , \24065 );
and \U$23863 ( \24241 , \24238 , \24240 );
xor \U$23864 ( \24242 , \24070 , \24072 );
and \U$23865 ( \24243 , \24240 , \24242 );
and \U$23866 ( \24244 , \24238 , \24242 );
or \U$23867 ( \24245 , \24241 , \24243 , \24244 );
xor \U$23868 ( \24246 , \24068 , \24073 );
xor \U$23869 ( \24247 , \24246 , \24076 );
and \U$23870 ( \24248 , \24245 , \24247 );
and \U$23871 ( \24249 , \24085 , \24248 );
xor \U$23872 ( \24250 , \24085 , \24248 );
xor \U$23873 ( \24251 , \24245 , \24247 );
xor \U$23874 ( \24252 , \23788 , \24102 );
xor \U$23875 ( \24253 , \24102 , \24103 );
not \U$23876 ( \24254 , \24253 );
and \U$23877 ( \24255 , \24252 , \24254 );
and \U$23878 ( \24256 , \21653 , \24255 );
not \U$23879 ( \24257 , \24256 );
xnor \U$23880 ( \24258 , \24257 , \24106 );
and \U$23881 ( \24259 , \21685 , \23933 );
and \U$23882 ( \24260 , \21667 , \23931 );
nor \U$23883 ( \24261 , \24259 , \24260 );
xnor \U$23884 ( \24262 , \24261 , \23791 );
and \U$23885 ( \24263 , \24258 , \24262 );
and \U$23886 ( \24264 , \21754 , \23637 );
and \U$23887 ( \24265 , \21706 , \23635 );
nor \U$23888 ( \24266 , \24264 , \24265 );
xnor \U$23889 ( \24267 , \24266 , \23500 );
and \U$23890 ( \24268 , \24262 , \24267 );
and \U$23891 ( \24269 , \24258 , \24267 );
or \U$23892 ( \24270 , \24263 , \24268 , \24269 );
and \U$23893 ( \24271 , \22126 , \22697 );
and \U$23894 ( \24272 , \22046 , \22695 );
nor \U$23895 ( \24273 , \24271 , \24272 );
xnor \U$23896 ( \24274 , \24273 , \22561 );
and \U$23897 ( \24275 , \22262 , \22497 );
and \U$23898 ( \24276 , \22200 , \22495 );
nor \U$23899 ( \24277 , \24275 , \24276 );
xnor \U$23900 ( \24278 , \24277 , \22419 );
and \U$23901 ( \24279 , \24274 , \24278 );
and \U$23902 ( \24280 , \22523 , \22333 );
and \U$23903 ( \24281 , \22325 , \22331 );
nor \U$23904 ( \24282 , \24280 , \24281 );
xnor \U$23905 ( \24283 , \24282 , \22239 );
and \U$23906 ( \24284 , \24278 , \24283 );
and \U$23907 ( \24285 , \24274 , \24283 );
or \U$23908 ( \24286 , \24279 , \24284 , \24285 );
and \U$23909 ( \24287 , \24270 , \24286 );
and \U$23910 ( \24288 , \21831 , \23431 );
and \U$23911 ( \24289 , \21762 , \23429 );
nor \U$23912 ( \24290 , \24288 , \24289 );
xnor \U$23913 ( \24291 , \24290 , \23279 );
and \U$23914 ( \24292 , \21890 , \23163 );
and \U$23915 ( \24293 , \21836 , \23161 );
nor \U$23916 ( \24294 , \24292 , \24293 );
xnor \U$23917 ( \24295 , \24294 , \23007 );
and \U$23918 ( \24296 , \24291 , \24295 );
and \U$23919 ( \24297 , \22018 , \22891 );
and \U$23920 ( \24298 , \21941 , \22889 );
nor \U$23921 ( \24299 , \24297 , \24298 );
xnor \U$23922 ( \24300 , \24299 , \22778 );
and \U$23923 ( \24301 , \24295 , \24300 );
and \U$23924 ( \24302 , \24291 , \24300 );
or \U$23925 ( \24303 , \24296 , \24301 , \24302 );
and \U$23926 ( \24304 , \24286 , \24303 );
and \U$23927 ( \24305 , \24270 , \24303 );
or \U$23928 ( \24306 , \24287 , \24304 , \24305 );
and \U$23929 ( \24307 , \23379 , \21815 );
and \U$23930 ( \24308 , \23136 , \21813 );
nor \U$23931 ( \24309 , \24307 , \24308 );
xnor \U$23932 ( \24310 , \24309 , \21774 );
and \U$23933 ( \24311 , \23570 , \21745 );
and \U$23934 ( \24312 , \23384 , \21743 );
nor \U$23935 ( \24313 , \24311 , \24312 );
xnor \U$23936 ( \24314 , \24313 , \21715 );
and \U$23937 ( \24315 , \24310 , \24314 );
and \U$23938 ( \24316 , \23978 , \21697 );
and \U$23939 ( \24317 , \23714 , \21695 );
nor \U$23940 ( \24318 , \24316 , \24317 );
xnor \U$23941 ( \24319 , \24318 , \21678 );
and \U$23942 ( \24320 , \24314 , \24319 );
and \U$23943 ( \24321 , \24310 , \24319 );
or \U$23944 ( \24322 , \24315 , \24320 , \24321 );
and \U$23945 ( \24323 , \22716 , \22163 );
and \U$23946 ( \24324 , \22611 , \22161 );
nor \U$23947 ( \24325 , \24323 , \24324 );
xnor \U$23948 ( \24326 , \24325 , \22091 );
and \U$23949 ( \24327 , \22837 , \22029 );
and \U$23950 ( \24328 , \22721 , \22027 );
nor \U$23951 ( \24329 , \24327 , \24328 );
xnor \U$23952 ( \24330 , \24329 , \21986 );
and \U$23953 ( \24331 , \24326 , \24330 );
and \U$23954 ( \24332 , \23128 , \21916 );
and \U$23955 ( \24333 , \22952 , \21914 );
nor \U$23956 ( \24334 , \24332 , \24333 );
xnor \U$23957 ( \24335 , \24334 , \21867 );
and \U$23958 ( \24336 , \24330 , \24335 );
and \U$23959 ( \24337 , \24326 , \24335 );
or \U$23960 ( \24338 , \24331 , \24336 , \24337 );
and \U$23961 ( \24339 , \24322 , \24338 );
and \U$23962 ( \24340 , \24177 , \21660 );
and \U$23963 ( \24341 , \24003 , \21658 );
nor \U$23964 ( \24342 , \24340 , \24341 );
xnor \U$23965 ( \24343 , \24342 , \21665 );
buf \U$23966 ( \24344 , RIc22a418_160);
and \U$23967 ( \24345 , \24344 , \21654 );
or \U$23968 ( \24346 , \24343 , \24345 );
and \U$23969 ( \24347 , \24338 , \24346 );
and \U$23970 ( \24348 , \24322 , \24346 );
or \U$23971 ( \24349 , \24339 , \24347 , \24348 );
and \U$23972 ( \24350 , \24306 , \24349 );
xor \U$23973 ( \24351 , \24143 , \24147 );
xor \U$23974 ( \24352 , \24351 , \24152 );
xor \U$23975 ( \24353 , \24159 , \24163 );
xor \U$23976 ( \24354 , \24353 , \24168 );
and \U$23977 ( \24355 , \24352 , \24354 );
xor \U$23978 ( \24356 , \24176 , \24178 );
and \U$23979 ( \24357 , \24354 , \24356 );
and \U$23980 ( \24358 , \24352 , \24356 );
or \U$23981 ( \24359 , \24355 , \24357 , \24358 );
and \U$23982 ( \24360 , \24349 , \24359 );
and \U$23983 ( \24361 , \24306 , \24359 );
or \U$23984 ( \24362 , \24350 , \24360 , \24361 );
xor \U$23985 ( \24363 , \24089 , \24093 );
xor \U$23986 ( \24364 , \24363 , \24098 );
xor \U$23987 ( \24365 , \24107 , \24111 );
xor \U$23988 ( \24366 , \24365 , \24116 );
and \U$23989 ( \24367 , \24364 , \24366 );
xor \U$23990 ( \24368 , \24124 , \24128 );
xor \U$23991 ( \24369 , \24368 , \24133 );
and \U$23992 ( \24370 , \24366 , \24369 );
and \U$23993 ( \24371 , \24364 , \24369 );
or \U$23994 ( \24372 , \24367 , \24370 , \24371 );
xor \U$23995 ( \24373 , \24197 , \24199 );
xor \U$23996 ( \24374 , \24373 , \24202 );
and \U$23997 ( \24375 , \24372 , \24374 );
xor \U$23998 ( \24376 , \24185 , \24187 );
xor \U$23999 ( \24377 , \24376 , \24189 );
and \U$24000 ( \24378 , \24374 , \24377 );
and \U$24001 ( \24379 , \24372 , \24377 );
or \U$24002 ( \24380 , \24375 , \24378 , \24379 );
and \U$24003 ( \24381 , \24362 , \24380 );
xor \U$24004 ( \24382 , \24101 , \24119 );
xor \U$24005 ( \24383 , \24382 , \24136 );
xor \U$24006 ( \24384 , \24155 , \24171 );
xor \U$24007 ( \24385 , \24384 , \24179 );
and \U$24008 ( \24386 , \24383 , \24385 );
and \U$24009 ( \24387 , \24380 , \24386 );
and \U$24010 ( \24388 , \24362 , \24386 );
or \U$24011 ( \24389 , \24381 , \24387 , \24388 );
xor \U$24012 ( \24390 , \24139 , \24182 );
xor \U$24013 ( \24391 , \24390 , \24192 );
xor \U$24014 ( \24392 , \24205 , \24207 );
xor \U$24015 ( \24393 , \24392 , \24210 );
and \U$24016 ( \24394 , \24391 , \24393 );
xor \U$24017 ( \24395 , \24216 , \24218 );
and \U$24018 ( \24396 , \24393 , \24395 );
and \U$24019 ( \24397 , \24391 , \24395 );
or \U$24020 ( \24398 , \24394 , \24396 , \24397 );
and \U$24021 ( \24399 , \24389 , \24398 );
xor \U$24022 ( \24400 , \24224 , \24226 );
xor \U$24023 ( \24401 , \24400 , \24229 );
and \U$24024 ( \24402 , \24398 , \24401 );
and \U$24025 ( \24403 , \24389 , \24401 );
or \U$24026 ( \24404 , \24399 , \24402 , \24403 );
xor \U$24027 ( \24405 , \24021 , \24039 );
xor \U$24028 ( \24406 , \24405 , \24049 );
and \U$24029 ( \24407 , \24404 , \24406 );
xor \U$24030 ( \24408 , \24222 , \24232 );
xor \U$24031 ( \24409 , \24408 , \24235 );
and \U$24032 ( \24410 , \24406 , \24409 );
and \U$24033 ( \24411 , \24404 , \24409 );
or \U$24034 ( \24412 , \24407 , \24410 , \24411 );
xor \U$24035 ( \24413 , \24238 , \24240 );
xor \U$24036 ( \24414 , \24413 , \24242 );
and \U$24037 ( \24415 , \24412 , \24414 );
and \U$24038 ( \24416 , \24251 , \24415 );
xor \U$24039 ( \24417 , \24251 , \24415 );
xor \U$24040 ( \24418 , \24412 , \24414 );
and \U$24041 ( \24419 , \21762 , \23637 );
and \U$24042 ( \24420 , \21754 , \23635 );
nor \U$24043 ( \24421 , \24419 , \24420 );
xnor \U$24044 ( \24422 , \24421 , \23500 );
and \U$24045 ( \24423 , \21836 , \23431 );
and \U$24046 ( \24424 , \21831 , \23429 );
nor \U$24047 ( \24425 , \24423 , \24424 );
xnor \U$24048 ( \24426 , \24425 , \23279 );
and \U$24049 ( \24427 , \24422 , \24426 );
and \U$24050 ( \24428 , \21941 , \23163 );
and \U$24051 ( \24429 , \21890 , \23161 );
nor \U$24052 ( \24430 , \24428 , \24429 );
xnor \U$24053 ( \24431 , \24430 , \23007 );
and \U$24054 ( \24432 , \24426 , \24431 );
and \U$24055 ( \24433 , \24422 , \24431 );
or \U$24056 ( \24434 , \24427 , \24432 , \24433 );
and \U$24057 ( \24435 , \22046 , \22891 );
and \U$24058 ( \24436 , \22018 , \22889 );
nor \U$24059 ( \24437 , \24435 , \24436 );
xnor \U$24060 ( \24438 , \24437 , \22778 );
and \U$24061 ( \24439 , \22200 , \22697 );
and \U$24062 ( \24440 , \22126 , \22695 );
nor \U$24063 ( \24441 , \24439 , \24440 );
xnor \U$24064 ( \24442 , \24441 , \22561 );
and \U$24065 ( \24443 , \24438 , \24442 );
and \U$24066 ( \24444 , \22325 , \22497 );
and \U$24067 ( \24445 , \22262 , \22495 );
nor \U$24068 ( \24446 , \24444 , \24445 );
xnor \U$24069 ( \24447 , \24446 , \22419 );
and \U$24070 ( \24448 , \24442 , \24447 );
and \U$24071 ( \24449 , \24438 , \24447 );
or \U$24072 ( \24450 , \24443 , \24448 , \24449 );
and \U$24073 ( \24451 , \24434 , \24450 );
buf \U$24074 ( \24452 , RIc226638_34);
buf \U$24075 ( \24453 , RIc2265c0_35);
and \U$24076 ( \24454 , \24452 , \24453 );
not \U$24077 ( \24455 , \24454 );
and \U$24078 ( \24456 , \24103 , \24455 );
not \U$24079 ( \24457 , \24456 );
and \U$24080 ( \24458 , \21667 , \24255 );
and \U$24081 ( \24459 , \21653 , \24253 );
nor \U$24082 ( \24460 , \24458 , \24459 );
xnor \U$24083 ( \24461 , \24460 , \24106 );
and \U$24084 ( \24462 , \24457 , \24461 );
and \U$24085 ( \24463 , \21706 , \23933 );
and \U$24086 ( \24464 , \21685 , \23931 );
nor \U$24087 ( \24465 , \24463 , \24464 );
xnor \U$24088 ( \24466 , \24465 , \23791 );
and \U$24089 ( \24467 , \24461 , \24466 );
and \U$24090 ( \24468 , \24457 , \24466 );
or \U$24091 ( \24469 , \24462 , \24467 , \24468 );
and \U$24092 ( \24470 , \24450 , \24469 );
and \U$24093 ( \24471 , \24434 , \24469 );
or \U$24094 ( \24472 , \24451 , \24470 , \24471 );
and \U$24095 ( \24473 , \24003 , \21697 );
and \U$24096 ( \24474 , \23978 , \21695 );
nor \U$24097 ( \24475 , \24473 , \24474 );
xnor \U$24098 ( \24476 , \24475 , \21678 );
and \U$24099 ( \24477 , \24344 , \21660 );
and \U$24100 ( \24478 , \24177 , \21658 );
nor \U$24101 ( \24479 , \24477 , \24478 );
xnor \U$24102 ( \24480 , \24479 , \21665 );
and \U$24103 ( \24481 , \24476 , \24480 );
buf \U$24104 ( \24482 , RIc22a490_161);
and \U$24105 ( \24483 , \24482 , \21654 );
and \U$24106 ( \24484 , \24480 , \24483 );
and \U$24107 ( \24485 , \24476 , \24483 );
or \U$24108 ( \24486 , \24481 , \24484 , \24485 );
and \U$24109 ( \24487 , \23136 , \21916 );
and \U$24110 ( \24488 , \23128 , \21914 );
nor \U$24111 ( \24489 , \24487 , \24488 );
xnor \U$24112 ( \24490 , \24489 , \21867 );
and \U$24113 ( \24491 , \23384 , \21815 );
and \U$24114 ( \24492 , \23379 , \21813 );
nor \U$24115 ( \24493 , \24491 , \24492 );
xnor \U$24116 ( \24494 , \24493 , \21774 );
and \U$24117 ( \24495 , \24490 , \24494 );
and \U$24118 ( \24496 , \23714 , \21745 );
and \U$24119 ( \24497 , \23570 , \21743 );
nor \U$24120 ( \24498 , \24496 , \24497 );
xnor \U$24121 ( \24499 , \24498 , \21715 );
and \U$24122 ( \24500 , \24494 , \24499 );
and \U$24123 ( \24501 , \24490 , \24499 );
or \U$24124 ( \24502 , \24495 , \24500 , \24501 );
and \U$24125 ( \24503 , \24486 , \24502 );
and \U$24126 ( \24504 , \22611 , \22333 );
and \U$24127 ( \24505 , \22523 , \22331 );
nor \U$24128 ( \24506 , \24504 , \24505 );
xnor \U$24129 ( \24507 , \24506 , \22239 );
and \U$24130 ( \24508 , \22721 , \22163 );
and \U$24131 ( \24509 , \22716 , \22161 );
nor \U$24132 ( \24510 , \24508 , \24509 );
xnor \U$24133 ( \24511 , \24510 , \22091 );
and \U$24134 ( \24512 , \24507 , \24511 );
and \U$24135 ( \24513 , \22952 , \22029 );
and \U$24136 ( \24514 , \22837 , \22027 );
nor \U$24137 ( \24515 , \24513 , \24514 );
xnor \U$24138 ( \24516 , \24515 , \21986 );
and \U$24139 ( \24517 , \24511 , \24516 );
and \U$24140 ( \24518 , \24507 , \24516 );
or \U$24141 ( \24519 , \24512 , \24517 , \24518 );
and \U$24142 ( \24520 , \24502 , \24519 );
and \U$24143 ( \24521 , \24486 , \24519 );
or \U$24144 ( \24522 , \24503 , \24520 , \24521 );
and \U$24145 ( \24523 , \24472 , \24522 );
xor \U$24146 ( \24524 , \24310 , \24314 );
xor \U$24147 ( \24525 , \24524 , \24319 );
xor \U$24148 ( \24526 , \24326 , \24330 );
xor \U$24149 ( \24527 , \24526 , \24335 );
and \U$24150 ( \24528 , \24525 , \24527 );
xnor \U$24151 ( \24529 , \24343 , \24345 );
and \U$24152 ( \24530 , \24527 , \24529 );
and \U$24153 ( \24531 , \24525 , \24529 );
or \U$24154 ( \24532 , \24528 , \24530 , \24531 );
and \U$24155 ( \24533 , \24522 , \24532 );
and \U$24156 ( \24534 , \24472 , \24532 );
or \U$24157 ( \24535 , \24523 , \24533 , \24534 );
xor \U$24158 ( \24536 , \24258 , \24262 );
xor \U$24159 ( \24537 , \24536 , \24267 );
xor \U$24160 ( \24538 , \24274 , \24278 );
xor \U$24161 ( \24539 , \24538 , \24283 );
and \U$24162 ( \24540 , \24537 , \24539 );
xor \U$24163 ( \24541 , \24291 , \24295 );
xor \U$24164 ( \24542 , \24541 , \24300 );
and \U$24165 ( \24543 , \24539 , \24542 );
and \U$24166 ( \24544 , \24537 , \24542 );
or \U$24167 ( \24545 , \24540 , \24543 , \24544 );
xor \U$24168 ( \24546 , \24364 , \24366 );
xor \U$24169 ( \24547 , \24546 , \24369 );
and \U$24170 ( \24548 , \24545 , \24547 );
xor \U$24171 ( \24549 , \24352 , \24354 );
xor \U$24172 ( \24550 , \24549 , \24356 );
and \U$24173 ( \24551 , \24547 , \24550 );
and \U$24174 ( \24552 , \24545 , \24550 );
or \U$24175 ( \24553 , \24548 , \24551 , \24552 );
and \U$24176 ( \24554 , \24535 , \24553 );
xor \U$24177 ( \24555 , \24270 , \24286 );
xor \U$24178 ( \24556 , \24555 , \24303 );
xor \U$24179 ( \24557 , \24322 , \24338 );
xor \U$24180 ( \24558 , \24557 , \24346 );
and \U$24181 ( \24559 , \24556 , \24558 );
and \U$24182 ( \24560 , \24553 , \24559 );
and \U$24183 ( \24561 , \24535 , \24559 );
or \U$24184 ( \24562 , \24554 , \24560 , \24561 );
xor \U$24185 ( \24563 , \24306 , \24349 );
xor \U$24186 ( \24564 , \24563 , \24359 );
xor \U$24187 ( \24565 , \24372 , \24374 );
xor \U$24188 ( \24566 , \24565 , \24377 );
and \U$24189 ( \24567 , \24564 , \24566 );
xor \U$24190 ( \24568 , \24383 , \24385 );
and \U$24191 ( \24569 , \24566 , \24568 );
and \U$24192 ( \24570 , \24564 , \24568 );
or \U$24193 ( \24571 , \24567 , \24569 , \24570 );
and \U$24194 ( \24572 , \24562 , \24571 );
xor \U$24195 ( \24573 , \24391 , \24393 );
xor \U$24196 ( \24574 , \24573 , \24395 );
and \U$24197 ( \24575 , \24571 , \24574 );
and \U$24198 ( \24576 , \24562 , \24574 );
or \U$24199 ( \24577 , \24572 , \24575 , \24576 );
xor \U$24200 ( \24578 , \24195 , \24213 );
xor \U$24201 ( \24579 , \24578 , \24219 );
and \U$24202 ( \24580 , \24577 , \24579 );
xor \U$24203 ( \24581 , \24389 , \24398 );
xor \U$24204 ( \24582 , \24581 , \24401 );
and \U$24205 ( \24583 , \24579 , \24582 );
and \U$24206 ( \24584 , \24577 , \24582 );
or \U$24207 ( \24585 , \24580 , \24583 , \24584 );
xor \U$24208 ( \24586 , \24404 , \24406 );
xor \U$24209 ( \24587 , \24586 , \24409 );
and \U$24210 ( \24588 , \24585 , \24587 );
and \U$24211 ( \24589 , \24418 , \24588 );
xor \U$24212 ( \24590 , \24418 , \24588 );
xor \U$24213 ( \24591 , \24585 , \24587 );
and \U$24214 ( \24592 , \24177 , \21697 );
and \U$24215 ( \24593 , \24003 , \21695 );
nor \U$24216 ( \24594 , \24592 , \24593 );
xnor \U$24217 ( \24595 , \24594 , \21678 );
and \U$24218 ( \24596 , \24482 , \21660 );
and \U$24219 ( \24597 , \24344 , \21658 );
nor \U$24220 ( \24598 , \24596 , \24597 );
xnor \U$24221 ( \24599 , \24598 , \21665 );
and \U$24222 ( \24600 , \24595 , \24599 );
buf \U$24223 ( \24601 , RIc22a508_162);
and \U$24224 ( \24602 , \24601 , \21654 );
and \U$24225 ( \24603 , \24599 , \24602 );
and \U$24226 ( \24604 , \24595 , \24602 );
or \U$24227 ( \24605 , \24600 , \24603 , \24604 );
and \U$24228 ( \24606 , \23379 , \21916 );
and \U$24229 ( \24607 , \23136 , \21914 );
nor \U$24230 ( \24608 , \24606 , \24607 );
xnor \U$24231 ( \24609 , \24608 , \21867 );
and \U$24232 ( \24610 , \23570 , \21815 );
and \U$24233 ( \24611 , \23384 , \21813 );
nor \U$24234 ( \24612 , \24610 , \24611 );
xnor \U$24235 ( \24613 , \24612 , \21774 );
and \U$24236 ( \24614 , \24609 , \24613 );
and \U$24237 ( \24615 , \23978 , \21745 );
and \U$24238 ( \24616 , \23714 , \21743 );
nor \U$24239 ( \24617 , \24615 , \24616 );
xnor \U$24240 ( \24618 , \24617 , \21715 );
and \U$24241 ( \24619 , \24613 , \24618 );
and \U$24242 ( \24620 , \24609 , \24618 );
or \U$24243 ( \24621 , \24614 , \24619 , \24620 );
and \U$24244 ( \24622 , \24605 , \24621 );
and \U$24245 ( \24623 , \22716 , \22333 );
and \U$24246 ( \24624 , \22611 , \22331 );
nor \U$24247 ( \24625 , \24623 , \24624 );
xnor \U$24248 ( \24626 , \24625 , \22239 );
and \U$24249 ( \24627 , \22837 , \22163 );
and \U$24250 ( \24628 , \22721 , \22161 );
nor \U$24251 ( \24629 , \24627 , \24628 );
xnor \U$24252 ( \24630 , \24629 , \22091 );
and \U$24253 ( \24631 , \24626 , \24630 );
and \U$24254 ( \24632 , \23128 , \22029 );
and \U$24255 ( \24633 , \22952 , \22027 );
nor \U$24256 ( \24634 , \24632 , \24633 );
xnor \U$24257 ( \24635 , \24634 , \21986 );
and \U$24258 ( \24636 , \24630 , \24635 );
and \U$24259 ( \24637 , \24626 , \24635 );
or \U$24260 ( \24638 , \24631 , \24636 , \24637 );
and \U$24261 ( \24639 , \24621 , \24638 );
and \U$24262 ( \24640 , \24605 , \24638 );
or \U$24263 ( \24641 , \24622 , \24639 , \24640 );
and \U$24264 ( \24642 , \21831 , \23637 );
and \U$24265 ( \24643 , \21762 , \23635 );
nor \U$24266 ( \24644 , \24642 , \24643 );
xnor \U$24267 ( \24645 , \24644 , \23500 );
and \U$24268 ( \24646 , \21890 , \23431 );
and \U$24269 ( \24647 , \21836 , \23429 );
nor \U$24270 ( \24648 , \24646 , \24647 );
xnor \U$24271 ( \24649 , \24648 , \23279 );
and \U$24272 ( \24650 , \24645 , \24649 );
and \U$24273 ( \24651 , \22018 , \23163 );
and \U$24274 ( \24652 , \21941 , \23161 );
nor \U$24275 ( \24653 , \24651 , \24652 );
xnor \U$24276 ( \24654 , \24653 , \23007 );
and \U$24277 ( \24655 , \24649 , \24654 );
and \U$24278 ( \24656 , \24645 , \24654 );
or \U$24279 ( \24657 , \24650 , \24655 , \24656 );
xor \U$24280 ( \24658 , \24103 , \24452 );
xor \U$24281 ( \24659 , \24452 , \24453 );
not \U$24282 ( \24660 , \24659 );
and \U$24283 ( \24661 , \24658 , \24660 );
and \U$24284 ( \24662 , \21653 , \24661 );
not \U$24285 ( \24663 , \24662 );
xnor \U$24286 ( \24664 , \24663 , \24456 );
and \U$24287 ( \24665 , \21685 , \24255 );
and \U$24288 ( \24666 , \21667 , \24253 );
nor \U$24289 ( \24667 , \24665 , \24666 );
xnor \U$24290 ( \24668 , \24667 , \24106 );
and \U$24291 ( \24669 , \24664 , \24668 );
and \U$24292 ( \24670 , \21754 , \23933 );
and \U$24293 ( \24671 , \21706 , \23931 );
nor \U$24294 ( \24672 , \24670 , \24671 );
xnor \U$24295 ( \24673 , \24672 , \23791 );
and \U$24296 ( \24674 , \24668 , \24673 );
and \U$24297 ( \24675 , \24664 , \24673 );
or \U$24298 ( \24676 , \24669 , \24674 , \24675 );
and \U$24299 ( \24677 , \24657 , \24676 );
and \U$24300 ( \24678 , \22126 , \22891 );
and \U$24301 ( \24679 , \22046 , \22889 );
nor \U$24302 ( \24680 , \24678 , \24679 );
xnor \U$24303 ( \24681 , \24680 , \22778 );
and \U$24304 ( \24682 , \22262 , \22697 );
and \U$24305 ( \24683 , \22200 , \22695 );
nor \U$24306 ( \24684 , \24682 , \24683 );
xnor \U$24307 ( \24685 , \24684 , \22561 );
and \U$24308 ( \24686 , \24681 , \24685 );
and \U$24309 ( \24687 , \22523 , \22497 );
and \U$24310 ( \24688 , \22325 , \22495 );
nor \U$24311 ( \24689 , \24687 , \24688 );
xnor \U$24312 ( \24690 , \24689 , \22419 );
and \U$24313 ( \24691 , \24685 , \24690 );
and \U$24314 ( \24692 , \24681 , \24690 );
or \U$24315 ( \24693 , \24686 , \24691 , \24692 );
and \U$24316 ( \24694 , \24676 , \24693 );
and \U$24317 ( \24695 , \24657 , \24693 );
or \U$24318 ( \24696 , \24677 , \24694 , \24695 );
and \U$24319 ( \24697 , \24641 , \24696 );
xor \U$24320 ( \24698 , \24476 , \24480 );
xor \U$24321 ( \24699 , \24698 , \24483 );
xor \U$24322 ( \24700 , \24490 , \24494 );
xor \U$24323 ( \24701 , \24700 , \24499 );
and \U$24324 ( \24702 , \24699 , \24701 );
xor \U$24325 ( \24703 , \24507 , \24511 );
xor \U$24326 ( \24704 , \24703 , \24516 );
and \U$24327 ( \24705 , \24701 , \24704 );
and \U$24328 ( \24706 , \24699 , \24704 );
or \U$24329 ( \24707 , \24702 , \24705 , \24706 );
and \U$24330 ( \24708 , \24696 , \24707 );
and \U$24331 ( \24709 , \24641 , \24707 );
or \U$24332 ( \24710 , \24697 , \24708 , \24709 );
xor \U$24333 ( \24711 , \24422 , \24426 );
xor \U$24334 ( \24712 , \24711 , \24431 );
xor \U$24335 ( \24713 , \24438 , \24442 );
xor \U$24336 ( \24714 , \24713 , \24447 );
and \U$24337 ( \24715 , \24712 , \24714 );
xor \U$24338 ( \24716 , \24457 , \24461 );
xor \U$24339 ( \24717 , \24716 , \24466 );
and \U$24340 ( \24718 , \24714 , \24717 );
and \U$24341 ( \24719 , \24712 , \24717 );
or \U$24342 ( \24720 , \24715 , \24718 , \24719 );
xor \U$24343 ( \24721 , \24537 , \24539 );
xor \U$24344 ( \24722 , \24721 , \24542 );
and \U$24345 ( \24723 , \24720 , \24722 );
xor \U$24346 ( \24724 , \24525 , \24527 );
xor \U$24347 ( \24725 , \24724 , \24529 );
and \U$24348 ( \24726 , \24722 , \24725 );
and \U$24349 ( \24727 , \24720 , \24725 );
or \U$24350 ( \24728 , \24723 , \24726 , \24727 );
and \U$24351 ( \24729 , \24710 , \24728 );
xor \U$24352 ( \24730 , \24434 , \24450 );
xor \U$24353 ( \24731 , \24730 , \24469 );
xor \U$24354 ( \24732 , \24486 , \24502 );
xor \U$24355 ( \24733 , \24732 , \24519 );
and \U$24356 ( \24734 , \24731 , \24733 );
and \U$24357 ( \24735 , \24728 , \24734 );
and \U$24358 ( \24736 , \24710 , \24734 );
or \U$24359 ( \24737 , \24729 , \24735 , \24736 );
xor \U$24360 ( \24738 , \24472 , \24522 );
xor \U$24361 ( \24739 , \24738 , \24532 );
xor \U$24362 ( \24740 , \24545 , \24547 );
xor \U$24363 ( \24741 , \24740 , \24550 );
and \U$24364 ( \24742 , \24739 , \24741 );
xor \U$24365 ( \24743 , \24556 , \24558 );
and \U$24366 ( \24744 , \24741 , \24743 );
and \U$24367 ( \24745 , \24739 , \24743 );
or \U$24368 ( \24746 , \24742 , \24744 , \24745 );
and \U$24369 ( \24747 , \24737 , \24746 );
xor \U$24370 ( \24748 , \24564 , \24566 );
xor \U$24371 ( \24749 , \24748 , \24568 );
and \U$24372 ( \24750 , \24746 , \24749 );
and \U$24373 ( \24751 , \24737 , \24749 );
or \U$24374 ( \24752 , \24747 , \24750 , \24751 );
xor \U$24375 ( \24753 , \24362 , \24380 );
xor \U$24376 ( \24754 , \24753 , \24386 );
and \U$24377 ( \24755 , \24752 , \24754 );
xor \U$24378 ( \24756 , \24562 , \24571 );
xor \U$24379 ( \24757 , \24756 , \24574 );
and \U$24380 ( \24758 , \24754 , \24757 );
and \U$24381 ( \24759 , \24752 , \24757 );
or \U$24382 ( \24760 , \24755 , \24758 , \24759 );
xor \U$24383 ( \24761 , \24577 , \24579 );
xor \U$24384 ( \24762 , \24761 , \24582 );
and \U$24385 ( \24763 , \24760 , \24762 );
and \U$24386 ( \24764 , \24591 , \24763 );
xor \U$24387 ( \24765 , \24591 , \24763 );
xor \U$24388 ( \24766 , \24760 , \24762 );
and \U$24389 ( \24767 , \22046 , \23163 );
and \U$24390 ( \24768 , \22018 , \23161 );
nor \U$24391 ( \24769 , \24767 , \24768 );
xnor \U$24392 ( \24770 , \24769 , \23007 );
and \U$24393 ( \24771 , \22200 , \22891 );
and \U$24394 ( \24772 , \22126 , \22889 );
nor \U$24395 ( \24773 , \24771 , \24772 );
xnor \U$24396 ( \24774 , \24773 , \22778 );
and \U$24397 ( \24775 , \24770 , \24774 );
and \U$24398 ( \24776 , \22325 , \22697 );
and \U$24399 ( \24777 , \22262 , \22695 );
nor \U$24400 ( \24778 , \24776 , \24777 );
xnor \U$24401 ( \24779 , \24778 , \22561 );
and \U$24402 ( \24780 , \24774 , \24779 );
and \U$24403 ( \24781 , \24770 , \24779 );
or \U$24404 ( \24782 , \24775 , \24780 , \24781 );
buf \U$24405 ( \24783 , RIc226548_36);
buf \U$24406 ( \24784 , RIc2264d0_37);
and \U$24407 ( \24785 , \24783 , \24784 );
not \U$24408 ( \24786 , \24785 );
and \U$24409 ( \24787 , \24453 , \24786 );
not \U$24410 ( \24788 , \24787 );
and \U$24411 ( \24789 , \21667 , \24661 );
and \U$24412 ( \24790 , \21653 , \24659 );
nor \U$24413 ( \24791 , \24789 , \24790 );
xnor \U$24414 ( \24792 , \24791 , \24456 );
and \U$24415 ( \24793 , \24788 , \24792 );
and \U$24416 ( \24794 , \21706 , \24255 );
and \U$24417 ( \24795 , \21685 , \24253 );
nor \U$24418 ( \24796 , \24794 , \24795 );
xnor \U$24419 ( \24797 , \24796 , \24106 );
and \U$24420 ( \24798 , \24792 , \24797 );
and \U$24421 ( \24799 , \24788 , \24797 );
or \U$24422 ( \24800 , \24793 , \24798 , \24799 );
and \U$24423 ( \24801 , \24782 , \24800 );
and \U$24424 ( \24802 , \21762 , \23933 );
and \U$24425 ( \24803 , \21754 , \23931 );
nor \U$24426 ( \24804 , \24802 , \24803 );
xnor \U$24427 ( \24805 , \24804 , \23791 );
and \U$24428 ( \24806 , \21836 , \23637 );
and \U$24429 ( \24807 , \21831 , \23635 );
nor \U$24430 ( \24808 , \24806 , \24807 );
xnor \U$24431 ( \24809 , \24808 , \23500 );
and \U$24432 ( \24810 , \24805 , \24809 );
and \U$24433 ( \24811 , \21941 , \23431 );
and \U$24434 ( \24812 , \21890 , \23429 );
nor \U$24435 ( \24813 , \24811 , \24812 );
xnor \U$24436 ( \24814 , \24813 , \23279 );
and \U$24437 ( \24815 , \24809 , \24814 );
and \U$24438 ( \24816 , \24805 , \24814 );
or \U$24439 ( \24817 , \24810 , \24815 , \24816 );
and \U$24440 ( \24818 , \24800 , \24817 );
and \U$24441 ( \24819 , \24782 , \24817 );
or \U$24442 ( \24820 , \24801 , \24818 , \24819 );
and \U$24443 ( \24821 , \24003 , \21745 );
and \U$24444 ( \24822 , \23978 , \21743 );
nor \U$24445 ( \24823 , \24821 , \24822 );
xnor \U$24446 ( \24824 , \24823 , \21715 );
and \U$24447 ( \24825 , \24344 , \21697 );
and \U$24448 ( \24826 , \24177 , \21695 );
nor \U$24449 ( \24827 , \24825 , \24826 );
xnor \U$24450 ( \24828 , \24827 , \21678 );
and \U$24451 ( \24829 , \24824 , \24828 );
and \U$24452 ( \24830 , \24601 , \21660 );
and \U$24453 ( \24831 , \24482 , \21658 );
nor \U$24454 ( \24832 , \24830 , \24831 );
xnor \U$24455 ( \24833 , \24832 , \21665 );
and \U$24456 ( \24834 , \24828 , \24833 );
and \U$24457 ( \24835 , \24824 , \24833 );
or \U$24458 ( \24836 , \24829 , \24834 , \24835 );
and \U$24459 ( \24837 , \22611 , \22497 );
and \U$24460 ( \24838 , \22523 , \22495 );
nor \U$24461 ( \24839 , \24837 , \24838 );
xnor \U$24462 ( \24840 , \24839 , \22419 );
and \U$24463 ( \24841 , \22721 , \22333 );
and \U$24464 ( \24842 , \22716 , \22331 );
nor \U$24465 ( \24843 , \24841 , \24842 );
xnor \U$24466 ( \24844 , \24843 , \22239 );
and \U$24467 ( \24845 , \24840 , \24844 );
and \U$24468 ( \24846 , \22952 , \22163 );
and \U$24469 ( \24847 , \22837 , \22161 );
nor \U$24470 ( \24848 , \24846 , \24847 );
xnor \U$24471 ( \24849 , \24848 , \22091 );
and \U$24472 ( \24850 , \24844 , \24849 );
and \U$24473 ( \24851 , \24840 , \24849 );
or \U$24474 ( \24852 , \24845 , \24850 , \24851 );
and \U$24475 ( \24853 , \24836 , \24852 );
and \U$24476 ( \24854 , \23136 , \22029 );
and \U$24477 ( \24855 , \23128 , \22027 );
nor \U$24478 ( \24856 , \24854 , \24855 );
xnor \U$24479 ( \24857 , \24856 , \21986 );
and \U$24480 ( \24858 , \23384 , \21916 );
and \U$24481 ( \24859 , \23379 , \21914 );
nor \U$24482 ( \24860 , \24858 , \24859 );
xnor \U$24483 ( \24861 , \24860 , \21867 );
and \U$24484 ( \24862 , \24857 , \24861 );
and \U$24485 ( \24863 , \23714 , \21815 );
and \U$24486 ( \24864 , \23570 , \21813 );
nor \U$24487 ( \24865 , \24863 , \24864 );
xnor \U$24488 ( \24866 , \24865 , \21774 );
and \U$24489 ( \24867 , \24861 , \24866 );
and \U$24490 ( \24868 , \24857 , \24866 );
or \U$24491 ( \24869 , \24862 , \24867 , \24868 );
and \U$24492 ( \24870 , \24852 , \24869 );
and \U$24493 ( \24871 , \24836 , \24869 );
or \U$24494 ( \24872 , \24853 , \24870 , \24871 );
and \U$24495 ( \24873 , \24820 , \24872 );
xor \U$24496 ( \24874 , \24595 , \24599 );
xor \U$24497 ( \24875 , \24874 , \24602 );
xor \U$24498 ( \24876 , \24609 , \24613 );
xor \U$24499 ( \24877 , \24876 , \24618 );
or \U$24500 ( \24878 , \24875 , \24877 );
and \U$24501 ( \24879 , \24872 , \24878 );
and \U$24502 ( \24880 , \24820 , \24878 );
or \U$24503 ( \24881 , \24873 , \24879 , \24880 );
xor \U$24504 ( \24882 , \24645 , \24649 );
xor \U$24505 ( \24883 , \24882 , \24654 );
xor \U$24506 ( \24884 , \24681 , \24685 );
xor \U$24507 ( \24885 , \24884 , \24690 );
and \U$24508 ( \24886 , \24883 , \24885 );
xor \U$24509 ( \24887 , \24626 , \24630 );
xor \U$24510 ( \24888 , \24887 , \24635 );
and \U$24511 ( \24889 , \24885 , \24888 );
and \U$24512 ( \24890 , \24883 , \24888 );
or \U$24513 ( \24891 , \24886 , \24889 , \24890 );
xor \U$24514 ( \24892 , \24699 , \24701 );
xor \U$24515 ( \24893 , \24892 , \24704 );
and \U$24516 ( \24894 , \24891 , \24893 );
xor \U$24517 ( \24895 , \24712 , \24714 );
xor \U$24518 ( \24896 , \24895 , \24717 );
and \U$24519 ( \24897 , \24893 , \24896 );
and \U$24520 ( \24898 , \24891 , \24896 );
or \U$24521 ( \24899 , \24894 , \24897 , \24898 );
and \U$24522 ( \24900 , \24881 , \24899 );
xor \U$24523 ( \24901 , \24605 , \24621 );
xor \U$24524 ( \24902 , \24901 , \24638 );
xor \U$24525 ( \24903 , \24657 , \24676 );
xor \U$24526 ( \24904 , \24903 , \24693 );
and \U$24527 ( \24905 , \24902 , \24904 );
and \U$24528 ( \24906 , \24899 , \24905 );
and \U$24529 ( \24907 , \24881 , \24905 );
or \U$24530 ( \24908 , \24900 , \24906 , \24907 );
xor \U$24531 ( \24909 , \24641 , \24696 );
xor \U$24532 ( \24910 , \24909 , \24707 );
xor \U$24533 ( \24911 , \24720 , \24722 );
xor \U$24534 ( \24912 , \24911 , \24725 );
and \U$24535 ( \24913 , \24910 , \24912 );
xor \U$24536 ( \24914 , \24731 , \24733 );
and \U$24537 ( \24915 , \24912 , \24914 );
and \U$24538 ( \24916 , \24910 , \24914 );
or \U$24539 ( \24917 , \24913 , \24915 , \24916 );
and \U$24540 ( \24918 , \24908 , \24917 );
xor \U$24541 ( \24919 , \24739 , \24741 );
xor \U$24542 ( \24920 , \24919 , \24743 );
and \U$24543 ( \24921 , \24917 , \24920 );
and \U$24544 ( \24922 , \24908 , \24920 );
or \U$24545 ( \24923 , \24918 , \24921 , \24922 );
xor \U$24546 ( \24924 , \24535 , \24553 );
xor \U$24547 ( \24925 , \24924 , \24559 );
and \U$24548 ( \24926 , \24923 , \24925 );
xor \U$24549 ( \24927 , \24737 , \24746 );
xor \U$24550 ( \24928 , \24927 , \24749 );
and \U$24551 ( \24929 , \24925 , \24928 );
and \U$24552 ( \24930 , \24923 , \24928 );
or \U$24553 ( \24931 , \24926 , \24929 , \24930 );
xor \U$24554 ( \24932 , \24752 , \24754 );
xor \U$24555 ( \24933 , \24932 , \24757 );
and \U$24556 ( \24934 , \24931 , \24933 );
and \U$24557 ( \24935 , \24766 , \24934 );
xor \U$24558 ( \24936 , \24766 , \24934 );
xor \U$24559 ( \24937 , \24931 , \24933 );
and \U$24560 ( \24938 , \22126 , \23163 );
and \U$24561 ( \24939 , \22046 , \23161 );
nor \U$24562 ( \24940 , \24938 , \24939 );
xnor \U$24563 ( \24941 , \24940 , \23007 );
and \U$24564 ( \24942 , \22262 , \22891 );
and \U$24565 ( \24943 , \22200 , \22889 );
nor \U$24566 ( \24944 , \24942 , \24943 );
xnor \U$24567 ( \24945 , \24944 , \22778 );
and \U$24568 ( \24946 , \24941 , \24945 );
and \U$24569 ( \24947 , \22523 , \22697 );
and \U$24570 ( \24948 , \22325 , \22695 );
nor \U$24571 ( \24949 , \24947 , \24948 );
xnor \U$24572 ( \24950 , \24949 , \22561 );
and \U$24573 ( \24951 , \24945 , \24950 );
and \U$24574 ( \24952 , \24941 , \24950 );
or \U$24575 ( \24953 , \24946 , \24951 , \24952 );
and \U$24576 ( \24954 , \21831 , \23933 );
and \U$24577 ( \24955 , \21762 , \23931 );
nor \U$24578 ( \24956 , \24954 , \24955 );
xnor \U$24579 ( \24957 , \24956 , \23791 );
and \U$24580 ( \24958 , \21890 , \23637 );
and \U$24581 ( \24959 , \21836 , \23635 );
nor \U$24582 ( \24960 , \24958 , \24959 );
xnor \U$24583 ( \24961 , \24960 , \23500 );
and \U$24584 ( \24962 , \24957 , \24961 );
and \U$24585 ( \24963 , \22018 , \23431 );
and \U$24586 ( \24964 , \21941 , \23429 );
nor \U$24587 ( \24965 , \24963 , \24964 );
xnor \U$24588 ( \24966 , \24965 , \23279 );
and \U$24589 ( \24967 , \24961 , \24966 );
and \U$24590 ( \24968 , \24957 , \24966 );
or \U$24591 ( \24969 , \24962 , \24967 , \24968 );
and \U$24592 ( \24970 , \24953 , \24969 );
xor \U$24593 ( \24971 , \24453 , \24783 );
xor \U$24594 ( \24972 , \24783 , \24784 );
not \U$24595 ( \24973 , \24972 );
and \U$24596 ( \24974 , \24971 , \24973 );
and \U$24597 ( \24975 , \21653 , \24974 );
not \U$24598 ( \24976 , \24975 );
xnor \U$24599 ( \24977 , \24976 , \24787 );
and \U$24600 ( \24978 , \21685 , \24661 );
and \U$24601 ( \24979 , \21667 , \24659 );
nor \U$24602 ( \24980 , \24978 , \24979 );
xnor \U$24603 ( \24981 , \24980 , \24456 );
and \U$24604 ( \24982 , \24977 , \24981 );
and \U$24605 ( \24983 , \21754 , \24255 );
and \U$24606 ( \24984 , \21706 , \24253 );
nor \U$24607 ( \24985 , \24983 , \24984 );
xnor \U$24608 ( \24986 , \24985 , \24106 );
and \U$24609 ( \24987 , \24981 , \24986 );
and \U$24610 ( \24988 , \24977 , \24986 );
or \U$24611 ( \24989 , \24982 , \24987 , \24988 );
and \U$24612 ( \24990 , \24969 , \24989 );
and \U$24613 ( \24991 , \24953 , \24989 );
or \U$24614 ( \24992 , \24970 , \24990 , \24991 );
and \U$24615 ( \24993 , \22716 , \22497 );
and \U$24616 ( \24994 , \22611 , \22495 );
nor \U$24617 ( \24995 , \24993 , \24994 );
xnor \U$24618 ( \24996 , \24995 , \22419 );
and \U$24619 ( \24997 , \22837 , \22333 );
and \U$24620 ( \24998 , \22721 , \22331 );
nor \U$24621 ( \24999 , \24997 , \24998 );
xnor \U$24622 ( \25000 , \24999 , \22239 );
and \U$24623 ( \25001 , \24996 , \25000 );
and \U$24624 ( \25002 , \23128 , \22163 );
and \U$24625 ( \25003 , \22952 , \22161 );
nor \U$24626 ( \25004 , \25002 , \25003 );
xnor \U$24627 ( \25005 , \25004 , \22091 );
and \U$24628 ( \25006 , \25000 , \25005 );
and \U$24629 ( \25007 , \24996 , \25005 );
or \U$24630 ( \25008 , \25001 , \25006 , \25007 );
and \U$24631 ( \25009 , \24177 , \21745 );
and \U$24632 ( \25010 , \24003 , \21743 );
nor \U$24633 ( \25011 , \25009 , \25010 );
xnor \U$24634 ( \25012 , \25011 , \21715 );
and \U$24635 ( \25013 , \24482 , \21697 );
and \U$24636 ( \25014 , \24344 , \21695 );
nor \U$24637 ( \25015 , \25013 , \25014 );
xnor \U$24638 ( \25016 , \25015 , \21678 );
and \U$24639 ( \25017 , \25012 , \25016 );
buf \U$24640 ( \25018 , RIc22a580_163);
and \U$24641 ( \25019 , \25018 , \21660 );
and \U$24642 ( \25020 , \24601 , \21658 );
nor \U$24643 ( \25021 , \25019 , \25020 );
xnor \U$24644 ( \25022 , \25021 , \21665 );
and \U$24645 ( \25023 , \25016 , \25022 );
and \U$24646 ( \25024 , \25012 , \25022 );
or \U$24647 ( \25025 , \25017 , \25023 , \25024 );
and \U$24648 ( \25026 , \25008 , \25025 );
and \U$24649 ( \25027 , \23379 , \22029 );
and \U$24650 ( \25028 , \23136 , \22027 );
nor \U$24651 ( \25029 , \25027 , \25028 );
xnor \U$24652 ( \25030 , \25029 , \21986 );
and \U$24653 ( \25031 , \23570 , \21916 );
and \U$24654 ( \25032 , \23384 , \21914 );
nor \U$24655 ( \25033 , \25031 , \25032 );
xnor \U$24656 ( \25034 , \25033 , \21867 );
and \U$24657 ( \25035 , \25030 , \25034 );
and \U$24658 ( \25036 , \23978 , \21815 );
and \U$24659 ( \25037 , \23714 , \21813 );
nor \U$24660 ( \25038 , \25036 , \25037 );
xnor \U$24661 ( \25039 , \25038 , \21774 );
and \U$24662 ( \25040 , \25034 , \25039 );
and \U$24663 ( \25041 , \25030 , \25039 );
or \U$24664 ( \25042 , \25035 , \25040 , \25041 );
and \U$24665 ( \25043 , \25025 , \25042 );
and \U$24666 ( \25044 , \25008 , \25042 );
or \U$24667 ( \25045 , \25026 , \25043 , \25044 );
and \U$24668 ( \25046 , \24992 , \25045 );
and \U$24669 ( \25047 , \25018 , \21654 );
xor \U$24670 ( \25048 , \24824 , \24828 );
xor \U$24671 ( \25049 , \25048 , \24833 );
and \U$24672 ( \25050 , \25047 , \25049 );
xor \U$24673 ( \25051 , \24857 , \24861 );
xor \U$24674 ( \25052 , \25051 , \24866 );
and \U$24675 ( \25053 , \25049 , \25052 );
and \U$24676 ( \25054 , \25047 , \25052 );
or \U$24677 ( \25055 , \25050 , \25053 , \25054 );
and \U$24678 ( \25056 , \25045 , \25055 );
and \U$24679 ( \25057 , \24992 , \25055 );
or \U$24680 ( \25058 , \25046 , \25056 , \25057 );
xor \U$24681 ( \25059 , \24770 , \24774 );
xor \U$24682 ( \25060 , \25059 , \24779 );
xor \U$24683 ( \25061 , \24840 , \24844 );
xor \U$24684 ( \25062 , \25061 , \24849 );
and \U$24685 ( \25063 , \25060 , \25062 );
xor \U$24686 ( \25064 , \24805 , \24809 );
xor \U$24687 ( \25065 , \25064 , \24814 );
and \U$24688 ( \25066 , \25062 , \25065 );
and \U$24689 ( \25067 , \25060 , \25065 );
or \U$24690 ( \25068 , \25063 , \25066 , \25067 );
xor \U$24691 ( \25069 , \24664 , \24668 );
xor \U$24692 ( \25070 , \25069 , \24673 );
and \U$24693 ( \25071 , \25068 , \25070 );
xor \U$24694 ( \25072 , \24883 , \24885 );
xor \U$24695 ( \25073 , \25072 , \24888 );
and \U$24696 ( \25074 , \25070 , \25073 );
and \U$24697 ( \25075 , \25068 , \25073 );
or \U$24698 ( \25076 , \25071 , \25074 , \25075 );
and \U$24699 ( \25077 , \25058 , \25076 );
xor \U$24700 ( \25078 , \24782 , \24800 );
xor \U$24701 ( \25079 , \25078 , \24817 );
xor \U$24702 ( \25080 , \24836 , \24852 );
xor \U$24703 ( \25081 , \25080 , \24869 );
and \U$24704 ( \25082 , \25079 , \25081 );
xnor \U$24705 ( \25083 , \24875 , \24877 );
and \U$24706 ( \25084 , \25081 , \25083 );
and \U$24707 ( \25085 , \25079 , \25083 );
or \U$24708 ( \25086 , \25082 , \25084 , \25085 );
and \U$24709 ( \25087 , \25076 , \25086 );
and \U$24710 ( \25088 , \25058 , \25086 );
or \U$24711 ( \25089 , \25077 , \25087 , \25088 );
xor \U$24712 ( \25090 , \24820 , \24872 );
xor \U$24713 ( \25091 , \25090 , \24878 );
xor \U$24714 ( \25092 , \24891 , \24893 );
xor \U$24715 ( \25093 , \25092 , \24896 );
and \U$24716 ( \25094 , \25091 , \25093 );
xor \U$24717 ( \25095 , \24902 , \24904 );
and \U$24718 ( \25096 , \25093 , \25095 );
and \U$24719 ( \25097 , \25091 , \25095 );
or \U$24720 ( \25098 , \25094 , \25096 , \25097 );
and \U$24721 ( \25099 , \25089 , \25098 );
xor \U$24722 ( \25100 , \24910 , \24912 );
xor \U$24723 ( \25101 , \25100 , \24914 );
and \U$24724 ( \25102 , \25098 , \25101 );
and \U$24725 ( \25103 , \25089 , \25101 );
or \U$24726 ( \25104 , \25099 , \25102 , \25103 );
xor \U$24727 ( \25105 , \24710 , \24728 );
xor \U$24728 ( \25106 , \25105 , \24734 );
and \U$24729 ( \25107 , \25104 , \25106 );
xor \U$24730 ( \25108 , \24908 , \24917 );
xor \U$24731 ( \25109 , \25108 , \24920 );
and \U$24732 ( \25110 , \25106 , \25109 );
and \U$24733 ( \25111 , \25104 , \25109 );
or \U$24734 ( \25112 , \25107 , \25110 , \25111 );
xor \U$24735 ( \25113 , \24923 , \24925 );
xor \U$24736 ( \25114 , \25113 , \24928 );
and \U$24737 ( \25115 , \25112 , \25114 );
and \U$24738 ( \25116 , \24937 , \25115 );
xor \U$24739 ( \25117 , \24937 , \25115 );
xor \U$24740 ( \25118 , \25112 , \25114 );
buf \U$24741 ( \25119 , RIc226458_38);
buf \U$24742 ( \25120 , RIc2263e0_39);
and \U$24743 ( \25121 , \25119 , \25120 );
not \U$24744 ( \25122 , \25121 );
and \U$24745 ( \25123 , \24784 , \25122 );
not \U$24746 ( \25124 , \25123 );
and \U$24747 ( \25125 , \21667 , \24974 );
and \U$24748 ( \25126 , \21653 , \24972 );
nor \U$24749 ( \25127 , \25125 , \25126 );
xnor \U$24750 ( \25128 , \25127 , \24787 );
and \U$24751 ( \25129 , \25124 , \25128 );
and \U$24752 ( \25130 , \21706 , \24661 );
and \U$24753 ( \25131 , \21685 , \24659 );
nor \U$24754 ( \25132 , \25130 , \25131 );
xnor \U$24755 ( \25133 , \25132 , \24456 );
and \U$24756 ( \25134 , \25128 , \25133 );
and \U$24757 ( \25135 , \25124 , \25133 );
or \U$24758 ( \25136 , \25129 , \25134 , \25135 );
and \U$24759 ( \25137 , \21762 , \24255 );
and \U$24760 ( \25138 , \21754 , \24253 );
nor \U$24761 ( \25139 , \25137 , \25138 );
xnor \U$24762 ( \25140 , \25139 , \24106 );
and \U$24763 ( \25141 , \21836 , \23933 );
and \U$24764 ( \25142 , \21831 , \23931 );
nor \U$24765 ( \25143 , \25141 , \25142 );
xnor \U$24766 ( \25144 , \25143 , \23791 );
and \U$24767 ( \25145 , \25140 , \25144 );
and \U$24768 ( \25146 , \21941 , \23637 );
and \U$24769 ( \25147 , \21890 , \23635 );
nor \U$24770 ( \25148 , \25146 , \25147 );
xnor \U$24771 ( \25149 , \25148 , \23500 );
and \U$24772 ( \25150 , \25144 , \25149 );
and \U$24773 ( \25151 , \25140 , \25149 );
or \U$24774 ( \25152 , \25145 , \25150 , \25151 );
and \U$24775 ( \25153 , \25136 , \25152 );
and \U$24776 ( \25154 , \22046 , \23431 );
and \U$24777 ( \25155 , \22018 , \23429 );
nor \U$24778 ( \25156 , \25154 , \25155 );
xnor \U$24779 ( \25157 , \25156 , \23279 );
and \U$24780 ( \25158 , \22200 , \23163 );
and \U$24781 ( \25159 , \22126 , \23161 );
nor \U$24782 ( \25160 , \25158 , \25159 );
xnor \U$24783 ( \25161 , \25160 , \23007 );
and \U$24784 ( \25162 , \25157 , \25161 );
and \U$24785 ( \25163 , \22325 , \22891 );
and \U$24786 ( \25164 , \22262 , \22889 );
nor \U$24787 ( \25165 , \25163 , \25164 );
xnor \U$24788 ( \25166 , \25165 , \22778 );
and \U$24789 ( \25167 , \25161 , \25166 );
and \U$24790 ( \25168 , \25157 , \25166 );
or \U$24791 ( \25169 , \25162 , \25167 , \25168 );
and \U$24792 ( \25170 , \25152 , \25169 );
and \U$24793 ( \25171 , \25136 , \25169 );
or \U$24794 ( \25172 , \25153 , \25170 , \25171 );
and \U$24795 ( \25173 , \23136 , \22163 );
and \U$24796 ( \25174 , \23128 , \22161 );
nor \U$24797 ( \25175 , \25173 , \25174 );
xnor \U$24798 ( \25176 , \25175 , \22091 );
and \U$24799 ( \25177 , \23384 , \22029 );
and \U$24800 ( \25178 , \23379 , \22027 );
nor \U$24801 ( \25179 , \25177 , \25178 );
xnor \U$24802 ( \25180 , \25179 , \21986 );
and \U$24803 ( \25181 , \25176 , \25180 );
and \U$24804 ( \25182 , \23714 , \21916 );
and \U$24805 ( \25183 , \23570 , \21914 );
nor \U$24806 ( \25184 , \25182 , \25183 );
xnor \U$24807 ( \25185 , \25184 , \21867 );
and \U$24808 ( \25186 , \25180 , \25185 );
and \U$24809 ( \25187 , \25176 , \25185 );
or \U$24810 ( \25188 , \25181 , \25186 , \25187 );
and \U$24811 ( \25189 , \22611 , \22697 );
and \U$24812 ( \25190 , \22523 , \22695 );
nor \U$24813 ( \25191 , \25189 , \25190 );
xnor \U$24814 ( \25192 , \25191 , \22561 );
and \U$24815 ( \25193 , \22721 , \22497 );
and \U$24816 ( \25194 , \22716 , \22495 );
nor \U$24817 ( \25195 , \25193 , \25194 );
xnor \U$24818 ( \25196 , \25195 , \22419 );
and \U$24819 ( \25197 , \25192 , \25196 );
and \U$24820 ( \25198 , \22952 , \22333 );
and \U$24821 ( \25199 , \22837 , \22331 );
nor \U$24822 ( \25200 , \25198 , \25199 );
xnor \U$24823 ( \25201 , \25200 , \22239 );
and \U$24824 ( \25202 , \25196 , \25201 );
and \U$24825 ( \25203 , \25192 , \25201 );
or \U$24826 ( \25204 , \25197 , \25202 , \25203 );
and \U$24827 ( \25205 , \25188 , \25204 );
and \U$24828 ( \25206 , \24003 , \21815 );
and \U$24829 ( \25207 , \23978 , \21813 );
nor \U$24830 ( \25208 , \25206 , \25207 );
xnor \U$24831 ( \25209 , \25208 , \21774 );
and \U$24832 ( \25210 , \24344 , \21745 );
and \U$24833 ( \25211 , \24177 , \21743 );
nor \U$24834 ( \25212 , \25210 , \25211 );
xnor \U$24835 ( \25213 , \25212 , \21715 );
and \U$24836 ( \25214 , \25209 , \25213 );
and \U$24837 ( \25215 , \24601 , \21697 );
and \U$24838 ( \25216 , \24482 , \21695 );
nor \U$24839 ( \25217 , \25215 , \25216 );
xnor \U$24840 ( \25218 , \25217 , \21678 );
and \U$24841 ( \25219 , \25213 , \25218 );
and \U$24842 ( \25220 , \25209 , \25218 );
or \U$24843 ( \25221 , \25214 , \25219 , \25220 );
and \U$24844 ( \25222 , \25204 , \25221 );
and \U$24845 ( \25223 , \25188 , \25221 );
or \U$24846 ( \25224 , \25205 , \25222 , \25223 );
and \U$24847 ( \25225 , \25172 , \25224 );
buf \U$24848 ( \25226 , RIc22a5f8_164);
and \U$24849 ( \25227 , \25226 , \21654 );
xor \U$24850 ( \25228 , \25012 , \25016 );
xor \U$24851 ( \25229 , \25228 , \25022 );
or \U$24852 ( \25230 , \25227 , \25229 );
and \U$24853 ( \25231 , \25224 , \25230 );
and \U$24854 ( \25232 , \25172 , \25230 );
or \U$24855 ( \25233 , \25225 , \25231 , \25232 );
xor \U$24856 ( \25234 , \24941 , \24945 );
xor \U$24857 ( \25235 , \25234 , \24950 );
xor \U$24858 ( \25236 , \24996 , \25000 );
xor \U$24859 ( \25237 , \25236 , \25005 );
and \U$24860 ( \25238 , \25235 , \25237 );
xor \U$24861 ( \25239 , \25030 , \25034 );
xor \U$24862 ( \25240 , \25239 , \25039 );
and \U$24863 ( \25241 , \25237 , \25240 );
and \U$24864 ( \25242 , \25235 , \25240 );
or \U$24865 ( \25243 , \25238 , \25241 , \25242 );
xor \U$24866 ( \25244 , \24788 , \24792 );
xor \U$24867 ( \25245 , \25244 , \24797 );
and \U$24868 ( \25246 , \25243 , \25245 );
xor \U$24869 ( \25247 , \25060 , \25062 );
xor \U$24870 ( \25248 , \25247 , \25065 );
and \U$24871 ( \25249 , \25245 , \25248 );
and \U$24872 ( \25250 , \25243 , \25248 );
or \U$24873 ( \25251 , \25246 , \25249 , \25250 );
and \U$24874 ( \25252 , \25233 , \25251 );
xor \U$24875 ( \25253 , \24953 , \24969 );
xor \U$24876 ( \25254 , \25253 , \24989 );
xor \U$24877 ( \25255 , \25008 , \25025 );
xor \U$24878 ( \25256 , \25255 , \25042 );
and \U$24879 ( \25257 , \25254 , \25256 );
xor \U$24880 ( \25258 , \25047 , \25049 );
xor \U$24881 ( \25259 , \25258 , \25052 );
and \U$24882 ( \25260 , \25256 , \25259 );
and \U$24883 ( \25261 , \25254 , \25259 );
or \U$24884 ( \25262 , \25257 , \25260 , \25261 );
and \U$24885 ( \25263 , \25251 , \25262 );
and \U$24886 ( \25264 , \25233 , \25262 );
or \U$24887 ( \25265 , \25252 , \25263 , \25264 );
xor \U$24888 ( \25266 , \24992 , \25045 );
xor \U$24889 ( \25267 , \25266 , \25055 );
xor \U$24890 ( \25268 , \25068 , \25070 );
xor \U$24891 ( \25269 , \25268 , \25073 );
and \U$24892 ( \25270 , \25267 , \25269 );
xor \U$24893 ( \25271 , \25079 , \25081 );
xor \U$24894 ( \25272 , \25271 , \25083 );
and \U$24895 ( \25273 , \25269 , \25272 );
and \U$24896 ( \25274 , \25267 , \25272 );
or \U$24897 ( \25275 , \25270 , \25273 , \25274 );
and \U$24898 ( \25276 , \25265 , \25275 );
xor \U$24899 ( \25277 , \25091 , \25093 );
xor \U$24900 ( \25278 , \25277 , \25095 );
and \U$24901 ( \25279 , \25275 , \25278 );
and \U$24902 ( \25280 , \25265 , \25278 );
or \U$24903 ( \25281 , \25276 , \25279 , \25280 );
xor \U$24904 ( \25282 , \24881 , \24899 );
xor \U$24905 ( \25283 , \25282 , \24905 );
and \U$24906 ( \25284 , \25281 , \25283 );
xor \U$24907 ( \25285 , \25089 , \25098 );
xor \U$24908 ( \25286 , \25285 , \25101 );
and \U$24909 ( \25287 , \25283 , \25286 );
and \U$24910 ( \25288 , \25281 , \25286 );
or \U$24911 ( \25289 , \25284 , \25287 , \25288 );
xor \U$24912 ( \25290 , \25104 , \25106 );
xor \U$24913 ( \25291 , \25290 , \25109 );
and \U$24914 ( \25292 , \25289 , \25291 );
and \U$24915 ( \25293 , \25118 , \25292 );
xor \U$24916 ( \25294 , \25118 , \25292 );
xor \U$24917 ( \25295 , \25289 , \25291 );
and \U$24918 ( \25296 , \22716 , \22697 );
and \U$24919 ( \25297 , \22611 , \22695 );
nor \U$24920 ( \25298 , \25296 , \25297 );
xnor \U$24921 ( \25299 , \25298 , \22561 );
and \U$24922 ( \25300 , \22837 , \22497 );
and \U$24923 ( \25301 , \22721 , \22495 );
nor \U$24924 ( \25302 , \25300 , \25301 );
xnor \U$24925 ( \25303 , \25302 , \22419 );
and \U$24926 ( \25304 , \25299 , \25303 );
and \U$24927 ( \25305 , \23128 , \22333 );
and \U$24928 ( \25306 , \22952 , \22331 );
nor \U$24929 ( \25307 , \25305 , \25306 );
xnor \U$24930 ( \25308 , \25307 , \22239 );
and \U$24931 ( \25309 , \25303 , \25308 );
and \U$24932 ( \25310 , \25299 , \25308 );
or \U$24933 ( \25311 , \25304 , \25309 , \25310 );
and \U$24934 ( \25312 , \23379 , \22163 );
and \U$24935 ( \25313 , \23136 , \22161 );
nor \U$24936 ( \25314 , \25312 , \25313 );
xnor \U$24937 ( \25315 , \25314 , \22091 );
and \U$24938 ( \25316 , \23570 , \22029 );
and \U$24939 ( \25317 , \23384 , \22027 );
nor \U$24940 ( \25318 , \25316 , \25317 );
xnor \U$24941 ( \25319 , \25318 , \21986 );
and \U$24942 ( \25320 , \25315 , \25319 );
and \U$24943 ( \25321 , \23978 , \21916 );
and \U$24944 ( \25322 , \23714 , \21914 );
nor \U$24945 ( \25323 , \25321 , \25322 );
xnor \U$24946 ( \25324 , \25323 , \21867 );
and \U$24947 ( \25325 , \25319 , \25324 );
and \U$24948 ( \25326 , \25315 , \25324 );
or \U$24949 ( \25327 , \25320 , \25325 , \25326 );
and \U$24950 ( \25328 , \25311 , \25327 );
and \U$24951 ( \25329 , \24177 , \21815 );
and \U$24952 ( \25330 , \24003 , \21813 );
nor \U$24953 ( \25331 , \25329 , \25330 );
xnor \U$24954 ( \25332 , \25331 , \21774 );
and \U$24955 ( \25333 , \24482 , \21745 );
and \U$24956 ( \25334 , \24344 , \21743 );
nor \U$24957 ( \25335 , \25333 , \25334 );
xnor \U$24958 ( \25336 , \25335 , \21715 );
and \U$24959 ( \25337 , \25332 , \25336 );
and \U$24960 ( \25338 , \25018 , \21697 );
and \U$24961 ( \25339 , \24601 , \21695 );
nor \U$24962 ( \25340 , \25338 , \25339 );
xnor \U$24963 ( \25341 , \25340 , \21678 );
and \U$24964 ( \25342 , \25336 , \25341 );
and \U$24965 ( \25343 , \25332 , \25341 );
or \U$24966 ( \25344 , \25337 , \25342 , \25343 );
and \U$24967 ( \25345 , \25327 , \25344 );
and \U$24968 ( \25346 , \25311 , \25344 );
or \U$24969 ( \25347 , \25328 , \25345 , \25346 );
buf \U$24970 ( \25348 , RIc22a670_165);
and \U$24971 ( \25349 , \25348 , \21660 );
and \U$24972 ( \25350 , \25226 , \21658 );
nor \U$24973 ( \25351 , \25349 , \25350 );
xnor \U$24974 ( \25352 , \25351 , \21665 );
buf \U$24975 ( \25353 , RIc22a6e8_166);
and \U$24976 ( \25354 , \25353 , \21654 );
or \U$24977 ( \25355 , \25352 , \25354 );
and \U$24978 ( \25356 , \25226 , \21660 );
and \U$24979 ( \25357 , \25018 , \21658 );
nor \U$24980 ( \25358 , \25356 , \25357 );
xnor \U$24981 ( \25359 , \25358 , \21665 );
and \U$24982 ( \25360 , \25355 , \25359 );
and \U$24983 ( \25361 , \25348 , \21654 );
and \U$24984 ( \25362 , \25359 , \25361 );
and \U$24985 ( \25363 , \25355 , \25361 );
or \U$24986 ( \25364 , \25360 , \25362 , \25363 );
and \U$24987 ( \25365 , \25347 , \25364 );
xor \U$24988 ( \25366 , \24784 , \25119 );
xor \U$24989 ( \25367 , \25119 , \25120 );
not \U$24990 ( \25368 , \25367 );
and \U$24991 ( \25369 , \25366 , \25368 );
and \U$24992 ( \25370 , \21653 , \25369 );
not \U$24993 ( \25371 , \25370 );
xnor \U$24994 ( \25372 , \25371 , \25123 );
and \U$24995 ( \25373 , \21685 , \24974 );
and \U$24996 ( \25374 , \21667 , \24972 );
nor \U$24997 ( \25375 , \25373 , \25374 );
xnor \U$24998 ( \25376 , \25375 , \24787 );
and \U$24999 ( \25377 , \25372 , \25376 );
and \U$25000 ( \25378 , \21754 , \24661 );
and \U$25001 ( \25379 , \21706 , \24659 );
nor \U$25002 ( \25380 , \25378 , \25379 );
xnor \U$25003 ( \25381 , \25380 , \24456 );
and \U$25004 ( \25382 , \25376 , \25381 );
and \U$25005 ( \25383 , \25372 , \25381 );
or \U$25006 ( \25384 , \25377 , \25382 , \25383 );
and \U$25007 ( \25385 , \21831 , \24255 );
and \U$25008 ( \25386 , \21762 , \24253 );
nor \U$25009 ( \25387 , \25385 , \25386 );
xnor \U$25010 ( \25388 , \25387 , \24106 );
and \U$25011 ( \25389 , \21890 , \23933 );
and \U$25012 ( \25390 , \21836 , \23931 );
nor \U$25013 ( \25391 , \25389 , \25390 );
xnor \U$25014 ( \25392 , \25391 , \23791 );
and \U$25015 ( \25393 , \25388 , \25392 );
and \U$25016 ( \25394 , \22018 , \23637 );
and \U$25017 ( \25395 , \21941 , \23635 );
nor \U$25018 ( \25396 , \25394 , \25395 );
xnor \U$25019 ( \25397 , \25396 , \23500 );
and \U$25020 ( \25398 , \25392 , \25397 );
and \U$25021 ( \25399 , \25388 , \25397 );
or \U$25022 ( \25400 , \25393 , \25398 , \25399 );
and \U$25023 ( \25401 , \25384 , \25400 );
and \U$25024 ( \25402 , \22126 , \23431 );
and \U$25025 ( \25403 , \22046 , \23429 );
nor \U$25026 ( \25404 , \25402 , \25403 );
xnor \U$25027 ( \25405 , \25404 , \23279 );
and \U$25028 ( \25406 , \22262 , \23163 );
and \U$25029 ( \25407 , \22200 , \23161 );
nor \U$25030 ( \25408 , \25406 , \25407 );
xnor \U$25031 ( \25409 , \25408 , \23007 );
and \U$25032 ( \25410 , \25405 , \25409 );
and \U$25033 ( \25411 , \22523 , \22891 );
and \U$25034 ( \25412 , \22325 , \22889 );
nor \U$25035 ( \25413 , \25411 , \25412 );
xnor \U$25036 ( \25414 , \25413 , \22778 );
and \U$25037 ( \25415 , \25409 , \25414 );
and \U$25038 ( \25416 , \25405 , \25414 );
or \U$25039 ( \25417 , \25410 , \25415 , \25416 );
and \U$25040 ( \25418 , \25400 , \25417 );
and \U$25041 ( \25419 , \25384 , \25417 );
or \U$25042 ( \25420 , \25401 , \25418 , \25419 );
and \U$25043 ( \25421 , \25364 , \25420 );
and \U$25044 ( \25422 , \25347 , \25420 );
or \U$25045 ( \25423 , \25365 , \25421 , \25422 );
xor \U$25046 ( \25424 , \25176 , \25180 );
xor \U$25047 ( \25425 , \25424 , \25185 );
xor \U$25048 ( \25426 , \25192 , \25196 );
xor \U$25049 ( \25427 , \25426 , \25201 );
and \U$25050 ( \25428 , \25425 , \25427 );
xor \U$25051 ( \25429 , \25209 , \25213 );
xor \U$25052 ( \25430 , \25429 , \25218 );
and \U$25053 ( \25431 , \25427 , \25430 );
and \U$25054 ( \25432 , \25425 , \25430 );
or \U$25055 ( \25433 , \25428 , \25431 , \25432 );
xor \U$25056 ( \25434 , \25124 , \25128 );
xor \U$25057 ( \25435 , \25434 , \25133 );
xor \U$25058 ( \25436 , \25140 , \25144 );
xor \U$25059 ( \25437 , \25436 , \25149 );
and \U$25060 ( \25438 , \25435 , \25437 );
xor \U$25061 ( \25439 , \25157 , \25161 );
xor \U$25062 ( \25440 , \25439 , \25166 );
and \U$25063 ( \25441 , \25437 , \25440 );
and \U$25064 ( \25442 , \25435 , \25440 );
or \U$25065 ( \25443 , \25438 , \25441 , \25442 );
and \U$25066 ( \25444 , \25433 , \25443 );
xor \U$25067 ( \25445 , \24957 , \24961 );
xor \U$25068 ( \25446 , \25445 , \24966 );
and \U$25069 ( \25447 , \25443 , \25446 );
and \U$25070 ( \25448 , \25433 , \25446 );
or \U$25071 ( \25449 , \25444 , \25447 , \25448 );
and \U$25072 ( \25450 , \25423 , \25449 );
xor \U$25073 ( \25451 , \24977 , \24981 );
xor \U$25074 ( \25452 , \25451 , \24986 );
xor \U$25075 ( \25453 , \25235 , \25237 );
xor \U$25076 ( \25454 , \25453 , \25240 );
and \U$25077 ( \25455 , \25452 , \25454 );
xnor \U$25078 ( \25456 , \25227 , \25229 );
and \U$25079 ( \25457 , \25454 , \25456 );
and \U$25080 ( \25458 , \25452 , \25456 );
or \U$25081 ( \25459 , \25455 , \25457 , \25458 );
and \U$25082 ( \25460 , \25449 , \25459 );
and \U$25083 ( \25461 , \25423 , \25459 );
or \U$25084 ( \25462 , \25450 , \25460 , \25461 );
xor \U$25085 ( \25463 , \25172 , \25224 );
xor \U$25086 ( \25464 , \25463 , \25230 );
xor \U$25087 ( \25465 , \25243 , \25245 );
xor \U$25088 ( \25466 , \25465 , \25248 );
and \U$25089 ( \25467 , \25464 , \25466 );
xor \U$25090 ( \25468 , \25254 , \25256 );
xor \U$25091 ( \25469 , \25468 , \25259 );
and \U$25092 ( \25470 , \25466 , \25469 );
and \U$25093 ( \25471 , \25464 , \25469 );
or \U$25094 ( \25472 , \25467 , \25470 , \25471 );
and \U$25095 ( \25473 , \25462 , \25472 );
xor \U$25096 ( \25474 , \25267 , \25269 );
xor \U$25097 ( \25475 , \25474 , \25272 );
and \U$25098 ( \25476 , \25472 , \25475 );
and \U$25099 ( \25477 , \25462 , \25475 );
or \U$25100 ( \25478 , \25473 , \25476 , \25477 );
xor \U$25101 ( \25479 , \25058 , \25076 );
xor \U$25102 ( \25480 , \25479 , \25086 );
and \U$25103 ( \25481 , \25478 , \25480 );
xor \U$25104 ( \25482 , \25265 , \25275 );
xor \U$25105 ( \25483 , \25482 , \25278 );
and \U$25106 ( \25484 , \25480 , \25483 );
and \U$25107 ( \25485 , \25478 , \25483 );
or \U$25108 ( \25486 , \25481 , \25484 , \25485 );
xor \U$25109 ( \25487 , \25281 , \25283 );
xor \U$25110 ( \25488 , \25487 , \25286 );
and \U$25111 ( \25489 , \25486 , \25488 );
and \U$25112 ( \25490 , \25295 , \25489 );
xor \U$25113 ( \25491 , \25295 , \25489 );
xor \U$25114 ( \25492 , \25486 , \25488 );
and \U$25115 ( \25493 , \23136 , \22333 );
and \U$25116 ( \25494 , \23128 , \22331 );
nor \U$25117 ( \25495 , \25493 , \25494 );
xnor \U$25118 ( \25496 , \25495 , \22239 );
and \U$25119 ( \25497 , \23384 , \22163 );
and \U$25120 ( \25498 , \23379 , \22161 );
nor \U$25121 ( \25499 , \25497 , \25498 );
xnor \U$25122 ( \25500 , \25499 , \22091 );
and \U$25123 ( \25501 , \25496 , \25500 );
and \U$25124 ( \25502 , \23714 , \22029 );
and \U$25125 ( \25503 , \23570 , \22027 );
nor \U$25126 ( \25504 , \25502 , \25503 );
xnor \U$25127 ( \25505 , \25504 , \21986 );
and \U$25128 ( \25506 , \25500 , \25505 );
and \U$25129 ( \25507 , \25496 , \25505 );
or \U$25130 ( \25508 , \25501 , \25506 , \25507 );
and \U$25131 ( \25509 , \22611 , \22891 );
and \U$25132 ( \25510 , \22523 , \22889 );
nor \U$25133 ( \25511 , \25509 , \25510 );
xnor \U$25134 ( \25512 , \25511 , \22778 );
and \U$25135 ( \25513 , \22721 , \22697 );
and \U$25136 ( \25514 , \22716 , \22695 );
nor \U$25137 ( \25515 , \25513 , \25514 );
xnor \U$25138 ( \25516 , \25515 , \22561 );
and \U$25139 ( \25517 , \25512 , \25516 );
and \U$25140 ( \25518 , \22952 , \22497 );
and \U$25141 ( \25519 , \22837 , \22495 );
nor \U$25142 ( \25520 , \25518 , \25519 );
xnor \U$25143 ( \25521 , \25520 , \22419 );
and \U$25144 ( \25522 , \25516 , \25521 );
and \U$25145 ( \25523 , \25512 , \25521 );
or \U$25146 ( \25524 , \25517 , \25522 , \25523 );
and \U$25147 ( \25525 , \25508 , \25524 );
and \U$25148 ( \25526 , \24003 , \21916 );
and \U$25149 ( \25527 , \23978 , \21914 );
nor \U$25150 ( \25528 , \25526 , \25527 );
xnor \U$25151 ( \25529 , \25528 , \21867 );
and \U$25152 ( \25530 , \24344 , \21815 );
and \U$25153 ( \25531 , \24177 , \21813 );
nor \U$25154 ( \25532 , \25530 , \25531 );
xnor \U$25155 ( \25533 , \25532 , \21774 );
and \U$25156 ( \25534 , \25529 , \25533 );
and \U$25157 ( \25535 , \24601 , \21745 );
and \U$25158 ( \25536 , \24482 , \21743 );
nor \U$25159 ( \25537 , \25535 , \25536 );
xnor \U$25160 ( \25538 , \25537 , \21715 );
and \U$25161 ( \25539 , \25533 , \25538 );
and \U$25162 ( \25540 , \25529 , \25538 );
or \U$25163 ( \25541 , \25534 , \25539 , \25540 );
and \U$25164 ( \25542 , \25524 , \25541 );
and \U$25165 ( \25543 , \25508 , \25541 );
or \U$25166 ( \25544 , \25525 , \25542 , \25543 );
buf \U$25167 ( \25545 , RIc226368_40);
buf \U$25168 ( \25546 , RIc2262f0_41);
and \U$25169 ( \25547 , \25545 , \25546 );
not \U$25170 ( \25548 , \25547 );
and \U$25171 ( \25549 , \25120 , \25548 );
not \U$25172 ( \25550 , \25549 );
and \U$25173 ( \25551 , \21667 , \25369 );
and \U$25174 ( \25552 , \21653 , \25367 );
nor \U$25175 ( \25553 , \25551 , \25552 );
xnor \U$25176 ( \25554 , \25553 , \25123 );
and \U$25177 ( \25555 , \25550 , \25554 );
and \U$25178 ( \25556 , \21706 , \24974 );
and \U$25179 ( \25557 , \21685 , \24972 );
nor \U$25180 ( \25558 , \25556 , \25557 );
xnor \U$25181 ( \25559 , \25558 , \24787 );
and \U$25182 ( \25560 , \25554 , \25559 );
and \U$25183 ( \25561 , \25550 , \25559 );
or \U$25184 ( \25562 , \25555 , \25560 , \25561 );
and \U$25185 ( \25563 , \21762 , \24661 );
and \U$25186 ( \25564 , \21754 , \24659 );
nor \U$25187 ( \25565 , \25563 , \25564 );
xnor \U$25188 ( \25566 , \25565 , \24456 );
and \U$25189 ( \25567 , \21836 , \24255 );
and \U$25190 ( \25568 , \21831 , \24253 );
nor \U$25191 ( \25569 , \25567 , \25568 );
xnor \U$25192 ( \25570 , \25569 , \24106 );
and \U$25193 ( \25571 , \25566 , \25570 );
and \U$25194 ( \25572 , \21941 , \23933 );
and \U$25195 ( \25573 , \21890 , \23931 );
nor \U$25196 ( \25574 , \25572 , \25573 );
xnor \U$25197 ( \25575 , \25574 , \23791 );
and \U$25198 ( \25576 , \25570 , \25575 );
and \U$25199 ( \25577 , \25566 , \25575 );
or \U$25200 ( \25578 , \25571 , \25576 , \25577 );
and \U$25201 ( \25579 , \25562 , \25578 );
and \U$25202 ( \25580 , \22046 , \23637 );
and \U$25203 ( \25581 , \22018 , \23635 );
nor \U$25204 ( \25582 , \25580 , \25581 );
xnor \U$25205 ( \25583 , \25582 , \23500 );
and \U$25206 ( \25584 , \22200 , \23431 );
and \U$25207 ( \25585 , \22126 , \23429 );
nor \U$25208 ( \25586 , \25584 , \25585 );
xnor \U$25209 ( \25587 , \25586 , \23279 );
and \U$25210 ( \25588 , \25583 , \25587 );
and \U$25211 ( \25589 , \22325 , \23163 );
and \U$25212 ( \25590 , \22262 , \23161 );
nor \U$25213 ( \25591 , \25589 , \25590 );
xnor \U$25214 ( \25592 , \25591 , \23007 );
and \U$25215 ( \25593 , \25587 , \25592 );
and \U$25216 ( \25594 , \25583 , \25592 );
or \U$25217 ( \25595 , \25588 , \25593 , \25594 );
and \U$25218 ( \25596 , \25578 , \25595 );
and \U$25219 ( \25597 , \25562 , \25595 );
or \U$25220 ( \25598 , \25579 , \25596 , \25597 );
and \U$25221 ( \25599 , \25544 , \25598 );
and \U$25222 ( \25600 , \25226 , \21697 );
and \U$25223 ( \25601 , \25018 , \21695 );
nor \U$25224 ( \25602 , \25600 , \25601 );
xnor \U$25225 ( \25603 , \25602 , \21678 );
and \U$25226 ( \25604 , \25353 , \21660 );
and \U$25227 ( \25605 , \25348 , \21658 );
nor \U$25228 ( \25606 , \25604 , \25605 );
xnor \U$25229 ( \25607 , \25606 , \21665 );
and \U$25230 ( \25608 , \25603 , \25607 );
buf \U$25231 ( \25609 , RIc22a760_167);
and \U$25232 ( \25610 , \25609 , \21654 );
and \U$25233 ( \25611 , \25607 , \25610 );
and \U$25234 ( \25612 , \25603 , \25610 );
or \U$25235 ( \25613 , \25608 , \25611 , \25612 );
xor \U$25236 ( \25614 , \25332 , \25336 );
xor \U$25237 ( \25615 , \25614 , \25341 );
and \U$25238 ( \25616 , \25613 , \25615 );
xnor \U$25239 ( \25617 , \25352 , \25354 );
and \U$25240 ( \25618 , \25615 , \25617 );
and \U$25241 ( \25619 , \25613 , \25617 );
or \U$25242 ( \25620 , \25616 , \25618 , \25619 );
and \U$25243 ( \25621 , \25598 , \25620 );
and \U$25244 ( \25622 , \25544 , \25620 );
or \U$25245 ( \25623 , \25599 , \25621 , \25622 );
xor \U$25246 ( \25624 , \25299 , \25303 );
xor \U$25247 ( \25625 , \25624 , \25308 );
xor \U$25248 ( \25626 , \25315 , \25319 );
xor \U$25249 ( \25627 , \25626 , \25324 );
and \U$25250 ( \25628 , \25625 , \25627 );
xor \U$25251 ( \25629 , \25405 , \25409 );
xor \U$25252 ( \25630 , \25629 , \25414 );
and \U$25253 ( \25631 , \25627 , \25630 );
and \U$25254 ( \25632 , \25625 , \25630 );
or \U$25255 ( \25633 , \25628 , \25631 , \25632 );
xor \U$25256 ( \25634 , \25372 , \25376 );
xor \U$25257 ( \25635 , \25634 , \25381 );
xor \U$25258 ( \25636 , \25388 , \25392 );
xor \U$25259 ( \25637 , \25636 , \25397 );
and \U$25260 ( \25638 , \25635 , \25637 );
and \U$25261 ( \25639 , \25633 , \25638 );
xor \U$25262 ( \25640 , \25435 , \25437 );
xor \U$25263 ( \25641 , \25640 , \25440 );
and \U$25264 ( \25642 , \25638 , \25641 );
and \U$25265 ( \25643 , \25633 , \25641 );
or \U$25266 ( \25644 , \25639 , \25642 , \25643 );
and \U$25267 ( \25645 , \25623 , \25644 );
xor \U$25268 ( \25646 , \25311 , \25327 );
xor \U$25269 ( \25647 , \25646 , \25344 );
xor \U$25270 ( \25648 , \25355 , \25359 );
xor \U$25271 ( \25649 , \25648 , \25361 );
and \U$25272 ( \25650 , \25647 , \25649 );
xor \U$25273 ( \25651 , \25425 , \25427 );
xor \U$25274 ( \25652 , \25651 , \25430 );
and \U$25275 ( \25653 , \25649 , \25652 );
and \U$25276 ( \25654 , \25647 , \25652 );
or \U$25277 ( \25655 , \25650 , \25653 , \25654 );
and \U$25278 ( \25656 , \25644 , \25655 );
and \U$25279 ( \25657 , \25623 , \25655 );
or \U$25280 ( \25658 , \25645 , \25656 , \25657 );
xor \U$25281 ( \25659 , \25136 , \25152 );
xor \U$25282 ( \25660 , \25659 , \25169 );
xor \U$25283 ( \25661 , \25188 , \25204 );
xor \U$25284 ( \25662 , \25661 , \25221 );
and \U$25285 ( \25663 , \25660 , \25662 );
xor \U$25286 ( \25664 , \25452 , \25454 );
xor \U$25287 ( \25665 , \25664 , \25456 );
and \U$25288 ( \25666 , \25662 , \25665 );
and \U$25289 ( \25667 , \25660 , \25665 );
or \U$25290 ( \25668 , \25663 , \25666 , \25667 );
and \U$25291 ( \25669 , \25658 , \25668 );
xor \U$25292 ( \25670 , \25464 , \25466 );
xor \U$25293 ( \25671 , \25670 , \25469 );
and \U$25294 ( \25672 , \25668 , \25671 );
and \U$25295 ( \25673 , \25658 , \25671 );
or \U$25296 ( \25674 , \25669 , \25672 , \25673 );
xor \U$25297 ( \25675 , \25233 , \25251 );
xor \U$25298 ( \25676 , \25675 , \25262 );
and \U$25299 ( \25677 , \25674 , \25676 );
xor \U$25300 ( \25678 , \25462 , \25472 );
xor \U$25301 ( \25679 , \25678 , \25475 );
and \U$25302 ( \25680 , \25676 , \25679 );
and \U$25303 ( \25681 , \25674 , \25679 );
or \U$25304 ( \25682 , \25677 , \25680 , \25681 );
xor \U$25305 ( \25683 , \25478 , \25480 );
xor \U$25306 ( \25684 , \25683 , \25483 );
and \U$25307 ( \25685 , \25682 , \25684 );
and \U$25308 ( \25686 , \25492 , \25685 );
xor \U$25309 ( \25687 , \25492 , \25685 );
xor \U$25310 ( \25688 , \25682 , \25684 );
xor \U$25311 ( \25689 , \25120 , \25545 );
xor \U$25312 ( \25690 , \25545 , \25546 );
not \U$25313 ( \25691 , \25690 );
and \U$25314 ( \25692 , \25689 , \25691 );
and \U$25315 ( \25693 , \21653 , \25692 );
not \U$25316 ( \25694 , \25693 );
xnor \U$25317 ( \25695 , \25694 , \25549 );
and \U$25318 ( \25696 , \21685 , \25369 );
and \U$25319 ( \25697 , \21667 , \25367 );
nor \U$25320 ( \25698 , \25696 , \25697 );
xnor \U$25321 ( \25699 , \25698 , \25123 );
and \U$25322 ( \25700 , \25695 , \25699 );
and \U$25323 ( \25701 , \21754 , \24974 );
and \U$25324 ( \25702 , \21706 , \24972 );
nor \U$25325 ( \25703 , \25701 , \25702 );
xnor \U$25326 ( \25704 , \25703 , \24787 );
and \U$25327 ( \25705 , \25699 , \25704 );
and \U$25328 ( \25706 , \25695 , \25704 );
or \U$25329 ( \25707 , \25700 , \25705 , \25706 );
and \U$25330 ( \25708 , \21831 , \24661 );
and \U$25331 ( \25709 , \21762 , \24659 );
nor \U$25332 ( \25710 , \25708 , \25709 );
xnor \U$25333 ( \25711 , \25710 , \24456 );
and \U$25334 ( \25712 , \21890 , \24255 );
and \U$25335 ( \25713 , \21836 , \24253 );
nor \U$25336 ( \25714 , \25712 , \25713 );
xnor \U$25337 ( \25715 , \25714 , \24106 );
and \U$25338 ( \25716 , \25711 , \25715 );
and \U$25339 ( \25717 , \22018 , \23933 );
and \U$25340 ( \25718 , \21941 , \23931 );
nor \U$25341 ( \25719 , \25717 , \25718 );
xnor \U$25342 ( \25720 , \25719 , \23791 );
and \U$25343 ( \25721 , \25715 , \25720 );
and \U$25344 ( \25722 , \25711 , \25720 );
or \U$25345 ( \25723 , \25716 , \25721 , \25722 );
and \U$25346 ( \25724 , \25707 , \25723 );
and \U$25347 ( \25725 , \22126 , \23637 );
and \U$25348 ( \25726 , \22046 , \23635 );
nor \U$25349 ( \25727 , \25725 , \25726 );
xnor \U$25350 ( \25728 , \25727 , \23500 );
and \U$25351 ( \25729 , \22262 , \23431 );
and \U$25352 ( \25730 , \22200 , \23429 );
nor \U$25353 ( \25731 , \25729 , \25730 );
xnor \U$25354 ( \25732 , \25731 , \23279 );
and \U$25355 ( \25733 , \25728 , \25732 );
and \U$25356 ( \25734 , \22523 , \23163 );
and \U$25357 ( \25735 , \22325 , \23161 );
nor \U$25358 ( \25736 , \25734 , \25735 );
xnor \U$25359 ( \25737 , \25736 , \23007 );
and \U$25360 ( \25738 , \25732 , \25737 );
and \U$25361 ( \25739 , \25728 , \25737 );
or \U$25362 ( \25740 , \25733 , \25738 , \25739 );
and \U$25363 ( \25741 , \25723 , \25740 );
and \U$25364 ( \25742 , \25707 , \25740 );
or \U$25365 ( \25743 , \25724 , \25741 , \25742 );
and \U$25366 ( \25744 , \24177 , \21916 );
and \U$25367 ( \25745 , \24003 , \21914 );
nor \U$25368 ( \25746 , \25744 , \25745 );
xnor \U$25369 ( \25747 , \25746 , \21867 );
and \U$25370 ( \25748 , \24482 , \21815 );
and \U$25371 ( \25749 , \24344 , \21813 );
nor \U$25372 ( \25750 , \25748 , \25749 );
xnor \U$25373 ( \25751 , \25750 , \21774 );
and \U$25374 ( \25752 , \25747 , \25751 );
and \U$25375 ( \25753 , \25018 , \21745 );
and \U$25376 ( \25754 , \24601 , \21743 );
nor \U$25377 ( \25755 , \25753 , \25754 );
xnor \U$25378 ( \25756 , \25755 , \21715 );
and \U$25379 ( \25757 , \25751 , \25756 );
and \U$25380 ( \25758 , \25747 , \25756 );
or \U$25381 ( \25759 , \25752 , \25757 , \25758 );
and \U$25382 ( \25760 , \22716 , \22891 );
and \U$25383 ( \25761 , \22611 , \22889 );
nor \U$25384 ( \25762 , \25760 , \25761 );
xnor \U$25385 ( \25763 , \25762 , \22778 );
and \U$25386 ( \25764 , \22837 , \22697 );
and \U$25387 ( \25765 , \22721 , \22695 );
nor \U$25388 ( \25766 , \25764 , \25765 );
xnor \U$25389 ( \25767 , \25766 , \22561 );
and \U$25390 ( \25768 , \25763 , \25767 );
and \U$25391 ( \25769 , \23128 , \22497 );
and \U$25392 ( \25770 , \22952 , \22495 );
nor \U$25393 ( \25771 , \25769 , \25770 );
xnor \U$25394 ( \25772 , \25771 , \22419 );
and \U$25395 ( \25773 , \25767 , \25772 );
and \U$25396 ( \25774 , \25763 , \25772 );
or \U$25397 ( \25775 , \25768 , \25773 , \25774 );
and \U$25398 ( \25776 , \25759 , \25775 );
and \U$25399 ( \25777 , \23379 , \22333 );
and \U$25400 ( \25778 , \23136 , \22331 );
nor \U$25401 ( \25779 , \25777 , \25778 );
xnor \U$25402 ( \25780 , \25779 , \22239 );
and \U$25403 ( \25781 , \23570 , \22163 );
and \U$25404 ( \25782 , \23384 , \22161 );
nor \U$25405 ( \25783 , \25781 , \25782 );
xnor \U$25406 ( \25784 , \25783 , \22091 );
and \U$25407 ( \25785 , \25780 , \25784 );
and \U$25408 ( \25786 , \23978 , \22029 );
and \U$25409 ( \25787 , \23714 , \22027 );
nor \U$25410 ( \25788 , \25786 , \25787 );
xnor \U$25411 ( \25789 , \25788 , \21986 );
and \U$25412 ( \25790 , \25784 , \25789 );
and \U$25413 ( \25791 , \25780 , \25789 );
or \U$25414 ( \25792 , \25785 , \25790 , \25791 );
and \U$25415 ( \25793 , \25775 , \25792 );
and \U$25416 ( \25794 , \25759 , \25792 );
or \U$25417 ( \25795 , \25776 , \25793 , \25794 );
and \U$25418 ( \25796 , \25743 , \25795 );
and \U$25419 ( \25797 , \25348 , \21697 );
and \U$25420 ( \25798 , \25226 , \21695 );
nor \U$25421 ( \25799 , \25797 , \25798 );
xnor \U$25422 ( \25800 , \25799 , \21678 );
and \U$25423 ( \25801 , \25609 , \21660 );
and \U$25424 ( \25802 , \25353 , \21658 );
nor \U$25425 ( \25803 , \25801 , \25802 );
xnor \U$25426 ( \25804 , \25803 , \21665 );
and \U$25427 ( \25805 , \25800 , \25804 );
buf \U$25428 ( \25806 , RIc22a7d8_168);
and \U$25429 ( \25807 , \25806 , \21654 );
and \U$25430 ( \25808 , \25804 , \25807 );
and \U$25431 ( \25809 , \25800 , \25807 );
or \U$25432 ( \25810 , \25805 , \25808 , \25809 );
xor \U$25433 ( \25811 , \25603 , \25607 );
xor \U$25434 ( \25812 , \25811 , \25610 );
and \U$25435 ( \25813 , \25810 , \25812 );
xor \U$25436 ( \25814 , \25529 , \25533 );
xor \U$25437 ( \25815 , \25814 , \25538 );
and \U$25438 ( \25816 , \25812 , \25815 );
and \U$25439 ( \25817 , \25810 , \25815 );
or \U$25440 ( \25818 , \25813 , \25816 , \25817 );
and \U$25441 ( \25819 , \25795 , \25818 );
and \U$25442 ( \25820 , \25743 , \25818 );
or \U$25443 ( \25821 , \25796 , \25819 , \25820 );
xor \U$25444 ( \25822 , \25508 , \25524 );
xor \U$25445 ( \25823 , \25822 , \25541 );
xor \U$25446 ( \25824 , \25562 , \25578 );
xor \U$25447 ( \25825 , \25824 , \25595 );
and \U$25448 ( \25826 , \25823 , \25825 );
xor \U$25449 ( \25827 , \25613 , \25615 );
xor \U$25450 ( \25828 , \25827 , \25617 );
and \U$25451 ( \25829 , \25825 , \25828 );
and \U$25452 ( \25830 , \25823 , \25828 );
or \U$25453 ( \25831 , \25826 , \25829 , \25830 );
and \U$25454 ( \25832 , \25821 , \25831 );
xor \U$25455 ( \25833 , \25496 , \25500 );
xor \U$25456 ( \25834 , \25833 , \25505 );
xor \U$25457 ( \25835 , \25512 , \25516 );
xor \U$25458 ( \25836 , \25835 , \25521 );
and \U$25459 ( \25837 , \25834 , \25836 );
xor \U$25460 ( \25838 , \25583 , \25587 );
xor \U$25461 ( \25839 , \25838 , \25592 );
and \U$25462 ( \25840 , \25836 , \25839 );
and \U$25463 ( \25841 , \25834 , \25839 );
or \U$25464 ( \25842 , \25837 , \25840 , \25841 );
xor \U$25465 ( \25843 , \25625 , \25627 );
xor \U$25466 ( \25844 , \25843 , \25630 );
and \U$25467 ( \25845 , \25842 , \25844 );
xor \U$25468 ( \25846 , \25635 , \25637 );
and \U$25469 ( \25847 , \25844 , \25846 );
and \U$25470 ( \25848 , \25842 , \25846 );
or \U$25471 ( \25849 , \25845 , \25847 , \25848 );
and \U$25472 ( \25850 , \25831 , \25849 );
and \U$25473 ( \25851 , \25821 , \25849 );
or \U$25474 ( \25852 , \25832 , \25850 , \25851 );
xor \U$25475 ( \25853 , \25384 , \25400 );
xor \U$25476 ( \25854 , \25853 , \25417 );
xor \U$25477 ( \25855 , \25633 , \25638 );
xor \U$25478 ( \25856 , \25855 , \25641 );
and \U$25479 ( \25857 , \25854 , \25856 );
xor \U$25480 ( \25858 , \25647 , \25649 );
xor \U$25481 ( \25859 , \25858 , \25652 );
and \U$25482 ( \25860 , \25856 , \25859 );
and \U$25483 ( \25861 , \25854 , \25859 );
or \U$25484 ( \25862 , \25857 , \25860 , \25861 );
and \U$25485 ( \25863 , \25852 , \25862 );
xor \U$25486 ( \25864 , \25433 , \25443 );
xor \U$25487 ( \25865 , \25864 , \25446 );
and \U$25488 ( \25866 , \25862 , \25865 );
and \U$25489 ( \25867 , \25852 , \25865 );
or \U$25490 ( \25868 , \25863 , \25866 , \25867 );
xor \U$25491 ( \25869 , \25347 , \25364 );
xor \U$25492 ( \25870 , \25869 , \25420 );
xor \U$25493 ( \25871 , \25623 , \25644 );
xor \U$25494 ( \25872 , \25871 , \25655 );
and \U$25495 ( \25873 , \25870 , \25872 );
xor \U$25496 ( \25874 , \25660 , \25662 );
xor \U$25497 ( \25875 , \25874 , \25665 );
and \U$25498 ( \25876 , \25872 , \25875 );
and \U$25499 ( \25877 , \25870 , \25875 );
or \U$25500 ( \25878 , \25873 , \25876 , \25877 );
and \U$25501 ( \25879 , \25868 , \25878 );
xor \U$25502 ( \25880 , \25423 , \25449 );
xor \U$25503 ( \25881 , \25880 , \25459 );
and \U$25504 ( \25882 , \25878 , \25881 );
and \U$25505 ( \25883 , \25868 , \25881 );
or \U$25506 ( \25884 , \25879 , \25882 , \25883 );
xor \U$25507 ( \25885 , \25674 , \25676 );
xor \U$25508 ( \25886 , \25885 , \25679 );
and \U$25509 ( \25887 , \25884 , \25886 );
and \U$25510 ( \25888 , \25688 , \25887 );
xor \U$25511 ( \25889 , \25688 , \25887 );
xor \U$25512 ( \25890 , \25884 , \25886 );
and \U$25513 ( \25891 , \22046 , \23933 );
and \U$25514 ( \25892 , \22018 , \23931 );
nor \U$25515 ( \25893 , \25891 , \25892 );
xnor \U$25516 ( \25894 , \25893 , \23791 );
and \U$25517 ( \25895 , \22200 , \23637 );
and \U$25518 ( \25896 , \22126 , \23635 );
nor \U$25519 ( \25897 , \25895 , \25896 );
xnor \U$25520 ( \25898 , \25897 , \23500 );
and \U$25521 ( \25899 , \25894 , \25898 );
and \U$25522 ( \25900 , \22325 , \23431 );
and \U$25523 ( \25901 , \22262 , \23429 );
nor \U$25524 ( \25902 , \25900 , \25901 );
xnor \U$25525 ( \25903 , \25902 , \23279 );
and \U$25526 ( \25904 , \25898 , \25903 );
and \U$25527 ( \25905 , \25894 , \25903 );
or \U$25528 ( \25906 , \25899 , \25904 , \25905 );
buf \U$25529 ( \25907 , RIc226278_42);
buf \U$25530 ( \25908 , RIc226200_43);
and \U$25531 ( \25909 , \25907 , \25908 );
not \U$25532 ( \25910 , \25909 );
and \U$25533 ( \25911 , \25546 , \25910 );
not \U$25534 ( \25912 , \25911 );
and \U$25535 ( \25913 , \21667 , \25692 );
and \U$25536 ( \25914 , \21653 , \25690 );
nor \U$25537 ( \25915 , \25913 , \25914 );
xnor \U$25538 ( \25916 , \25915 , \25549 );
and \U$25539 ( \25917 , \25912 , \25916 );
and \U$25540 ( \25918 , \21706 , \25369 );
and \U$25541 ( \25919 , \21685 , \25367 );
nor \U$25542 ( \25920 , \25918 , \25919 );
xnor \U$25543 ( \25921 , \25920 , \25123 );
and \U$25544 ( \25922 , \25916 , \25921 );
and \U$25545 ( \25923 , \25912 , \25921 );
or \U$25546 ( \25924 , \25917 , \25922 , \25923 );
and \U$25547 ( \25925 , \25906 , \25924 );
and \U$25548 ( \25926 , \21762 , \24974 );
and \U$25549 ( \25927 , \21754 , \24972 );
nor \U$25550 ( \25928 , \25926 , \25927 );
xnor \U$25551 ( \25929 , \25928 , \24787 );
and \U$25552 ( \25930 , \21836 , \24661 );
and \U$25553 ( \25931 , \21831 , \24659 );
nor \U$25554 ( \25932 , \25930 , \25931 );
xnor \U$25555 ( \25933 , \25932 , \24456 );
and \U$25556 ( \25934 , \25929 , \25933 );
and \U$25557 ( \25935 , \21941 , \24255 );
and \U$25558 ( \25936 , \21890 , \24253 );
nor \U$25559 ( \25937 , \25935 , \25936 );
xnor \U$25560 ( \25938 , \25937 , \24106 );
and \U$25561 ( \25939 , \25933 , \25938 );
and \U$25562 ( \25940 , \25929 , \25938 );
or \U$25563 ( \25941 , \25934 , \25939 , \25940 );
and \U$25564 ( \25942 , \25924 , \25941 );
and \U$25565 ( \25943 , \25906 , \25941 );
or \U$25566 ( \25944 , \25925 , \25942 , \25943 );
and \U$25567 ( \25945 , \24003 , \22029 );
and \U$25568 ( \25946 , \23978 , \22027 );
nor \U$25569 ( \25947 , \25945 , \25946 );
xnor \U$25570 ( \25948 , \25947 , \21986 );
and \U$25571 ( \25949 , \24344 , \21916 );
and \U$25572 ( \25950 , \24177 , \21914 );
nor \U$25573 ( \25951 , \25949 , \25950 );
xnor \U$25574 ( \25952 , \25951 , \21867 );
and \U$25575 ( \25953 , \25948 , \25952 );
and \U$25576 ( \25954 , \24601 , \21815 );
and \U$25577 ( \25955 , \24482 , \21813 );
nor \U$25578 ( \25956 , \25954 , \25955 );
xnor \U$25579 ( \25957 , \25956 , \21774 );
and \U$25580 ( \25958 , \25952 , \25957 );
and \U$25581 ( \25959 , \25948 , \25957 );
or \U$25582 ( \25960 , \25953 , \25958 , \25959 );
and \U$25583 ( \25961 , \22611 , \23163 );
and \U$25584 ( \25962 , \22523 , \23161 );
nor \U$25585 ( \25963 , \25961 , \25962 );
xnor \U$25586 ( \25964 , \25963 , \23007 );
and \U$25587 ( \25965 , \22721 , \22891 );
and \U$25588 ( \25966 , \22716 , \22889 );
nor \U$25589 ( \25967 , \25965 , \25966 );
xnor \U$25590 ( \25968 , \25967 , \22778 );
and \U$25591 ( \25969 , \25964 , \25968 );
and \U$25592 ( \25970 , \22952 , \22697 );
and \U$25593 ( \25971 , \22837 , \22695 );
nor \U$25594 ( \25972 , \25970 , \25971 );
xnor \U$25595 ( \25973 , \25972 , \22561 );
and \U$25596 ( \25974 , \25968 , \25973 );
and \U$25597 ( \25975 , \25964 , \25973 );
or \U$25598 ( \25976 , \25969 , \25974 , \25975 );
and \U$25599 ( \25977 , \25960 , \25976 );
and \U$25600 ( \25978 , \23136 , \22497 );
and \U$25601 ( \25979 , \23128 , \22495 );
nor \U$25602 ( \25980 , \25978 , \25979 );
xnor \U$25603 ( \25981 , \25980 , \22419 );
and \U$25604 ( \25982 , \23384 , \22333 );
and \U$25605 ( \25983 , \23379 , \22331 );
nor \U$25606 ( \25984 , \25982 , \25983 );
xnor \U$25607 ( \25985 , \25984 , \22239 );
and \U$25608 ( \25986 , \25981 , \25985 );
and \U$25609 ( \25987 , \23714 , \22163 );
and \U$25610 ( \25988 , \23570 , \22161 );
nor \U$25611 ( \25989 , \25987 , \25988 );
xnor \U$25612 ( \25990 , \25989 , \22091 );
and \U$25613 ( \25991 , \25985 , \25990 );
and \U$25614 ( \25992 , \25981 , \25990 );
or \U$25615 ( \25993 , \25986 , \25991 , \25992 );
and \U$25616 ( \25994 , \25976 , \25993 );
and \U$25617 ( \25995 , \25960 , \25993 );
or \U$25618 ( \25996 , \25977 , \25994 , \25995 );
and \U$25619 ( \25997 , \25944 , \25996 );
and \U$25620 ( \25998 , \25226 , \21745 );
and \U$25621 ( \25999 , \25018 , \21743 );
nor \U$25622 ( \26000 , \25998 , \25999 );
xnor \U$25623 ( \26001 , \26000 , \21715 );
and \U$25624 ( \26002 , \25353 , \21697 );
and \U$25625 ( \26003 , \25348 , \21695 );
nor \U$25626 ( \26004 , \26002 , \26003 );
xnor \U$25627 ( \26005 , \26004 , \21678 );
and \U$25628 ( \26006 , \26001 , \26005 );
and \U$25629 ( \26007 , \25806 , \21660 );
and \U$25630 ( \26008 , \25609 , \21658 );
nor \U$25631 ( \26009 , \26007 , \26008 );
xnor \U$25632 ( \26010 , \26009 , \21665 );
and \U$25633 ( \26011 , \26005 , \26010 );
and \U$25634 ( \26012 , \26001 , \26010 );
or \U$25635 ( \26013 , \26006 , \26011 , \26012 );
xor \U$25636 ( \26014 , \25800 , \25804 );
xor \U$25637 ( \26015 , \26014 , \25807 );
or \U$25638 ( \26016 , \26013 , \26015 );
and \U$25639 ( \26017 , \25996 , \26016 );
and \U$25640 ( \26018 , \25944 , \26016 );
or \U$25641 ( \26019 , \25997 , \26017 , \26018 );
xor \U$25642 ( \26020 , \25747 , \25751 );
xor \U$25643 ( \26021 , \26020 , \25756 );
xor \U$25644 ( \26022 , \25763 , \25767 );
xor \U$25645 ( \26023 , \26022 , \25772 );
and \U$25646 ( \26024 , \26021 , \26023 );
xor \U$25647 ( \26025 , \25780 , \25784 );
xor \U$25648 ( \26026 , \26025 , \25789 );
and \U$25649 ( \26027 , \26023 , \26026 );
and \U$25650 ( \26028 , \26021 , \26026 );
or \U$25651 ( \26029 , \26024 , \26027 , \26028 );
xor \U$25652 ( \26030 , \25695 , \25699 );
xor \U$25653 ( \26031 , \26030 , \25704 );
xor \U$25654 ( \26032 , \25711 , \25715 );
xor \U$25655 ( \26033 , \26032 , \25720 );
and \U$25656 ( \26034 , \26031 , \26033 );
xor \U$25657 ( \26035 , \25728 , \25732 );
xor \U$25658 ( \26036 , \26035 , \25737 );
and \U$25659 ( \26037 , \26033 , \26036 );
and \U$25660 ( \26038 , \26031 , \26036 );
or \U$25661 ( \26039 , \26034 , \26037 , \26038 );
and \U$25662 ( \26040 , \26029 , \26039 );
xor \U$25663 ( \26041 , \25566 , \25570 );
xor \U$25664 ( \26042 , \26041 , \25575 );
and \U$25665 ( \26043 , \26039 , \26042 );
and \U$25666 ( \26044 , \26029 , \26042 );
or \U$25667 ( \26045 , \26040 , \26043 , \26044 );
and \U$25668 ( \26046 , \26019 , \26045 );
xor \U$25669 ( \26047 , \25550 , \25554 );
xor \U$25670 ( \26048 , \26047 , \25559 );
xor \U$25671 ( \26049 , \25834 , \25836 );
xor \U$25672 ( \26050 , \26049 , \25839 );
and \U$25673 ( \26051 , \26048 , \26050 );
xor \U$25674 ( \26052 , \25810 , \25812 );
xor \U$25675 ( \26053 , \26052 , \25815 );
and \U$25676 ( \26054 , \26050 , \26053 );
and \U$25677 ( \26055 , \26048 , \26053 );
or \U$25678 ( \26056 , \26051 , \26054 , \26055 );
and \U$25679 ( \26057 , \26045 , \26056 );
and \U$25680 ( \26058 , \26019 , \26056 );
or \U$25681 ( \26059 , \26046 , \26057 , \26058 );
xor \U$25682 ( \26060 , \25743 , \25795 );
xor \U$25683 ( \26061 , \26060 , \25818 );
xor \U$25684 ( \26062 , \25823 , \25825 );
xor \U$25685 ( \26063 , \26062 , \25828 );
and \U$25686 ( \26064 , \26061 , \26063 );
xor \U$25687 ( \26065 , \25842 , \25844 );
xor \U$25688 ( \26066 , \26065 , \25846 );
and \U$25689 ( \26067 , \26063 , \26066 );
and \U$25690 ( \26068 , \26061 , \26066 );
or \U$25691 ( \26069 , \26064 , \26067 , \26068 );
and \U$25692 ( \26070 , \26059 , \26069 );
xor \U$25693 ( \26071 , \25544 , \25598 );
xor \U$25694 ( \26072 , \26071 , \25620 );
and \U$25695 ( \26073 , \26069 , \26072 );
and \U$25696 ( \26074 , \26059 , \26072 );
or \U$25697 ( \26075 , \26070 , \26073 , \26074 );
xor \U$25698 ( \26076 , \25821 , \25831 );
xor \U$25699 ( \26077 , \26076 , \25849 );
xor \U$25700 ( \26078 , \25854 , \25856 );
xor \U$25701 ( \26079 , \26078 , \25859 );
and \U$25702 ( \26080 , \26077 , \26079 );
and \U$25703 ( \26081 , \26075 , \26080 );
xor \U$25704 ( \26082 , \25870 , \25872 );
xor \U$25705 ( \26083 , \26082 , \25875 );
and \U$25706 ( \26084 , \26080 , \26083 );
and \U$25707 ( \26085 , \26075 , \26083 );
or \U$25708 ( \26086 , \26081 , \26084 , \26085 );
xor \U$25709 ( \26087 , \25868 , \25878 );
xor \U$25710 ( \26088 , \26087 , \25881 );
and \U$25711 ( \26089 , \26086 , \26088 );
xor \U$25712 ( \26090 , \25658 , \25668 );
xor \U$25713 ( \26091 , \26090 , \25671 );
and \U$25714 ( \26092 , \26088 , \26091 );
and \U$25715 ( \26093 , \26086 , \26091 );
or \U$25716 ( \26094 , \26089 , \26092 , \26093 );
and \U$25717 ( \26095 , \25890 , \26094 );
xor \U$25718 ( \26096 , \25890 , \26094 );
xor \U$25719 ( \26097 , \26086 , \26088 );
xor \U$25720 ( \26098 , \26097 , \26091 );
and \U$25721 ( \26099 , \25348 , \21745 );
and \U$25722 ( \26100 , \25226 , \21743 );
nor \U$25723 ( \26101 , \26099 , \26100 );
xnor \U$25724 ( \26102 , \26101 , \21715 );
and \U$25725 ( \26103 , \25609 , \21697 );
and \U$25726 ( \26104 , \25353 , \21695 );
nor \U$25727 ( \26105 , \26103 , \26104 );
xnor \U$25728 ( \26106 , \26105 , \21678 );
and \U$25729 ( \26107 , \26102 , \26106 );
buf \U$25730 ( \26108 , RIc22a850_169);
and \U$25731 ( \26109 , \26108 , \21660 );
and \U$25732 ( \26110 , \25806 , \21658 );
nor \U$25733 ( \26111 , \26109 , \26110 );
xnor \U$25734 ( \26112 , \26111 , \21665 );
and \U$25735 ( \26113 , \26106 , \26112 );
and \U$25736 ( \26114 , \26102 , \26112 );
or \U$25737 ( \26115 , \26107 , \26113 , \26114 );
buf \U$25738 ( \26116 , RIc22a8c8_170);
and \U$25739 ( \26117 , \26116 , \21654 );
buf \U$25740 ( \26118 , \26117 );
and \U$25741 ( \26119 , \26115 , \26118 );
and \U$25742 ( \26120 , \26108 , \21654 );
and \U$25743 ( \26121 , \26118 , \26120 );
and \U$25744 ( \26122 , \26115 , \26120 );
or \U$25745 ( \26123 , \26119 , \26121 , \26122 );
and \U$25746 ( \26124 , \22126 , \23933 );
and \U$25747 ( \26125 , \22046 , \23931 );
nor \U$25748 ( \26126 , \26124 , \26125 );
xnor \U$25749 ( \26127 , \26126 , \23791 );
and \U$25750 ( \26128 , \22262 , \23637 );
and \U$25751 ( \26129 , \22200 , \23635 );
nor \U$25752 ( \26130 , \26128 , \26129 );
xnor \U$25753 ( \26131 , \26130 , \23500 );
and \U$25754 ( \26132 , \26127 , \26131 );
and \U$25755 ( \26133 , \22523 , \23431 );
and \U$25756 ( \26134 , \22325 , \23429 );
nor \U$25757 ( \26135 , \26133 , \26134 );
xnor \U$25758 ( \26136 , \26135 , \23279 );
and \U$25759 ( \26137 , \26131 , \26136 );
and \U$25760 ( \26138 , \26127 , \26136 );
or \U$25761 ( \26139 , \26132 , \26137 , \26138 );
xor \U$25762 ( \26140 , \25546 , \25907 );
xor \U$25763 ( \26141 , \25907 , \25908 );
not \U$25764 ( \26142 , \26141 );
and \U$25765 ( \26143 , \26140 , \26142 );
and \U$25766 ( \26144 , \21653 , \26143 );
not \U$25767 ( \26145 , \26144 );
xnor \U$25768 ( \26146 , \26145 , \25911 );
and \U$25769 ( \26147 , \21685 , \25692 );
and \U$25770 ( \26148 , \21667 , \25690 );
nor \U$25771 ( \26149 , \26147 , \26148 );
xnor \U$25772 ( \26150 , \26149 , \25549 );
and \U$25773 ( \26151 , \26146 , \26150 );
and \U$25774 ( \26152 , \21754 , \25369 );
and \U$25775 ( \26153 , \21706 , \25367 );
nor \U$25776 ( \26154 , \26152 , \26153 );
xnor \U$25777 ( \26155 , \26154 , \25123 );
and \U$25778 ( \26156 , \26150 , \26155 );
and \U$25779 ( \26157 , \26146 , \26155 );
or \U$25780 ( \26158 , \26151 , \26156 , \26157 );
and \U$25781 ( \26159 , \26139 , \26158 );
and \U$25782 ( \26160 , \21831 , \24974 );
and \U$25783 ( \26161 , \21762 , \24972 );
nor \U$25784 ( \26162 , \26160 , \26161 );
xnor \U$25785 ( \26163 , \26162 , \24787 );
and \U$25786 ( \26164 , \21890 , \24661 );
and \U$25787 ( \26165 , \21836 , \24659 );
nor \U$25788 ( \26166 , \26164 , \26165 );
xnor \U$25789 ( \26167 , \26166 , \24456 );
and \U$25790 ( \26168 , \26163 , \26167 );
and \U$25791 ( \26169 , \22018 , \24255 );
and \U$25792 ( \26170 , \21941 , \24253 );
nor \U$25793 ( \26171 , \26169 , \26170 );
xnor \U$25794 ( \26172 , \26171 , \24106 );
and \U$25795 ( \26173 , \26167 , \26172 );
and \U$25796 ( \26174 , \26163 , \26172 );
or \U$25797 ( \26175 , \26168 , \26173 , \26174 );
and \U$25798 ( \26176 , \26158 , \26175 );
and \U$25799 ( \26177 , \26139 , \26175 );
or \U$25800 ( \26178 , \26159 , \26176 , \26177 );
and \U$25801 ( \26179 , \26123 , \26178 );
and \U$25802 ( \26180 , \24177 , \22029 );
and \U$25803 ( \26181 , \24003 , \22027 );
nor \U$25804 ( \26182 , \26180 , \26181 );
xnor \U$25805 ( \26183 , \26182 , \21986 );
and \U$25806 ( \26184 , \24482 , \21916 );
and \U$25807 ( \26185 , \24344 , \21914 );
nor \U$25808 ( \26186 , \26184 , \26185 );
xnor \U$25809 ( \26187 , \26186 , \21867 );
and \U$25810 ( \26188 , \26183 , \26187 );
and \U$25811 ( \26189 , \25018 , \21815 );
and \U$25812 ( \26190 , \24601 , \21813 );
nor \U$25813 ( \26191 , \26189 , \26190 );
xnor \U$25814 ( \26192 , \26191 , \21774 );
and \U$25815 ( \26193 , \26187 , \26192 );
and \U$25816 ( \26194 , \26183 , \26192 );
or \U$25817 ( \26195 , \26188 , \26193 , \26194 );
and \U$25818 ( \26196 , \23379 , \22497 );
and \U$25819 ( \26197 , \23136 , \22495 );
nor \U$25820 ( \26198 , \26196 , \26197 );
xnor \U$25821 ( \26199 , \26198 , \22419 );
and \U$25822 ( \26200 , \23570 , \22333 );
and \U$25823 ( \26201 , \23384 , \22331 );
nor \U$25824 ( \26202 , \26200 , \26201 );
xnor \U$25825 ( \26203 , \26202 , \22239 );
and \U$25826 ( \26204 , \26199 , \26203 );
and \U$25827 ( \26205 , \23978 , \22163 );
and \U$25828 ( \26206 , \23714 , \22161 );
nor \U$25829 ( \26207 , \26205 , \26206 );
xnor \U$25830 ( \26208 , \26207 , \22091 );
and \U$25831 ( \26209 , \26203 , \26208 );
and \U$25832 ( \26210 , \26199 , \26208 );
or \U$25833 ( \26211 , \26204 , \26209 , \26210 );
and \U$25834 ( \26212 , \26195 , \26211 );
and \U$25835 ( \26213 , \22716 , \23163 );
and \U$25836 ( \26214 , \22611 , \23161 );
nor \U$25837 ( \26215 , \26213 , \26214 );
xnor \U$25838 ( \26216 , \26215 , \23007 );
and \U$25839 ( \26217 , \22837 , \22891 );
and \U$25840 ( \26218 , \22721 , \22889 );
nor \U$25841 ( \26219 , \26217 , \26218 );
xnor \U$25842 ( \26220 , \26219 , \22778 );
and \U$25843 ( \26221 , \26216 , \26220 );
and \U$25844 ( \26222 , \23128 , \22697 );
and \U$25845 ( \26223 , \22952 , \22695 );
nor \U$25846 ( \26224 , \26222 , \26223 );
xnor \U$25847 ( \26225 , \26224 , \22561 );
and \U$25848 ( \26226 , \26220 , \26225 );
and \U$25849 ( \26227 , \26216 , \26225 );
or \U$25850 ( \26228 , \26221 , \26226 , \26227 );
and \U$25851 ( \26229 , \26211 , \26228 );
and \U$25852 ( \26230 , \26195 , \26228 );
or \U$25853 ( \26231 , \26212 , \26229 , \26230 );
and \U$25854 ( \26232 , \26178 , \26231 );
and \U$25855 ( \26233 , \26123 , \26231 );
or \U$25856 ( \26234 , \26179 , \26232 , \26233 );
xor \U$25857 ( \26235 , \25948 , \25952 );
xor \U$25858 ( \26236 , \26235 , \25957 );
xor \U$25859 ( \26237 , \25981 , \25985 );
xor \U$25860 ( \26238 , \26237 , \25990 );
and \U$25861 ( \26239 , \26236 , \26238 );
xor \U$25862 ( \26240 , \26001 , \26005 );
xor \U$25863 ( \26241 , \26240 , \26010 );
and \U$25864 ( \26242 , \26238 , \26241 );
and \U$25865 ( \26243 , \26236 , \26241 );
or \U$25866 ( \26244 , \26239 , \26242 , \26243 );
xor \U$25867 ( \26245 , \25894 , \25898 );
xor \U$25868 ( \26246 , \26245 , \25903 );
xor \U$25869 ( \26247 , \25964 , \25968 );
xor \U$25870 ( \26248 , \26247 , \25973 );
and \U$25871 ( \26249 , \26246 , \26248 );
xor \U$25872 ( \26250 , \25929 , \25933 );
xor \U$25873 ( \26251 , \26250 , \25938 );
and \U$25874 ( \26252 , \26248 , \26251 );
and \U$25875 ( \26253 , \26246 , \26251 );
or \U$25876 ( \26254 , \26249 , \26252 , \26253 );
and \U$25877 ( \26255 , \26244 , \26254 );
xor \U$25878 ( \26256 , \26031 , \26033 );
xor \U$25879 ( \26257 , \26256 , \26036 );
and \U$25880 ( \26258 , \26254 , \26257 );
and \U$25881 ( \26259 , \26244 , \26257 );
or \U$25882 ( \26260 , \26255 , \26258 , \26259 );
and \U$25883 ( \26261 , \26234 , \26260 );
xor \U$25884 ( \26262 , \25960 , \25976 );
xor \U$25885 ( \26263 , \26262 , \25993 );
xor \U$25886 ( \26264 , \26021 , \26023 );
xor \U$25887 ( \26265 , \26264 , \26026 );
and \U$25888 ( \26266 , \26263 , \26265 );
xnor \U$25889 ( \26267 , \26013 , \26015 );
and \U$25890 ( \26268 , \26265 , \26267 );
and \U$25891 ( \26269 , \26263 , \26267 );
or \U$25892 ( \26270 , \26266 , \26268 , \26269 );
and \U$25893 ( \26271 , \26260 , \26270 );
and \U$25894 ( \26272 , \26234 , \26270 );
or \U$25895 ( \26273 , \26261 , \26271 , \26272 );
xor \U$25896 ( \26274 , \25707 , \25723 );
xor \U$25897 ( \26275 , \26274 , \25740 );
xor \U$25898 ( \26276 , \25759 , \25775 );
xor \U$25899 ( \26277 , \26276 , \25792 );
and \U$25900 ( \26278 , \26275 , \26277 );
xor \U$25901 ( \26279 , \26048 , \26050 );
xor \U$25902 ( \26280 , \26279 , \26053 );
and \U$25903 ( \26281 , \26277 , \26280 );
and \U$25904 ( \26282 , \26275 , \26280 );
or \U$25905 ( \26283 , \26278 , \26281 , \26282 );
and \U$25906 ( \26284 , \26273 , \26283 );
xor \U$25907 ( \26285 , \26061 , \26063 );
xor \U$25908 ( \26286 , \26285 , \26066 );
and \U$25909 ( \26287 , \26283 , \26286 );
and \U$25910 ( \26288 , \26273 , \26286 );
or \U$25911 ( \26289 , \26284 , \26287 , \26288 );
xor \U$25912 ( \26290 , \26059 , \26069 );
xor \U$25913 ( \26291 , \26290 , \26072 );
and \U$25914 ( \26292 , \26289 , \26291 );
xor \U$25915 ( \26293 , \26077 , \26079 );
and \U$25916 ( \26294 , \26291 , \26293 );
and \U$25917 ( \26295 , \26289 , \26293 );
or \U$25918 ( \26296 , \26292 , \26294 , \26295 );
xor \U$25919 ( \26297 , \25852 , \25862 );
xor \U$25920 ( \26298 , \26297 , \25865 );
and \U$25921 ( \26299 , \26296 , \26298 );
xor \U$25922 ( \26300 , \26075 , \26080 );
xor \U$25923 ( \26301 , \26300 , \26083 );
and \U$25924 ( \26302 , \26298 , \26301 );
and \U$25925 ( \26303 , \26296 , \26301 );
or \U$25926 ( \26304 , \26299 , \26302 , \26303 );
and \U$25927 ( \26305 , \26098 , \26304 );
xor \U$25928 ( \26306 , \26098 , \26304 );
xor \U$25929 ( \26307 , \26296 , \26298 );
xor \U$25930 ( \26308 , \26307 , \26301 );
and \U$25931 ( \26309 , \22046 , \24255 );
and \U$25932 ( \26310 , \22018 , \24253 );
nor \U$25933 ( \26311 , \26309 , \26310 );
xnor \U$25934 ( \26312 , \26311 , \24106 );
and \U$25935 ( \26313 , \22200 , \23933 );
and \U$25936 ( \26314 , \22126 , \23931 );
nor \U$25937 ( \26315 , \26313 , \26314 );
xnor \U$25938 ( \26316 , \26315 , \23791 );
and \U$25939 ( \26317 , \26312 , \26316 );
and \U$25940 ( \26318 , \22325 , \23637 );
and \U$25941 ( \26319 , \22262 , \23635 );
nor \U$25942 ( \26320 , \26318 , \26319 );
xnor \U$25943 ( \26321 , \26320 , \23500 );
and \U$25944 ( \26322 , \26316 , \26321 );
and \U$25945 ( \26323 , \26312 , \26321 );
or \U$25946 ( \26324 , \26317 , \26322 , \26323 );
buf \U$25947 ( \26325 , RIc226188_44);
buf \U$25948 ( \26326 , RIc226110_45);
and \U$25949 ( \26327 , \26325 , \26326 );
not \U$25950 ( \26328 , \26327 );
and \U$25951 ( \26329 , \25908 , \26328 );
not \U$25952 ( \26330 , \26329 );
and \U$25953 ( \26331 , \21667 , \26143 );
and \U$25954 ( \26332 , \21653 , \26141 );
nor \U$25955 ( \26333 , \26331 , \26332 );
xnor \U$25956 ( \26334 , \26333 , \25911 );
and \U$25957 ( \26335 , \26330 , \26334 );
and \U$25958 ( \26336 , \21706 , \25692 );
and \U$25959 ( \26337 , \21685 , \25690 );
nor \U$25960 ( \26338 , \26336 , \26337 );
xnor \U$25961 ( \26339 , \26338 , \25549 );
and \U$25962 ( \26340 , \26334 , \26339 );
and \U$25963 ( \26341 , \26330 , \26339 );
or \U$25964 ( \26342 , \26335 , \26340 , \26341 );
and \U$25965 ( \26343 , \26324 , \26342 );
and \U$25966 ( \26344 , \21762 , \25369 );
and \U$25967 ( \26345 , \21754 , \25367 );
nor \U$25968 ( \26346 , \26344 , \26345 );
xnor \U$25969 ( \26347 , \26346 , \25123 );
and \U$25970 ( \26348 , \21836 , \24974 );
and \U$25971 ( \26349 , \21831 , \24972 );
nor \U$25972 ( \26350 , \26348 , \26349 );
xnor \U$25973 ( \26351 , \26350 , \24787 );
and \U$25974 ( \26352 , \26347 , \26351 );
and \U$25975 ( \26353 , \21941 , \24661 );
and \U$25976 ( \26354 , \21890 , \24659 );
nor \U$25977 ( \26355 , \26353 , \26354 );
xnor \U$25978 ( \26356 , \26355 , \24456 );
and \U$25979 ( \26357 , \26351 , \26356 );
and \U$25980 ( \26358 , \26347 , \26356 );
or \U$25981 ( \26359 , \26352 , \26357 , \26358 );
and \U$25982 ( \26360 , \26342 , \26359 );
and \U$25983 ( \26361 , \26324 , \26359 );
or \U$25984 ( \26362 , \26343 , \26360 , \26361 );
and \U$25985 ( \26363 , \22611 , \23431 );
and \U$25986 ( \26364 , \22523 , \23429 );
nor \U$25987 ( \26365 , \26363 , \26364 );
xnor \U$25988 ( \26366 , \26365 , \23279 );
and \U$25989 ( \26367 , \22721 , \23163 );
and \U$25990 ( \26368 , \22716 , \23161 );
nor \U$25991 ( \26369 , \26367 , \26368 );
xnor \U$25992 ( \26370 , \26369 , \23007 );
and \U$25993 ( \26371 , \26366 , \26370 );
and \U$25994 ( \26372 , \22952 , \22891 );
and \U$25995 ( \26373 , \22837 , \22889 );
nor \U$25996 ( \26374 , \26372 , \26373 );
xnor \U$25997 ( \26375 , \26374 , \22778 );
and \U$25998 ( \26376 , \26370 , \26375 );
and \U$25999 ( \26377 , \26366 , \26375 );
or \U$26000 ( \26378 , \26371 , \26376 , \26377 );
and \U$26001 ( \26379 , \24003 , \22163 );
and \U$26002 ( \26380 , \23978 , \22161 );
nor \U$26003 ( \26381 , \26379 , \26380 );
xnor \U$26004 ( \26382 , \26381 , \22091 );
and \U$26005 ( \26383 , \24344 , \22029 );
and \U$26006 ( \26384 , \24177 , \22027 );
nor \U$26007 ( \26385 , \26383 , \26384 );
xnor \U$26008 ( \26386 , \26385 , \21986 );
and \U$26009 ( \26387 , \26382 , \26386 );
and \U$26010 ( \26388 , \24601 , \21916 );
and \U$26011 ( \26389 , \24482 , \21914 );
nor \U$26012 ( \26390 , \26388 , \26389 );
xnor \U$26013 ( \26391 , \26390 , \21867 );
and \U$26014 ( \26392 , \26386 , \26391 );
and \U$26015 ( \26393 , \26382 , \26391 );
or \U$26016 ( \26394 , \26387 , \26392 , \26393 );
and \U$26017 ( \26395 , \26378 , \26394 );
and \U$26018 ( \26396 , \23136 , \22697 );
and \U$26019 ( \26397 , \23128 , \22695 );
nor \U$26020 ( \26398 , \26396 , \26397 );
xnor \U$26021 ( \26399 , \26398 , \22561 );
and \U$26022 ( \26400 , \23384 , \22497 );
and \U$26023 ( \26401 , \23379 , \22495 );
nor \U$26024 ( \26402 , \26400 , \26401 );
xnor \U$26025 ( \26403 , \26402 , \22419 );
and \U$26026 ( \26404 , \26399 , \26403 );
and \U$26027 ( \26405 , \23714 , \22333 );
and \U$26028 ( \26406 , \23570 , \22331 );
nor \U$26029 ( \26407 , \26405 , \26406 );
xnor \U$26030 ( \26408 , \26407 , \22239 );
and \U$26031 ( \26409 , \26403 , \26408 );
and \U$26032 ( \26410 , \26399 , \26408 );
or \U$26033 ( \26411 , \26404 , \26409 , \26410 );
and \U$26034 ( \26412 , \26394 , \26411 );
and \U$26035 ( \26413 , \26378 , \26411 );
or \U$26036 ( \26414 , \26395 , \26412 , \26413 );
and \U$26037 ( \26415 , \26362 , \26414 );
and \U$26038 ( \26416 , \25226 , \21815 );
and \U$26039 ( \26417 , \25018 , \21813 );
nor \U$26040 ( \26418 , \26416 , \26417 );
xnor \U$26041 ( \26419 , \26418 , \21774 );
and \U$26042 ( \26420 , \25353 , \21745 );
and \U$26043 ( \26421 , \25348 , \21743 );
nor \U$26044 ( \26422 , \26420 , \26421 );
xnor \U$26045 ( \26423 , \26422 , \21715 );
and \U$26046 ( \26424 , \26419 , \26423 );
and \U$26047 ( \26425 , \25806 , \21697 );
and \U$26048 ( \26426 , \25609 , \21695 );
nor \U$26049 ( \26427 , \26425 , \26426 );
xnor \U$26050 ( \26428 , \26427 , \21678 );
and \U$26051 ( \26429 , \26423 , \26428 );
and \U$26052 ( \26430 , \26419 , \26428 );
or \U$26053 ( \26431 , \26424 , \26429 , \26430 );
xor \U$26054 ( \26432 , \26102 , \26106 );
xor \U$26055 ( \26433 , \26432 , \26112 );
and \U$26056 ( \26434 , \26431 , \26433 );
not \U$26057 ( \26435 , \26117 );
and \U$26058 ( \26436 , \26433 , \26435 );
and \U$26059 ( \26437 , \26431 , \26435 );
or \U$26060 ( \26438 , \26434 , \26436 , \26437 );
and \U$26061 ( \26439 , \26414 , \26438 );
and \U$26062 ( \26440 , \26362 , \26438 );
or \U$26063 ( \26441 , \26415 , \26439 , \26440 );
xor \U$26064 ( \26442 , \26183 , \26187 );
xor \U$26065 ( \26443 , \26442 , \26192 );
xor \U$26066 ( \26444 , \26199 , \26203 );
xor \U$26067 ( \26445 , \26444 , \26208 );
and \U$26068 ( \26446 , \26443 , \26445 );
xor \U$26069 ( \26447 , \26216 , \26220 );
xor \U$26070 ( \26448 , \26447 , \26225 );
and \U$26071 ( \26449 , \26445 , \26448 );
and \U$26072 ( \26450 , \26443 , \26448 );
or \U$26073 ( \26451 , \26446 , \26449 , \26450 );
xor \U$26074 ( \26452 , \26127 , \26131 );
xor \U$26075 ( \26453 , \26452 , \26136 );
xor \U$26076 ( \26454 , \26146 , \26150 );
xor \U$26077 ( \26455 , \26454 , \26155 );
and \U$26078 ( \26456 , \26453 , \26455 );
xor \U$26079 ( \26457 , \26163 , \26167 );
xor \U$26080 ( \26458 , \26457 , \26172 );
and \U$26081 ( \26459 , \26455 , \26458 );
and \U$26082 ( \26460 , \26453 , \26458 );
or \U$26083 ( \26461 , \26456 , \26459 , \26460 );
and \U$26084 ( \26462 , \26451 , \26461 );
xor \U$26085 ( \26463 , \25912 , \25916 );
xor \U$26086 ( \26464 , \26463 , \25921 );
and \U$26087 ( \26465 , \26461 , \26464 );
and \U$26088 ( \26466 , \26451 , \26464 );
or \U$26089 ( \26467 , \26462 , \26465 , \26466 );
and \U$26090 ( \26468 , \26441 , \26467 );
xor \U$26091 ( \26469 , \26115 , \26118 );
xor \U$26092 ( \26470 , \26469 , \26120 );
xor \U$26093 ( \26471 , \26236 , \26238 );
xor \U$26094 ( \26472 , \26471 , \26241 );
and \U$26095 ( \26473 , \26470 , \26472 );
xor \U$26096 ( \26474 , \26246 , \26248 );
xor \U$26097 ( \26475 , \26474 , \26251 );
and \U$26098 ( \26476 , \26472 , \26475 );
and \U$26099 ( \26477 , \26470 , \26475 );
or \U$26100 ( \26478 , \26473 , \26476 , \26477 );
and \U$26101 ( \26479 , \26467 , \26478 );
and \U$26102 ( \26480 , \26441 , \26478 );
or \U$26103 ( \26481 , \26468 , \26479 , \26480 );
xor \U$26104 ( \26482 , \25906 , \25924 );
xor \U$26105 ( \26483 , \26482 , \25941 );
xor \U$26106 ( \26484 , \26244 , \26254 );
xor \U$26107 ( \26485 , \26484 , \26257 );
and \U$26108 ( \26486 , \26483 , \26485 );
xor \U$26109 ( \26487 , \26263 , \26265 );
xor \U$26110 ( \26488 , \26487 , \26267 );
and \U$26111 ( \26489 , \26485 , \26488 );
and \U$26112 ( \26490 , \26483 , \26488 );
or \U$26113 ( \26491 , \26486 , \26489 , \26490 );
and \U$26114 ( \26492 , \26481 , \26491 );
xor \U$26115 ( \26493 , \26029 , \26039 );
xor \U$26116 ( \26494 , \26493 , \26042 );
and \U$26117 ( \26495 , \26491 , \26494 );
and \U$26118 ( \26496 , \26481 , \26494 );
or \U$26119 ( \26497 , \26492 , \26495 , \26496 );
xor \U$26120 ( \26498 , \25944 , \25996 );
xor \U$26121 ( \26499 , \26498 , \26016 );
xor \U$26122 ( \26500 , \26234 , \26260 );
xor \U$26123 ( \26501 , \26500 , \26270 );
and \U$26124 ( \26502 , \26499 , \26501 );
xor \U$26125 ( \26503 , \26275 , \26277 );
xor \U$26126 ( \26504 , \26503 , \26280 );
and \U$26127 ( \26505 , \26501 , \26504 );
and \U$26128 ( \26506 , \26499 , \26504 );
or \U$26129 ( \26507 , \26502 , \26505 , \26506 );
and \U$26130 ( \26508 , \26497 , \26507 );
xor \U$26131 ( \26509 , \26019 , \26045 );
xor \U$26132 ( \26510 , \26509 , \26056 );
and \U$26133 ( \26511 , \26507 , \26510 );
and \U$26134 ( \26512 , \26497 , \26510 );
or \U$26135 ( \26513 , \26508 , \26511 , \26512 );
xor \U$26136 ( \26514 , \25908 , \26325 );
xor \U$26137 ( \26515 , \26325 , \26326 );
not \U$26138 ( \26516 , \26515 );
and \U$26139 ( \26517 , \26514 , \26516 );
and \U$26140 ( \26518 , \21653 , \26517 );
not \U$26141 ( \26519 , \26518 );
xnor \U$26142 ( \26520 , \26519 , \26329 );
and \U$26143 ( \26521 , \21685 , \26143 );
and \U$26144 ( \26522 , \21667 , \26141 );
nor \U$26145 ( \26523 , \26521 , \26522 );
xnor \U$26146 ( \26524 , \26523 , \25911 );
and \U$26147 ( \26525 , \26520 , \26524 );
and \U$26148 ( \26526 , \21754 , \25692 );
and \U$26149 ( \26527 , \21706 , \25690 );
nor \U$26150 ( \26528 , \26526 , \26527 );
xnor \U$26151 ( \26529 , \26528 , \25549 );
and \U$26152 ( \26530 , \26524 , \26529 );
and \U$26153 ( \26531 , \26520 , \26529 );
or \U$26154 ( \26532 , \26525 , \26530 , \26531 );
and \U$26155 ( \26533 , \22126 , \24255 );
and \U$26156 ( \26534 , \22046 , \24253 );
nor \U$26157 ( \26535 , \26533 , \26534 );
xnor \U$26158 ( \26536 , \26535 , \24106 );
and \U$26159 ( \26537 , \22262 , \23933 );
and \U$26160 ( \26538 , \22200 , \23931 );
nor \U$26161 ( \26539 , \26537 , \26538 );
xnor \U$26162 ( \26540 , \26539 , \23791 );
and \U$26163 ( \26541 , \26536 , \26540 );
and \U$26164 ( \26542 , \22523 , \23637 );
and \U$26165 ( \26543 , \22325 , \23635 );
nor \U$26166 ( \26544 , \26542 , \26543 );
xnor \U$26167 ( \26545 , \26544 , \23500 );
and \U$26168 ( \26546 , \26540 , \26545 );
and \U$26169 ( \26547 , \26536 , \26545 );
or \U$26170 ( \26548 , \26541 , \26546 , \26547 );
and \U$26171 ( \26549 , \26532 , \26548 );
and \U$26172 ( \26550 , \21831 , \25369 );
and \U$26173 ( \26551 , \21762 , \25367 );
nor \U$26174 ( \26552 , \26550 , \26551 );
xnor \U$26175 ( \26553 , \26552 , \25123 );
and \U$26176 ( \26554 , \21890 , \24974 );
and \U$26177 ( \26555 , \21836 , \24972 );
nor \U$26178 ( \26556 , \26554 , \26555 );
xnor \U$26179 ( \26557 , \26556 , \24787 );
and \U$26180 ( \26558 , \26553 , \26557 );
and \U$26181 ( \26559 , \22018 , \24661 );
and \U$26182 ( \26560 , \21941 , \24659 );
nor \U$26183 ( \26561 , \26559 , \26560 );
xnor \U$26184 ( \26562 , \26561 , \24456 );
and \U$26185 ( \26563 , \26557 , \26562 );
and \U$26186 ( \26564 , \26553 , \26562 );
or \U$26187 ( \26565 , \26558 , \26563 , \26564 );
and \U$26188 ( \26566 , \26548 , \26565 );
and \U$26189 ( \26567 , \26532 , \26565 );
or \U$26190 ( \26568 , \26549 , \26566 , \26567 );
and \U$26191 ( \26569 , \25348 , \21815 );
and \U$26192 ( \26570 , \25226 , \21813 );
nor \U$26193 ( \26571 , \26569 , \26570 );
xnor \U$26194 ( \26572 , \26571 , \21774 );
and \U$26195 ( \26573 , \25609 , \21745 );
and \U$26196 ( \26574 , \25353 , \21743 );
nor \U$26197 ( \26575 , \26573 , \26574 );
xnor \U$26198 ( \26576 , \26575 , \21715 );
and \U$26199 ( \26577 , \26572 , \26576 );
and \U$26200 ( \26578 , \26108 , \21697 );
and \U$26201 ( \26579 , \25806 , \21695 );
nor \U$26202 ( \26580 , \26578 , \26579 );
xnor \U$26203 ( \26581 , \26580 , \21678 );
and \U$26204 ( \26582 , \26576 , \26581 );
and \U$26205 ( \26583 , \26572 , \26581 );
or \U$26206 ( \26584 , \26577 , \26582 , \26583 );
buf \U$26207 ( \26585 , RIc22a940_171);
and \U$26208 ( \26586 , \26585 , \21660 );
and \U$26209 ( \26587 , \26116 , \21658 );
nor \U$26210 ( \26588 , \26586 , \26587 );
xnor \U$26211 ( \26589 , \26588 , \21665 );
buf \U$26212 ( \26590 , RIc22a9b8_172);
and \U$26213 ( \26591 , \26590 , \21654 );
or \U$26214 ( \26592 , \26589 , \26591 );
and \U$26215 ( \26593 , \26584 , \26592 );
and \U$26216 ( \26594 , \26116 , \21660 );
and \U$26217 ( \26595 , \26108 , \21658 );
nor \U$26218 ( \26596 , \26594 , \26595 );
xnor \U$26219 ( \26597 , \26596 , \21665 );
and \U$26220 ( \26598 , \26592 , \26597 );
and \U$26221 ( \26599 , \26584 , \26597 );
or \U$26222 ( \26600 , \26593 , \26598 , \26599 );
and \U$26223 ( \26601 , \26568 , \26600 );
and \U$26224 ( \26602 , \22716 , \23431 );
and \U$26225 ( \26603 , \22611 , \23429 );
nor \U$26226 ( \26604 , \26602 , \26603 );
xnor \U$26227 ( \26605 , \26604 , \23279 );
and \U$26228 ( \26606 , \22837 , \23163 );
and \U$26229 ( \26607 , \22721 , \23161 );
nor \U$26230 ( \26608 , \26606 , \26607 );
xnor \U$26231 ( \26609 , \26608 , \23007 );
and \U$26232 ( \26610 , \26605 , \26609 );
and \U$26233 ( \26611 , \23128 , \22891 );
and \U$26234 ( \26612 , \22952 , \22889 );
nor \U$26235 ( \26613 , \26611 , \26612 );
xnor \U$26236 ( \26614 , \26613 , \22778 );
and \U$26237 ( \26615 , \26609 , \26614 );
and \U$26238 ( \26616 , \26605 , \26614 );
or \U$26239 ( \26617 , \26610 , \26615 , \26616 );
and \U$26240 ( \26618 , \23379 , \22697 );
and \U$26241 ( \26619 , \23136 , \22695 );
nor \U$26242 ( \26620 , \26618 , \26619 );
xnor \U$26243 ( \26621 , \26620 , \22561 );
and \U$26244 ( \26622 , \23570 , \22497 );
and \U$26245 ( \26623 , \23384 , \22495 );
nor \U$26246 ( \26624 , \26622 , \26623 );
xnor \U$26247 ( \26625 , \26624 , \22419 );
and \U$26248 ( \26626 , \26621 , \26625 );
and \U$26249 ( \26627 , \23978 , \22333 );
and \U$26250 ( \26628 , \23714 , \22331 );
nor \U$26251 ( \26629 , \26627 , \26628 );
xnor \U$26252 ( \26630 , \26629 , \22239 );
and \U$26253 ( \26631 , \26625 , \26630 );
and \U$26254 ( \26632 , \26621 , \26630 );
or \U$26255 ( \26633 , \26626 , \26631 , \26632 );
and \U$26256 ( \26634 , \26617 , \26633 );
and \U$26257 ( \26635 , \24177 , \22163 );
and \U$26258 ( \26636 , \24003 , \22161 );
nor \U$26259 ( \26637 , \26635 , \26636 );
xnor \U$26260 ( \26638 , \26637 , \22091 );
and \U$26261 ( \26639 , \24482 , \22029 );
and \U$26262 ( \26640 , \24344 , \22027 );
nor \U$26263 ( \26641 , \26639 , \26640 );
xnor \U$26264 ( \26642 , \26641 , \21986 );
and \U$26265 ( \26643 , \26638 , \26642 );
and \U$26266 ( \26644 , \25018 , \21916 );
and \U$26267 ( \26645 , \24601 , \21914 );
nor \U$26268 ( \26646 , \26644 , \26645 );
xnor \U$26269 ( \26647 , \26646 , \21867 );
and \U$26270 ( \26648 , \26642 , \26647 );
and \U$26271 ( \26649 , \26638 , \26647 );
or \U$26272 ( \26650 , \26643 , \26648 , \26649 );
and \U$26273 ( \26651 , \26633 , \26650 );
and \U$26274 ( \26652 , \26617 , \26650 );
or \U$26275 ( \26653 , \26634 , \26651 , \26652 );
and \U$26276 ( \26654 , \26600 , \26653 );
and \U$26277 ( \26655 , \26568 , \26653 );
or \U$26278 ( \26656 , \26601 , \26654 , \26655 );
and \U$26279 ( \26657 , \26585 , \21654 );
xor \U$26280 ( \26658 , \26419 , \26423 );
xor \U$26281 ( \26659 , \26658 , \26428 );
and \U$26282 ( \26660 , \26657 , \26659 );
xor \U$26283 ( \26661 , \26382 , \26386 );
xor \U$26284 ( \26662 , \26661 , \26391 );
and \U$26285 ( \26663 , \26659 , \26662 );
and \U$26286 ( \26664 , \26657 , \26662 );
or \U$26287 ( \26665 , \26660 , \26663 , \26664 );
xor \U$26288 ( \26666 , \26366 , \26370 );
xor \U$26289 ( \26667 , \26666 , \26375 );
xor \U$26290 ( \26668 , \26312 , \26316 );
xor \U$26291 ( \26669 , \26668 , \26321 );
and \U$26292 ( \26670 , \26667 , \26669 );
xor \U$26293 ( \26671 , \26399 , \26403 );
xor \U$26294 ( \26672 , \26671 , \26408 );
and \U$26295 ( \26673 , \26669 , \26672 );
and \U$26296 ( \26674 , \26667 , \26672 );
or \U$26297 ( \26675 , \26670 , \26673 , \26674 );
and \U$26298 ( \26676 , \26665 , \26675 );
xor \U$26299 ( \26677 , \26453 , \26455 );
xor \U$26300 ( \26678 , \26677 , \26458 );
and \U$26301 ( \26679 , \26675 , \26678 );
and \U$26302 ( \26680 , \26665 , \26678 );
or \U$26303 ( \26681 , \26676 , \26679 , \26680 );
and \U$26304 ( \26682 , \26656 , \26681 );
xor \U$26305 ( \26683 , \26378 , \26394 );
xor \U$26306 ( \26684 , \26683 , \26411 );
xor \U$26307 ( \26685 , \26443 , \26445 );
xor \U$26308 ( \26686 , \26685 , \26448 );
and \U$26309 ( \26687 , \26684 , \26686 );
xor \U$26310 ( \26688 , \26431 , \26433 );
xor \U$26311 ( \26689 , \26688 , \26435 );
and \U$26312 ( \26690 , \26686 , \26689 );
and \U$26313 ( \26691 , \26684 , \26689 );
or \U$26314 ( \26692 , \26687 , \26690 , \26691 );
and \U$26315 ( \26693 , \26681 , \26692 );
and \U$26316 ( \26694 , \26656 , \26692 );
or \U$26317 ( \26695 , \26682 , \26693 , \26694 );
xor \U$26318 ( \26696 , \26139 , \26158 );
xor \U$26319 ( \26697 , \26696 , \26175 );
xor \U$26320 ( \26698 , \26195 , \26211 );
xor \U$26321 ( \26699 , \26698 , \26228 );
and \U$26322 ( \26700 , \26697 , \26699 );
xor \U$26323 ( \26701 , \26470 , \26472 );
xor \U$26324 ( \26702 , \26701 , \26475 );
and \U$26325 ( \26703 , \26699 , \26702 );
and \U$26326 ( \26704 , \26697 , \26702 );
or \U$26327 ( \26705 , \26700 , \26703 , \26704 );
and \U$26328 ( \26706 , \26695 , \26705 );
xor \U$26329 ( \26707 , \26123 , \26178 );
xor \U$26330 ( \26708 , \26707 , \26231 );
and \U$26331 ( \26709 , \26705 , \26708 );
and \U$26332 ( \26710 , \26695 , \26708 );
or \U$26333 ( \26711 , \26706 , \26709 , \26710 );
xor \U$26334 ( \26712 , \26481 , \26491 );
xor \U$26335 ( \26713 , \26712 , \26494 );
and \U$26336 ( \26714 , \26711 , \26713 );
xor \U$26337 ( \26715 , \26499 , \26501 );
xor \U$26338 ( \26716 , \26715 , \26504 );
and \U$26339 ( \26717 , \26713 , \26716 );
and \U$26340 ( \26718 , \26711 , \26716 );
or \U$26341 ( \26719 , \26714 , \26717 , \26718 );
xor \U$26342 ( \26720 , \26497 , \26507 );
xor \U$26343 ( \26721 , \26720 , \26510 );
and \U$26344 ( \26722 , \26719 , \26721 );
xor \U$26345 ( \26723 , \26273 , \26283 );
xor \U$26346 ( \26724 , \26723 , \26286 );
and \U$26347 ( \26725 , \26721 , \26724 );
and \U$26348 ( \26726 , \26719 , \26724 );
or \U$26349 ( \26727 , \26722 , \26725 , \26726 );
and \U$26350 ( \26728 , \26513 , \26727 );
xor \U$26351 ( \26729 , \26289 , \26291 );
xor \U$26352 ( \26730 , \26729 , \26293 );
and \U$26353 ( \26731 , \26727 , \26730 );
and \U$26354 ( \26732 , \26513 , \26730 );
or \U$26355 ( \26733 , \26728 , \26731 , \26732 );
and \U$26356 ( \26734 , \26308 , \26733 );
xor \U$26357 ( \26735 , \26308 , \26733 );
xor \U$26358 ( \26736 , \26513 , \26727 );
xor \U$26359 ( \26737 , \26736 , \26730 );
buf \U$26360 ( \26738 , RIc226098_46);
buf \U$26361 ( \26739 , RIc226020_47);
and \U$26362 ( \26740 , \26738 , \26739 );
not \U$26363 ( \26741 , \26740 );
and \U$26364 ( \26742 , \26326 , \26741 );
not \U$26365 ( \26743 , \26742 );
and \U$26366 ( \26744 , \21667 , \26517 );
and \U$26367 ( \26745 , \21653 , \26515 );
nor \U$26368 ( \26746 , \26744 , \26745 );
xnor \U$26369 ( \26747 , \26746 , \26329 );
and \U$26370 ( \26748 , \26743 , \26747 );
and \U$26371 ( \26749 , \21706 , \26143 );
and \U$26372 ( \26750 , \21685 , \26141 );
nor \U$26373 ( \26751 , \26749 , \26750 );
xnor \U$26374 ( \26752 , \26751 , \25911 );
and \U$26375 ( \26753 , \26747 , \26752 );
and \U$26376 ( \26754 , \26743 , \26752 );
or \U$26377 ( \26755 , \26748 , \26753 , \26754 );
and \U$26378 ( \26756 , \21762 , \25692 );
and \U$26379 ( \26757 , \21754 , \25690 );
nor \U$26380 ( \26758 , \26756 , \26757 );
xnor \U$26381 ( \26759 , \26758 , \25549 );
and \U$26382 ( \26760 , \21836 , \25369 );
and \U$26383 ( \26761 , \21831 , \25367 );
nor \U$26384 ( \26762 , \26760 , \26761 );
xnor \U$26385 ( \26763 , \26762 , \25123 );
and \U$26386 ( \26764 , \26759 , \26763 );
and \U$26387 ( \26765 , \21941 , \24974 );
and \U$26388 ( \26766 , \21890 , \24972 );
nor \U$26389 ( \26767 , \26765 , \26766 );
xnor \U$26390 ( \26768 , \26767 , \24787 );
and \U$26391 ( \26769 , \26763 , \26768 );
and \U$26392 ( \26770 , \26759 , \26768 );
or \U$26393 ( \26771 , \26764 , \26769 , \26770 );
and \U$26394 ( \26772 , \26755 , \26771 );
and \U$26395 ( \26773 , \22046 , \24661 );
and \U$26396 ( \26774 , \22018 , \24659 );
nor \U$26397 ( \26775 , \26773 , \26774 );
xnor \U$26398 ( \26776 , \26775 , \24456 );
and \U$26399 ( \26777 , \22200 , \24255 );
and \U$26400 ( \26778 , \22126 , \24253 );
nor \U$26401 ( \26779 , \26777 , \26778 );
xnor \U$26402 ( \26780 , \26779 , \24106 );
and \U$26403 ( \26781 , \26776 , \26780 );
and \U$26404 ( \26782 , \22325 , \23933 );
and \U$26405 ( \26783 , \22262 , \23931 );
nor \U$26406 ( \26784 , \26782 , \26783 );
xnor \U$26407 ( \26785 , \26784 , \23791 );
and \U$26408 ( \26786 , \26780 , \26785 );
and \U$26409 ( \26787 , \26776 , \26785 );
or \U$26410 ( \26788 , \26781 , \26786 , \26787 );
and \U$26411 ( \26789 , \26771 , \26788 );
and \U$26412 ( \26790 , \26755 , \26788 );
or \U$26413 ( \26791 , \26772 , \26789 , \26790 );
and \U$26414 ( \26792 , \22611 , \23637 );
and \U$26415 ( \26793 , \22523 , \23635 );
nor \U$26416 ( \26794 , \26792 , \26793 );
xnor \U$26417 ( \26795 , \26794 , \23500 );
and \U$26418 ( \26796 , \22721 , \23431 );
and \U$26419 ( \26797 , \22716 , \23429 );
nor \U$26420 ( \26798 , \26796 , \26797 );
xnor \U$26421 ( \26799 , \26798 , \23279 );
and \U$26422 ( \26800 , \26795 , \26799 );
and \U$26423 ( \26801 , \22952 , \23163 );
and \U$26424 ( \26802 , \22837 , \23161 );
nor \U$26425 ( \26803 , \26801 , \26802 );
xnor \U$26426 ( \26804 , \26803 , \23007 );
and \U$26427 ( \26805 , \26799 , \26804 );
and \U$26428 ( \26806 , \26795 , \26804 );
or \U$26429 ( \26807 , \26800 , \26805 , \26806 );
and \U$26430 ( \26808 , \23136 , \22891 );
and \U$26431 ( \26809 , \23128 , \22889 );
nor \U$26432 ( \26810 , \26808 , \26809 );
xnor \U$26433 ( \26811 , \26810 , \22778 );
and \U$26434 ( \26812 , \23384 , \22697 );
and \U$26435 ( \26813 , \23379 , \22695 );
nor \U$26436 ( \26814 , \26812 , \26813 );
xnor \U$26437 ( \26815 , \26814 , \22561 );
and \U$26438 ( \26816 , \26811 , \26815 );
and \U$26439 ( \26817 , \23714 , \22497 );
and \U$26440 ( \26818 , \23570 , \22495 );
nor \U$26441 ( \26819 , \26817 , \26818 );
xnor \U$26442 ( \26820 , \26819 , \22419 );
and \U$26443 ( \26821 , \26815 , \26820 );
and \U$26444 ( \26822 , \26811 , \26820 );
or \U$26445 ( \26823 , \26816 , \26821 , \26822 );
and \U$26446 ( \26824 , \26807 , \26823 );
and \U$26447 ( \26825 , \24003 , \22333 );
and \U$26448 ( \26826 , \23978 , \22331 );
nor \U$26449 ( \26827 , \26825 , \26826 );
xnor \U$26450 ( \26828 , \26827 , \22239 );
and \U$26451 ( \26829 , \24344 , \22163 );
and \U$26452 ( \26830 , \24177 , \22161 );
nor \U$26453 ( \26831 , \26829 , \26830 );
xnor \U$26454 ( \26832 , \26831 , \22091 );
and \U$26455 ( \26833 , \26828 , \26832 );
and \U$26456 ( \26834 , \24601 , \22029 );
and \U$26457 ( \26835 , \24482 , \22027 );
nor \U$26458 ( \26836 , \26834 , \26835 );
xnor \U$26459 ( \26837 , \26836 , \21986 );
and \U$26460 ( \26838 , \26832 , \26837 );
and \U$26461 ( \26839 , \26828 , \26837 );
or \U$26462 ( \26840 , \26833 , \26838 , \26839 );
and \U$26463 ( \26841 , \26823 , \26840 );
and \U$26464 ( \26842 , \26807 , \26840 );
or \U$26465 ( \26843 , \26824 , \26841 , \26842 );
and \U$26466 ( \26844 , \26791 , \26843 );
and \U$26467 ( \26845 , \26116 , \21697 );
and \U$26468 ( \26846 , \26108 , \21695 );
nor \U$26469 ( \26847 , \26845 , \26846 );
xnor \U$26470 ( \26848 , \26847 , \21678 );
and \U$26471 ( \26849 , \26590 , \21660 );
and \U$26472 ( \26850 , \26585 , \21658 );
nor \U$26473 ( \26851 , \26849 , \26850 );
xnor \U$26474 ( \26852 , \26851 , \21665 );
and \U$26475 ( \26853 , \26848 , \26852 );
buf \U$26476 ( \26854 , RIc22aa30_173);
and \U$26477 ( \26855 , \26854 , \21654 );
and \U$26478 ( \26856 , \26852 , \26855 );
and \U$26479 ( \26857 , \26848 , \26855 );
or \U$26480 ( \26858 , \26853 , \26856 , \26857 );
and \U$26481 ( \26859 , \25226 , \21916 );
and \U$26482 ( \26860 , \25018 , \21914 );
nor \U$26483 ( \26861 , \26859 , \26860 );
xnor \U$26484 ( \26862 , \26861 , \21867 );
and \U$26485 ( \26863 , \25353 , \21815 );
and \U$26486 ( \26864 , \25348 , \21813 );
nor \U$26487 ( \26865 , \26863 , \26864 );
xnor \U$26488 ( \26866 , \26865 , \21774 );
and \U$26489 ( \26867 , \26862 , \26866 );
and \U$26490 ( \26868 , \25806 , \21745 );
and \U$26491 ( \26869 , \25609 , \21743 );
nor \U$26492 ( \26870 , \26868 , \26869 );
xnor \U$26493 ( \26871 , \26870 , \21715 );
and \U$26494 ( \26872 , \26866 , \26871 );
and \U$26495 ( \26873 , \26862 , \26871 );
or \U$26496 ( \26874 , \26867 , \26872 , \26873 );
and \U$26497 ( \26875 , \26858 , \26874 );
xnor \U$26498 ( \26876 , \26589 , \26591 );
and \U$26499 ( \26877 , \26874 , \26876 );
and \U$26500 ( \26878 , \26858 , \26876 );
or \U$26501 ( \26879 , \26875 , \26877 , \26878 );
and \U$26502 ( \26880 , \26843 , \26879 );
and \U$26503 ( \26881 , \26791 , \26879 );
or \U$26504 ( \26882 , \26844 , \26880 , \26881 );
xor \U$26505 ( \26883 , \26572 , \26576 );
xor \U$26506 ( \26884 , \26883 , \26581 );
xor \U$26507 ( \26885 , \26621 , \26625 );
xor \U$26508 ( \26886 , \26885 , \26630 );
and \U$26509 ( \26887 , \26884 , \26886 );
xor \U$26510 ( \26888 , \26638 , \26642 );
xor \U$26511 ( \26889 , \26888 , \26647 );
and \U$26512 ( \26890 , \26886 , \26889 );
and \U$26513 ( \26891 , \26884 , \26889 );
or \U$26514 ( \26892 , \26887 , \26890 , \26891 );
xor \U$26515 ( \26893 , \26605 , \26609 );
xor \U$26516 ( \26894 , \26893 , \26614 );
xor \U$26517 ( \26895 , \26536 , \26540 );
xor \U$26518 ( \26896 , \26895 , \26545 );
and \U$26519 ( \26897 , \26894 , \26896 );
xor \U$26520 ( \26898 , \26553 , \26557 );
xor \U$26521 ( \26899 , \26898 , \26562 );
and \U$26522 ( \26900 , \26896 , \26899 );
and \U$26523 ( \26901 , \26894 , \26899 );
or \U$26524 ( \26902 , \26897 , \26900 , \26901 );
and \U$26525 ( \26903 , \26892 , \26902 );
xor \U$26526 ( \26904 , \26347 , \26351 );
xor \U$26527 ( \26905 , \26904 , \26356 );
and \U$26528 ( \26906 , \26902 , \26905 );
and \U$26529 ( \26907 , \26892 , \26905 );
or \U$26530 ( \26908 , \26903 , \26906 , \26907 );
and \U$26531 ( \26909 , \26882 , \26908 );
xor \U$26532 ( \26910 , \26330 , \26334 );
xor \U$26533 ( \26911 , \26910 , \26339 );
xor \U$26534 ( \26912 , \26657 , \26659 );
xor \U$26535 ( \26913 , \26912 , \26662 );
and \U$26536 ( \26914 , \26911 , \26913 );
xor \U$26537 ( \26915 , \26667 , \26669 );
xor \U$26538 ( \26916 , \26915 , \26672 );
and \U$26539 ( \26917 , \26913 , \26916 );
and \U$26540 ( \26918 , \26911 , \26916 );
or \U$26541 ( \26919 , \26914 , \26917 , \26918 );
and \U$26542 ( \26920 , \26908 , \26919 );
and \U$26543 ( \26921 , \26882 , \26919 );
or \U$26544 ( \26922 , \26909 , \26920 , \26921 );
xor \U$26545 ( \26923 , \26532 , \26548 );
xor \U$26546 ( \26924 , \26923 , \26565 );
xor \U$26547 ( \26925 , \26584 , \26592 );
xor \U$26548 ( \26926 , \26925 , \26597 );
and \U$26549 ( \26927 , \26924 , \26926 );
xor \U$26550 ( \26928 , \26617 , \26633 );
xor \U$26551 ( \26929 , \26928 , \26650 );
and \U$26552 ( \26930 , \26926 , \26929 );
and \U$26553 ( \26931 , \26924 , \26929 );
or \U$26554 ( \26932 , \26927 , \26930 , \26931 );
xor \U$26555 ( \26933 , \26324 , \26342 );
xor \U$26556 ( \26934 , \26933 , \26359 );
and \U$26557 ( \26935 , \26932 , \26934 );
xor \U$26558 ( \26936 , \26684 , \26686 );
xor \U$26559 ( \26937 , \26936 , \26689 );
and \U$26560 ( \26938 , \26934 , \26937 );
and \U$26561 ( \26939 , \26932 , \26937 );
or \U$26562 ( \26940 , \26935 , \26938 , \26939 );
and \U$26563 ( \26941 , \26922 , \26940 );
xor \U$26564 ( \26942 , \26451 , \26461 );
xor \U$26565 ( \26943 , \26942 , \26464 );
and \U$26566 ( \26944 , \26940 , \26943 );
and \U$26567 ( \26945 , \26922 , \26943 );
or \U$26568 ( \26946 , \26941 , \26944 , \26945 );
xor \U$26569 ( \26947 , \26362 , \26414 );
xor \U$26570 ( \26948 , \26947 , \26438 );
xor \U$26571 ( \26949 , \26656 , \26681 );
xor \U$26572 ( \26950 , \26949 , \26692 );
and \U$26573 ( \26951 , \26948 , \26950 );
xor \U$26574 ( \26952 , \26697 , \26699 );
xor \U$26575 ( \26953 , \26952 , \26702 );
and \U$26576 ( \26954 , \26950 , \26953 );
and \U$26577 ( \26955 , \26948 , \26953 );
or \U$26578 ( \26956 , \26951 , \26954 , \26955 );
and \U$26579 ( \26957 , \26946 , \26956 );
xor \U$26580 ( \26958 , \26483 , \26485 );
xor \U$26581 ( \26959 , \26958 , \26488 );
and \U$26582 ( \26960 , \26956 , \26959 );
and \U$26583 ( \26961 , \26946 , \26959 );
or \U$26584 ( \26962 , \26957 , \26960 , \26961 );
xor \U$26585 ( \26963 , \26441 , \26467 );
xor \U$26586 ( \26964 , \26963 , \26478 );
xor \U$26587 ( \26965 , \26695 , \26705 );
xor \U$26588 ( \26966 , \26965 , \26708 );
and \U$26589 ( \26967 , \26964 , \26966 );
and \U$26590 ( \26968 , \26962 , \26967 );
xor \U$26591 ( \26969 , \26711 , \26713 );
xor \U$26592 ( \26970 , \26969 , \26716 );
and \U$26593 ( \26971 , \26967 , \26970 );
and \U$26594 ( \26972 , \26962 , \26970 );
or \U$26595 ( \26973 , \26968 , \26971 , \26972 );
xor \U$26596 ( \26974 , \26719 , \26721 );
xor \U$26597 ( \26975 , \26974 , \26724 );
and \U$26598 ( \26976 , \26973 , \26975 );
and \U$26599 ( \26977 , \26737 , \26976 );
xor \U$26600 ( \26978 , \26737 , \26976 );
xor \U$26601 ( \26979 , \26973 , \26975 );
xor \U$26602 ( \26980 , \26326 , \26738 );
xor \U$26603 ( \26981 , \26738 , \26739 );
not \U$26604 ( \26982 , \26981 );
and \U$26605 ( \26983 , \26980 , \26982 );
and \U$26606 ( \26984 , \21653 , \26983 );
not \U$26607 ( \26985 , \26984 );
xnor \U$26608 ( \26986 , \26985 , \26742 );
and \U$26609 ( \26987 , \21685 , \26517 );
and \U$26610 ( \26988 , \21667 , \26515 );
nor \U$26611 ( \26989 , \26987 , \26988 );
xnor \U$26612 ( \26990 , \26989 , \26329 );
and \U$26613 ( \26991 , \26986 , \26990 );
and \U$26614 ( \26992 , \21754 , \26143 );
and \U$26615 ( \26993 , \21706 , \26141 );
nor \U$26616 ( \26994 , \26992 , \26993 );
xnor \U$26617 ( \26995 , \26994 , \25911 );
and \U$26618 ( \26996 , \26990 , \26995 );
and \U$26619 ( \26997 , \26986 , \26995 );
or \U$26620 ( \26998 , \26991 , \26996 , \26997 );
and \U$26621 ( \26999 , \21831 , \25692 );
and \U$26622 ( \27000 , \21762 , \25690 );
nor \U$26623 ( \27001 , \26999 , \27000 );
xnor \U$26624 ( \27002 , \27001 , \25549 );
and \U$26625 ( \27003 , \21890 , \25369 );
and \U$26626 ( \27004 , \21836 , \25367 );
nor \U$26627 ( \27005 , \27003 , \27004 );
xnor \U$26628 ( \27006 , \27005 , \25123 );
and \U$26629 ( \27007 , \27002 , \27006 );
and \U$26630 ( \27008 , \22018 , \24974 );
and \U$26631 ( \27009 , \21941 , \24972 );
nor \U$26632 ( \27010 , \27008 , \27009 );
xnor \U$26633 ( \27011 , \27010 , \24787 );
and \U$26634 ( \27012 , \27006 , \27011 );
and \U$26635 ( \27013 , \27002 , \27011 );
or \U$26636 ( \27014 , \27007 , \27012 , \27013 );
and \U$26637 ( \27015 , \26998 , \27014 );
and \U$26638 ( \27016 , \22126 , \24661 );
and \U$26639 ( \27017 , \22046 , \24659 );
nor \U$26640 ( \27018 , \27016 , \27017 );
xnor \U$26641 ( \27019 , \27018 , \24456 );
and \U$26642 ( \27020 , \22262 , \24255 );
and \U$26643 ( \27021 , \22200 , \24253 );
nor \U$26644 ( \27022 , \27020 , \27021 );
xnor \U$26645 ( \27023 , \27022 , \24106 );
and \U$26646 ( \27024 , \27019 , \27023 );
and \U$26647 ( \27025 , \22523 , \23933 );
and \U$26648 ( \27026 , \22325 , \23931 );
nor \U$26649 ( \27027 , \27025 , \27026 );
xnor \U$26650 ( \27028 , \27027 , \23791 );
and \U$26651 ( \27029 , \27023 , \27028 );
and \U$26652 ( \27030 , \27019 , \27028 );
or \U$26653 ( \27031 , \27024 , \27029 , \27030 );
and \U$26654 ( \27032 , \27014 , \27031 );
and \U$26655 ( \27033 , \26998 , \27031 );
or \U$26656 ( \27034 , \27015 , \27032 , \27033 );
and \U$26657 ( \27035 , \22716 , \23637 );
and \U$26658 ( \27036 , \22611 , \23635 );
nor \U$26659 ( \27037 , \27035 , \27036 );
xnor \U$26660 ( \27038 , \27037 , \23500 );
and \U$26661 ( \27039 , \22837 , \23431 );
and \U$26662 ( \27040 , \22721 , \23429 );
nor \U$26663 ( \27041 , \27039 , \27040 );
xnor \U$26664 ( \27042 , \27041 , \23279 );
and \U$26665 ( \27043 , \27038 , \27042 );
and \U$26666 ( \27044 , \23128 , \23163 );
and \U$26667 ( \27045 , \22952 , \23161 );
nor \U$26668 ( \27046 , \27044 , \27045 );
xnor \U$26669 ( \27047 , \27046 , \23007 );
and \U$26670 ( \27048 , \27042 , \27047 );
and \U$26671 ( \27049 , \27038 , \27047 );
or \U$26672 ( \27050 , \27043 , \27048 , \27049 );
and \U$26673 ( \27051 , \23379 , \22891 );
and \U$26674 ( \27052 , \23136 , \22889 );
nor \U$26675 ( \27053 , \27051 , \27052 );
xnor \U$26676 ( \27054 , \27053 , \22778 );
and \U$26677 ( \27055 , \23570 , \22697 );
and \U$26678 ( \27056 , \23384 , \22695 );
nor \U$26679 ( \27057 , \27055 , \27056 );
xnor \U$26680 ( \27058 , \27057 , \22561 );
and \U$26681 ( \27059 , \27054 , \27058 );
and \U$26682 ( \27060 , \23978 , \22497 );
and \U$26683 ( \27061 , \23714 , \22495 );
nor \U$26684 ( \27062 , \27060 , \27061 );
xnor \U$26685 ( \27063 , \27062 , \22419 );
and \U$26686 ( \27064 , \27058 , \27063 );
and \U$26687 ( \27065 , \27054 , \27063 );
or \U$26688 ( \27066 , \27059 , \27064 , \27065 );
and \U$26689 ( \27067 , \27050 , \27066 );
and \U$26690 ( \27068 , \24177 , \22333 );
and \U$26691 ( \27069 , \24003 , \22331 );
nor \U$26692 ( \27070 , \27068 , \27069 );
xnor \U$26693 ( \27071 , \27070 , \22239 );
and \U$26694 ( \27072 , \24482 , \22163 );
and \U$26695 ( \27073 , \24344 , \22161 );
nor \U$26696 ( \27074 , \27072 , \27073 );
xnor \U$26697 ( \27075 , \27074 , \22091 );
and \U$26698 ( \27076 , \27071 , \27075 );
and \U$26699 ( \27077 , \25018 , \22029 );
and \U$26700 ( \27078 , \24601 , \22027 );
nor \U$26701 ( \27079 , \27077 , \27078 );
xnor \U$26702 ( \27080 , \27079 , \21986 );
and \U$26703 ( \27081 , \27075 , \27080 );
and \U$26704 ( \27082 , \27071 , \27080 );
or \U$26705 ( \27083 , \27076 , \27081 , \27082 );
and \U$26706 ( \27084 , \27066 , \27083 );
and \U$26707 ( \27085 , \27050 , \27083 );
or \U$26708 ( \27086 , \27067 , \27084 , \27085 );
and \U$26709 ( \27087 , \27034 , \27086 );
and \U$26710 ( \27088 , \25348 , \21916 );
and \U$26711 ( \27089 , \25226 , \21914 );
nor \U$26712 ( \27090 , \27088 , \27089 );
xnor \U$26713 ( \27091 , \27090 , \21867 );
and \U$26714 ( \27092 , \25609 , \21815 );
and \U$26715 ( \27093 , \25353 , \21813 );
nor \U$26716 ( \27094 , \27092 , \27093 );
xnor \U$26717 ( \27095 , \27094 , \21774 );
and \U$26718 ( \27096 , \27091 , \27095 );
and \U$26719 ( \27097 , \26108 , \21745 );
and \U$26720 ( \27098 , \25806 , \21743 );
nor \U$26721 ( \27099 , \27097 , \27098 );
xnor \U$26722 ( \27100 , \27099 , \21715 );
and \U$26723 ( \27101 , \27095 , \27100 );
and \U$26724 ( \27102 , \27091 , \27100 );
or \U$26725 ( \27103 , \27096 , \27101 , \27102 );
and \U$26726 ( \27104 , \26585 , \21697 );
and \U$26727 ( \27105 , \26116 , \21695 );
nor \U$26728 ( \27106 , \27104 , \27105 );
xnor \U$26729 ( \27107 , \27106 , \21678 );
and \U$26730 ( \27108 , \26854 , \21660 );
and \U$26731 ( \27109 , \26590 , \21658 );
nor \U$26732 ( \27110 , \27108 , \27109 );
xnor \U$26733 ( \27111 , \27110 , \21665 );
and \U$26734 ( \27112 , \27107 , \27111 );
buf \U$26735 ( \27113 , RIc22aaa8_174);
and \U$26736 ( \27114 , \27113 , \21654 );
and \U$26737 ( \27115 , \27111 , \27114 );
and \U$26738 ( \27116 , \27107 , \27114 );
or \U$26739 ( \27117 , \27112 , \27115 , \27116 );
and \U$26740 ( \27118 , \27103 , \27117 );
xor \U$26741 ( \27119 , \26848 , \26852 );
xor \U$26742 ( \27120 , \27119 , \26855 );
and \U$26743 ( \27121 , \27117 , \27120 );
and \U$26744 ( \27122 , \27103 , \27120 );
or \U$26745 ( \27123 , \27118 , \27121 , \27122 );
and \U$26746 ( \27124 , \27086 , \27123 );
and \U$26747 ( \27125 , \27034 , \27123 );
or \U$26748 ( \27126 , \27087 , \27124 , \27125 );
xor \U$26749 ( \27127 , \26795 , \26799 );
xor \U$26750 ( \27128 , \27127 , \26804 );
xor \U$26751 ( \27129 , \26759 , \26763 );
xor \U$26752 ( \27130 , \27129 , \26768 );
and \U$26753 ( \27131 , \27128 , \27130 );
xor \U$26754 ( \27132 , \26776 , \26780 );
xor \U$26755 ( \27133 , \27132 , \26785 );
and \U$26756 ( \27134 , \27130 , \27133 );
and \U$26757 ( \27135 , \27128 , \27133 );
or \U$26758 ( \27136 , \27131 , \27134 , \27135 );
xor \U$26759 ( \27137 , \26811 , \26815 );
xor \U$26760 ( \27138 , \27137 , \26820 );
xor \U$26761 ( \27139 , \26828 , \26832 );
xor \U$26762 ( \27140 , \27139 , \26837 );
and \U$26763 ( \27141 , \27138 , \27140 );
xor \U$26764 ( \27142 , \26862 , \26866 );
xor \U$26765 ( \27143 , \27142 , \26871 );
and \U$26766 ( \27144 , \27140 , \27143 );
and \U$26767 ( \27145 , \27138 , \27143 );
or \U$26768 ( \27146 , \27141 , \27144 , \27145 );
and \U$26769 ( \27147 , \27136 , \27146 );
xor \U$26770 ( \27148 , \26520 , \26524 );
xor \U$26771 ( \27149 , \27148 , \26529 );
and \U$26772 ( \27150 , \27146 , \27149 );
and \U$26773 ( \27151 , \27136 , \27149 );
or \U$26774 ( \27152 , \27147 , \27150 , \27151 );
and \U$26775 ( \27153 , \27126 , \27152 );
xor \U$26776 ( \27154 , \26884 , \26886 );
xor \U$26777 ( \27155 , \27154 , \26889 );
xor \U$26778 ( \27156 , \26894 , \26896 );
xor \U$26779 ( \27157 , \27156 , \26899 );
and \U$26780 ( \27158 , \27155 , \27157 );
xor \U$26781 ( \27159 , \26858 , \26874 );
xor \U$26782 ( \27160 , \27159 , \26876 );
and \U$26783 ( \27161 , \27157 , \27160 );
and \U$26784 ( \27162 , \27155 , \27160 );
or \U$26785 ( \27163 , \27158 , \27161 , \27162 );
and \U$26786 ( \27164 , \27152 , \27163 );
and \U$26787 ( \27165 , \27126 , \27163 );
or \U$26788 ( \27166 , \27153 , \27164 , \27165 );
xor \U$26789 ( \27167 , \26892 , \26902 );
xor \U$26790 ( \27168 , \27167 , \26905 );
xor \U$26791 ( \27169 , \26924 , \26926 );
xor \U$26792 ( \27170 , \27169 , \26929 );
and \U$26793 ( \27171 , \27168 , \27170 );
xor \U$26794 ( \27172 , \26911 , \26913 );
xor \U$26795 ( \27173 , \27172 , \26916 );
and \U$26796 ( \27174 , \27170 , \27173 );
and \U$26797 ( \27175 , \27168 , \27173 );
or \U$26798 ( \27176 , \27171 , \27174 , \27175 );
and \U$26799 ( \27177 , \27166 , \27176 );
xor \U$26800 ( \27178 , \26665 , \26675 );
xor \U$26801 ( \27179 , \27178 , \26678 );
and \U$26802 ( \27180 , \27176 , \27179 );
and \U$26803 ( \27181 , \27166 , \27179 );
or \U$26804 ( \27182 , \27177 , \27180 , \27181 );
xor \U$26805 ( \27183 , \26568 , \26600 );
xor \U$26806 ( \27184 , \27183 , \26653 );
xor \U$26807 ( \27185 , \26882 , \26908 );
xor \U$26808 ( \27186 , \27185 , \26919 );
and \U$26809 ( \27187 , \27184 , \27186 );
xor \U$26810 ( \27188 , \26932 , \26934 );
xor \U$26811 ( \27189 , \27188 , \26937 );
and \U$26812 ( \27190 , \27186 , \27189 );
and \U$26813 ( \27191 , \27184 , \27189 );
or \U$26814 ( \27192 , \27187 , \27190 , \27191 );
and \U$26815 ( \27193 , \27182 , \27192 );
xor \U$26816 ( \27194 , \26948 , \26950 );
xor \U$26817 ( \27195 , \27194 , \26953 );
and \U$26818 ( \27196 , \27192 , \27195 );
and \U$26819 ( \27197 , \27182 , \27195 );
or \U$26820 ( \27198 , \27193 , \27196 , \27197 );
xor \U$26821 ( \27199 , \26946 , \26956 );
xor \U$26822 ( \27200 , \27199 , \26959 );
and \U$26823 ( \27201 , \27198 , \27200 );
xor \U$26824 ( \27202 , \26964 , \26966 );
and \U$26825 ( \27203 , \27200 , \27202 );
and \U$26826 ( \27204 , \27198 , \27202 );
or \U$26827 ( \27205 , \27201 , \27203 , \27204 );
xor \U$26828 ( \27206 , \26962 , \26967 );
xor \U$26829 ( \27207 , \27206 , \26970 );
and \U$26830 ( \27208 , \27205 , \27207 );
and \U$26831 ( \27209 , \26979 , \27208 );
xor \U$26832 ( \27210 , \26979 , \27208 );
xor \U$26833 ( \27211 , \27205 , \27207 );
and \U$26834 ( \27212 , \21762 , \26143 );
and \U$26835 ( \27213 , \21754 , \26141 );
nor \U$26836 ( \27214 , \27212 , \27213 );
xnor \U$26837 ( \27215 , \27214 , \25911 );
and \U$26838 ( \27216 , \21836 , \25692 );
and \U$26839 ( \27217 , \21831 , \25690 );
nor \U$26840 ( \27218 , \27216 , \27217 );
xnor \U$26841 ( \27219 , \27218 , \25549 );
and \U$26842 ( \27220 , \27215 , \27219 );
and \U$26843 ( \27221 , \21941 , \25369 );
and \U$26844 ( \27222 , \21890 , \25367 );
nor \U$26845 ( \27223 , \27221 , \27222 );
xnor \U$26846 ( \27224 , \27223 , \25123 );
and \U$26847 ( \27225 , \27219 , \27224 );
and \U$26848 ( \27226 , \27215 , \27224 );
or \U$26849 ( \27227 , \27220 , \27225 , \27226 );
buf \U$26850 ( \27228 , RIc225fa8_48);
buf \U$26851 ( \27229 , RIc225f30_49);
and \U$26852 ( \27230 , \27228 , \27229 );
not \U$26853 ( \27231 , \27230 );
and \U$26854 ( \27232 , \26739 , \27231 );
not \U$26855 ( \27233 , \27232 );
and \U$26856 ( \27234 , \21667 , \26983 );
and \U$26857 ( \27235 , \21653 , \26981 );
nor \U$26858 ( \27236 , \27234 , \27235 );
xnor \U$26859 ( \27237 , \27236 , \26742 );
and \U$26860 ( \27238 , \27233 , \27237 );
and \U$26861 ( \27239 , \21706 , \26517 );
and \U$26862 ( \27240 , \21685 , \26515 );
nor \U$26863 ( \27241 , \27239 , \27240 );
xnor \U$26864 ( \27242 , \27241 , \26329 );
and \U$26865 ( \27243 , \27237 , \27242 );
and \U$26866 ( \27244 , \27233 , \27242 );
or \U$26867 ( \27245 , \27238 , \27243 , \27244 );
and \U$26868 ( \27246 , \27227 , \27245 );
and \U$26869 ( \27247 , \22046 , \24974 );
and \U$26870 ( \27248 , \22018 , \24972 );
nor \U$26871 ( \27249 , \27247 , \27248 );
xnor \U$26872 ( \27250 , \27249 , \24787 );
and \U$26873 ( \27251 , \22200 , \24661 );
and \U$26874 ( \27252 , \22126 , \24659 );
nor \U$26875 ( \27253 , \27251 , \27252 );
xnor \U$26876 ( \27254 , \27253 , \24456 );
and \U$26877 ( \27255 , \27250 , \27254 );
and \U$26878 ( \27256 , \22325 , \24255 );
and \U$26879 ( \27257 , \22262 , \24253 );
nor \U$26880 ( \27258 , \27256 , \27257 );
xnor \U$26881 ( \27259 , \27258 , \24106 );
and \U$26882 ( \27260 , \27254 , \27259 );
and \U$26883 ( \27261 , \27250 , \27259 );
or \U$26884 ( \27262 , \27255 , \27260 , \27261 );
and \U$26885 ( \27263 , \27245 , \27262 );
and \U$26886 ( \27264 , \27227 , \27262 );
or \U$26887 ( \27265 , \27246 , \27263 , \27264 );
and \U$26888 ( \27266 , \24003 , \22497 );
and \U$26889 ( \27267 , \23978 , \22495 );
nor \U$26890 ( \27268 , \27266 , \27267 );
xnor \U$26891 ( \27269 , \27268 , \22419 );
and \U$26892 ( \27270 , \24344 , \22333 );
and \U$26893 ( \27271 , \24177 , \22331 );
nor \U$26894 ( \27272 , \27270 , \27271 );
xnor \U$26895 ( \27273 , \27272 , \22239 );
and \U$26896 ( \27274 , \27269 , \27273 );
and \U$26897 ( \27275 , \24601 , \22163 );
and \U$26898 ( \27276 , \24482 , \22161 );
nor \U$26899 ( \27277 , \27275 , \27276 );
xnor \U$26900 ( \27278 , \27277 , \22091 );
and \U$26901 ( \27279 , \27273 , \27278 );
and \U$26902 ( \27280 , \27269 , \27278 );
or \U$26903 ( \27281 , \27274 , \27279 , \27280 );
and \U$26904 ( \27282 , \23136 , \23163 );
and \U$26905 ( \27283 , \23128 , \23161 );
nor \U$26906 ( \27284 , \27282 , \27283 );
xnor \U$26907 ( \27285 , \27284 , \23007 );
and \U$26908 ( \27286 , \23384 , \22891 );
and \U$26909 ( \27287 , \23379 , \22889 );
nor \U$26910 ( \27288 , \27286 , \27287 );
xnor \U$26911 ( \27289 , \27288 , \22778 );
and \U$26912 ( \27290 , \27285 , \27289 );
and \U$26913 ( \27291 , \23714 , \22697 );
and \U$26914 ( \27292 , \23570 , \22695 );
nor \U$26915 ( \27293 , \27291 , \27292 );
xnor \U$26916 ( \27294 , \27293 , \22561 );
and \U$26917 ( \27295 , \27289 , \27294 );
and \U$26918 ( \27296 , \27285 , \27294 );
or \U$26919 ( \27297 , \27290 , \27295 , \27296 );
and \U$26920 ( \27298 , \27281 , \27297 );
and \U$26921 ( \27299 , \22611 , \23933 );
and \U$26922 ( \27300 , \22523 , \23931 );
nor \U$26923 ( \27301 , \27299 , \27300 );
xnor \U$26924 ( \27302 , \27301 , \23791 );
and \U$26925 ( \27303 , \22721 , \23637 );
and \U$26926 ( \27304 , \22716 , \23635 );
nor \U$26927 ( \27305 , \27303 , \27304 );
xnor \U$26928 ( \27306 , \27305 , \23500 );
and \U$26929 ( \27307 , \27302 , \27306 );
and \U$26930 ( \27308 , \22952 , \23431 );
and \U$26931 ( \27309 , \22837 , \23429 );
nor \U$26932 ( \27310 , \27308 , \27309 );
xnor \U$26933 ( \27311 , \27310 , \23279 );
and \U$26934 ( \27312 , \27306 , \27311 );
and \U$26935 ( \27313 , \27302 , \27311 );
or \U$26936 ( \27314 , \27307 , \27312 , \27313 );
and \U$26937 ( \27315 , \27297 , \27314 );
and \U$26938 ( \27316 , \27281 , \27314 );
or \U$26939 ( \27317 , \27298 , \27315 , \27316 );
and \U$26940 ( \27318 , \27265 , \27317 );
and \U$26941 ( \27319 , \25226 , \22029 );
and \U$26942 ( \27320 , \25018 , \22027 );
nor \U$26943 ( \27321 , \27319 , \27320 );
xnor \U$26944 ( \27322 , \27321 , \21986 );
and \U$26945 ( \27323 , \25353 , \21916 );
and \U$26946 ( \27324 , \25348 , \21914 );
nor \U$26947 ( \27325 , \27323 , \27324 );
xnor \U$26948 ( \27326 , \27325 , \21867 );
and \U$26949 ( \27327 , \27322 , \27326 );
and \U$26950 ( \27328 , \25806 , \21815 );
and \U$26951 ( \27329 , \25609 , \21813 );
nor \U$26952 ( \27330 , \27328 , \27329 );
xnor \U$26953 ( \27331 , \27330 , \21774 );
and \U$26954 ( \27332 , \27326 , \27331 );
and \U$26955 ( \27333 , \27322 , \27331 );
or \U$26956 ( \27334 , \27327 , \27332 , \27333 );
and \U$26957 ( \27335 , \26116 , \21745 );
and \U$26958 ( \27336 , \26108 , \21743 );
nor \U$26959 ( \27337 , \27335 , \27336 );
xnor \U$26960 ( \27338 , \27337 , \21715 );
and \U$26961 ( \27339 , \26590 , \21697 );
and \U$26962 ( \27340 , \26585 , \21695 );
nor \U$26963 ( \27341 , \27339 , \27340 );
xnor \U$26964 ( \27342 , \27341 , \21678 );
and \U$26965 ( \27343 , \27338 , \27342 );
and \U$26966 ( \27344 , \27113 , \21660 );
and \U$26967 ( \27345 , \26854 , \21658 );
nor \U$26968 ( \27346 , \27344 , \27345 );
xnor \U$26969 ( \27347 , \27346 , \21665 );
and \U$26970 ( \27348 , \27342 , \27347 );
and \U$26971 ( \27349 , \27338 , \27347 );
or \U$26972 ( \27350 , \27343 , \27348 , \27349 );
or \U$26973 ( \27351 , \27334 , \27350 );
and \U$26974 ( \27352 , \27317 , \27351 );
and \U$26975 ( \27353 , \27265 , \27351 );
or \U$26976 ( \27354 , \27318 , \27352 , \27353 );
xor \U$26977 ( \27355 , \27038 , \27042 );
xor \U$26978 ( \27356 , \27355 , \27047 );
xor \U$26979 ( \27357 , \27054 , \27058 );
xor \U$26980 ( \27358 , \27357 , \27063 );
and \U$26981 ( \27359 , \27356 , \27358 );
xor \U$26982 ( \27360 , \27019 , \27023 );
xor \U$26983 ( \27361 , \27360 , \27028 );
and \U$26984 ( \27362 , \27358 , \27361 );
and \U$26985 ( \27363 , \27356 , \27361 );
or \U$26986 ( \27364 , \27359 , \27362 , \27363 );
xor \U$26987 ( \27365 , \27071 , \27075 );
xor \U$26988 ( \27366 , \27365 , \27080 );
xor \U$26989 ( \27367 , \27091 , \27095 );
xor \U$26990 ( \27368 , \27367 , \27100 );
and \U$26991 ( \27369 , \27366 , \27368 );
xor \U$26992 ( \27370 , \27107 , \27111 );
xor \U$26993 ( \27371 , \27370 , \27114 );
and \U$26994 ( \27372 , \27368 , \27371 );
and \U$26995 ( \27373 , \27366 , \27371 );
or \U$26996 ( \27374 , \27369 , \27372 , \27373 );
and \U$26997 ( \27375 , \27364 , \27374 );
xor \U$26998 ( \27376 , \26986 , \26990 );
xor \U$26999 ( \27377 , \27376 , \26995 );
xor \U$27000 ( \27378 , \27002 , \27006 );
xor \U$27001 ( \27379 , \27378 , \27011 );
and \U$27002 ( \27380 , \27377 , \27379 );
and \U$27003 ( \27381 , \27374 , \27380 );
and \U$27004 ( \27382 , \27364 , \27380 );
or \U$27005 ( \27383 , \27375 , \27381 , \27382 );
and \U$27006 ( \27384 , \27354 , \27383 );
xor \U$27007 ( \27385 , \26743 , \26747 );
xor \U$27008 ( \27386 , \27385 , \26752 );
xor \U$27009 ( \27387 , \27128 , \27130 );
xor \U$27010 ( \27388 , \27387 , \27133 );
and \U$27011 ( \27389 , \27386 , \27388 );
xor \U$27012 ( \27390 , \27138 , \27140 );
xor \U$27013 ( \27391 , \27390 , \27143 );
and \U$27014 ( \27392 , \27388 , \27391 );
and \U$27015 ( \27393 , \27386 , \27391 );
or \U$27016 ( \27394 , \27389 , \27392 , \27393 );
and \U$27017 ( \27395 , \27383 , \27394 );
and \U$27018 ( \27396 , \27354 , \27394 );
or \U$27019 ( \27397 , \27384 , \27395 , \27396 );
xor \U$27020 ( \27398 , \26998 , \27014 );
xor \U$27021 ( \27399 , \27398 , \27031 );
xor \U$27022 ( \27400 , \27050 , \27066 );
xor \U$27023 ( \27401 , \27400 , \27083 );
and \U$27024 ( \27402 , \27399 , \27401 );
xor \U$27025 ( \27403 , \27103 , \27117 );
xor \U$27026 ( \27404 , \27403 , \27120 );
and \U$27027 ( \27405 , \27401 , \27404 );
and \U$27028 ( \27406 , \27399 , \27404 );
or \U$27029 ( \27407 , \27402 , \27405 , \27406 );
xor \U$27030 ( \27408 , \26755 , \26771 );
xor \U$27031 ( \27409 , \27408 , \26788 );
and \U$27032 ( \27410 , \27407 , \27409 );
xor \U$27033 ( \27411 , \26807 , \26823 );
xor \U$27034 ( \27412 , \27411 , \26840 );
and \U$27035 ( \27413 , \27409 , \27412 );
and \U$27036 ( \27414 , \27407 , \27412 );
or \U$27037 ( \27415 , \27410 , \27413 , \27414 );
and \U$27038 ( \27416 , \27397 , \27415 );
xor \U$27039 ( \27417 , \27034 , \27086 );
xor \U$27040 ( \27418 , \27417 , \27123 );
xor \U$27041 ( \27419 , \27136 , \27146 );
xor \U$27042 ( \27420 , \27419 , \27149 );
and \U$27043 ( \27421 , \27418 , \27420 );
xor \U$27044 ( \27422 , \27155 , \27157 );
xor \U$27045 ( \27423 , \27422 , \27160 );
and \U$27046 ( \27424 , \27420 , \27423 );
and \U$27047 ( \27425 , \27418 , \27423 );
or \U$27048 ( \27426 , \27421 , \27424 , \27425 );
and \U$27049 ( \27427 , \27415 , \27426 );
and \U$27050 ( \27428 , \27397 , \27426 );
or \U$27051 ( \27429 , \27416 , \27427 , \27428 );
xor \U$27052 ( \27430 , \26791 , \26843 );
xor \U$27053 ( \27431 , \27430 , \26879 );
xor \U$27054 ( \27432 , \27126 , \27152 );
xor \U$27055 ( \27433 , \27432 , \27163 );
and \U$27056 ( \27434 , \27431 , \27433 );
xor \U$27057 ( \27435 , \27168 , \27170 );
xor \U$27058 ( \27436 , \27435 , \27173 );
and \U$27059 ( \27437 , \27433 , \27436 );
and \U$27060 ( \27438 , \27431 , \27436 );
or \U$27061 ( \27439 , \27434 , \27437 , \27438 );
and \U$27062 ( \27440 , \27429 , \27439 );
xor \U$27063 ( \27441 , \27184 , \27186 );
xor \U$27064 ( \27442 , \27441 , \27189 );
and \U$27065 ( \27443 , \27439 , \27442 );
and \U$27066 ( \27444 , \27429 , \27442 );
or \U$27067 ( \27445 , \27440 , \27443 , \27444 );
xor \U$27068 ( \27446 , \26922 , \26940 );
xor \U$27069 ( \27447 , \27446 , \26943 );
and \U$27070 ( \27448 , \27445 , \27447 );
xor \U$27071 ( \27449 , \27182 , \27192 );
xor \U$27072 ( \27450 , \27449 , \27195 );
and \U$27073 ( \27451 , \27447 , \27450 );
and \U$27074 ( \27452 , \27445 , \27450 );
or \U$27075 ( \27453 , \27448 , \27451 , \27452 );
xor \U$27076 ( \27454 , \27198 , \27200 );
xor \U$27077 ( \27455 , \27454 , \27202 );
and \U$27078 ( \27456 , \27453 , \27455 );
and \U$27079 ( \27457 , \27211 , \27456 );
xor \U$27080 ( \27458 , \27211 , \27456 );
xor \U$27081 ( \27459 , \27453 , \27455 );
and \U$27082 ( \27460 , \25348 , \22029 );
and \U$27083 ( \27461 , \25226 , \22027 );
nor \U$27084 ( \27462 , \27460 , \27461 );
xnor \U$27085 ( \27463 , \27462 , \21986 );
and \U$27086 ( \27464 , \25609 , \21916 );
and \U$27087 ( \27465 , \25353 , \21914 );
nor \U$27088 ( \27466 , \27464 , \27465 );
xnor \U$27089 ( \27467 , \27466 , \21867 );
and \U$27090 ( \27468 , \27463 , \27467 );
and \U$27091 ( \27469 , \26108 , \21815 );
and \U$27092 ( \27470 , \25806 , \21813 );
nor \U$27093 ( \27471 , \27469 , \27470 );
xnor \U$27094 ( \27472 , \27471 , \21774 );
and \U$27095 ( \27473 , \27467 , \27472 );
and \U$27096 ( \27474 , \27463 , \27472 );
or \U$27097 ( \27475 , \27468 , \27473 , \27474 );
and \U$27098 ( \27476 , \26585 , \21745 );
and \U$27099 ( \27477 , \26116 , \21743 );
nor \U$27100 ( \27478 , \27476 , \27477 );
xnor \U$27101 ( \27479 , \27478 , \21715 );
and \U$27102 ( \27480 , \26854 , \21697 );
and \U$27103 ( \27481 , \26590 , \21695 );
nor \U$27104 ( \27482 , \27480 , \27481 );
xnor \U$27105 ( \27483 , \27482 , \21678 );
and \U$27106 ( \27484 , \27479 , \27483 );
buf \U$27107 ( \27485 , RIc22ab20_175);
and \U$27108 ( \27486 , \27485 , \21660 );
and \U$27109 ( \27487 , \27113 , \21658 );
nor \U$27110 ( \27488 , \27486 , \27487 );
xnor \U$27111 ( \27489 , \27488 , \21665 );
and \U$27112 ( \27490 , \27483 , \27489 );
and \U$27113 ( \27491 , \27479 , \27489 );
or \U$27114 ( \27492 , \27484 , \27490 , \27491 );
and \U$27115 ( \27493 , \27475 , \27492 );
buf \U$27116 ( \27494 , RIc22ab98_176);
and \U$27117 ( \27495 , \27494 , \21654 );
buf \U$27118 ( \27496 , \27495 );
and \U$27119 ( \27497 , \27492 , \27496 );
and \U$27120 ( \27498 , \27475 , \27496 );
or \U$27121 ( \27499 , \27493 , \27497 , \27498 );
and \U$27122 ( \27500 , \23379 , \23163 );
and \U$27123 ( \27501 , \23136 , \23161 );
nor \U$27124 ( \27502 , \27500 , \27501 );
xnor \U$27125 ( \27503 , \27502 , \23007 );
and \U$27126 ( \27504 , \23570 , \22891 );
and \U$27127 ( \27505 , \23384 , \22889 );
nor \U$27128 ( \27506 , \27504 , \27505 );
xnor \U$27129 ( \27507 , \27506 , \22778 );
and \U$27130 ( \27508 , \27503 , \27507 );
and \U$27131 ( \27509 , \23978 , \22697 );
and \U$27132 ( \27510 , \23714 , \22695 );
nor \U$27133 ( \27511 , \27509 , \27510 );
xnor \U$27134 ( \27512 , \27511 , \22561 );
and \U$27135 ( \27513 , \27507 , \27512 );
and \U$27136 ( \27514 , \27503 , \27512 );
or \U$27137 ( \27515 , \27508 , \27513 , \27514 );
and \U$27138 ( \27516 , \22716 , \23933 );
and \U$27139 ( \27517 , \22611 , \23931 );
nor \U$27140 ( \27518 , \27516 , \27517 );
xnor \U$27141 ( \27519 , \27518 , \23791 );
and \U$27142 ( \27520 , \22837 , \23637 );
and \U$27143 ( \27521 , \22721 , \23635 );
nor \U$27144 ( \27522 , \27520 , \27521 );
xnor \U$27145 ( \27523 , \27522 , \23500 );
and \U$27146 ( \27524 , \27519 , \27523 );
and \U$27147 ( \27525 , \23128 , \23431 );
and \U$27148 ( \27526 , \22952 , \23429 );
nor \U$27149 ( \27527 , \27525 , \27526 );
xnor \U$27150 ( \27528 , \27527 , \23279 );
and \U$27151 ( \27529 , \27523 , \27528 );
and \U$27152 ( \27530 , \27519 , \27528 );
or \U$27153 ( \27531 , \27524 , \27529 , \27530 );
and \U$27154 ( \27532 , \27515 , \27531 );
and \U$27155 ( \27533 , \24177 , \22497 );
and \U$27156 ( \27534 , \24003 , \22495 );
nor \U$27157 ( \27535 , \27533 , \27534 );
xnor \U$27158 ( \27536 , \27535 , \22419 );
and \U$27159 ( \27537 , \24482 , \22333 );
and \U$27160 ( \27538 , \24344 , \22331 );
nor \U$27161 ( \27539 , \27537 , \27538 );
xnor \U$27162 ( \27540 , \27539 , \22239 );
and \U$27163 ( \27541 , \27536 , \27540 );
and \U$27164 ( \27542 , \25018 , \22163 );
and \U$27165 ( \27543 , \24601 , \22161 );
nor \U$27166 ( \27544 , \27542 , \27543 );
xnor \U$27167 ( \27545 , \27544 , \22091 );
and \U$27168 ( \27546 , \27540 , \27545 );
and \U$27169 ( \27547 , \27536 , \27545 );
or \U$27170 ( \27548 , \27541 , \27546 , \27547 );
and \U$27171 ( \27549 , \27531 , \27548 );
and \U$27172 ( \27550 , \27515 , \27548 );
or \U$27173 ( \27551 , \27532 , \27549 , \27550 );
and \U$27174 ( \27552 , \27499 , \27551 );
and \U$27175 ( \27553 , \21831 , \26143 );
and \U$27176 ( \27554 , \21762 , \26141 );
nor \U$27177 ( \27555 , \27553 , \27554 );
xnor \U$27178 ( \27556 , \27555 , \25911 );
and \U$27179 ( \27557 , \21890 , \25692 );
and \U$27180 ( \27558 , \21836 , \25690 );
nor \U$27181 ( \27559 , \27557 , \27558 );
xnor \U$27182 ( \27560 , \27559 , \25549 );
and \U$27183 ( \27561 , \27556 , \27560 );
and \U$27184 ( \27562 , \22018 , \25369 );
and \U$27185 ( \27563 , \21941 , \25367 );
nor \U$27186 ( \27564 , \27562 , \27563 );
xnor \U$27187 ( \27565 , \27564 , \25123 );
and \U$27188 ( \27566 , \27560 , \27565 );
and \U$27189 ( \27567 , \27556 , \27565 );
or \U$27190 ( \27568 , \27561 , \27566 , \27567 );
xor \U$27191 ( \27569 , \26739 , \27228 );
xor \U$27192 ( \27570 , \27228 , \27229 );
not \U$27193 ( \27571 , \27570 );
and \U$27194 ( \27572 , \27569 , \27571 );
and \U$27195 ( \27573 , \21653 , \27572 );
not \U$27196 ( \27574 , \27573 );
xnor \U$27197 ( \27575 , \27574 , \27232 );
and \U$27198 ( \27576 , \21685 , \26983 );
and \U$27199 ( \27577 , \21667 , \26981 );
nor \U$27200 ( \27578 , \27576 , \27577 );
xnor \U$27201 ( \27579 , \27578 , \26742 );
and \U$27202 ( \27580 , \27575 , \27579 );
and \U$27203 ( \27581 , \21754 , \26517 );
and \U$27204 ( \27582 , \21706 , \26515 );
nor \U$27205 ( \27583 , \27581 , \27582 );
xnor \U$27206 ( \27584 , \27583 , \26329 );
and \U$27207 ( \27585 , \27579 , \27584 );
and \U$27208 ( \27586 , \27575 , \27584 );
or \U$27209 ( \27587 , \27580 , \27585 , \27586 );
and \U$27210 ( \27588 , \27568 , \27587 );
and \U$27211 ( \27589 , \22126 , \24974 );
and \U$27212 ( \27590 , \22046 , \24972 );
nor \U$27213 ( \27591 , \27589 , \27590 );
xnor \U$27214 ( \27592 , \27591 , \24787 );
and \U$27215 ( \27593 , \22262 , \24661 );
and \U$27216 ( \27594 , \22200 , \24659 );
nor \U$27217 ( \27595 , \27593 , \27594 );
xnor \U$27218 ( \27596 , \27595 , \24456 );
and \U$27219 ( \27597 , \27592 , \27596 );
and \U$27220 ( \27598 , \22523 , \24255 );
and \U$27221 ( \27599 , \22325 , \24253 );
nor \U$27222 ( \27600 , \27598 , \27599 );
xnor \U$27223 ( \27601 , \27600 , \24106 );
and \U$27224 ( \27602 , \27596 , \27601 );
and \U$27225 ( \27603 , \27592 , \27601 );
or \U$27226 ( \27604 , \27597 , \27602 , \27603 );
and \U$27227 ( \27605 , \27587 , \27604 );
and \U$27228 ( \27606 , \27568 , \27604 );
or \U$27229 ( \27607 , \27588 , \27605 , \27606 );
and \U$27230 ( \27608 , \27551 , \27607 );
and \U$27231 ( \27609 , \27499 , \27607 );
or \U$27232 ( \27610 , \27552 , \27608 , \27609 );
xor \U$27233 ( \27611 , \27215 , \27219 );
xor \U$27234 ( \27612 , \27611 , \27224 );
xor \U$27235 ( \27613 , \27233 , \27237 );
xor \U$27236 ( \27614 , \27613 , \27242 );
and \U$27237 ( \27615 , \27612 , \27614 );
xor \U$27238 ( \27616 , \27250 , \27254 );
xor \U$27239 ( \27617 , \27616 , \27259 );
and \U$27240 ( \27618 , \27614 , \27617 );
and \U$27241 ( \27619 , \27612 , \27617 );
or \U$27242 ( \27620 , \27615 , \27618 , \27619 );
xor \U$27243 ( \27621 , \27269 , \27273 );
xor \U$27244 ( \27622 , \27621 , \27278 );
xor \U$27245 ( \27623 , \27285 , \27289 );
xor \U$27246 ( \27624 , \27623 , \27294 );
and \U$27247 ( \27625 , \27622 , \27624 );
xor \U$27248 ( \27626 , \27302 , \27306 );
xor \U$27249 ( \27627 , \27626 , \27311 );
and \U$27250 ( \27628 , \27624 , \27627 );
and \U$27251 ( \27629 , \27622 , \27627 );
or \U$27252 ( \27630 , \27625 , \27628 , \27629 );
and \U$27253 ( \27631 , \27620 , \27630 );
and \U$27254 ( \27632 , \27485 , \21654 );
xor \U$27255 ( \27633 , \27322 , \27326 );
xor \U$27256 ( \27634 , \27633 , \27331 );
and \U$27257 ( \27635 , \27632 , \27634 );
xor \U$27258 ( \27636 , \27338 , \27342 );
xor \U$27259 ( \27637 , \27636 , \27347 );
and \U$27260 ( \27638 , \27634 , \27637 );
and \U$27261 ( \27639 , \27632 , \27637 );
or \U$27262 ( \27640 , \27635 , \27638 , \27639 );
and \U$27263 ( \27641 , \27630 , \27640 );
and \U$27264 ( \27642 , \27620 , \27640 );
or \U$27265 ( \27643 , \27631 , \27641 , \27642 );
and \U$27266 ( \27644 , \27610 , \27643 );
xor \U$27267 ( \27645 , \27356 , \27358 );
xor \U$27268 ( \27646 , \27645 , \27361 );
xor \U$27269 ( \27647 , \27366 , \27368 );
xor \U$27270 ( \27648 , \27647 , \27371 );
and \U$27271 ( \27649 , \27646 , \27648 );
xor \U$27272 ( \27650 , \27377 , \27379 );
and \U$27273 ( \27651 , \27648 , \27650 );
and \U$27274 ( \27652 , \27646 , \27650 );
or \U$27275 ( \27653 , \27649 , \27651 , \27652 );
and \U$27276 ( \27654 , \27643 , \27653 );
and \U$27277 ( \27655 , \27610 , \27653 );
or \U$27278 ( \27656 , \27644 , \27654 , \27655 );
xor \U$27279 ( \27657 , \27227 , \27245 );
xor \U$27280 ( \27658 , \27657 , \27262 );
xor \U$27281 ( \27659 , \27281 , \27297 );
xor \U$27282 ( \27660 , \27659 , \27314 );
and \U$27283 ( \27661 , \27658 , \27660 );
xnor \U$27284 ( \27662 , \27334 , \27350 );
and \U$27285 ( \27663 , \27660 , \27662 );
and \U$27286 ( \27664 , \27658 , \27662 );
or \U$27287 ( \27665 , \27661 , \27663 , \27664 );
xor \U$27288 ( \27666 , \27386 , \27388 );
xor \U$27289 ( \27667 , \27666 , \27391 );
and \U$27290 ( \27668 , \27665 , \27667 );
xor \U$27291 ( \27669 , \27399 , \27401 );
xor \U$27292 ( \27670 , \27669 , \27404 );
and \U$27293 ( \27671 , \27667 , \27670 );
and \U$27294 ( \27672 , \27665 , \27670 );
or \U$27295 ( \27673 , \27668 , \27671 , \27672 );
and \U$27296 ( \27674 , \27656 , \27673 );
xor \U$27297 ( \27675 , \27265 , \27317 );
xor \U$27298 ( \27676 , \27675 , \27351 );
xor \U$27299 ( \27677 , \27364 , \27374 );
xor \U$27300 ( \27678 , \27677 , \27380 );
and \U$27301 ( \27679 , \27676 , \27678 );
and \U$27302 ( \27680 , \27673 , \27679 );
and \U$27303 ( \27681 , \27656 , \27679 );
or \U$27304 ( \27682 , \27674 , \27680 , \27681 );
xor \U$27305 ( \27683 , \27354 , \27383 );
xor \U$27306 ( \27684 , \27683 , \27394 );
xor \U$27307 ( \27685 , \27407 , \27409 );
xor \U$27308 ( \27686 , \27685 , \27412 );
and \U$27309 ( \27687 , \27684 , \27686 );
xor \U$27310 ( \27688 , \27418 , \27420 );
xor \U$27311 ( \27689 , \27688 , \27423 );
and \U$27312 ( \27690 , \27686 , \27689 );
and \U$27313 ( \27691 , \27684 , \27689 );
or \U$27314 ( \27692 , \27687 , \27690 , \27691 );
and \U$27315 ( \27693 , \27682 , \27692 );
xor \U$27316 ( \27694 , \27431 , \27433 );
xor \U$27317 ( \27695 , \27694 , \27436 );
and \U$27318 ( \27696 , \27692 , \27695 );
and \U$27319 ( \27697 , \27682 , \27695 );
or \U$27320 ( \27698 , \27693 , \27696 , \27697 );
xor \U$27321 ( \27699 , \27166 , \27176 );
xor \U$27322 ( \27700 , \27699 , \27179 );
and \U$27323 ( \27701 , \27698 , \27700 );
xor \U$27324 ( \27702 , \27429 , \27439 );
xor \U$27325 ( \27703 , \27702 , \27442 );
and \U$27326 ( \27704 , \27700 , \27703 );
and \U$27327 ( \27705 , \27698 , \27703 );
or \U$27328 ( \27706 , \27701 , \27704 , \27705 );
xor \U$27329 ( \27707 , \27445 , \27447 );
xor \U$27330 ( \27708 , \27707 , \27450 );
and \U$27331 ( \27709 , \27706 , \27708 );
and \U$27332 ( \27710 , \27459 , \27709 );
xor \U$27333 ( \27711 , \27459 , \27709 );
xor \U$27334 ( \27712 , \27706 , \27708 );
xor \U$27335 ( \27713 , \27503 , \27507 );
xor \U$27336 ( \27714 , \27713 , \27512 );
xor \U$27337 ( \27715 , \27519 , \27523 );
xor \U$27338 ( \27716 , \27715 , \27528 );
and \U$27339 ( \27717 , \27714 , \27716 );
xor \U$27340 ( \27718 , \27536 , \27540 );
xor \U$27341 ( \27719 , \27718 , \27545 );
and \U$27342 ( \27720 , \27716 , \27719 );
and \U$27343 ( \27721 , \27714 , \27719 );
or \U$27344 ( \27722 , \27717 , \27720 , \27721 );
xor \U$27345 ( \27723 , \27556 , \27560 );
xor \U$27346 ( \27724 , \27723 , \27565 );
xor \U$27347 ( \27725 , \27575 , \27579 );
xor \U$27348 ( \27726 , \27725 , \27584 );
and \U$27349 ( \27727 , \27724 , \27726 );
xor \U$27350 ( \27728 , \27592 , \27596 );
xor \U$27351 ( \27729 , \27728 , \27601 );
and \U$27352 ( \27730 , \27726 , \27729 );
and \U$27353 ( \27731 , \27724 , \27729 );
or \U$27354 ( \27732 , \27727 , \27730 , \27731 );
and \U$27355 ( \27733 , \27722 , \27732 );
xor \U$27356 ( \27734 , \27463 , \27467 );
xor \U$27357 ( \27735 , \27734 , \27472 );
xor \U$27358 ( \27736 , \27479 , \27483 );
xor \U$27359 ( \27737 , \27736 , \27489 );
and \U$27360 ( \27738 , \27735 , \27737 );
not \U$27361 ( \27739 , \27495 );
and \U$27362 ( \27740 , \27737 , \27739 );
and \U$27363 ( \27741 , \27735 , \27739 );
or \U$27364 ( \27742 , \27738 , \27740 , \27741 );
and \U$27365 ( \27743 , \27732 , \27742 );
and \U$27366 ( \27744 , \27722 , \27742 );
or \U$27367 ( \27745 , \27733 , \27743 , \27744 );
and \U$27368 ( \27746 , \21762 , \26517 );
and \U$27369 ( \27747 , \21754 , \26515 );
nor \U$27370 ( \27748 , \27746 , \27747 );
xnor \U$27371 ( \27749 , \27748 , \26329 );
and \U$27372 ( \27750 , \21836 , \26143 );
and \U$27373 ( \27751 , \21831 , \26141 );
nor \U$27374 ( \27752 , \27750 , \27751 );
xnor \U$27375 ( \27753 , \27752 , \25911 );
and \U$27376 ( \27754 , \27749 , \27753 );
and \U$27377 ( \27755 , \21941 , \25692 );
and \U$27378 ( \27756 , \21890 , \25690 );
nor \U$27379 ( \27757 , \27755 , \27756 );
xnor \U$27380 ( \27758 , \27757 , \25549 );
and \U$27381 ( \27759 , \27753 , \27758 );
and \U$27382 ( \27760 , \27749 , \27758 );
or \U$27383 ( \27761 , \27754 , \27759 , \27760 );
buf \U$27384 ( \27762 , RIc225eb8_50);
buf \U$27385 ( \27763 , RIc225e40_51);
and \U$27386 ( \27764 , \27762 , \27763 );
not \U$27387 ( \27765 , \27764 );
and \U$27388 ( \27766 , \27229 , \27765 );
not \U$27389 ( \27767 , \27766 );
and \U$27390 ( \27768 , \21667 , \27572 );
and \U$27391 ( \27769 , \21653 , \27570 );
nor \U$27392 ( \27770 , \27768 , \27769 );
xnor \U$27393 ( \27771 , \27770 , \27232 );
and \U$27394 ( \27772 , \27767 , \27771 );
and \U$27395 ( \27773 , \21706 , \26983 );
and \U$27396 ( \27774 , \21685 , \26981 );
nor \U$27397 ( \27775 , \27773 , \27774 );
xnor \U$27398 ( \27776 , \27775 , \26742 );
and \U$27399 ( \27777 , \27771 , \27776 );
and \U$27400 ( \27778 , \27767 , \27776 );
or \U$27401 ( \27779 , \27772 , \27777 , \27778 );
and \U$27402 ( \27780 , \27761 , \27779 );
and \U$27403 ( \27781 , \22046 , \25369 );
and \U$27404 ( \27782 , \22018 , \25367 );
nor \U$27405 ( \27783 , \27781 , \27782 );
xnor \U$27406 ( \27784 , \27783 , \25123 );
and \U$27407 ( \27785 , \22200 , \24974 );
and \U$27408 ( \27786 , \22126 , \24972 );
nor \U$27409 ( \27787 , \27785 , \27786 );
xnor \U$27410 ( \27788 , \27787 , \24787 );
and \U$27411 ( \27789 , \27784 , \27788 );
and \U$27412 ( \27790 , \22325 , \24661 );
and \U$27413 ( \27791 , \22262 , \24659 );
nor \U$27414 ( \27792 , \27790 , \27791 );
xnor \U$27415 ( \27793 , \27792 , \24456 );
and \U$27416 ( \27794 , \27788 , \27793 );
and \U$27417 ( \27795 , \27784 , \27793 );
or \U$27418 ( \27796 , \27789 , \27794 , \27795 );
and \U$27419 ( \27797 , \27779 , \27796 );
and \U$27420 ( \27798 , \27761 , \27796 );
or \U$27421 ( \27799 , \27780 , \27797 , \27798 );
and \U$27422 ( \27800 , \25226 , \22163 );
and \U$27423 ( \27801 , \25018 , \22161 );
nor \U$27424 ( \27802 , \27800 , \27801 );
xnor \U$27425 ( \27803 , \27802 , \22091 );
and \U$27426 ( \27804 , \25353 , \22029 );
and \U$27427 ( \27805 , \25348 , \22027 );
nor \U$27428 ( \27806 , \27804 , \27805 );
xnor \U$27429 ( \27807 , \27806 , \21986 );
and \U$27430 ( \27808 , \27803 , \27807 );
and \U$27431 ( \27809 , \25806 , \21916 );
and \U$27432 ( \27810 , \25609 , \21914 );
nor \U$27433 ( \27811 , \27809 , \27810 );
xnor \U$27434 ( \27812 , \27811 , \21867 );
and \U$27435 ( \27813 , \27807 , \27812 );
and \U$27436 ( \27814 , \27803 , \27812 );
or \U$27437 ( \27815 , \27808 , \27813 , \27814 );
and \U$27438 ( \27816 , \26116 , \21815 );
and \U$27439 ( \27817 , \26108 , \21813 );
nor \U$27440 ( \27818 , \27816 , \27817 );
xnor \U$27441 ( \27819 , \27818 , \21774 );
and \U$27442 ( \27820 , \26590 , \21745 );
and \U$27443 ( \27821 , \26585 , \21743 );
nor \U$27444 ( \27822 , \27820 , \27821 );
xnor \U$27445 ( \27823 , \27822 , \21715 );
and \U$27446 ( \27824 , \27819 , \27823 );
and \U$27447 ( \27825 , \27113 , \21697 );
and \U$27448 ( \27826 , \26854 , \21695 );
nor \U$27449 ( \27827 , \27825 , \27826 );
xnor \U$27450 ( \27828 , \27827 , \21678 );
and \U$27451 ( \27829 , \27823 , \27828 );
and \U$27452 ( \27830 , \27819 , \27828 );
or \U$27453 ( \27831 , \27824 , \27829 , \27830 );
and \U$27454 ( \27832 , \27815 , \27831 );
and \U$27455 ( \27833 , \27494 , \21660 );
and \U$27456 ( \27834 , \27485 , \21658 );
nor \U$27457 ( \27835 , \27833 , \27834 );
xnor \U$27458 ( \27836 , \27835 , \21665 );
buf \U$27459 ( \27837 , RIc22ac10_177);
and \U$27460 ( \27838 , \27837 , \21654 );
and \U$27461 ( \27839 , \27836 , \27838 );
and \U$27462 ( \27840 , \27831 , \27839 );
and \U$27463 ( \27841 , \27815 , \27839 );
or \U$27464 ( \27842 , \27832 , \27840 , \27841 );
and \U$27465 ( \27843 , \27799 , \27842 );
and \U$27466 ( \27844 , \22611 , \24255 );
and \U$27467 ( \27845 , \22523 , \24253 );
nor \U$27468 ( \27846 , \27844 , \27845 );
xnor \U$27469 ( \27847 , \27846 , \24106 );
and \U$27470 ( \27848 , \22721 , \23933 );
and \U$27471 ( \27849 , \22716 , \23931 );
nor \U$27472 ( \27850 , \27848 , \27849 );
xnor \U$27473 ( \27851 , \27850 , \23791 );
and \U$27474 ( \27852 , \27847 , \27851 );
and \U$27475 ( \27853 , \22952 , \23637 );
and \U$27476 ( \27854 , \22837 , \23635 );
nor \U$27477 ( \27855 , \27853 , \27854 );
xnor \U$27478 ( \27856 , \27855 , \23500 );
and \U$27479 ( \27857 , \27851 , \27856 );
and \U$27480 ( \27858 , \27847 , \27856 );
or \U$27481 ( \27859 , \27852 , \27857 , \27858 );
and \U$27482 ( \27860 , \23136 , \23431 );
and \U$27483 ( \27861 , \23128 , \23429 );
nor \U$27484 ( \27862 , \27860 , \27861 );
xnor \U$27485 ( \27863 , \27862 , \23279 );
and \U$27486 ( \27864 , \23384 , \23163 );
and \U$27487 ( \27865 , \23379 , \23161 );
nor \U$27488 ( \27866 , \27864 , \27865 );
xnor \U$27489 ( \27867 , \27866 , \23007 );
and \U$27490 ( \27868 , \27863 , \27867 );
and \U$27491 ( \27869 , \23714 , \22891 );
and \U$27492 ( \27870 , \23570 , \22889 );
nor \U$27493 ( \27871 , \27869 , \27870 );
xnor \U$27494 ( \27872 , \27871 , \22778 );
and \U$27495 ( \27873 , \27867 , \27872 );
and \U$27496 ( \27874 , \27863 , \27872 );
or \U$27497 ( \27875 , \27868 , \27873 , \27874 );
and \U$27498 ( \27876 , \27859 , \27875 );
and \U$27499 ( \27877 , \24003 , \22697 );
and \U$27500 ( \27878 , \23978 , \22695 );
nor \U$27501 ( \27879 , \27877 , \27878 );
xnor \U$27502 ( \27880 , \27879 , \22561 );
and \U$27503 ( \27881 , \24344 , \22497 );
and \U$27504 ( \27882 , \24177 , \22495 );
nor \U$27505 ( \27883 , \27881 , \27882 );
xnor \U$27506 ( \27884 , \27883 , \22419 );
and \U$27507 ( \27885 , \27880 , \27884 );
and \U$27508 ( \27886 , \24601 , \22333 );
and \U$27509 ( \27887 , \24482 , \22331 );
nor \U$27510 ( \27888 , \27886 , \27887 );
xnor \U$27511 ( \27889 , \27888 , \22239 );
and \U$27512 ( \27890 , \27884 , \27889 );
and \U$27513 ( \27891 , \27880 , \27889 );
or \U$27514 ( \27892 , \27885 , \27890 , \27891 );
and \U$27515 ( \27893 , \27875 , \27892 );
and \U$27516 ( \27894 , \27859 , \27892 );
or \U$27517 ( \27895 , \27876 , \27893 , \27894 );
and \U$27518 ( \27896 , \27842 , \27895 );
and \U$27519 ( \27897 , \27799 , \27895 );
or \U$27520 ( \27898 , \27843 , \27896 , \27897 );
and \U$27521 ( \27899 , \27745 , \27898 );
xor \U$27522 ( \27900 , \27612 , \27614 );
xor \U$27523 ( \27901 , \27900 , \27617 );
xor \U$27524 ( \27902 , \27622 , \27624 );
xor \U$27525 ( \27903 , \27902 , \27627 );
and \U$27526 ( \27904 , \27901 , \27903 );
xor \U$27527 ( \27905 , \27632 , \27634 );
xor \U$27528 ( \27906 , \27905 , \27637 );
and \U$27529 ( \27907 , \27903 , \27906 );
and \U$27530 ( \27908 , \27901 , \27906 );
or \U$27531 ( \27909 , \27904 , \27907 , \27908 );
and \U$27532 ( \27910 , \27898 , \27909 );
and \U$27533 ( \27911 , \27745 , \27909 );
or \U$27534 ( \27912 , \27899 , \27910 , \27911 );
xor \U$27535 ( \27913 , \27475 , \27492 );
xor \U$27536 ( \27914 , \27913 , \27496 );
xor \U$27537 ( \27915 , \27515 , \27531 );
xor \U$27538 ( \27916 , \27915 , \27548 );
and \U$27539 ( \27917 , \27914 , \27916 );
xor \U$27540 ( \27918 , \27568 , \27587 );
xor \U$27541 ( \27919 , \27918 , \27604 );
and \U$27542 ( \27920 , \27916 , \27919 );
and \U$27543 ( \27921 , \27914 , \27919 );
or \U$27544 ( \27922 , \27917 , \27920 , \27921 );
xor \U$27545 ( \27923 , \27658 , \27660 );
xor \U$27546 ( \27924 , \27923 , \27662 );
and \U$27547 ( \27925 , \27922 , \27924 );
xor \U$27548 ( \27926 , \27646 , \27648 );
xor \U$27549 ( \27927 , \27926 , \27650 );
and \U$27550 ( \27928 , \27924 , \27927 );
and \U$27551 ( \27929 , \27922 , \27927 );
or \U$27552 ( \27930 , \27925 , \27928 , \27929 );
and \U$27553 ( \27931 , \27912 , \27930 );
xor \U$27554 ( \27932 , \27499 , \27551 );
xor \U$27555 ( \27933 , \27932 , \27607 );
xor \U$27556 ( \27934 , \27620 , \27630 );
xor \U$27557 ( \27935 , \27934 , \27640 );
and \U$27558 ( \27936 , \27933 , \27935 );
and \U$27559 ( \27937 , \27930 , \27936 );
and \U$27560 ( \27938 , \27912 , \27936 );
or \U$27561 ( \27939 , \27931 , \27937 , \27938 );
xor \U$27562 ( \27940 , \27610 , \27643 );
xor \U$27563 ( \27941 , \27940 , \27653 );
xor \U$27564 ( \27942 , \27665 , \27667 );
xor \U$27565 ( \27943 , \27942 , \27670 );
and \U$27566 ( \27944 , \27941 , \27943 );
xor \U$27567 ( \27945 , \27676 , \27678 );
and \U$27568 ( \27946 , \27943 , \27945 );
and \U$27569 ( \27947 , \27941 , \27945 );
or \U$27570 ( \27948 , \27944 , \27946 , \27947 );
and \U$27571 ( \27949 , \27939 , \27948 );
xor \U$27572 ( \27950 , \27684 , \27686 );
xor \U$27573 ( \27951 , \27950 , \27689 );
and \U$27574 ( \27952 , \27948 , \27951 );
and \U$27575 ( \27953 , \27939 , \27951 );
or \U$27576 ( \27954 , \27949 , \27952 , \27953 );
xor \U$27577 ( \27955 , \27397 , \27415 );
xor \U$27578 ( \27956 , \27955 , \27426 );
and \U$27579 ( \27957 , \27954 , \27956 );
xor \U$27580 ( \27958 , \27682 , \27692 );
xor \U$27581 ( \27959 , \27958 , \27695 );
and \U$27582 ( \27960 , \27956 , \27959 );
and \U$27583 ( \27961 , \27954 , \27959 );
or \U$27584 ( \27962 , \27957 , \27960 , \27961 );
xor \U$27585 ( \27963 , \27698 , \27700 );
xor \U$27586 ( \27964 , \27963 , \27703 );
and \U$27587 ( \27965 , \27962 , \27964 );
and \U$27588 ( \27966 , \27712 , \27965 );
xor \U$27589 ( \27967 , \27712 , \27965 );
xor \U$27590 ( \27968 , \27962 , \27964 );
xor \U$27591 ( \27969 , \27847 , \27851 );
xor \U$27592 ( \27970 , \27969 , \27856 );
xor \U$27593 ( \27971 , \27863 , \27867 );
xor \U$27594 ( \27972 , \27971 , \27872 );
and \U$27595 ( \27973 , \27970 , \27972 );
xor \U$27596 ( \27974 , \27880 , \27884 );
xor \U$27597 ( \27975 , \27974 , \27889 );
and \U$27598 ( \27976 , \27972 , \27975 );
and \U$27599 ( \27977 , \27970 , \27975 );
or \U$27600 ( \27978 , \27973 , \27976 , \27977 );
xor \U$27601 ( \27979 , \27749 , \27753 );
xor \U$27602 ( \27980 , \27979 , \27758 );
xor \U$27603 ( \27981 , \27767 , \27771 );
xor \U$27604 ( \27982 , \27981 , \27776 );
and \U$27605 ( \27983 , \27980 , \27982 );
xor \U$27606 ( \27984 , \27784 , \27788 );
xor \U$27607 ( \27985 , \27984 , \27793 );
and \U$27608 ( \27986 , \27982 , \27985 );
and \U$27609 ( \27987 , \27980 , \27985 );
or \U$27610 ( \27988 , \27983 , \27986 , \27987 );
and \U$27611 ( \27989 , \27978 , \27988 );
xor \U$27612 ( \27990 , \27803 , \27807 );
xor \U$27613 ( \27991 , \27990 , \27812 );
xor \U$27614 ( \27992 , \27819 , \27823 );
xor \U$27615 ( \27993 , \27992 , \27828 );
and \U$27616 ( \27994 , \27991 , \27993 );
xor \U$27617 ( \27995 , \27836 , \27838 );
and \U$27618 ( \27996 , \27993 , \27995 );
and \U$27619 ( \27997 , \27991 , \27995 );
or \U$27620 ( \27998 , \27994 , \27996 , \27997 );
and \U$27621 ( \27999 , \27988 , \27998 );
and \U$27622 ( \28000 , \27978 , \27998 );
or \U$27623 ( \28001 , \27989 , \27999 , \28000 );
and \U$27624 ( \28002 , \25348 , \22163 );
and \U$27625 ( \28003 , \25226 , \22161 );
nor \U$27626 ( \28004 , \28002 , \28003 );
xnor \U$27627 ( \28005 , \28004 , \22091 );
and \U$27628 ( \28006 , \25609 , \22029 );
and \U$27629 ( \28007 , \25353 , \22027 );
nor \U$27630 ( \28008 , \28006 , \28007 );
xnor \U$27631 ( \28009 , \28008 , \21986 );
and \U$27632 ( \28010 , \28005 , \28009 );
and \U$27633 ( \28011 , \26108 , \21916 );
and \U$27634 ( \28012 , \25806 , \21914 );
nor \U$27635 ( \28013 , \28011 , \28012 );
xnor \U$27636 ( \28014 , \28013 , \21867 );
and \U$27637 ( \28015 , \28009 , \28014 );
and \U$27638 ( \28016 , \28005 , \28014 );
or \U$27639 ( \28017 , \28010 , \28015 , \28016 );
and \U$27640 ( \28018 , \26585 , \21815 );
and \U$27641 ( \28019 , \26116 , \21813 );
nor \U$27642 ( \28020 , \28018 , \28019 );
xnor \U$27643 ( \28021 , \28020 , \21774 );
and \U$27644 ( \28022 , \26854 , \21745 );
and \U$27645 ( \28023 , \26590 , \21743 );
nor \U$27646 ( \28024 , \28022 , \28023 );
xnor \U$27647 ( \28025 , \28024 , \21715 );
and \U$27648 ( \28026 , \28021 , \28025 );
and \U$27649 ( \28027 , \27485 , \21697 );
and \U$27650 ( \28028 , \27113 , \21695 );
nor \U$27651 ( \28029 , \28027 , \28028 );
xnor \U$27652 ( \28030 , \28029 , \21678 );
and \U$27653 ( \28031 , \28025 , \28030 );
and \U$27654 ( \28032 , \28021 , \28030 );
or \U$27655 ( \28033 , \28026 , \28031 , \28032 );
and \U$27656 ( \28034 , \28017 , \28033 );
and \U$27657 ( \28035 , \27837 , \21660 );
and \U$27658 ( \28036 , \27494 , \21658 );
nor \U$27659 ( \28037 , \28035 , \28036 );
xnor \U$27660 ( \28038 , \28037 , \21665 );
buf \U$27661 ( \28039 , RIc22ac88_178);
and \U$27662 ( \28040 , \28039 , \21654 );
or \U$27663 ( \28041 , \28038 , \28040 );
and \U$27664 ( \28042 , \28033 , \28041 );
and \U$27665 ( \28043 , \28017 , \28041 );
or \U$27666 ( \28044 , \28034 , \28042 , \28043 );
and \U$27667 ( \28045 , \22126 , \25369 );
and \U$27668 ( \28046 , \22046 , \25367 );
nor \U$27669 ( \28047 , \28045 , \28046 );
xnor \U$27670 ( \28048 , \28047 , \25123 );
and \U$27671 ( \28049 , \22262 , \24974 );
and \U$27672 ( \28050 , \22200 , \24972 );
nor \U$27673 ( \28051 , \28049 , \28050 );
xnor \U$27674 ( \28052 , \28051 , \24787 );
and \U$27675 ( \28053 , \28048 , \28052 );
and \U$27676 ( \28054 , \22523 , \24661 );
and \U$27677 ( \28055 , \22325 , \24659 );
nor \U$27678 ( \28056 , \28054 , \28055 );
xnor \U$27679 ( \28057 , \28056 , \24456 );
and \U$27680 ( \28058 , \28052 , \28057 );
and \U$27681 ( \28059 , \28048 , \28057 );
or \U$27682 ( \28060 , \28053 , \28058 , \28059 );
and \U$27683 ( \28061 , \21831 , \26517 );
and \U$27684 ( \28062 , \21762 , \26515 );
nor \U$27685 ( \28063 , \28061 , \28062 );
xnor \U$27686 ( \28064 , \28063 , \26329 );
and \U$27687 ( \28065 , \21890 , \26143 );
and \U$27688 ( \28066 , \21836 , \26141 );
nor \U$27689 ( \28067 , \28065 , \28066 );
xnor \U$27690 ( \28068 , \28067 , \25911 );
and \U$27691 ( \28069 , \28064 , \28068 );
and \U$27692 ( \28070 , \22018 , \25692 );
and \U$27693 ( \28071 , \21941 , \25690 );
nor \U$27694 ( \28072 , \28070 , \28071 );
xnor \U$27695 ( \28073 , \28072 , \25549 );
and \U$27696 ( \28074 , \28068 , \28073 );
and \U$27697 ( \28075 , \28064 , \28073 );
or \U$27698 ( \28076 , \28069 , \28074 , \28075 );
and \U$27699 ( \28077 , \28060 , \28076 );
xor \U$27700 ( \28078 , \27229 , \27762 );
xor \U$27701 ( \28079 , \27762 , \27763 );
not \U$27702 ( \28080 , \28079 );
and \U$27703 ( \28081 , \28078 , \28080 );
and \U$27704 ( \28082 , \21653 , \28081 );
not \U$27705 ( \28083 , \28082 );
xnor \U$27706 ( \28084 , \28083 , \27766 );
and \U$27707 ( \28085 , \21685 , \27572 );
and \U$27708 ( \28086 , \21667 , \27570 );
nor \U$27709 ( \28087 , \28085 , \28086 );
xnor \U$27710 ( \28088 , \28087 , \27232 );
and \U$27711 ( \28089 , \28084 , \28088 );
and \U$27712 ( \28090 , \21754 , \26983 );
and \U$27713 ( \28091 , \21706 , \26981 );
nor \U$27714 ( \28092 , \28090 , \28091 );
xnor \U$27715 ( \28093 , \28092 , \26742 );
and \U$27716 ( \28094 , \28088 , \28093 );
and \U$27717 ( \28095 , \28084 , \28093 );
or \U$27718 ( \28096 , \28089 , \28094 , \28095 );
and \U$27719 ( \28097 , \28076 , \28096 );
and \U$27720 ( \28098 , \28060 , \28096 );
or \U$27721 ( \28099 , \28077 , \28097 , \28098 );
and \U$27722 ( \28100 , \28044 , \28099 );
and \U$27723 ( \28101 , \23379 , \23431 );
and \U$27724 ( \28102 , \23136 , \23429 );
nor \U$27725 ( \28103 , \28101 , \28102 );
xnor \U$27726 ( \28104 , \28103 , \23279 );
and \U$27727 ( \28105 , \23570 , \23163 );
and \U$27728 ( \28106 , \23384 , \23161 );
nor \U$27729 ( \28107 , \28105 , \28106 );
xnor \U$27730 ( \28108 , \28107 , \23007 );
and \U$27731 ( \28109 , \28104 , \28108 );
and \U$27732 ( \28110 , \23978 , \22891 );
and \U$27733 ( \28111 , \23714 , \22889 );
nor \U$27734 ( \28112 , \28110 , \28111 );
xnor \U$27735 ( \28113 , \28112 , \22778 );
and \U$27736 ( \28114 , \28108 , \28113 );
and \U$27737 ( \28115 , \28104 , \28113 );
or \U$27738 ( \28116 , \28109 , \28114 , \28115 );
and \U$27739 ( \28117 , \24177 , \22697 );
and \U$27740 ( \28118 , \24003 , \22695 );
nor \U$27741 ( \28119 , \28117 , \28118 );
xnor \U$27742 ( \28120 , \28119 , \22561 );
and \U$27743 ( \28121 , \24482 , \22497 );
and \U$27744 ( \28122 , \24344 , \22495 );
nor \U$27745 ( \28123 , \28121 , \28122 );
xnor \U$27746 ( \28124 , \28123 , \22419 );
and \U$27747 ( \28125 , \28120 , \28124 );
and \U$27748 ( \28126 , \25018 , \22333 );
and \U$27749 ( \28127 , \24601 , \22331 );
nor \U$27750 ( \28128 , \28126 , \28127 );
xnor \U$27751 ( \28129 , \28128 , \22239 );
and \U$27752 ( \28130 , \28124 , \28129 );
and \U$27753 ( \28131 , \28120 , \28129 );
or \U$27754 ( \28132 , \28125 , \28130 , \28131 );
and \U$27755 ( \28133 , \28116 , \28132 );
and \U$27756 ( \28134 , \22716 , \24255 );
and \U$27757 ( \28135 , \22611 , \24253 );
nor \U$27758 ( \28136 , \28134 , \28135 );
xnor \U$27759 ( \28137 , \28136 , \24106 );
and \U$27760 ( \28138 , \22837 , \23933 );
and \U$27761 ( \28139 , \22721 , \23931 );
nor \U$27762 ( \28140 , \28138 , \28139 );
xnor \U$27763 ( \28141 , \28140 , \23791 );
and \U$27764 ( \28142 , \28137 , \28141 );
and \U$27765 ( \28143 , \23128 , \23637 );
and \U$27766 ( \28144 , \22952 , \23635 );
nor \U$27767 ( \28145 , \28143 , \28144 );
xnor \U$27768 ( \28146 , \28145 , \23500 );
and \U$27769 ( \28147 , \28141 , \28146 );
and \U$27770 ( \28148 , \28137 , \28146 );
or \U$27771 ( \28149 , \28142 , \28147 , \28148 );
and \U$27772 ( \28150 , \28132 , \28149 );
and \U$27773 ( \28151 , \28116 , \28149 );
or \U$27774 ( \28152 , \28133 , \28150 , \28151 );
and \U$27775 ( \28153 , \28099 , \28152 );
and \U$27776 ( \28154 , \28044 , \28152 );
or \U$27777 ( \28155 , \28100 , \28153 , \28154 );
and \U$27778 ( \28156 , \28001 , \28155 );
xor \U$27779 ( \28157 , \27714 , \27716 );
xor \U$27780 ( \28158 , \28157 , \27719 );
xor \U$27781 ( \28159 , \27724 , \27726 );
xor \U$27782 ( \28160 , \28159 , \27729 );
and \U$27783 ( \28161 , \28158 , \28160 );
xor \U$27784 ( \28162 , \27735 , \27737 );
xor \U$27785 ( \28163 , \28162 , \27739 );
and \U$27786 ( \28164 , \28160 , \28163 );
and \U$27787 ( \28165 , \28158 , \28163 );
or \U$27788 ( \28166 , \28161 , \28164 , \28165 );
and \U$27789 ( \28167 , \28155 , \28166 );
and \U$27790 ( \28168 , \28001 , \28166 );
or \U$27791 ( \28169 , \28156 , \28167 , \28168 );
xor \U$27792 ( \28170 , \27761 , \27779 );
xor \U$27793 ( \28171 , \28170 , \27796 );
xor \U$27794 ( \28172 , \27815 , \27831 );
xor \U$27795 ( \28173 , \28172 , \27839 );
and \U$27796 ( \28174 , \28171 , \28173 );
xor \U$27797 ( \28175 , \27859 , \27875 );
xor \U$27798 ( \28176 , \28175 , \27892 );
and \U$27799 ( \28177 , \28173 , \28176 );
and \U$27800 ( \28178 , \28171 , \28176 );
or \U$27801 ( \28179 , \28174 , \28177 , \28178 );
xor \U$27802 ( \28180 , \27914 , \27916 );
xor \U$27803 ( \28181 , \28180 , \27919 );
and \U$27804 ( \28182 , \28179 , \28181 );
xor \U$27805 ( \28183 , \27901 , \27903 );
xor \U$27806 ( \28184 , \28183 , \27906 );
and \U$27807 ( \28185 , \28181 , \28184 );
and \U$27808 ( \28186 , \28179 , \28184 );
or \U$27809 ( \28187 , \28182 , \28185 , \28186 );
and \U$27810 ( \28188 , \28169 , \28187 );
xor \U$27811 ( \28189 , \27722 , \27732 );
xor \U$27812 ( \28190 , \28189 , \27742 );
xor \U$27813 ( \28191 , \27799 , \27842 );
xor \U$27814 ( \28192 , \28191 , \27895 );
and \U$27815 ( \28193 , \28190 , \28192 );
and \U$27816 ( \28194 , \28187 , \28193 );
and \U$27817 ( \28195 , \28169 , \28193 );
or \U$27818 ( \28196 , \28188 , \28194 , \28195 );
xor \U$27819 ( \28197 , \27745 , \27898 );
xor \U$27820 ( \28198 , \28197 , \27909 );
xor \U$27821 ( \28199 , \27922 , \27924 );
xor \U$27822 ( \28200 , \28199 , \27927 );
and \U$27823 ( \28201 , \28198 , \28200 );
xor \U$27824 ( \28202 , \27933 , \27935 );
and \U$27825 ( \28203 , \28200 , \28202 );
and \U$27826 ( \28204 , \28198 , \28202 );
or \U$27827 ( \28205 , \28201 , \28203 , \28204 );
and \U$27828 ( \28206 , \28196 , \28205 );
xor \U$27829 ( \28207 , \27941 , \27943 );
xor \U$27830 ( \28208 , \28207 , \27945 );
and \U$27831 ( \28209 , \28205 , \28208 );
and \U$27832 ( \28210 , \28196 , \28208 );
or \U$27833 ( \28211 , \28206 , \28209 , \28210 );
xor \U$27834 ( \28212 , \27656 , \27673 );
xor \U$27835 ( \28213 , \28212 , \27679 );
and \U$27836 ( \28214 , \28211 , \28213 );
xor \U$27837 ( \28215 , \27939 , \27948 );
xor \U$27838 ( \28216 , \28215 , \27951 );
and \U$27839 ( \28217 , \28213 , \28216 );
and \U$27840 ( \28218 , \28211 , \28216 );
or \U$27841 ( \28219 , \28214 , \28217 , \28218 );
xor \U$27842 ( \28220 , \27954 , \27956 );
xor \U$27843 ( \28221 , \28220 , \27959 );
and \U$27844 ( \28222 , \28219 , \28221 );
and \U$27845 ( \28223 , \27968 , \28222 );
xor \U$27846 ( \28224 , \27968 , \28222 );
xor \U$27847 ( \28225 , \28219 , \28221 );
and \U$27848 ( \28226 , \22611 , \24661 );
and \U$27849 ( \28227 , \22523 , \24659 );
nor \U$27850 ( \28228 , \28226 , \28227 );
xnor \U$27851 ( \28229 , \28228 , \24456 );
and \U$27852 ( \28230 , \22721 , \24255 );
and \U$27853 ( \28231 , \22716 , \24253 );
nor \U$27854 ( \28232 , \28230 , \28231 );
xnor \U$27855 ( \28233 , \28232 , \24106 );
and \U$27856 ( \28234 , \28229 , \28233 );
and \U$27857 ( \28235 , \22952 , \23933 );
and \U$27858 ( \28236 , \22837 , \23931 );
nor \U$27859 ( \28237 , \28235 , \28236 );
xnor \U$27860 ( \28238 , \28237 , \23791 );
and \U$27861 ( \28239 , \28233 , \28238 );
and \U$27862 ( \28240 , \28229 , \28238 );
or \U$27863 ( \28241 , \28234 , \28239 , \28240 );
and \U$27864 ( \28242 , \23136 , \23637 );
and \U$27865 ( \28243 , \23128 , \23635 );
nor \U$27866 ( \28244 , \28242 , \28243 );
xnor \U$27867 ( \28245 , \28244 , \23500 );
and \U$27868 ( \28246 , \23384 , \23431 );
and \U$27869 ( \28247 , \23379 , \23429 );
nor \U$27870 ( \28248 , \28246 , \28247 );
xnor \U$27871 ( \28249 , \28248 , \23279 );
and \U$27872 ( \28250 , \28245 , \28249 );
and \U$27873 ( \28251 , \23714 , \23163 );
and \U$27874 ( \28252 , \23570 , \23161 );
nor \U$27875 ( \28253 , \28251 , \28252 );
xnor \U$27876 ( \28254 , \28253 , \23007 );
and \U$27877 ( \28255 , \28249 , \28254 );
and \U$27878 ( \28256 , \28245 , \28254 );
or \U$27879 ( \28257 , \28250 , \28255 , \28256 );
and \U$27880 ( \28258 , \28241 , \28257 );
and \U$27881 ( \28259 , \24003 , \22891 );
and \U$27882 ( \28260 , \23978 , \22889 );
nor \U$27883 ( \28261 , \28259 , \28260 );
xnor \U$27884 ( \28262 , \28261 , \22778 );
and \U$27885 ( \28263 , \24344 , \22697 );
and \U$27886 ( \28264 , \24177 , \22695 );
nor \U$27887 ( \28265 , \28263 , \28264 );
xnor \U$27888 ( \28266 , \28265 , \22561 );
and \U$27889 ( \28267 , \28262 , \28266 );
and \U$27890 ( \28268 , \24601 , \22497 );
and \U$27891 ( \28269 , \24482 , \22495 );
nor \U$27892 ( \28270 , \28268 , \28269 );
xnor \U$27893 ( \28271 , \28270 , \22419 );
and \U$27894 ( \28272 , \28266 , \28271 );
and \U$27895 ( \28273 , \28262 , \28271 );
or \U$27896 ( \28274 , \28267 , \28272 , \28273 );
and \U$27897 ( \28275 , \28257 , \28274 );
and \U$27898 ( \28276 , \28241 , \28274 );
or \U$27899 ( \28277 , \28258 , \28275 , \28276 );
and \U$27900 ( \28278 , \21762 , \26983 );
and \U$27901 ( \28279 , \21754 , \26981 );
nor \U$27902 ( \28280 , \28278 , \28279 );
xnor \U$27903 ( \28281 , \28280 , \26742 );
and \U$27904 ( \28282 , \21836 , \26517 );
and \U$27905 ( \28283 , \21831 , \26515 );
nor \U$27906 ( \28284 , \28282 , \28283 );
xnor \U$27907 ( \28285 , \28284 , \26329 );
and \U$27908 ( \28286 , \28281 , \28285 );
and \U$27909 ( \28287 , \21941 , \26143 );
and \U$27910 ( \28288 , \21890 , \26141 );
nor \U$27911 ( \28289 , \28287 , \28288 );
xnor \U$27912 ( \28290 , \28289 , \25911 );
and \U$27913 ( \28291 , \28285 , \28290 );
and \U$27914 ( \28292 , \28281 , \28290 );
or \U$27915 ( \28293 , \28286 , \28291 , \28292 );
and \U$27916 ( \28294 , \22046 , \25692 );
and \U$27917 ( \28295 , \22018 , \25690 );
nor \U$27918 ( \28296 , \28294 , \28295 );
xnor \U$27919 ( \28297 , \28296 , \25549 );
and \U$27920 ( \28298 , \22200 , \25369 );
and \U$27921 ( \28299 , \22126 , \25367 );
nor \U$27922 ( \28300 , \28298 , \28299 );
xnor \U$27923 ( \28301 , \28300 , \25123 );
and \U$27924 ( \28302 , \28297 , \28301 );
and \U$27925 ( \28303 , \22325 , \24974 );
and \U$27926 ( \28304 , \22262 , \24972 );
nor \U$27927 ( \28305 , \28303 , \28304 );
xnor \U$27928 ( \28306 , \28305 , \24787 );
and \U$27929 ( \28307 , \28301 , \28306 );
and \U$27930 ( \28308 , \28297 , \28306 );
or \U$27931 ( \28309 , \28302 , \28307 , \28308 );
and \U$27932 ( \28310 , \28293 , \28309 );
buf \U$27933 ( \28311 , RIc225dc8_52);
buf \U$27934 ( \28312 , RIc225d50_53);
and \U$27935 ( \28313 , \28311 , \28312 );
not \U$27936 ( \28314 , \28313 );
and \U$27937 ( \28315 , \27763 , \28314 );
not \U$27938 ( \28316 , \28315 );
and \U$27939 ( \28317 , \21667 , \28081 );
and \U$27940 ( \28318 , \21653 , \28079 );
nor \U$27941 ( \28319 , \28317 , \28318 );
xnor \U$27942 ( \28320 , \28319 , \27766 );
and \U$27943 ( \28321 , \28316 , \28320 );
and \U$27944 ( \28322 , \21706 , \27572 );
and \U$27945 ( \28323 , \21685 , \27570 );
nor \U$27946 ( \28324 , \28322 , \28323 );
xnor \U$27947 ( \28325 , \28324 , \27232 );
and \U$27948 ( \28326 , \28320 , \28325 );
and \U$27949 ( \28327 , \28316 , \28325 );
or \U$27950 ( \28328 , \28321 , \28326 , \28327 );
and \U$27951 ( \28329 , \28309 , \28328 );
and \U$27952 ( \28330 , \28293 , \28328 );
or \U$27953 ( \28331 , \28310 , \28329 , \28330 );
and \U$27954 ( \28332 , \28277 , \28331 );
and \U$27955 ( \28333 , \27494 , \21697 );
and \U$27956 ( \28334 , \27485 , \21695 );
nor \U$27957 ( \28335 , \28333 , \28334 );
xnor \U$27958 ( \28336 , \28335 , \21678 );
and \U$27959 ( \28337 , \28039 , \21660 );
and \U$27960 ( \28338 , \27837 , \21658 );
nor \U$27961 ( \28339 , \28337 , \28338 );
xnor \U$27962 ( \28340 , \28339 , \21665 );
and \U$27963 ( \28341 , \28336 , \28340 );
buf \U$27964 ( \28342 , RIc22ad00_179);
and \U$27965 ( \28343 , \28342 , \21654 );
and \U$27966 ( \28344 , \28340 , \28343 );
and \U$27967 ( \28345 , \28336 , \28343 );
or \U$27968 ( \28346 , \28341 , \28344 , \28345 );
and \U$27969 ( \28347 , \25226 , \22333 );
and \U$27970 ( \28348 , \25018 , \22331 );
nor \U$27971 ( \28349 , \28347 , \28348 );
xnor \U$27972 ( \28350 , \28349 , \22239 );
and \U$27973 ( \28351 , \25353 , \22163 );
and \U$27974 ( \28352 , \25348 , \22161 );
nor \U$27975 ( \28353 , \28351 , \28352 );
xnor \U$27976 ( \28354 , \28353 , \22091 );
and \U$27977 ( \28355 , \28350 , \28354 );
and \U$27978 ( \28356 , \25806 , \22029 );
and \U$27979 ( \28357 , \25609 , \22027 );
nor \U$27980 ( \28358 , \28356 , \28357 );
xnor \U$27981 ( \28359 , \28358 , \21986 );
and \U$27982 ( \28360 , \28354 , \28359 );
and \U$27983 ( \28361 , \28350 , \28359 );
or \U$27984 ( \28362 , \28355 , \28360 , \28361 );
and \U$27985 ( \28363 , \28346 , \28362 );
and \U$27986 ( \28364 , \26116 , \21916 );
and \U$27987 ( \28365 , \26108 , \21914 );
nor \U$27988 ( \28366 , \28364 , \28365 );
xnor \U$27989 ( \28367 , \28366 , \21867 );
and \U$27990 ( \28368 , \26590 , \21815 );
and \U$27991 ( \28369 , \26585 , \21813 );
nor \U$27992 ( \28370 , \28368 , \28369 );
xnor \U$27993 ( \28371 , \28370 , \21774 );
and \U$27994 ( \28372 , \28367 , \28371 );
and \U$27995 ( \28373 , \27113 , \21745 );
and \U$27996 ( \28374 , \26854 , \21743 );
nor \U$27997 ( \28375 , \28373 , \28374 );
xnor \U$27998 ( \28376 , \28375 , \21715 );
and \U$27999 ( \28377 , \28371 , \28376 );
and \U$28000 ( \28378 , \28367 , \28376 );
or \U$28001 ( \28379 , \28372 , \28377 , \28378 );
and \U$28002 ( \28380 , \28362 , \28379 );
and \U$28003 ( \28381 , \28346 , \28379 );
or \U$28004 ( \28382 , \28363 , \28380 , \28381 );
and \U$28005 ( \28383 , \28331 , \28382 );
and \U$28006 ( \28384 , \28277 , \28382 );
or \U$28007 ( \28385 , \28332 , \28383 , \28384 );
xor \U$28008 ( \28386 , \28104 , \28108 );
xor \U$28009 ( \28387 , \28386 , \28113 );
xor \U$28010 ( \28388 , \28120 , \28124 );
xor \U$28011 ( \28389 , \28388 , \28129 );
and \U$28012 ( \28390 , \28387 , \28389 );
xor \U$28013 ( \28391 , \28137 , \28141 );
xor \U$28014 ( \28392 , \28391 , \28146 );
and \U$28015 ( \28393 , \28389 , \28392 );
and \U$28016 ( \28394 , \28387 , \28392 );
or \U$28017 ( \28395 , \28390 , \28393 , \28394 );
xor \U$28018 ( \28396 , \28048 , \28052 );
xor \U$28019 ( \28397 , \28396 , \28057 );
xor \U$28020 ( \28398 , \28064 , \28068 );
xor \U$28021 ( \28399 , \28398 , \28073 );
and \U$28022 ( \28400 , \28397 , \28399 );
xor \U$28023 ( \28401 , \28084 , \28088 );
xor \U$28024 ( \28402 , \28401 , \28093 );
and \U$28025 ( \28403 , \28399 , \28402 );
and \U$28026 ( \28404 , \28397 , \28402 );
or \U$28027 ( \28405 , \28400 , \28403 , \28404 );
and \U$28028 ( \28406 , \28395 , \28405 );
xor \U$28029 ( \28407 , \28005 , \28009 );
xor \U$28030 ( \28408 , \28407 , \28014 );
xor \U$28031 ( \28409 , \28021 , \28025 );
xor \U$28032 ( \28410 , \28409 , \28030 );
and \U$28033 ( \28411 , \28408 , \28410 );
xnor \U$28034 ( \28412 , \28038 , \28040 );
and \U$28035 ( \28413 , \28410 , \28412 );
and \U$28036 ( \28414 , \28408 , \28412 );
or \U$28037 ( \28415 , \28411 , \28413 , \28414 );
and \U$28038 ( \28416 , \28405 , \28415 );
and \U$28039 ( \28417 , \28395 , \28415 );
or \U$28040 ( \28418 , \28406 , \28416 , \28417 );
and \U$28041 ( \28419 , \28385 , \28418 );
xor \U$28042 ( \28420 , \27970 , \27972 );
xor \U$28043 ( \28421 , \28420 , \27975 );
xor \U$28044 ( \28422 , \27980 , \27982 );
xor \U$28045 ( \28423 , \28422 , \27985 );
and \U$28046 ( \28424 , \28421 , \28423 );
xor \U$28047 ( \28425 , \27991 , \27993 );
xor \U$28048 ( \28426 , \28425 , \27995 );
and \U$28049 ( \28427 , \28423 , \28426 );
and \U$28050 ( \28428 , \28421 , \28426 );
or \U$28051 ( \28429 , \28424 , \28427 , \28428 );
and \U$28052 ( \28430 , \28418 , \28429 );
and \U$28053 ( \28431 , \28385 , \28429 );
or \U$28054 ( \28432 , \28419 , \28430 , \28431 );
xor \U$28055 ( \28433 , \28017 , \28033 );
xor \U$28056 ( \28434 , \28433 , \28041 );
xor \U$28057 ( \28435 , \28060 , \28076 );
xor \U$28058 ( \28436 , \28435 , \28096 );
and \U$28059 ( \28437 , \28434 , \28436 );
xor \U$28060 ( \28438 , \28116 , \28132 );
xor \U$28061 ( \28439 , \28438 , \28149 );
and \U$28062 ( \28440 , \28436 , \28439 );
and \U$28063 ( \28441 , \28434 , \28439 );
or \U$28064 ( \28442 , \28437 , \28440 , \28441 );
xor \U$28065 ( \28443 , \28171 , \28173 );
xor \U$28066 ( \28444 , \28443 , \28176 );
and \U$28067 ( \28445 , \28442 , \28444 );
xor \U$28068 ( \28446 , \28158 , \28160 );
xor \U$28069 ( \28447 , \28446 , \28163 );
and \U$28070 ( \28448 , \28444 , \28447 );
and \U$28071 ( \28449 , \28442 , \28447 );
or \U$28072 ( \28450 , \28445 , \28448 , \28449 );
and \U$28073 ( \28451 , \28432 , \28450 );
xor \U$28074 ( \28452 , \27978 , \27988 );
xor \U$28075 ( \28453 , \28452 , \27998 );
xor \U$28076 ( \28454 , \28044 , \28099 );
xor \U$28077 ( \28455 , \28454 , \28152 );
and \U$28078 ( \28456 , \28453 , \28455 );
and \U$28079 ( \28457 , \28450 , \28456 );
and \U$28080 ( \28458 , \28432 , \28456 );
or \U$28081 ( \28459 , \28451 , \28457 , \28458 );
xor \U$28082 ( \28460 , \28001 , \28155 );
xor \U$28083 ( \28461 , \28460 , \28166 );
xor \U$28084 ( \28462 , \28179 , \28181 );
xor \U$28085 ( \28463 , \28462 , \28184 );
and \U$28086 ( \28464 , \28461 , \28463 );
xor \U$28087 ( \28465 , \28190 , \28192 );
and \U$28088 ( \28466 , \28463 , \28465 );
and \U$28089 ( \28467 , \28461 , \28465 );
or \U$28090 ( \28468 , \28464 , \28466 , \28467 );
and \U$28091 ( \28469 , \28459 , \28468 );
xor \U$28092 ( \28470 , \28198 , \28200 );
xor \U$28093 ( \28471 , \28470 , \28202 );
and \U$28094 ( \28472 , \28468 , \28471 );
and \U$28095 ( \28473 , \28459 , \28471 );
or \U$28096 ( \28474 , \28469 , \28472 , \28473 );
xor \U$28097 ( \28475 , \27912 , \27930 );
xor \U$28098 ( \28476 , \28475 , \27936 );
and \U$28099 ( \28477 , \28474 , \28476 );
xor \U$28100 ( \28478 , \28196 , \28205 );
xor \U$28101 ( \28479 , \28478 , \28208 );
and \U$28102 ( \28480 , \28476 , \28479 );
and \U$28103 ( \28481 , \28474 , \28479 );
or \U$28104 ( \28482 , \28477 , \28480 , \28481 );
xor \U$28105 ( \28483 , \28211 , \28213 );
xor \U$28106 ( \28484 , \28483 , \28216 );
and \U$28107 ( \28485 , \28482 , \28484 );
and \U$28108 ( \28486 , \28225 , \28485 );
xor \U$28109 ( \28487 , \28225 , \28485 );
xor \U$28110 ( \28488 , \28482 , \28484 );
and \U$28111 ( \28489 , \25348 , \22333 );
and \U$28112 ( \28490 , \25226 , \22331 );
nor \U$28113 ( \28491 , \28489 , \28490 );
xnor \U$28114 ( \28492 , \28491 , \22239 );
and \U$28115 ( \28493 , \25609 , \22163 );
and \U$28116 ( \28494 , \25353 , \22161 );
nor \U$28117 ( \28495 , \28493 , \28494 );
xnor \U$28118 ( \28496 , \28495 , \22091 );
and \U$28119 ( \28497 , \28492 , \28496 );
and \U$28120 ( \28498 , \26108 , \22029 );
and \U$28121 ( \28499 , \25806 , \22027 );
nor \U$28122 ( \28500 , \28498 , \28499 );
xnor \U$28123 ( \28501 , \28500 , \21986 );
and \U$28124 ( \28502 , \28496 , \28501 );
and \U$28125 ( \28503 , \28492 , \28501 );
or \U$28126 ( \28504 , \28497 , \28502 , \28503 );
and \U$28127 ( \28505 , \27837 , \21697 );
and \U$28128 ( \28506 , \27494 , \21695 );
nor \U$28129 ( \28507 , \28505 , \28506 );
xnor \U$28130 ( \28508 , \28507 , \21678 );
and \U$28131 ( \28509 , \28342 , \21660 );
and \U$28132 ( \28510 , \28039 , \21658 );
nor \U$28133 ( \28511 , \28509 , \28510 );
xnor \U$28134 ( \28512 , \28511 , \21665 );
and \U$28135 ( \28513 , \28508 , \28512 );
buf \U$28136 ( \28514 , RIc22ad78_180);
and \U$28137 ( \28515 , \28514 , \21654 );
and \U$28138 ( \28516 , \28512 , \28515 );
and \U$28139 ( \28517 , \28508 , \28515 );
or \U$28140 ( \28518 , \28513 , \28516 , \28517 );
and \U$28141 ( \28519 , \28504 , \28518 );
and \U$28142 ( \28520 , \26585 , \21916 );
and \U$28143 ( \28521 , \26116 , \21914 );
nor \U$28144 ( \28522 , \28520 , \28521 );
xnor \U$28145 ( \28523 , \28522 , \21867 );
and \U$28146 ( \28524 , \26854 , \21815 );
and \U$28147 ( \28525 , \26590 , \21813 );
nor \U$28148 ( \28526 , \28524 , \28525 );
xnor \U$28149 ( \28527 , \28526 , \21774 );
and \U$28150 ( \28528 , \28523 , \28527 );
and \U$28151 ( \28529 , \27485 , \21745 );
and \U$28152 ( \28530 , \27113 , \21743 );
nor \U$28153 ( \28531 , \28529 , \28530 );
xnor \U$28154 ( \28532 , \28531 , \21715 );
and \U$28155 ( \28533 , \28527 , \28532 );
and \U$28156 ( \28534 , \28523 , \28532 );
or \U$28157 ( \28535 , \28528 , \28533 , \28534 );
and \U$28158 ( \28536 , \28518 , \28535 );
and \U$28159 ( \28537 , \28504 , \28535 );
or \U$28160 ( \28538 , \28519 , \28536 , \28537 );
and \U$28161 ( \28539 , \21831 , \26983 );
and \U$28162 ( \28540 , \21762 , \26981 );
nor \U$28163 ( \28541 , \28539 , \28540 );
xnor \U$28164 ( \28542 , \28541 , \26742 );
and \U$28165 ( \28543 , \21890 , \26517 );
and \U$28166 ( \28544 , \21836 , \26515 );
nor \U$28167 ( \28545 , \28543 , \28544 );
xnor \U$28168 ( \28546 , \28545 , \26329 );
and \U$28169 ( \28547 , \28542 , \28546 );
and \U$28170 ( \28548 , \22018 , \26143 );
and \U$28171 ( \28549 , \21941 , \26141 );
nor \U$28172 ( \28550 , \28548 , \28549 );
xnor \U$28173 ( \28551 , \28550 , \25911 );
and \U$28174 ( \28552 , \28546 , \28551 );
and \U$28175 ( \28553 , \28542 , \28551 );
or \U$28176 ( \28554 , \28547 , \28552 , \28553 );
and \U$28177 ( \28555 , \22126 , \25692 );
and \U$28178 ( \28556 , \22046 , \25690 );
nor \U$28179 ( \28557 , \28555 , \28556 );
xnor \U$28180 ( \28558 , \28557 , \25549 );
and \U$28181 ( \28559 , \22262 , \25369 );
and \U$28182 ( \28560 , \22200 , \25367 );
nor \U$28183 ( \28561 , \28559 , \28560 );
xnor \U$28184 ( \28562 , \28561 , \25123 );
and \U$28185 ( \28563 , \28558 , \28562 );
and \U$28186 ( \28564 , \22523 , \24974 );
and \U$28187 ( \28565 , \22325 , \24972 );
nor \U$28188 ( \28566 , \28564 , \28565 );
xnor \U$28189 ( \28567 , \28566 , \24787 );
and \U$28190 ( \28568 , \28562 , \28567 );
and \U$28191 ( \28569 , \28558 , \28567 );
or \U$28192 ( \28570 , \28563 , \28568 , \28569 );
and \U$28193 ( \28571 , \28554 , \28570 );
xor \U$28194 ( \28572 , \27763 , \28311 );
xor \U$28195 ( \28573 , \28311 , \28312 );
not \U$28196 ( \28574 , \28573 );
and \U$28197 ( \28575 , \28572 , \28574 );
and \U$28198 ( \28576 , \21653 , \28575 );
not \U$28199 ( \28577 , \28576 );
xnor \U$28200 ( \28578 , \28577 , \28315 );
and \U$28201 ( \28579 , \21685 , \28081 );
and \U$28202 ( \28580 , \21667 , \28079 );
nor \U$28203 ( \28581 , \28579 , \28580 );
xnor \U$28204 ( \28582 , \28581 , \27766 );
and \U$28205 ( \28583 , \28578 , \28582 );
and \U$28206 ( \28584 , \21754 , \27572 );
and \U$28207 ( \28585 , \21706 , \27570 );
nor \U$28208 ( \28586 , \28584 , \28585 );
xnor \U$28209 ( \28587 , \28586 , \27232 );
and \U$28210 ( \28588 , \28582 , \28587 );
and \U$28211 ( \28589 , \28578 , \28587 );
or \U$28212 ( \28590 , \28583 , \28588 , \28589 );
and \U$28213 ( \28591 , \28570 , \28590 );
and \U$28214 ( \28592 , \28554 , \28590 );
or \U$28215 ( \28593 , \28571 , \28591 , \28592 );
and \U$28216 ( \28594 , \28538 , \28593 );
and \U$28217 ( \28595 , \22716 , \24661 );
and \U$28218 ( \28596 , \22611 , \24659 );
nor \U$28219 ( \28597 , \28595 , \28596 );
xnor \U$28220 ( \28598 , \28597 , \24456 );
and \U$28221 ( \28599 , \22837 , \24255 );
and \U$28222 ( \28600 , \22721 , \24253 );
nor \U$28223 ( \28601 , \28599 , \28600 );
xnor \U$28224 ( \28602 , \28601 , \24106 );
and \U$28225 ( \28603 , \28598 , \28602 );
and \U$28226 ( \28604 , \23128 , \23933 );
and \U$28227 ( \28605 , \22952 , \23931 );
nor \U$28228 ( \28606 , \28604 , \28605 );
xnor \U$28229 ( \28607 , \28606 , \23791 );
and \U$28230 ( \28608 , \28602 , \28607 );
and \U$28231 ( \28609 , \28598 , \28607 );
or \U$28232 ( \28610 , \28603 , \28608 , \28609 );
and \U$28233 ( \28611 , \23379 , \23637 );
and \U$28234 ( \28612 , \23136 , \23635 );
nor \U$28235 ( \28613 , \28611 , \28612 );
xnor \U$28236 ( \28614 , \28613 , \23500 );
and \U$28237 ( \28615 , \23570 , \23431 );
and \U$28238 ( \28616 , \23384 , \23429 );
nor \U$28239 ( \28617 , \28615 , \28616 );
xnor \U$28240 ( \28618 , \28617 , \23279 );
and \U$28241 ( \28619 , \28614 , \28618 );
and \U$28242 ( \28620 , \23978 , \23163 );
and \U$28243 ( \28621 , \23714 , \23161 );
nor \U$28244 ( \28622 , \28620 , \28621 );
xnor \U$28245 ( \28623 , \28622 , \23007 );
and \U$28246 ( \28624 , \28618 , \28623 );
and \U$28247 ( \28625 , \28614 , \28623 );
or \U$28248 ( \28626 , \28619 , \28624 , \28625 );
and \U$28249 ( \28627 , \28610 , \28626 );
and \U$28250 ( \28628 , \24177 , \22891 );
and \U$28251 ( \28629 , \24003 , \22889 );
nor \U$28252 ( \28630 , \28628 , \28629 );
xnor \U$28253 ( \28631 , \28630 , \22778 );
and \U$28254 ( \28632 , \24482 , \22697 );
and \U$28255 ( \28633 , \24344 , \22695 );
nor \U$28256 ( \28634 , \28632 , \28633 );
xnor \U$28257 ( \28635 , \28634 , \22561 );
and \U$28258 ( \28636 , \28631 , \28635 );
and \U$28259 ( \28637 , \25018 , \22497 );
and \U$28260 ( \28638 , \24601 , \22495 );
nor \U$28261 ( \28639 , \28637 , \28638 );
xnor \U$28262 ( \28640 , \28639 , \22419 );
and \U$28263 ( \28641 , \28635 , \28640 );
and \U$28264 ( \28642 , \28631 , \28640 );
or \U$28265 ( \28643 , \28636 , \28641 , \28642 );
and \U$28266 ( \28644 , \28626 , \28643 );
and \U$28267 ( \28645 , \28610 , \28643 );
or \U$28268 ( \28646 , \28627 , \28644 , \28645 );
and \U$28269 ( \28647 , \28593 , \28646 );
and \U$28270 ( \28648 , \28538 , \28646 );
or \U$28271 ( \28649 , \28594 , \28647 , \28648 );
xor \U$28272 ( \28650 , \28336 , \28340 );
xor \U$28273 ( \28651 , \28650 , \28343 );
xor \U$28274 ( \28652 , \28350 , \28354 );
xor \U$28275 ( \28653 , \28652 , \28359 );
and \U$28276 ( \28654 , \28651 , \28653 );
xor \U$28277 ( \28655 , \28367 , \28371 );
xor \U$28278 ( \28656 , \28655 , \28376 );
and \U$28279 ( \28657 , \28653 , \28656 );
and \U$28280 ( \28658 , \28651 , \28656 );
or \U$28281 ( \28659 , \28654 , \28657 , \28658 );
xor \U$28282 ( \28660 , \28229 , \28233 );
xor \U$28283 ( \28661 , \28660 , \28238 );
xor \U$28284 ( \28662 , \28245 , \28249 );
xor \U$28285 ( \28663 , \28662 , \28254 );
and \U$28286 ( \28664 , \28661 , \28663 );
xor \U$28287 ( \28665 , \28262 , \28266 );
xor \U$28288 ( \28666 , \28665 , \28271 );
and \U$28289 ( \28667 , \28663 , \28666 );
and \U$28290 ( \28668 , \28661 , \28666 );
or \U$28291 ( \28669 , \28664 , \28667 , \28668 );
and \U$28292 ( \28670 , \28659 , \28669 );
xor \U$28293 ( \28671 , \28281 , \28285 );
xor \U$28294 ( \28672 , \28671 , \28290 );
xor \U$28295 ( \28673 , \28297 , \28301 );
xor \U$28296 ( \28674 , \28673 , \28306 );
and \U$28297 ( \28675 , \28672 , \28674 );
xor \U$28298 ( \28676 , \28316 , \28320 );
xor \U$28299 ( \28677 , \28676 , \28325 );
and \U$28300 ( \28678 , \28674 , \28677 );
and \U$28301 ( \28679 , \28672 , \28677 );
or \U$28302 ( \28680 , \28675 , \28678 , \28679 );
and \U$28303 ( \28681 , \28669 , \28680 );
and \U$28304 ( \28682 , \28659 , \28680 );
or \U$28305 ( \28683 , \28670 , \28681 , \28682 );
and \U$28306 ( \28684 , \28649 , \28683 );
xor \U$28307 ( \28685 , \28387 , \28389 );
xor \U$28308 ( \28686 , \28685 , \28392 );
xor \U$28309 ( \28687 , \28397 , \28399 );
xor \U$28310 ( \28688 , \28687 , \28402 );
and \U$28311 ( \28689 , \28686 , \28688 );
xor \U$28312 ( \28690 , \28408 , \28410 );
xor \U$28313 ( \28691 , \28690 , \28412 );
and \U$28314 ( \28692 , \28688 , \28691 );
and \U$28315 ( \28693 , \28686 , \28691 );
or \U$28316 ( \28694 , \28689 , \28692 , \28693 );
and \U$28317 ( \28695 , \28683 , \28694 );
and \U$28318 ( \28696 , \28649 , \28694 );
or \U$28319 ( \28697 , \28684 , \28695 , \28696 );
xor \U$28320 ( \28698 , \28241 , \28257 );
xor \U$28321 ( \28699 , \28698 , \28274 );
xor \U$28322 ( \28700 , \28293 , \28309 );
xor \U$28323 ( \28701 , \28700 , \28328 );
and \U$28324 ( \28702 , \28699 , \28701 );
xor \U$28325 ( \28703 , \28346 , \28362 );
xor \U$28326 ( \28704 , \28703 , \28379 );
and \U$28327 ( \28705 , \28701 , \28704 );
and \U$28328 ( \28706 , \28699 , \28704 );
or \U$28329 ( \28707 , \28702 , \28705 , \28706 );
xor \U$28330 ( \28708 , \28434 , \28436 );
xor \U$28331 ( \28709 , \28708 , \28439 );
and \U$28332 ( \28710 , \28707 , \28709 );
xor \U$28333 ( \28711 , \28421 , \28423 );
xor \U$28334 ( \28712 , \28711 , \28426 );
and \U$28335 ( \28713 , \28709 , \28712 );
and \U$28336 ( \28714 , \28707 , \28712 );
or \U$28337 ( \28715 , \28710 , \28713 , \28714 );
and \U$28338 ( \28716 , \28697 , \28715 );
xor \U$28339 ( \28717 , \28277 , \28331 );
xor \U$28340 ( \28718 , \28717 , \28382 );
xor \U$28341 ( \28719 , \28395 , \28405 );
xor \U$28342 ( \28720 , \28719 , \28415 );
and \U$28343 ( \28721 , \28718 , \28720 );
and \U$28344 ( \28722 , \28715 , \28721 );
and \U$28345 ( \28723 , \28697 , \28721 );
or \U$28346 ( \28724 , \28716 , \28722 , \28723 );
xor \U$28347 ( \28725 , \28385 , \28418 );
xor \U$28348 ( \28726 , \28725 , \28429 );
xor \U$28349 ( \28727 , \28442 , \28444 );
xor \U$28350 ( \28728 , \28727 , \28447 );
and \U$28351 ( \28729 , \28726 , \28728 );
xor \U$28352 ( \28730 , \28453 , \28455 );
and \U$28353 ( \28731 , \28728 , \28730 );
and \U$28354 ( \28732 , \28726 , \28730 );
or \U$28355 ( \28733 , \28729 , \28731 , \28732 );
and \U$28356 ( \28734 , \28724 , \28733 );
xor \U$28357 ( \28735 , \28461 , \28463 );
xor \U$28358 ( \28736 , \28735 , \28465 );
and \U$28359 ( \28737 , \28733 , \28736 );
and \U$28360 ( \28738 , \28724 , \28736 );
or \U$28361 ( \28739 , \28734 , \28737 , \28738 );
xor \U$28362 ( \28740 , \28169 , \28187 );
xor \U$28363 ( \28741 , \28740 , \28193 );
and \U$28364 ( \28742 , \28739 , \28741 );
xor \U$28365 ( \28743 , \28459 , \28468 );
xor \U$28366 ( \28744 , \28743 , \28471 );
and \U$28367 ( \28745 , \28741 , \28744 );
and \U$28368 ( \28746 , \28739 , \28744 );
or \U$28369 ( \28747 , \28742 , \28745 , \28746 );
xor \U$28370 ( \28748 , \28474 , \28476 );
xor \U$28371 ( \28749 , \28748 , \28479 );
and \U$28372 ( \28750 , \28747 , \28749 );
and \U$28373 ( \28751 , \28488 , \28750 );
xor \U$28374 ( \28752 , \28488 , \28750 );
xor \U$28375 ( \28753 , \28747 , \28749 );
xor \U$28376 ( \28754 , \28542 , \28546 );
xor \U$28377 ( \28755 , \28754 , \28551 );
xor \U$28378 ( \28756 , \28598 , \28602 );
xor \U$28379 ( \28757 , \28756 , \28607 );
and \U$28380 ( \28758 , \28755 , \28757 );
xor \U$28381 ( \28759 , \28558 , \28562 );
xor \U$28382 ( \28760 , \28759 , \28567 );
and \U$28383 ( \28761 , \28757 , \28760 );
and \U$28384 ( \28762 , \28755 , \28760 );
or \U$28385 ( \28763 , \28758 , \28761 , \28762 );
xor \U$28386 ( \28764 , \28614 , \28618 );
xor \U$28387 ( \28765 , \28764 , \28623 );
xor \U$28388 ( \28766 , \28492 , \28496 );
xor \U$28389 ( \28767 , \28766 , \28501 );
and \U$28390 ( \28768 , \28765 , \28767 );
xor \U$28391 ( \28769 , \28631 , \28635 );
xor \U$28392 ( \28770 , \28769 , \28640 );
and \U$28393 ( \28771 , \28767 , \28770 );
and \U$28394 ( \28772 , \28765 , \28770 );
or \U$28395 ( \28773 , \28768 , \28771 , \28772 );
and \U$28396 ( \28774 , \28763 , \28773 );
xor \U$28397 ( \28775 , \28508 , \28512 );
xor \U$28398 ( \28776 , \28775 , \28515 );
xor \U$28399 ( \28777 , \28523 , \28527 );
xor \U$28400 ( \28778 , \28777 , \28532 );
or \U$28401 ( \28779 , \28776 , \28778 );
and \U$28402 ( \28780 , \28773 , \28779 );
and \U$28403 ( \28781 , \28763 , \28779 );
or \U$28404 ( \28782 , \28774 , \28780 , \28781 );
and \U$28405 ( \28783 , \23136 , \23933 );
and \U$28406 ( \28784 , \23128 , \23931 );
nor \U$28407 ( \28785 , \28783 , \28784 );
xnor \U$28408 ( \28786 , \28785 , \23791 );
and \U$28409 ( \28787 , \23384 , \23637 );
and \U$28410 ( \28788 , \23379 , \23635 );
nor \U$28411 ( \28789 , \28787 , \28788 );
xnor \U$28412 ( \28790 , \28789 , \23500 );
and \U$28413 ( \28791 , \28786 , \28790 );
and \U$28414 ( \28792 , \23714 , \23431 );
and \U$28415 ( \28793 , \23570 , \23429 );
nor \U$28416 ( \28794 , \28792 , \28793 );
xnor \U$28417 ( \28795 , \28794 , \23279 );
and \U$28418 ( \28796 , \28790 , \28795 );
and \U$28419 ( \28797 , \28786 , \28795 );
or \U$28420 ( \28798 , \28791 , \28796 , \28797 );
and \U$28421 ( \28799 , \22611 , \24974 );
and \U$28422 ( \28800 , \22523 , \24972 );
nor \U$28423 ( \28801 , \28799 , \28800 );
xnor \U$28424 ( \28802 , \28801 , \24787 );
and \U$28425 ( \28803 , \22721 , \24661 );
and \U$28426 ( \28804 , \22716 , \24659 );
nor \U$28427 ( \28805 , \28803 , \28804 );
xnor \U$28428 ( \28806 , \28805 , \24456 );
and \U$28429 ( \28807 , \28802 , \28806 );
and \U$28430 ( \28808 , \22952 , \24255 );
and \U$28431 ( \28809 , \22837 , \24253 );
nor \U$28432 ( \28810 , \28808 , \28809 );
xnor \U$28433 ( \28811 , \28810 , \24106 );
and \U$28434 ( \28812 , \28806 , \28811 );
and \U$28435 ( \28813 , \28802 , \28811 );
or \U$28436 ( \28814 , \28807 , \28812 , \28813 );
and \U$28437 ( \28815 , \28798 , \28814 );
and \U$28438 ( \28816 , \24003 , \23163 );
and \U$28439 ( \28817 , \23978 , \23161 );
nor \U$28440 ( \28818 , \28816 , \28817 );
xnor \U$28441 ( \28819 , \28818 , \23007 );
and \U$28442 ( \28820 , \24344 , \22891 );
and \U$28443 ( \28821 , \24177 , \22889 );
nor \U$28444 ( \28822 , \28820 , \28821 );
xnor \U$28445 ( \28823 , \28822 , \22778 );
and \U$28446 ( \28824 , \28819 , \28823 );
and \U$28447 ( \28825 , \24601 , \22697 );
and \U$28448 ( \28826 , \24482 , \22695 );
nor \U$28449 ( \28827 , \28825 , \28826 );
xnor \U$28450 ( \28828 , \28827 , \22561 );
and \U$28451 ( \28829 , \28823 , \28828 );
and \U$28452 ( \28830 , \28819 , \28828 );
or \U$28453 ( \28831 , \28824 , \28829 , \28830 );
and \U$28454 ( \28832 , \28814 , \28831 );
and \U$28455 ( \28833 , \28798 , \28831 );
or \U$28456 ( \28834 , \28815 , \28832 , \28833 );
and \U$28457 ( \28835 , \21762 , \27572 );
and \U$28458 ( \28836 , \21754 , \27570 );
nor \U$28459 ( \28837 , \28835 , \28836 );
xnor \U$28460 ( \28838 , \28837 , \27232 );
and \U$28461 ( \28839 , \21836 , \26983 );
and \U$28462 ( \28840 , \21831 , \26981 );
nor \U$28463 ( \28841 , \28839 , \28840 );
xnor \U$28464 ( \28842 , \28841 , \26742 );
and \U$28465 ( \28843 , \28838 , \28842 );
and \U$28466 ( \28844 , \21941 , \26517 );
and \U$28467 ( \28845 , \21890 , \26515 );
nor \U$28468 ( \28846 , \28844 , \28845 );
xnor \U$28469 ( \28847 , \28846 , \26329 );
and \U$28470 ( \28848 , \28842 , \28847 );
and \U$28471 ( \28849 , \28838 , \28847 );
or \U$28472 ( \28850 , \28843 , \28848 , \28849 );
buf \U$28473 ( \28851 , RIc225cd8_54);
buf \U$28474 ( \28852 , RIc225c60_55);
and \U$28475 ( \28853 , \28851 , \28852 );
not \U$28476 ( \28854 , \28853 );
and \U$28477 ( \28855 , \28312 , \28854 );
not \U$28478 ( \28856 , \28855 );
and \U$28479 ( \28857 , \21667 , \28575 );
and \U$28480 ( \28858 , \21653 , \28573 );
nor \U$28481 ( \28859 , \28857 , \28858 );
xnor \U$28482 ( \28860 , \28859 , \28315 );
and \U$28483 ( \28861 , \28856 , \28860 );
and \U$28484 ( \28862 , \21706 , \28081 );
and \U$28485 ( \28863 , \21685 , \28079 );
nor \U$28486 ( \28864 , \28862 , \28863 );
xnor \U$28487 ( \28865 , \28864 , \27766 );
and \U$28488 ( \28866 , \28860 , \28865 );
and \U$28489 ( \28867 , \28856 , \28865 );
or \U$28490 ( \28868 , \28861 , \28866 , \28867 );
and \U$28491 ( \28869 , \28850 , \28868 );
and \U$28492 ( \28870 , \22046 , \26143 );
and \U$28493 ( \28871 , \22018 , \26141 );
nor \U$28494 ( \28872 , \28870 , \28871 );
xnor \U$28495 ( \28873 , \28872 , \25911 );
and \U$28496 ( \28874 , \22200 , \25692 );
and \U$28497 ( \28875 , \22126 , \25690 );
nor \U$28498 ( \28876 , \28874 , \28875 );
xnor \U$28499 ( \28877 , \28876 , \25549 );
and \U$28500 ( \28878 , \28873 , \28877 );
and \U$28501 ( \28879 , \22325 , \25369 );
and \U$28502 ( \28880 , \22262 , \25367 );
nor \U$28503 ( \28881 , \28879 , \28880 );
xnor \U$28504 ( \28882 , \28881 , \25123 );
and \U$28505 ( \28883 , \28877 , \28882 );
and \U$28506 ( \28884 , \28873 , \28882 );
or \U$28507 ( \28885 , \28878 , \28883 , \28884 );
and \U$28508 ( \28886 , \28868 , \28885 );
and \U$28509 ( \28887 , \28850 , \28885 );
or \U$28510 ( \28888 , \28869 , \28886 , \28887 );
and \U$28511 ( \28889 , \28834 , \28888 );
and \U$28512 ( \28890 , \25226 , \22497 );
and \U$28513 ( \28891 , \25018 , \22495 );
nor \U$28514 ( \28892 , \28890 , \28891 );
xnor \U$28515 ( \28893 , \28892 , \22419 );
and \U$28516 ( \28894 , \25353 , \22333 );
and \U$28517 ( \28895 , \25348 , \22331 );
nor \U$28518 ( \28896 , \28894 , \28895 );
xnor \U$28519 ( \28897 , \28896 , \22239 );
and \U$28520 ( \28898 , \28893 , \28897 );
and \U$28521 ( \28899 , \25806 , \22163 );
and \U$28522 ( \28900 , \25609 , \22161 );
nor \U$28523 ( \28901 , \28899 , \28900 );
xnor \U$28524 ( \28902 , \28901 , \22091 );
and \U$28525 ( \28903 , \28897 , \28902 );
and \U$28526 ( \28904 , \28893 , \28902 );
or \U$28527 ( \28905 , \28898 , \28903 , \28904 );
and \U$28528 ( \28906 , \26116 , \22029 );
and \U$28529 ( \28907 , \26108 , \22027 );
nor \U$28530 ( \28908 , \28906 , \28907 );
xnor \U$28531 ( \28909 , \28908 , \21986 );
and \U$28532 ( \28910 , \26590 , \21916 );
and \U$28533 ( \28911 , \26585 , \21914 );
nor \U$28534 ( \28912 , \28910 , \28911 );
xnor \U$28535 ( \28913 , \28912 , \21867 );
and \U$28536 ( \28914 , \28909 , \28913 );
and \U$28537 ( \28915 , \27113 , \21815 );
and \U$28538 ( \28916 , \26854 , \21813 );
nor \U$28539 ( \28917 , \28915 , \28916 );
xnor \U$28540 ( \28918 , \28917 , \21774 );
and \U$28541 ( \28919 , \28913 , \28918 );
and \U$28542 ( \28920 , \28909 , \28918 );
or \U$28543 ( \28921 , \28914 , \28919 , \28920 );
and \U$28544 ( \28922 , \28905 , \28921 );
and \U$28545 ( \28923 , \27494 , \21745 );
and \U$28546 ( \28924 , \27485 , \21743 );
nor \U$28547 ( \28925 , \28923 , \28924 );
xnor \U$28548 ( \28926 , \28925 , \21715 );
and \U$28549 ( \28927 , \28039 , \21697 );
and \U$28550 ( \28928 , \27837 , \21695 );
nor \U$28551 ( \28929 , \28927 , \28928 );
xnor \U$28552 ( \28930 , \28929 , \21678 );
and \U$28553 ( \28931 , \28926 , \28930 );
and \U$28554 ( \28932 , \28514 , \21660 );
and \U$28555 ( \28933 , \28342 , \21658 );
nor \U$28556 ( \28934 , \28932 , \28933 );
xnor \U$28557 ( \28935 , \28934 , \21665 );
and \U$28558 ( \28936 , \28930 , \28935 );
and \U$28559 ( \28937 , \28926 , \28935 );
or \U$28560 ( \28938 , \28931 , \28936 , \28937 );
and \U$28561 ( \28939 , \28921 , \28938 );
and \U$28562 ( \28940 , \28905 , \28938 );
or \U$28563 ( \28941 , \28922 , \28939 , \28940 );
and \U$28564 ( \28942 , \28888 , \28941 );
and \U$28565 ( \28943 , \28834 , \28941 );
or \U$28566 ( \28944 , \28889 , \28942 , \28943 );
and \U$28567 ( \28945 , \28782 , \28944 );
xor \U$28568 ( \28946 , \28651 , \28653 );
xor \U$28569 ( \28947 , \28946 , \28656 );
xor \U$28570 ( \28948 , \28661 , \28663 );
xor \U$28571 ( \28949 , \28948 , \28666 );
and \U$28572 ( \28950 , \28947 , \28949 );
xor \U$28573 ( \28951 , \28672 , \28674 );
xor \U$28574 ( \28952 , \28951 , \28677 );
and \U$28575 ( \28953 , \28949 , \28952 );
and \U$28576 ( \28954 , \28947 , \28952 );
or \U$28577 ( \28955 , \28950 , \28953 , \28954 );
and \U$28578 ( \28956 , \28944 , \28955 );
and \U$28579 ( \28957 , \28782 , \28955 );
or \U$28580 ( \28958 , \28945 , \28956 , \28957 );
xor \U$28581 ( \28959 , \28504 , \28518 );
xor \U$28582 ( \28960 , \28959 , \28535 );
xor \U$28583 ( \28961 , \28554 , \28570 );
xor \U$28584 ( \28962 , \28961 , \28590 );
and \U$28585 ( \28963 , \28960 , \28962 );
xor \U$28586 ( \28964 , \28610 , \28626 );
xor \U$28587 ( \28965 , \28964 , \28643 );
and \U$28588 ( \28966 , \28962 , \28965 );
and \U$28589 ( \28967 , \28960 , \28965 );
or \U$28590 ( \28968 , \28963 , \28966 , \28967 );
xor \U$28591 ( \28969 , \28699 , \28701 );
xor \U$28592 ( \28970 , \28969 , \28704 );
and \U$28593 ( \28971 , \28968 , \28970 );
xor \U$28594 ( \28972 , \28686 , \28688 );
xor \U$28595 ( \28973 , \28972 , \28691 );
and \U$28596 ( \28974 , \28970 , \28973 );
and \U$28597 ( \28975 , \28968 , \28973 );
or \U$28598 ( \28976 , \28971 , \28974 , \28975 );
and \U$28599 ( \28977 , \28958 , \28976 );
xor \U$28600 ( \28978 , \28538 , \28593 );
xor \U$28601 ( \28979 , \28978 , \28646 );
xor \U$28602 ( \28980 , \28659 , \28669 );
xor \U$28603 ( \28981 , \28980 , \28680 );
and \U$28604 ( \28982 , \28979 , \28981 );
and \U$28605 ( \28983 , \28976 , \28982 );
and \U$28606 ( \28984 , \28958 , \28982 );
or \U$28607 ( \28985 , \28977 , \28983 , \28984 );
xor \U$28608 ( \28986 , \28649 , \28683 );
xor \U$28609 ( \28987 , \28986 , \28694 );
xor \U$28610 ( \28988 , \28707 , \28709 );
xor \U$28611 ( \28989 , \28988 , \28712 );
and \U$28612 ( \28990 , \28987 , \28989 );
xor \U$28613 ( \28991 , \28718 , \28720 );
and \U$28614 ( \28992 , \28989 , \28991 );
and \U$28615 ( \28993 , \28987 , \28991 );
or \U$28616 ( \28994 , \28990 , \28992 , \28993 );
and \U$28617 ( \28995 , \28985 , \28994 );
xor \U$28618 ( \28996 , \28726 , \28728 );
xor \U$28619 ( \28997 , \28996 , \28730 );
and \U$28620 ( \28998 , \28994 , \28997 );
and \U$28621 ( \28999 , \28985 , \28997 );
or \U$28622 ( \29000 , \28995 , \28998 , \28999 );
xor \U$28623 ( \29001 , \28432 , \28450 );
xor \U$28624 ( \29002 , \29001 , \28456 );
and \U$28625 ( \29003 , \29000 , \29002 );
xor \U$28626 ( \29004 , \28724 , \28733 );
xor \U$28627 ( \29005 , \29004 , \28736 );
and \U$28628 ( \29006 , \29002 , \29005 );
and \U$28629 ( \29007 , \29000 , \29005 );
or \U$28630 ( \29008 , \29003 , \29006 , \29007 );
xor \U$28631 ( \29009 , \28739 , \28741 );
xor \U$28632 ( \29010 , \29009 , \28744 );
and \U$28633 ( \29011 , \29008 , \29010 );
and \U$28634 ( \29012 , \28753 , \29011 );
xor \U$28635 ( \29013 , \28753 , \29011 );
xor \U$28636 ( \29014 , \29008 , \29010 );
and \U$28637 ( \29015 , \25348 , \22497 );
and \U$28638 ( \29016 , \25226 , \22495 );
nor \U$28639 ( \29017 , \29015 , \29016 );
xnor \U$28640 ( \29018 , \29017 , \22419 );
and \U$28641 ( \29019 , \25609 , \22333 );
and \U$28642 ( \29020 , \25353 , \22331 );
nor \U$28643 ( \29021 , \29019 , \29020 );
xnor \U$28644 ( \29022 , \29021 , \22239 );
and \U$28645 ( \29023 , \29018 , \29022 );
and \U$28646 ( \29024 , \26108 , \22163 );
and \U$28647 ( \29025 , \25806 , \22161 );
nor \U$28648 ( \29026 , \29024 , \29025 );
xnor \U$28649 ( \29027 , \29026 , \22091 );
and \U$28650 ( \29028 , \29022 , \29027 );
and \U$28651 ( \29029 , \29018 , \29027 );
or \U$28652 ( \29030 , \29023 , \29028 , \29029 );
and \U$28653 ( \29031 , \27837 , \21745 );
and \U$28654 ( \29032 , \27494 , \21743 );
nor \U$28655 ( \29033 , \29031 , \29032 );
xnor \U$28656 ( \29034 , \29033 , \21715 );
and \U$28657 ( \29035 , \28342 , \21697 );
and \U$28658 ( \29036 , \28039 , \21695 );
nor \U$28659 ( \29037 , \29035 , \29036 );
xnor \U$28660 ( \29038 , \29037 , \21678 );
and \U$28661 ( \29039 , \29034 , \29038 );
buf \U$28662 ( \29040 , RIc22adf0_181);
and \U$28663 ( \29041 , \29040 , \21660 );
and \U$28664 ( \29042 , \28514 , \21658 );
nor \U$28665 ( \29043 , \29041 , \29042 );
xnor \U$28666 ( \29044 , \29043 , \21665 );
and \U$28667 ( \29045 , \29038 , \29044 );
and \U$28668 ( \29046 , \29034 , \29044 );
or \U$28669 ( \29047 , \29039 , \29045 , \29046 );
and \U$28670 ( \29048 , \29030 , \29047 );
and \U$28671 ( \29049 , \26585 , \22029 );
and \U$28672 ( \29050 , \26116 , \22027 );
nor \U$28673 ( \29051 , \29049 , \29050 );
xnor \U$28674 ( \29052 , \29051 , \21986 );
and \U$28675 ( \29053 , \26854 , \21916 );
and \U$28676 ( \29054 , \26590 , \21914 );
nor \U$28677 ( \29055 , \29053 , \29054 );
xnor \U$28678 ( \29056 , \29055 , \21867 );
and \U$28679 ( \29057 , \29052 , \29056 );
and \U$28680 ( \29058 , \27485 , \21815 );
and \U$28681 ( \29059 , \27113 , \21813 );
nor \U$28682 ( \29060 , \29058 , \29059 );
xnor \U$28683 ( \29061 , \29060 , \21774 );
and \U$28684 ( \29062 , \29056 , \29061 );
and \U$28685 ( \29063 , \29052 , \29061 );
or \U$28686 ( \29064 , \29057 , \29062 , \29063 );
and \U$28687 ( \29065 , \29047 , \29064 );
and \U$28688 ( \29066 , \29030 , \29064 );
or \U$28689 ( \29067 , \29048 , \29065 , \29066 );
and \U$28690 ( \29068 , \21831 , \27572 );
and \U$28691 ( \29069 , \21762 , \27570 );
nor \U$28692 ( \29070 , \29068 , \29069 );
xnor \U$28693 ( \29071 , \29070 , \27232 );
and \U$28694 ( \29072 , \21890 , \26983 );
and \U$28695 ( \29073 , \21836 , \26981 );
nor \U$28696 ( \29074 , \29072 , \29073 );
xnor \U$28697 ( \29075 , \29074 , \26742 );
and \U$28698 ( \29076 , \29071 , \29075 );
and \U$28699 ( \29077 , \22018 , \26517 );
and \U$28700 ( \29078 , \21941 , \26515 );
nor \U$28701 ( \29079 , \29077 , \29078 );
xnor \U$28702 ( \29080 , \29079 , \26329 );
and \U$28703 ( \29081 , \29075 , \29080 );
and \U$28704 ( \29082 , \29071 , \29080 );
or \U$28705 ( \29083 , \29076 , \29081 , \29082 );
and \U$28706 ( \29084 , \22126 , \26143 );
and \U$28707 ( \29085 , \22046 , \26141 );
nor \U$28708 ( \29086 , \29084 , \29085 );
xnor \U$28709 ( \29087 , \29086 , \25911 );
and \U$28710 ( \29088 , \22262 , \25692 );
and \U$28711 ( \29089 , \22200 , \25690 );
nor \U$28712 ( \29090 , \29088 , \29089 );
xnor \U$28713 ( \29091 , \29090 , \25549 );
and \U$28714 ( \29092 , \29087 , \29091 );
and \U$28715 ( \29093 , \22523 , \25369 );
and \U$28716 ( \29094 , \22325 , \25367 );
nor \U$28717 ( \29095 , \29093 , \29094 );
xnor \U$28718 ( \29096 , \29095 , \25123 );
and \U$28719 ( \29097 , \29091 , \29096 );
and \U$28720 ( \29098 , \29087 , \29096 );
or \U$28721 ( \29099 , \29092 , \29097 , \29098 );
and \U$28722 ( \29100 , \29083 , \29099 );
xor \U$28723 ( \29101 , \28312 , \28851 );
xor \U$28724 ( \29102 , \28851 , \28852 );
not \U$28725 ( \29103 , \29102 );
and \U$28726 ( \29104 , \29101 , \29103 );
and \U$28727 ( \29105 , \21653 , \29104 );
not \U$28728 ( \29106 , \29105 );
xnor \U$28729 ( \29107 , \29106 , \28855 );
and \U$28730 ( \29108 , \21685 , \28575 );
and \U$28731 ( \29109 , \21667 , \28573 );
nor \U$28732 ( \29110 , \29108 , \29109 );
xnor \U$28733 ( \29111 , \29110 , \28315 );
and \U$28734 ( \29112 , \29107 , \29111 );
and \U$28735 ( \29113 , \21754 , \28081 );
and \U$28736 ( \29114 , \21706 , \28079 );
nor \U$28737 ( \29115 , \29113 , \29114 );
xnor \U$28738 ( \29116 , \29115 , \27766 );
and \U$28739 ( \29117 , \29111 , \29116 );
and \U$28740 ( \29118 , \29107 , \29116 );
or \U$28741 ( \29119 , \29112 , \29117 , \29118 );
and \U$28742 ( \29120 , \29099 , \29119 );
and \U$28743 ( \29121 , \29083 , \29119 );
or \U$28744 ( \29122 , \29100 , \29120 , \29121 );
and \U$28745 ( \29123 , \29067 , \29122 );
and \U$28746 ( \29124 , \24177 , \23163 );
and \U$28747 ( \29125 , \24003 , \23161 );
nor \U$28748 ( \29126 , \29124 , \29125 );
xnor \U$28749 ( \29127 , \29126 , \23007 );
and \U$28750 ( \29128 , \24482 , \22891 );
and \U$28751 ( \29129 , \24344 , \22889 );
nor \U$28752 ( \29130 , \29128 , \29129 );
xnor \U$28753 ( \29131 , \29130 , \22778 );
and \U$28754 ( \29132 , \29127 , \29131 );
and \U$28755 ( \29133 , \25018 , \22697 );
and \U$28756 ( \29134 , \24601 , \22695 );
nor \U$28757 ( \29135 , \29133 , \29134 );
xnor \U$28758 ( \29136 , \29135 , \22561 );
and \U$28759 ( \29137 , \29131 , \29136 );
and \U$28760 ( \29138 , \29127 , \29136 );
or \U$28761 ( \29139 , \29132 , \29137 , \29138 );
and \U$28762 ( \29140 , \22716 , \24974 );
and \U$28763 ( \29141 , \22611 , \24972 );
nor \U$28764 ( \29142 , \29140 , \29141 );
xnor \U$28765 ( \29143 , \29142 , \24787 );
and \U$28766 ( \29144 , \22837 , \24661 );
and \U$28767 ( \29145 , \22721 , \24659 );
nor \U$28768 ( \29146 , \29144 , \29145 );
xnor \U$28769 ( \29147 , \29146 , \24456 );
and \U$28770 ( \29148 , \29143 , \29147 );
and \U$28771 ( \29149 , \23128 , \24255 );
and \U$28772 ( \29150 , \22952 , \24253 );
nor \U$28773 ( \29151 , \29149 , \29150 );
xnor \U$28774 ( \29152 , \29151 , \24106 );
and \U$28775 ( \29153 , \29147 , \29152 );
and \U$28776 ( \29154 , \29143 , \29152 );
or \U$28777 ( \29155 , \29148 , \29153 , \29154 );
and \U$28778 ( \29156 , \29139 , \29155 );
and \U$28779 ( \29157 , \23379 , \23933 );
and \U$28780 ( \29158 , \23136 , \23931 );
nor \U$28781 ( \29159 , \29157 , \29158 );
xnor \U$28782 ( \29160 , \29159 , \23791 );
and \U$28783 ( \29161 , \23570 , \23637 );
and \U$28784 ( \29162 , \23384 , \23635 );
nor \U$28785 ( \29163 , \29161 , \29162 );
xnor \U$28786 ( \29164 , \29163 , \23500 );
and \U$28787 ( \29165 , \29160 , \29164 );
and \U$28788 ( \29166 , \23978 , \23431 );
and \U$28789 ( \29167 , \23714 , \23429 );
nor \U$28790 ( \29168 , \29166 , \29167 );
xnor \U$28791 ( \29169 , \29168 , \23279 );
and \U$28792 ( \29170 , \29164 , \29169 );
and \U$28793 ( \29171 , \29160 , \29169 );
or \U$28794 ( \29172 , \29165 , \29170 , \29171 );
and \U$28795 ( \29173 , \29155 , \29172 );
and \U$28796 ( \29174 , \29139 , \29172 );
or \U$28797 ( \29175 , \29156 , \29173 , \29174 );
and \U$28798 ( \29176 , \29122 , \29175 );
and \U$28799 ( \29177 , \29067 , \29175 );
or \U$28800 ( \29178 , \29123 , \29176 , \29177 );
xor \U$28801 ( \29179 , \28838 , \28842 );
xor \U$28802 ( \29180 , \29179 , \28847 );
xor \U$28803 ( \29181 , \28802 , \28806 );
xor \U$28804 ( \29182 , \29181 , \28811 );
and \U$28805 ( \29183 , \29180 , \29182 );
xor \U$28806 ( \29184 , \28873 , \28877 );
xor \U$28807 ( \29185 , \29184 , \28882 );
and \U$28808 ( \29186 , \29182 , \29185 );
and \U$28809 ( \29187 , \29180 , \29185 );
or \U$28810 ( \29188 , \29183 , \29186 , \29187 );
and \U$28811 ( \29189 , \29040 , \21654 );
xor \U$28812 ( \29190 , \28909 , \28913 );
xor \U$28813 ( \29191 , \29190 , \28918 );
and \U$28814 ( \29192 , \29189 , \29191 );
xor \U$28815 ( \29193 , \28926 , \28930 );
xor \U$28816 ( \29194 , \29193 , \28935 );
and \U$28817 ( \29195 , \29191 , \29194 );
and \U$28818 ( \29196 , \29189 , \29194 );
or \U$28819 ( \29197 , \29192 , \29195 , \29196 );
and \U$28820 ( \29198 , \29188 , \29197 );
xor \U$28821 ( \29199 , \28893 , \28897 );
xor \U$28822 ( \29200 , \29199 , \28902 );
xor \U$28823 ( \29201 , \28786 , \28790 );
xor \U$28824 ( \29202 , \29201 , \28795 );
and \U$28825 ( \29203 , \29200 , \29202 );
xor \U$28826 ( \29204 , \28819 , \28823 );
xor \U$28827 ( \29205 , \29204 , \28828 );
and \U$28828 ( \29206 , \29202 , \29205 );
and \U$28829 ( \29207 , \29200 , \29205 );
or \U$28830 ( \29208 , \29203 , \29206 , \29207 );
and \U$28831 ( \29209 , \29197 , \29208 );
and \U$28832 ( \29210 , \29188 , \29208 );
or \U$28833 ( \29211 , \29198 , \29209 , \29210 );
and \U$28834 ( \29212 , \29178 , \29211 );
xor \U$28835 ( \29213 , \28578 , \28582 );
xor \U$28836 ( \29214 , \29213 , \28587 );
xor \U$28837 ( \29215 , \28755 , \28757 );
xor \U$28838 ( \29216 , \29215 , \28760 );
and \U$28839 ( \29217 , \29214 , \29216 );
xor \U$28840 ( \29218 , \28765 , \28767 );
xor \U$28841 ( \29219 , \29218 , \28770 );
and \U$28842 ( \29220 , \29216 , \29219 );
and \U$28843 ( \29221 , \29214 , \29219 );
or \U$28844 ( \29222 , \29217 , \29220 , \29221 );
and \U$28845 ( \29223 , \29211 , \29222 );
and \U$28846 ( \29224 , \29178 , \29222 );
or \U$28847 ( \29225 , \29212 , \29223 , \29224 );
xor \U$28848 ( \29226 , \28798 , \28814 );
xor \U$28849 ( \29227 , \29226 , \28831 );
xor \U$28850 ( \29228 , \28905 , \28921 );
xor \U$28851 ( \29229 , \29228 , \28938 );
and \U$28852 ( \29230 , \29227 , \29229 );
xnor \U$28853 ( \29231 , \28776 , \28778 );
and \U$28854 ( \29232 , \29229 , \29231 );
and \U$28855 ( \29233 , \29227 , \29231 );
or \U$28856 ( \29234 , \29230 , \29232 , \29233 );
xor \U$28857 ( \29235 , \28960 , \28962 );
xor \U$28858 ( \29236 , \29235 , \28965 );
and \U$28859 ( \29237 , \29234 , \29236 );
xor \U$28860 ( \29238 , \28947 , \28949 );
xor \U$28861 ( \29239 , \29238 , \28952 );
and \U$28862 ( \29240 , \29236 , \29239 );
and \U$28863 ( \29241 , \29234 , \29239 );
or \U$28864 ( \29242 , \29237 , \29240 , \29241 );
and \U$28865 ( \29243 , \29225 , \29242 );
xor \U$28866 ( \29244 , \28763 , \28773 );
xor \U$28867 ( \29245 , \29244 , \28779 );
xor \U$28868 ( \29246 , \28834 , \28888 );
xor \U$28869 ( \29247 , \29246 , \28941 );
and \U$28870 ( \29248 , \29245 , \29247 );
and \U$28871 ( \29249 , \29242 , \29248 );
and \U$28872 ( \29250 , \29225 , \29248 );
or \U$28873 ( \29251 , \29243 , \29249 , \29250 );
xor \U$28874 ( \29252 , \28782 , \28944 );
xor \U$28875 ( \29253 , \29252 , \28955 );
xor \U$28876 ( \29254 , \28968 , \28970 );
xor \U$28877 ( \29255 , \29254 , \28973 );
and \U$28878 ( \29256 , \29253 , \29255 );
xor \U$28879 ( \29257 , \28979 , \28981 );
and \U$28880 ( \29258 , \29255 , \29257 );
and \U$28881 ( \29259 , \29253 , \29257 );
or \U$28882 ( \29260 , \29256 , \29258 , \29259 );
and \U$28883 ( \29261 , \29251 , \29260 );
xor \U$28884 ( \29262 , \28987 , \28989 );
xor \U$28885 ( \29263 , \29262 , \28991 );
and \U$28886 ( \29264 , \29260 , \29263 );
and \U$28887 ( \29265 , \29251 , \29263 );
or \U$28888 ( \29266 , \29261 , \29264 , \29265 );
xor \U$28889 ( \29267 , \28697 , \28715 );
xor \U$28890 ( \29268 , \29267 , \28721 );
and \U$28891 ( \29269 , \29266 , \29268 );
xor \U$28892 ( \29270 , \28985 , \28994 );
xor \U$28893 ( \29271 , \29270 , \28997 );
and \U$28894 ( \29272 , \29268 , \29271 );
and \U$28895 ( \29273 , \29266 , \29271 );
or \U$28896 ( \29274 , \29269 , \29272 , \29273 );
xor \U$28897 ( \29275 , \29000 , \29002 );
xor \U$28898 ( \29276 , \29275 , \29005 );
and \U$28899 ( \29277 , \29274 , \29276 );
and \U$28900 ( \29278 , \29014 , \29277 );
xor \U$28901 ( \29279 , \29014 , \29277 );
xor \U$28902 ( \29280 , \29274 , \29276 );
and \U$28903 ( \29281 , \24003 , \23431 );
and \U$28904 ( \29282 , \23978 , \23429 );
nor \U$28905 ( \29283 , \29281 , \29282 );
xnor \U$28906 ( \29284 , \29283 , \23279 );
and \U$28907 ( \29285 , \24344 , \23163 );
and \U$28908 ( \29286 , \24177 , \23161 );
nor \U$28909 ( \29287 , \29285 , \29286 );
xnor \U$28910 ( \29288 , \29287 , \23007 );
and \U$28911 ( \29289 , \29284 , \29288 );
and \U$28912 ( \29290 , \24601 , \22891 );
and \U$28913 ( \29291 , \24482 , \22889 );
nor \U$28914 ( \29292 , \29290 , \29291 );
xnor \U$28915 ( \29293 , \29292 , \22778 );
and \U$28916 ( \29294 , \29288 , \29293 );
and \U$28917 ( \29295 , \29284 , \29293 );
or \U$28918 ( \29296 , \29289 , \29294 , \29295 );
and \U$28919 ( \29297 , \22611 , \25369 );
and \U$28920 ( \29298 , \22523 , \25367 );
nor \U$28921 ( \29299 , \29297 , \29298 );
xnor \U$28922 ( \29300 , \29299 , \25123 );
and \U$28923 ( \29301 , \22721 , \24974 );
and \U$28924 ( \29302 , \22716 , \24972 );
nor \U$28925 ( \29303 , \29301 , \29302 );
xnor \U$28926 ( \29304 , \29303 , \24787 );
and \U$28927 ( \29305 , \29300 , \29304 );
and \U$28928 ( \29306 , \22952 , \24661 );
and \U$28929 ( \29307 , \22837 , \24659 );
nor \U$28930 ( \29308 , \29306 , \29307 );
xnor \U$28931 ( \29309 , \29308 , \24456 );
and \U$28932 ( \29310 , \29304 , \29309 );
and \U$28933 ( \29311 , \29300 , \29309 );
or \U$28934 ( \29312 , \29305 , \29310 , \29311 );
and \U$28935 ( \29313 , \29296 , \29312 );
and \U$28936 ( \29314 , \23136 , \24255 );
and \U$28937 ( \29315 , \23128 , \24253 );
nor \U$28938 ( \29316 , \29314 , \29315 );
xnor \U$28939 ( \29317 , \29316 , \24106 );
and \U$28940 ( \29318 , \23384 , \23933 );
and \U$28941 ( \29319 , \23379 , \23931 );
nor \U$28942 ( \29320 , \29318 , \29319 );
xnor \U$28943 ( \29321 , \29320 , \23791 );
and \U$28944 ( \29322 , \29317 , \29321 );
and \U$28945 ( \29323 , \23714 , \23637 );
and \U$28946 ( \29324 , \23570 , \23635 );
nor \U$28947 ( \29325 , \29323 , \29324 );
xnor \U$28948 ( \29326 , \29325 , \23500 );
and \U$28949 ( \29327 , \29321 , \29326 );
and \U$28950 ( \29328 , \29317 , \29326 );
or \U$28951 ( \29329 , \29322 , \29327 , \29328 );
and \U$28952 ( \29330 , \29312 , \29329 );
and \U$28953 ( \29331 , \29296 , \29329 );
or \U$28954 ( \29332 , \29313 , \29330 , \29331 );
and \U$28955 ( \29333 , \22046 , \26517 );
and \U$28956 ( \29334 , \22018 , \26515 );
nor \U$28957 ( \29335 , \29333 , \29334 );
xnor \U$28958 ( \29336 , \29335 , \26329 );
and \U$28959 ( \29337 , \22200 , \26143 );
and \U$28960 ( \29338 , \22126 , \26141 );
nor \U$28961 ( \29339 , \29337 , \29338 );
xnor \U$28962 ( \29340 , \29339 , \25911 );
and \U$28963 ( \29341 , \29336 , \29340 );
and \U$28964 ( \29342 , \22325 , \25692 );
and \U$28965 ( \29343 , \22262 , \25690 );
nor \U$28966 ( \29344 , \29342 , \29343 );
xnor \U$28967 ( \29345 , \29344 , \25549 );
and \U$28968 ( \29346 , \29340 , \29345 );
and \U$28969 ( \29347 , \29336 , \29345 );
or \U$28970 ( \29348 , \29341 , \29346 , \29347 );
buf \U$28971 ( \29349 , RIc225be8_56);
buf \U$28972 ( \29350 , RIc225b70_57);
and \U$28973 ( \29351 , \29349 , \29350 );
not \U$28974 ( \29352 , \29351 );
and \U$28975 ( \29353 , \28852 , \29352 );
not \U$28976 ( \29354 , \29353 );
and \U$28977 ( \29355 , \21667 , \29104 );
and \U$28978 ( \29356 , \21653 , \29102 );
nor \U$28979 ( \29357 , \29355 , \29356 );
xnor \U$28980 ( \29358 , \29357 , \28855 );
and \U$28981 ( \29359 , \29354 , \29358 );
and \U$28982 ( \29360 , \21706 , \28575 );
and \U$28983 ( \29361 , \21685 , \28573 );
nor \U$28984 ( \29362 , \29360 , \29361 );
xnor \U$28985 ( \29363 , \29362 , \28315 );
and \U$28986 ( \29364 , \29358 , \29363 );
and \U$28987 ( \29365 , \29354 , \29363 );
or \U$28988 ( \29366 , \29359 , \29364 , \29365 );
and \U$28989 ( \29367 , \29348 , \29366 );
and \U$28990 ( \29368 , \21762 , \28081 );
and \U$28991 ( \29369 , \21754 , \28079 );
nor \U$28992 ( \29370 , \29368 , \29369 );
xnor \U$28993 ( \29371 , \29370 , \27766 );
and \U$28994 ( \29372 , \21836 , \27572 );
and \U$28995 ( \29373 , \21831 , \27570 );
nor \U$28996 ( \29374 , \29372 , \29373 );
xnor \U$28997 ( \29375 , \29374 , \27232 );
and \U$28998 ( \29376 , \29371 , \29375 );
and \U$28999 ( \29377 , \21941 , \26983 );
and \U$29000 ( \29378 , \21890 , \26981 );
nor \U$29001 ( \29379 , \29377 , \29378 );
xnor \U$29002 ( \29380 , \29379 , \26742 );
and \U$29003 ( \29381 , \29375 , \29380 );
and \U$29004 ( \29382 , \29371 , \29380 );
or \U$29005 ( \29383 , \29376 , \29381 , \29382 );
and \U$29006 ( \29384 , \29366 , \29383 );
and \U$29007 ( \29385 , \29348 , \29383 );
or \U$29008 ( \29386 , \29367 , \29384 , \29385 );
and \U$29009 ( \29387 , \29332 , \29386 );
and \U$29010 ( \29388 , \26116 , \22163 );
and \U$29011 ( \29389 , \26108 , \22161 );
nor \U$29012 ( \29390 , \29388 , \29389 );
xnor \U$29013 ( \29391 , \29390 , \22091 );
and \U$29014 ( \29392 , \26590 , \22029 );
and \U$29015 ( \29393 , \26585 , \22027 );
nor \U$29016 ( \29394 , \29392 , \29393 );
xnor \U$29017 ( \29395 , \29394 , \21986 );
and \U$29018 ( \29396 , \29391 , \29395 );
and \U$29019 ( \29397 , \27113 , \21916 );
and \U$29020 ( \29398 , \26854 , \21914 );
nor \U$29021 ( \29399 , \29397 , \29398 );
xnor \U$29022 ( \29400 , \29399 , \21867 );
and \U$29023 ( \29401 , \29395 , \29400 );
and \U$29024 ( \29402 , \29391 , \29400 );
or \U$29025 ( \29403 , \29396 , \29401 , \29402 );
and \U$29026 ( \29404 , \27494 , \21815 );
and \U$29027 ( \29405 , \27485 , \21813 );
nor \U$29028 ( \29406 , \29404 , \29405 );
xnor \U$29029 ( \29407 , \29406 , \21774 );
and \U$29030 ( \29408 , \28039 , \21745 );
and \U$29031 ( \29409 , \27837 , \21743 );
nor \U$29032 ( \29410 , \29408 , \29409 );
xnor \U$29033 ( \29411 , \29410 , \21715 );
and \U$29034 ( \29412 , \29407 , \29411 );
and \U$29035 ( \29413 , \28514 , \21697 );
and \U$29036 ( \29414 , \28342 , \21695 );
nor \U$29037 ( \29415 , \29413 , \29414 );
xnor \U$29038 ( \29416 , \29415 , \21678 );
and \U$29039 ( \29417 , \29411 , \29416 );
and \U$29040 ( \29418 , \29407 , \29416 );
or \U$29041 ( \29419 , \29412 , \29417 , \29418 );
and \U$29042 ( \29420 , \29403 , \29419 );
and \U$29043 ( \29421 , \25226 , \22697 );
and \U$29044 ( \29422 , \25018 , \22695 );
nor \U$29045 ( \29423 , \29421 , \29422 );
xnor \U$29046 ( \29424 , \29423 , \22561 );
and \U$29047 ( \29425 , \25353 , \22497 );
and \U$29048 ( \29426 , \25348 , \22495 );
nor \U$29049 ( \29427 , \29425 , \29426 );
xnor \U$29050 ( \29428 , \29427 , \22419 );
and \U$29051 ( \29429 , \29424 , \29428 );
and \U$29052 ( \29430 , \25806 , \22333 );
and \U$29053 ( \29431 , \25609 , \22331 );
nor \U$29054 ( \29432 , \29430 , \29431 );
xnor \U$29055 ( \29433 , \29432 , \22239 );
and \U$29056 ( \29434 , \29428 , \29433 );
and \U$29057 ( \29435 , \29424 , \29433 );
or \U$29058 ( \29436 , \29429 , \29434 , \29435 );
and \U$29059 ( \29437 , \29419 , \29436 );
and \U$29060 ( \29438 , \29403 , \29436 );
or \U$29061 ( \29439 , \29420 , \29437 , \29438 );
and \U$29062 ( \29440 , \29386 , \29439 );
and \U$29063 ( \29441 , \29332 , \29439 );
or \U$29064 ( \29442 , \29387 , \29440 , \29441 );
xor \U$29065 ( \29443 , \29018 , \29022 );
xor \U$29066 ( \29444 , \29443 , \29027 );
xor \U$29067 ( \29445 , \29127 , \29131 );
xor \U$29068 ( \29446 , \29445 , \29136 );
and \U$29069 ( \29447 , \29444 , \29446 );
xor \U$29070 ( \29448 , \29052 , \29056 );
xor \U$29071 ( \29449 , \29448 , \29061 );
and \U$29072 ( \29450 , \29446 , \29449 );
and \U$29073 ( \29451 , \29444 , \29449 );
or \U$29074 ( \29452 , \29447 , \29450 , \29451 );
xor \U$29075 ( \29453 , \29087 , \29091 );
xor \U$29076 ( \29454 , \29453 , \29096 );
xor \U$29077 ( \29455 , \29143 , \29147 );
xor \U$29078 ( \29456 , \29455 , \29152 );
and \U$29079 ( \29457 , \29454 , \29456 );
xor \U$29080 ( \29458 , \29160 , \29164 );
xor \U$29081 ( \29459 , \29458 , \29169 );
and \U$29082 ( \29460 , \29456 , \29459 );
and \U$29083 ( \29461 , \29454 , \29459 );
or \U$29084 ( \29462 , \29457 , \29460 , \29461 );
and \U$29085 ( \29463 , \29452 , \29462 );
buf \U$29086 ( \29464 , RIc22ae68_182);
and \U$29087 ( \29465 , \29464 , \21654 );
xor \U$29088 ( \29466 , \29034 , \29038 );
xor \U$29089 ( \29467 , \29466 , \29044 );
or \U$29090 ( \29468 , \29465 , \29467 );
and \U$29091 ( \29469 , \29462 , \29468 );
and \U$29092 ( \29470 , \29452 , \29468 );
or \U$29093 ( \29471 , \29463 , \29469 , \29470 );
and \U$29094 ( \29472 , \29442 , \29471 );
xor \U$29095 ( \29473 , \28856 , \28860 );
xor \U$29096 ( \29474 , \29473 , \28865 );
xor \U$29097 ( \29475 , \29180 , \29182 );
xor \U$29098 ( \29476 , \29475 , \29185 );
and \U$29099 ( \29477 , \29474 , \29476 );
xor \U$29100 ( \29478 , \29200 , \29202 );
xor \U$29101 ( \29479 , \29478 , \29205 );
and \U$29102 ( \29480 , \29476 , \29479 );
and \U$29103 ( \29481 , \29474 , \29479 );
or \U$29104 ( \29482 , \29477 , \29480 , \29481 );
and \U$29105 ( \29483 , \29471 , \29482 );
and \U$29106 ( \29484 , \29442 , \29482 );
or \U$29107 ( \29485 , \29472 , \29483 , \29484 );
xor \U$29108 ( \29486 , \29067 , \29122 );
xor \U$29109 ( \29487 , \29486 , \29175 );
xor \U$29110 ( \29488 , \29188 , \29197 );
xor \U$29111 ( \29489 , \29488 , \29208 );
and \U$29112 ( \29490 , \29487 , \29489 );
xor \U$29113 ( \29491 , \29214 , \29216 );
xor \U$29114 ( \29492 , \29491 , \29219 );
and \U$29115 ( \29493 , \29489 , \29492 );
and \U$29116 ( \29494 , \29487 , \29492 );
or \U$29117 ( \29495 , \29490 , \29493 , \29494 );
and \U$29118 ( \29496 , \29485 , \29495 );
xor \U$29119 ( \29497 , \29030 , \29047 );
xor \U$29120 ( \29498 , \29497 , \29064 );
xor \U$29121 ( \29499 , \29139 , \29155 );
xor \U$29122 ( \29500 , \29499 , \29172 );
and \U$29123 ( \29501 , \29498 , \29500 );
xor \U$29124 ( \29502 , \29189 , \29191 );
xor \U$29125 ( \29503 , \29502 , \29194 );
and \U$29126 ( \29504 , \29500 , \29503 );
and \U$29127 ( \29505 , \29498 , \29503 );
or \U$29128 ( \29506 , \29501 , \29504 , \29505 );
xor \U$29129 ( \29507 , \28850 , \28868 );
xor \U$29130 ( \29508 , \29507 , \28885 );
and \U$29131 ( \29509 , \29506 , \29508 );
xor \U$29132 ( \29510 , \29227 , \29229 );
xor \U$29133 ( \29511 , \29510 , \29231 );
and \U$29134 ( \29512 , \29508 , \29511 );
and \U$29135 ( \29513 , \29506 , \29511 );
or \U$29136 ( \29514 , \29509 , \29512 , \29513 );
and \U$29137 ( \29515 , \29495 , \29514 );
and \U$29138 ( \29516 , \29485 , \29514 );
or \U$29139 ( \29517 , \29496 , \29515 , \29516 );
xor \U$29140 ( \29518 , \29178 , \29211 );
xor \U$29141 ( \29519 , \29518 , \29222 );
xor \U$29142 ( \29520 , \29234 , \29236 );
xor \U$29143 ( \29521 , \29520 , \29239 );
and \U$29144 ( \29522 , \29519 , \29521 );
xor \U$29145 ( \29523 , \29245 , \29247 );
and \U$29146 ( \29524 , \29521 , \29523 );
and \U$29147 ( \29525 , \29519 , \29523 );
or \U$29148 ( \29526 , \29522 , \29524 , \29525 );
and \U$29149 ( \29527 , \29517 , \29526 );
xor \U$29150 ( \29528 , \29253 , \29255 );
xor \U$29151 ( \29529 , \29528 , \29257 );
and \U$29152 ( \29530 , \29526 , \29529 );
and \U$29153 ( \29531 , \29517 , \29529 );
or \U$29154 ( \29532 , \29527 , \29530 , \29531 );
xor \U$29155 ( \29533 , \28958 , \28976 );
xor \U$29156 ( \29534 , \29533 , \28982 );
and \U$29157 ( \29535 , \29532 , \29534 );
xor \U$29158 ( \29536 , \29251 , \29260 );
xor \U$29159 ( \29537 , \29536 , \29263 );
and \U$29160 ( \29538 , \29534 , \29537 );
and \U$29161 ( \29539 , \29532 , \29537 );
or \U$29162 ( \29540 , \29535 , \29538 , \29539 );
xor \U$29163 ( \29541 , \29266 , \29268 );
xor \U$29164 ( \29542 , \29541 , \29271 );
and \U$29165 ( \29543 , \29540 , \29542 );
and \U$29166 ( \29544 , \29280 , \29543 );
xor \U$29167 ( \29545 , \29280 , \29543 );
xor \U$29168 ( \29546 , \29540 , \29542 );
and \U$29169 ( \29547 , \23379 , \24255 );
and \U$29170 ( \29548 , \23136 , \24253 );
nor \U$29171 ( \29549 , \29547 , \29548 );
xnor \U$29172 ( \29550 , \29549 , \24106 );
and \U$29173 ( \29551 , \23570 , \23933 );
and \U$29174 ( \29552 , \23384 , \23931 );
nor \U$29175 ( \29553 , \29551 , \29552 );
xnor \U$29176 ( \29554 , \29553 , \23791 );
and \U$29177 ( \29555 , \29550 , \29554 );
and \U$29178 ( \29556 , \23978 , \23637 );
and \U$29179 ( \29557 , \23714 , \23635 );
nor \U$29180 ( \29558 , \29556 , \29557 );
xnor \U$29181 ( \29559 , \29558 , \23500 );
and \U$29182 ( \29560 , \29554 , \29559 );
and \U$29183 ( \29561 , \29550 , \29559 );
or \U$29184 ( \29562 , \29555 , \29560 , \29561 );
and \U$29185 ( \29563 , \24177 , \23431 );
and \U$29186 ( \29564 , \24003 , \23429 );
nor \U$29187 ( \29565 , \29563 , \29564 );
xnor \U$29188 ( \29566 , \29565 , \23279 );
and \U$29189 ( \29567 , \24482 , \23163 );
and \U$29190 ( \29568 , \24344 , \23161 );
nor \U$29191 ( \29569 , \29567 , \29568 );
xnor \U$29192 ( \29570 , \29569 , \23007 );
and \U$29193 ( \29571 , \29566 , \29570 );
and \U$29194 ( \29572 , \25018 , \22891 );
and \U$29195 ( \29573 , \24601 , \22889 );
nor \U$29196 ( \29574 , \29572 , \29573 );
xnor \U$29197 ( \29575 , \29574 , \22778 );
and \U$29198 ( \29576 , \29570 , \29575 );
and \U$29199 ( \29577 , \29566 , \29575 );
or \U$29200 ( \29578 , \29571 , \29576 , \29577 );
and \U$29201 ( \29579 , \29562 , \29578 );
and \U$29202 ( \29580 , \22716 , \25369 );
and \U$29203 ( \29581 , \22611 , \25367 );
nor \U$29204 ( \29582 , \29580 , \29581 );
xnor \U$29205 ( \29583 , \29582 , \25123 );
and \U$29206 ( \29584 , \22837 , \24974 );
and \U$29207 ( \29585 , \22721 , \24972 );
nor \U$29208 ( \29586 , \29584 , \29585 );
xnor \U$29209 ( \29587 , \29586 , \24787 );
and \U$29210 ( \29588 , \29583 , \29587 );
and \U$29211 ( \29589 , \23128 , \24661 );
and \U$29212 ( \29590 , \22952 , \24659 );
nor \U$29213 ( \29591 , \29589 , \29590 );
xnor \U$29214 ( \29592 , \29591 , \24456 );
and \U$29215 ( \29593 , \29587 , \29592 );
and \U$29216 ( \29594 , \29583 , \29592 );
or \U$29217 ( \29595 , \29588 , \29593 , \29594 );
and \U$29218 ( \29596 , \29578 , \29595 );
and \U$29219 ( \29597 , \29562 , \29595 );
or \U$29220 ( \29598 , \29579 , \29596 , \29597 );
and \U$29221 ( \29599 , \26585 , \22163 );
and \U$29222 ( \29600 , \26116 , \22161 );
nor \U$29223 ( \29601 , \29599 , \29600 );
xnor \U$29224 ( \29602 , \29601 , \22091 );
and \U$29225 ( \29603 , \26854 , \22029 );
and \U$29226 ( \29604 , \26590 , \22027 );
nor \U$29227 ( \29605 , \29603 , \29604 );
xnor \U$29228 ( \29606 , \29605 , \21986 );
and \U$29229 ( \29607 , \29602 , \29606 );
and \U$29230 ( \29608 , \27485 , \21916 );
and \U$29231 ( \29609 , \27113 , \21914 );
nor \U$29232 ( \29610 , \29608 , \29609 );
xnor \U$29233 ( \29611 , \29610 , \21867 );
and \U$29234 ( \29612 , \29606 , \29611 );
and \U$29235 ( \29613 , \29602 , \29611 );
or \U$29236 ( \29614 , \29607 , \29612 , \29613 );
and \U$29237 ( \29615 , \25348 , \22697 );
and \U$29238 ( \29616 , \25226 , \22695 );
nor \U$29239 ( \29617 , \29615 , \29616 );
xnor \U$29240 ( \29618 , \29617 , \22561 );
and \U$29241 ( \29619 , \25609 , \22497 );
and \U$29242 ( \29620 , \25353 , \22495 );
nor \U$29243 ( \29621 , \29619 , \29620 );
xnor \U$29244 ( \29622 , \29621 , \22419 );
and \U$29245 ( \29623 , \29618 , \29622 );
and \U$29246 ( \29624 , \26108 , \22333 );
and \U$29247 ( \29625 , \25806 , \22331 );
nor \U$29248 ( \29626 , \29624 , \29625 );
xnor \U$29249 ( \29627 , \29626 , \22239 );
and \U$29250 ( \29628 , \29622 , \29627 );
and \U$29251 ( \29629 , \29618 , \29627 );
or \U$29252 ( \29630 , \29623 , \29628 , \29629 );
and \U$29253 ( \29631 , \29614 , \29630 );
and \U$29254 ( \29632 , \27837 , \21815 );
and \U$29255 ( \29633 , \27494 , \21813 );
nor \U$29256 ( \29634 , \29632 , \29633 );
xnor \U$29257 ( \29635 , \29634 , \21774 );
and \U$29258 ( \29636 , \28342 , \21745 );
and \U$29259 ( \29637 , \28039 , \21743 );
nor \U$29260 ( \29638 , \29636 , \29637 );
xnor \U$29261 ( \29639 , \29638 , \21715 );
and \U$29262 ( \29640 , \29635 , \29639 );
and \U$29263 ( \29641 , \29040 , \21697 );
and \U$29264 ( \29642 , \28514 , \21695 );
nor \U$29265 ( \29643 , \29641 , \29642 );
xnor \U$29266 ( \29644 , \29643 , \21678 );
and \U$29267 ( \29645 , \29639 , \29644 );
and \U$29268 ( \29646 , \29635 , \29644 );
or \U$29269 ( \29647 , \29640 , \29645 , \29646 );
and \U$29270 ( \29648 , \29630 , \29647 );
and \U$29271 ( \29649 , \29614 , \29647 );
or \U$29272 ( \29650 , \29631 , \29648 , \29649 );
and \U$29273 ( \29651 , \29598 , \29650 );
and \U$29274 ( \29652 , \22126 , \26517 );
and \U$29275 ( \29653 , \22046 , \26515 );
nor \U$29276 ( \29654 , \29652 , \29653 );
xnor \U$29277 ( \29655 , \29654 , \26329 );
and \U$29278 ( \29656 , \22262 , \26143 );
and \U$29279 ( \29657 , \22200 , \26141 );
nor \U$29280 ( \29658 , \29656 , \29657 );
xnor \U$29281 ( \29659 , \29658 , \25911 );
and \U$29282 ( \29660 , \29655 , \29659 );
and \U$29283 ( \29661 , \22523 , \25692 );
and \U$29284 ( \29662 , \22325 , \25690 );
nor \U$29285 ( \29663 , \29661 , \29662 );
xnor \U$29286 ( \29664 , \29663 , \25549 );
and \U$29287 ( \29665 , \29659 , \29664 );
and \U$29288 ( \29666 , \29655 , \29664 );
or \U$29289 ( \29667 , \29660 , \29665 , \29666 );
xor \U$29290 ( \29668 , \28852 , \29349 );
xor \U$29291 ( \29669 , \29349 , \29350 );
not \U$29292 ( \29670 , \29669 );
and \U$29293 ( \29671 , \29668 , \29670 );
and \U$29294 ( \29672 , \21653 , \29671 );
not \U$29295 ( \29673 , \29672 );
xnor \U$29296 ( \29674 , \29673 , \29353 );
and \U$29297 ( \29675 , \21685 , \29104 );
and \U$29298 ( \29676 , \21667 , \29102 );
nor \U$29299 ( \29677 , \29675 , \29676 );
xnor \U$29300 ( \29678 , \29677 , \28855 );
and \U$29301 ( \29679 , \29674 , \29678 );
and \U$29302 ( \29680 , \21754 , \28575 );
and \U$29303 ( \29681 , \21706 , \28573 );
nor \U$29304 ( \29682 , \29680 , \29681 );
xnor \U$29305 ( \29683 , \29682 , \28315 );
and \U$29306 ( \29684 , \29678 , \29683 );
and \U$29307 ( \29685 , \29674 , \29683 );
or \U$29308 ( \29686 , \29679 , \29684 , \29685 );
and \U$29309 ( \29687 , \29667 , \29686 );
and \U$29310 ( \29688 , \21831 , \28081 );
and \U$29311 ( \29689 , \21762 , \28079 );
nor \U$29312 ( \29690 , \29688 , \29689 );
xnor \U$29313 ( \29691 , \29690 , \27766 );
and \U$29314 ( \29692 , \21890 , \27572 );
and \U$29315 ( \29693 , \21836 , \27570 );
nor \U$29316 ( \29694 , \29692 , \29693 );
xnor \U$29317 ( \29695 , \29694 , \27232 );
and \U$29318 ( \29696 , \29691 , \29695 );
and \U$29319 ( \29697 , \22018 , \26983 );
and \U$29320 ( \29698 , \21941 , \26981 );
nor \U$29321 ( \29699 , \29697 , \29698 );
xnor \U$29322 ( \29700 , \29699 , \26742 );
and \U$29323 ( \29701 , \29695 , \29700 );
and \U$29324 ( \29702 , \29691 , \29700 );
or \U$29325 ( \29703 , \29696 , \29701 , \29702 );
and \U$29326 ( \29704 , \29686 , \29703 );
and \U$29327 ( \29705 , \29667 , \29703 );
or \U$29328 ( \29706 , \29687 , \29704 , \29705 );
and \U$29329 ( \29707 , \29650 , \29706 );
and \U$29330 ( \29708 , \29598 , \29706 );
or \U$29331 ( \29709 , \29651 , \29707 , \29708 );
buf \U$29332 ( \29710 , RIc22aee0_183);
and \U$29333 ( \29711 , \29710 , \21660 );
and \U$29334 ( \29712 , \29464 , \21658 );
nor \U$29335 ( \29713 , \29711 , \29712 );
xnor \U$29336 ( \29714 , \29713 , \21665 );
buf \U$29337 ( \29715 , RIc22af58_184);
and \U$29338 ( \29716 , \29715 , \21654 );
or \U$29339 ( \29717 , \29714 , \29716 );
and \U$29340 ( \29718 , \29464 , \21660 );
and \U$29341 ( \29719 , \29040 , \21658 );
nor \U$29342 ( \29720 , \29718 , \29719 );
xnor \U$29343 ( \29721 , \29720 , \21665 );
and \U$29344 ( \29722 , \29717 , \29721 );
and \U$29345 ( \29723 , \29710 , \21654 );
and \U$29346 ( \29724 , \29721 , \29723 );
and \U$29347 ( \29725 , \29717 , \29723 );
or \U$29348 ( \29726 , \29722 , \29724 , \29725 );
xor \U$29349 ( \29727 , \29391 , \29395 );
xor \U$29350 ( \29728 , \29727 , \29400 );
xor \U$29351 ( \29729 , \29407 , \29411 );
xor \U$29352 ( \29730 , \29729 , \29416 );
and \U$29353 ( \29731 , \29728 , \29730 );
xor \U$29354 ( \29732 , \29424 , \29428 );
xor \U$29355 ( \29733 , \29732 , \29433 );
and \U$29356 ( \29734 , \29730 , \29733 );
and \U$29357 ( \29735 , \29728 , \29733 );
or \U$29358 ( \29736 , \29731 , \29734 , \29735 );
and \U$29359 ( \29737 , \29726 , \29736 );
xor \U$29360 ( \29738 , \29284 , \29288 );
xor \U$29361 ( \29739 , \29738 , \29293 );
xor \U$29362 ( \29740 , \29300 , \29304 );
xor \U$29363 ( \29741 , \29740 , \29309 );
and \U$29364 ( \29742 , \29739 , \29741 );
xor \U$29365 ( \29743 , \29317 , \29321 );
xor \U$29366 ( \29744 , \29743 , \29326 );
and \U$29367 ( \29745 , \29741 , \29744 );
and \U$29368 ( \29746 , \29739 , \29744 );
or \U$29369 ( \29747 , \29742 , \29745 , \29746 );
and \U$29370 ( \29748 , \29736 , \29747 );
and \U$29371 ( \29749 , \29726 , \29747 );
or \U$29372 ( \29750 , \29737 , \29748 , \29749 );
and \U$29373 ( \29751 , \29709 , \29750 );
xor \U$29374 ( \29752 , \29336 , \29340 );
xor \U$29375 ( \29753 , \29752 , \29345 );
xor \U$29376 ( \29754 , \29354 , \29358 );
xor \U$29377 ( \29755 , \29754 , \29363 );
and \U$29378 ( \29756 , \29753 , \29755 );
xor \U$29379 ( \29757 , \29371 , \29375 );
xor \U$29380 ( \29758 , \29757 , \29380 );
and \U$29381 ( \29759 , \29755 , \29758 );
and \U$29382 ( \29760 , \29753 , \29758 );
or \U$29383 ( \29761 , \29756 , \29759 , \29760 );
xor \U$29384 ( \29762 , \29071 , \29075 );
xor \U$29385 ( \29763 , \29762 , \29080 );
and \U$29386 ( \29764 , \29761 , \29763 );
xor \U$29387 ( \29765 , \29107 , \29111 );
xor \U$29388 ( \29766 , \29765 , \29116 );
and \U$29389 ( \29767 , \29763 , \29766 );
and \U$29390 ( \29768 , \29761 , \29766 );
or \U$29391 ( \29769 , \29764 , \29767 , \29768 );
and \U$29392 ( \29770 , \29750 , \29769 );
and \U$29393 ( \29771 , \29709 , \29769 );
or \U$29394 ( \29772 , \29751 , \29770 , \29771 );
xor \U$29395 ( \29773 , \29296 , \29312 );
xor \U$29396 ( \29774 , \29773 , \29329 );
xor \U$29397 ( \29775 , \29348 , \29366 );
xor \U$29398 ( \29776 , \29775 , \29383 );
and \U$29399 ( \29777 , \29774 , \29776 );
xor \U$29400 ( \29778 , \29403 , \29419 );
xor \U$29401 ( \29779 , \29778 , \29436 );
and \U$29402 ( \29780 , \29776 , \29779 );
and \U$29403 ( \29781 , \29774 , \29779 );
or \U$29404 ( \29782 , \29777 , \29780 , \29781 );
xor \U$29405 ( \29783 , \29444 , \29446 );
xor \U$29406 ( \29784 , \29783 , \29449 );
xor \U$29407 ( \29785 , \29454 , \29456 );
xor \U$29408 ( \29786 , \29785 , \29459 );
and \U$29409 ( \29787 , \29784 , \29786 );
xnor \U$29410 ( \29788 , \29465 , \29467 );
and \U$29411 ( \29789 , \29786 , \29788 );
and \U$29412 ( \29790 , \29784 , \29788 );
or \U$29413 ( \29791 , \29787 , \29789 , \29790 );
and \U$29414 ( \29792 , \29782 , \29791 );
xor \U$29415 ( \29793 , \29083 , \29099 );
xor \U$29416 ( \29794 , \29793 , \29119 );
and \U$29417 ( \29795 , \29791 , \29794 );
and \U$29418 ( \29796 , \29782 , \29794 );
or \U$29419 ( \29797 , \29792 , \29795 , \29796 );
and \U$29420 ( \29798 , \29772 , \29797 );
xor \U$29421 ( \29799 , \29452 , \29462 );
xor \U$29422 ( \29800 , \29799 , \29468 );
xor \U$29423 ( \29801 , \29498 , \29500 );
xor \U$29424 ( \29802 , \29801 , \29503 );
and \U$29425 ( \29803 , \29800 , \29802 );
xor \U$29426 ( \29804 , \29474 , \29476 );
xor \U$29427 ( \29805 , \29804 , \29479 );
and \U$29428 ( \29806 , \29802 , \29805 );
and \U$29429 ( \29807 , \29800 , \29805 );
or \U$29430 ( \29808 , \29803 , \29806 , \29807 );
and \U$29431 ( \29809 , \29797 , \29808 );
and \U$29432 ( \29810 , \29772 , \29808 );
or \U$29433 ( \29811 , \29798 , \29809 , \29810 );
xor \U$29434 ( \29812 , \29442 , \29471 );
xor \U$29435 ( \29813 , \29812 , \29482 );
xor \U$29436 ( \29814 , \29487 , \29489 );
xor \U$29437 ( \29815 , \29814 , \29492 );
and \U$29438 ( \29816 , \29813 , \29815 );
xor \U$29439 ( \29817 , \29506 , \29508 );
xor \U$29440 ( \29818 , \29817 , \29511 );
and \U$29441 ( \29819 , \29815 , \29818 );
and \U$29442 ( \29820 , \29813 , \29818 );
or \U$29443 ( \29821 , \29816 , \29819 , \29820 );
and \U$29444 ( \29822 , \29811 , \29821 );
xor \U$29445 ( \29823 , \29519 , \29521 );
xor \U$29446 ( \29824 , \29823 , \29523 );
and \U$29447 ( \29825 , \29821 , \29824 );
and \U$29448 ( \29826 , \29811 , \29824 );
or \U$29449 ( \29827 , \29822 , \29825 , \29826 );
xor \U$29450 ( \29828 , \29225 , \29242 );
xor \U$29451 ( \29829 , \29828 , \29248 );
and \U$29452 ( \29830 , \29827 , \29829 );
xor \U$29453 ( \29831 , \29517 , \29526 );
xor \U$29454 ( \29832 , \29831 , \29529 );
and \U$29455 ( \29833 , \29829 , \29832 );
and \U$29456 ( \29834 , \29827 , \29832 );
or \U$29457 ( \29835 , \29830 , \29833 , \29834 );
xor \U$29458 ( \29836 , \29532 , \29534 );
xor \U$29459 ( \29837 , \29836 , \29537 );
and \U$29460 ( \29838 , \29835 , \29837 );
and \U$29461 ( \29839 , \29546 , \29838 );
xor \U$29462 ( \29840 , \29546 , \29838 );
xor \U$29463 ( \29841 , \29835 , \29837 );
and \U$29464 ( \29842 , \21762 , \28575 );
and \U$29465 ( \29843 , \21754 , \28573 );
nor \U$29466 ( \29844 , \29842 , \29843 );
xnor \U$29467 ( \29845 , \29844 , \28315 );
and \U$29468 ( \29846 , \21836 , \28081 );
and \U$29469 ( \29847 , \21831 , \28079 );
nor \U$29470 ( \29848 , \29846 , \29847 );
xnor \U$29471 ( \29849 , \29848 , \27766 );
and \U$29472 ( \29850 , \29845 , \29849 );
and \U$29473 ( \29851 , \21941 , \27572 );
and \U$29474 ( \29852 , \21890 , \27570 );
nor \U$29475 ( \29853 , \29851 , \29852 );
xnor \U$29476 ( \29854 , \29853 , \27232 );
and \U$29477 ( \29855 , \29849 , \29854 );
and \U$29478 ( \29856 , \29845 , \29854 );
or \U$29479 ( \29857 , \29850 , \29855 , \29856 );
buf \U$29480 ( \29858 , RIc225af8_58);
buf \U$29481 ( \29859 , RIc225a80_59);
and \U$29482 ( \29860 , \29858 , \29859 );
not \U$29483 ( \29861 , \29860 );
and \U$29484 ( \29862 , \29350 , \29861 );
not \U$29485 ( \29863 , \29862 );
and \U$29486 ( \29864 , \21667 , \29671 );
and \U$29487 ( \29865 , \21653 , \29669 );
nor \U$29488 ( \29866 , \29864 , \29865 );
xnor \U$29489 ( \29867 , \29866 , \29353 );
and \U$29490 ( \29868 , \29863 , \29867 );
and \U$29491 ( \29869 , \21706 , \29104 );
and \U$29492 ( \29870 , \21685 , \29102 );
nor \U$29493 ( \29871 , \29869 , \29870 );
xnor \U$29494 ( \29872 , \29871 , \28855 );
and \U$29495 ( \29873 , \29867 , \29872 );
and \U$29496 ( \29874 , \29863 , \29872 );
or \U$29497 ( \29875 , \29868 , \29873 , \29874 );
and \U$29498 ( \29876 , \29857 , \29875 );
and \U$29499 ( \29877 , \22046 , \26983 );
and \U$29500 ( \29878 , \22018 , \26981 );
nor \U$29501 ( \29879 , \29877 , \29878 );
xnor \U$29502 ( \29880 , \29879 , \26742 );
and \U$29503 ( \29881 , \22200 , \26517 );
and \U$29504 ( \29882 , \22126 , \26515 );
nor \U$29505 ( \29883 , \29881 , \29882 );
xnor \U$29506 ( \29884 , \29883 , \26329 );
and \U$29507 ( \29885 , \29880 , \29884 );
and \U$29508 ( \29886 , \22325 , \26143 );
and \U$29509 ( \29887 , \22262 , \26141 );
nor \U$29510 ( \29888 , \29886 , \29887 );
xnor \U$29511 ( \29889 , \29888 , \25911 );
and \U$29512 ( \29890 , \29884 , \29889 );
and \U$29513 ( \29891 , \29880 , \29889 );
or \U$29514 ( \29892 , \29885 , \29890 , \29891 );
and \U$29515 ( \29893 , \29875 , \29892 );
and \U$29516 ( \29894 , \29857 , \29892 );
or \U$29517 ( \29895 , \29876 , \29893 , \29894 );
and \U$29518 ( \29896 , \24003 , \23637 );
and \U$29519 ( \29897 , \23978 , \23635 );
nor \U$29520 ( \29898 , \29896 , \29897 );
xnor \U$29521 ( \29899 , \29898 , \23500 );
and \U$29522 ( \29900 , \24344 , \23431 );
and \U$29523 ( \29901 , \24177 , \23429 );
nor \U$29524 ( \29902 , \29900 , \29901 );
xnor \U$29525 ( \29903 , \29902 , \23279 );
and \U$29526 ( \29904 , \29899 , \29903 );
and \U$29527 ( \29905 , \24601 , \23163 );
and \U$29528 ( \29906 , \24482 , \23161 );
nor \U$29529 ( \29907 , \29905 , \29906 );
xnor \U$29530 ( \29908 , \29907 , \23007 );
and \U$29531 ( \29909 , \29903 , \29908 );
and \U$29532 ( \29910 , \29899 , \29908 );
or \U$29533 ( \29911 , \29904 , \29909 , \29910 );
and \U$29534 ( \29912 , \23136 , \24661 );
and \U$29535 ( \29913 , \23128 , \24659 );
nor \U$29536 ( \29914 , \29912 , \29913 );
xnor \U$29537 ( \29915 , \29914 , \24456 );
and \U$29538 ( \29916 , \23384 , \24255 );
and \U$29539 ( \29917 , \23379 , \24253 );
nor \U$29540 ( \29918 , \29916 , \29917 );
xnor \U$29541 ( \29919 , \29918 , \24106 );
and \U$29542 ( \29920 , \29915 , \29919 );
and \U$29543 ( \29921 , \23714 , \23933 );
and \U$29544 ( \29922 , \23570 , \23931 );
nor \U$29545 ( \29923 , \29921 , \29922 );
xnor \U$29546 ( \29924 , \29923 , \23791 );
and \U$29547 ( \29925 , \29919 , \29924 );
and \U$29548 ( \29926 , \29915 , \29924 );
or \U$29549 ( \29927 , \29920 , \29925 , \29926 );
and \U$29550 ( \29928 , \29911 , \29927 );
and \U$29551 ( \29929 , \22611 , \25692 );
and \U$29552 ( \29930 , \22523 , \25690 );
nor \U$29553 ( \29931 , \29929 , \29930 );
xnor \U$29554 ( \29932 , \29931 , \25549 );
and \U$29555 ( \29933 , \22721 , \25369 );
and \U$29556 ( \29934 , \22716 , \25367 );
nor \U$29557 ( \29935 , \29933 , \29934 );
xnor \U$29558 ( \29936 , \29935 , \25123 );
and \U$29559 ( \29937 , \29932 , \29936 );
and \U$29560 ( \29938 , \22952 , \24974 );
and \U$29561 ( \29939 , \22837 , \24972 );
nor \U$29562 ( \29940 , \29938 , \29939 );
xnor \U$29563 ( \29941 , \29940 , \24787 );
and \U$29564 ( \29942 , \29936 , \29941 );
and \U$29565 ( \29943 , \29932 , \29941 );
or \U$29566 ( \29944 , \29937 , \29942 , \29943 );
and \U$29567 ( \29945 , \29927 , \29944 );
and \U$29568 ( \29946 , \29911 , \29944 );
or \U$29569 ( \29947 , \29928 , \29945 , \29946 );
and \U$29570 ( \29948 , \29895 , \29947 );
and \U$29571 ( \29949 , \26116 , \22333 );
and \U$29572 ( \29950 , \26108 , \22331 );
nor \U$29573 ( \29951 , \29949 , \29950 );
xnor \U$29574 ( \29952 , \29951 , \22239 );
and \U$29575 ( \29953 , \26590 , \22163 );
and \U$29576 ( \29954 , \26585 , \22161 );
nor \U$29577 ( \29955 , \29953 , \29954 );
xnor \U$29578 ( \29956 , \29955 , \22091 );
and \U$29579 ( \29957 , \29952 , \29956 );
and \U$29580 ( \29958 , \27113 , \22029 );
and \U$29581 ( \29959 , \26854 , \22027 );
nor \U$29582 ( \29960 , \29958 , \29959 );
xnor \U$29583 ( \29961 , \29960 , \21986 );
and \U$29584 ( \29962 , \29956 , \29961 );
and \U$29585 ( \29963 , \29952 , \29961 );
or \U$29586 ( \29964 , \29957 , \29962 , \29963 );
and \U$29587 ( \29965 , \25226 , \22891 );
and \U$29588 ( \29966 , \25018 , \22889 );
nor \U$29589 ( \29967 , \29965 , \29966 );
xnor \U$29590 ( \29968 , \29967 , \22778 );
and \U$29591 ( \29969 , \25353 , \22697 );
and \U$29592 ( \29970 , \25348 , \22695 );
nor \U$29593 ( \29971 , \29969 , \29970 );
xnor \U$29594 ( \29972 , \29971 , \22561 );
and \U$29595 ( \29973 , \29968 , \29972 );
and \U$29596 ( \29974 , \25806 , \22497 );
and \U$29597 ( \29975 , \25609 , \22495 );
nor \U$29598 ( \29976 , \29974 , \29975 );
xnor \U$29599 ( \29977 , \29976 , \22419 );
and \U$29600 ( \29978 , \29972 , \29977 );
and \U$29601 ( \29979 , \29968 , \29977 );
or \U$29602 ( \29980 , \29973 , \29978 , \29979 );
and \U$29603 ( \29981 , \29964 , \29980 );
and \U$29604 ( \29982 , \27494 , \21916 );
and \U$29605 ( \29983 , \27485 , \21914 );
nor \U$29606 ( \29984 , \29982 , \29983 );
xnor \U$29607 ( \29985 , \29984 , \21867 );
and \U$29608 ( \29986 , \28039 , \21815 );
and \U$29609 ( \29987 , \27837 , \21813 );
nor \U$29610 ( \29988 , \29986 , \29987 );
xnor \U$29611 ( \29989 , \29988 , \21774 );
and \U$29612 ( \29990 , \29985 , \29989 );
and \U$29613 ( \29991 , \28514 , \21745 );
and \U$29614 ( \29992 , \28342 , \21743 );
nor \U$29615 ( \29993 , \29991 , \29992 );
xnor \U$29616 ( \29994 , \29993 , \21715 );
and \U$29617 ( \29995 , \29989 , \29994 );
and \U$29618 ( \29996 , \29985 , \29994 );
or \U$29619 ( \29997 , \29990 , \29995 , \29996 );
and \U$29620 ( \29998 , \29980 , \29997 );
and \U$29621 ( \29999 , \29964 , \29997 );
or \U$29622 ( \30000 , \29981 , \29998 , \29999 );
and \U$29623 ( \30001 , \29947 , \30000 );
and \U$29624 ( \30002 , \29895 , \30000 );
or \U$29625 ( \30003 , \29948 , \30001 , \30002 );
xor \U$29626 ( \30004 , \29550 , \29554 );
xor \U$29627 ( \30005 , \30004 , \29559 );
xor \U$29628 ( \30006 , \29655 , \29659 );
xor \U$29629 ( \30007 , \30006 , \29664 );
and \U$29630 ( \30008 , \30005 , \30007 );
xor \U$29631 ( \30009 , \29583 , \29587 );
xor \U$29632 ( \30010 , \30009 , \29592 );
and \U$29633 ( \30011 , \30007 , \30010 );
and \U$29634 ( \30012 , \30005 , \30010 );
or \U$29635 ( \30013 , \30008 , \30011 , \30012 );
xor \U$29636 ( \30014 , \29566 , \29570 );
xor \U$29637 ( \30015 , \30014 , \29575 );
xor \U$29638 ( \30016 , \29602 , \29606 );
xor \U$29639 ( \30017 , \30016 , \29611 );
and \U$29640 ( \30018 , \30015 , \30017 );
xor \U$29641 ( \30019 , \29618 , \29622 );
xor \U$29642 ( \30020 , \30019 , \29627 );
and \U$29643 ( \30021 , \30017 , \30020 );
and \U$29644 ( \30022 , \30015 , \30020 );
or \U$29645 ( \30023 , \30018 , \30021 , \30022 );
and \U$29646 ( \30024 , \30013 , \30023 );
and \U$29647 ( \30025 , \29464 , \21697 );
and \U$29648 ( \30026 , \29040 , \21695 );
nor \U$29649 ( \30027 , \30025 , \30026 );
xnor \U$29650 ( \30028 , \30027 , \21678 );
and \U$29651 ( \30029 , \29715 , \21660 );
and \U$29652 ( \30030 , \29710 , \21658 );
nor \U$29653 ( \30031 , \30029 , \30030 );
xnor \U$29654 ( \30032 , \30031 , \21665 );
and \U$29655 ( \30033 , \30028 , \30032 );
buf \U$29656 ( \30034 , RIc22afd0_185);
and \U$29657 ( \30035 , \30034 , \21654 );
and \U$29658 ( \30036 , \30032 , \30035 );
and \U$29659 ( \30037 , \30028 , \30035 );
or \U$29660 ( \30038 , \30033 , \30036 , \30037 );
xor \U$29661 ( \30039 , \29635 , \29639 );
xor \U$29662 ( \30040 , \30039 , \29644 );
and \U$29663 ( \30041 , \30038 , \30040 );
xnor \U$29664 ( \30042 , \29714 , \29716 );
and \U$29665 ( \30043 , \30040 , \30042 );
and \U$29666 ( \30044 , \30038 , \30042 );
or \U$29667 ( \30045 , \30041 , \30043 , \30044 );
and \U$29668 ( \30046 , \30023 , \30045 );
and \U$29669 ( \30047 , \30013 , \30045 );
or \U$29670 ( \30048 , \30024 , \30046 , \30047 );
and \U$29671 ( \30049 , \30003 , \30048 );
xor \U$29672 ( \30050 , \29728 , \29730 );
xor \U$29673 ( \30051 , \30050 , \29733 );
xor \U$29674 ( \30052 , \29739 , \29741 );
xor \U$29675 ( \30053 , \30052 , \29744 );
and \U$29676 ( \30054 , \30051 , \30053 );
xor \U$29677 ( \30055 , \29753 , \29755 );
xor \U$29678 ( \30056 , \30055 , \29758 );
and \U$29679 ( \30057 , \30053 , \30056 );
and \U$29680 ( \30058 , \30051 , \30056 );
or \U$29681 ( \30059 , \30054 , \30057 , \30058 );
and \U$29682 ( \30060 , \30048 , \30059 );
and \U$29683 ( \30061 , \30003 , \30059 );
or \U$29684 ( \30062 , \30049 , \30060 , \30061 );
xor \U$29685 ( \30063 , \29598 , \29650 );
xor \U$29686 ( \30064 , \30063 , \29706 );
xor \U$29687 ( \30065 , \29726 , \29736 );
xor \U$29688 ( \30066 , \30065 , \29747 );
and \U$29689 ( \30067 , \30064 , \30066 );
xor \U$29690 ( \30068 , \29761 , \29763 );
xor \U$29691 ( \30069 , \30068 , \29766 );
and \U$29692 ( \30070 , \30066 , \30069 );
and \U$29693 ( \30071 , \30064 , \30069 );
or \U$29694 ( \30072 , \30067 , \30070 , \30071 );
and \U$29695 ( \30073 , \30062 , \30072 );
xor \U$29696 ( \30074 , \29562 , \29578 );
xor \U$29697 ( \30075 , \30074 , \29595 );
xor \U$29698 ( \30076 , \29614 , \29630 );
xor \U$29699 ( \30077 , \30076 , \29647 );
and \U$29700 ( \30078 , \30075 , \30077 );
xor \U$29701 ( \30079 , \29717 , \29721 );
xor \U$29702 ( \30080 , \30079 , \29723 );
and \U$29703 ( \30081 , \30077 , \30080 );
and \U$29704 ( \30082 , \30075 , \30080 );
or \U$29705 ( \30083 , \30078 , \30081 , \30082 );
xor \U$29706 ( \30084 , \29774 , \29776 );
xor \U$29707 ( \30085 , \30084 , \29779 );
and \U$29708 ( \30086 , \30083 , \30085 );
xor \U$29709 ( \30087 , \29784 , \29786 );
xor \U$29710 ( \30088 , \30087 , \29788 );
and \U$29711 ( \30089 , \30085 , \30088 );
and \U$29712 ( \30090 , \30083 , \30088 );
or \U$29713 ( \30091 , \30086 , \30089 , \30090 );
and \U$29714 ( \30092 , \30072 , \30091 );
and \U$29715 ( \30093 , \30062 , \30091 );
or \U$29716 ( \30094 , \30073 , \30092 , \30093 );
xor \U$29717 ( \30095 , \29332 , \29386 );
xor \U$29718 ( \30096 , \30095 , \29439 );
xor \U$29719 ( \30097 , \29782 , \29791 );
xor \U$29720 ( \30098 , \30097 , \29794 );
and \U$29721 ( \30099 , \30096 , \30098 );
xor \U$29722 ( \30100 , \29800 , \29802 );
xor \U$29723 ( \30101 , \30100 , \29805 );
and \U$29724 ( \30102 , \30098 , \30101 );
and \U$29725 ( \30103 , \30096 , \30101 );
or \U$29726 ( \30104 , \30099 , \30102 , \30103 );
and \U$29727 ( \30105 , \30094 , \30104 );
xor \U$29728 ( \30106 , \29813 , \29815 );
xor \U$29729 ( \30107 , \30106 , \29818 );
and \U$29730 ( \30108 , \30104 , \30107 );
and \U$29731 ( \30109 , \30094 , \30107 );
or \U$29732 ( \30110 , \30105 , \30108 , \30109 );
xor \U$29733 ( \30111 , \29485 , \29495 );
xor \U$29734 ( \30112 , \30111 , \29514 );
and \U$29735 ( \30113 , \30110 , \30112 );
xor \U$29736 ( \30114 , \29811 , \29821 );
xor \U$29737 ( \30115 , \30114 , \29824 );
and \U$29738 ( \30116 , \30112 , \30115 );
and \U$29739 ( \30117 , \30110 , \30115 );
or \U$29740 ( \30118 , \30113 , \30116 , \30117 );
xor \U$29741 ( \30119 , \29827 , \29829 );
xor \U$29742 ( \30120 , \30119 , \29832 );
and \U$29743 ( \30121 , \30118 , \30120 );
and \U$29744 ( \30122 , \29841 , \30121 );
xor \U$29745 ( \30123 , \29841 , \30121 );
xor \U$29746 ( \30124 , \30118 , \30120 );
and \U$29747 ( \30125 , \24177 , \23637 );
and \U$29748 ( \30126 , \24003 , \23635 );
nor \U$29749 ( \30127 , \30125 , \30126 );
xnor \U$29750 ( \30128 , \30127 , \23500 );
and \U$29751 ( \30129 , \24482 , \23431 );
and \U$29752 ( \30130 , \24344 , \23429 );
nor \U$29753 ( \30131 , \30129 , \30130 );
xnor \U$29754 ( \30132 , \30131 , \23279 );
and \U$29755 ( \30133 , \30128 , \30132 );
and \U$29756 ( \30134 , \25018 , \23163 );
and \U$29757 ( \30135 , \24601 , \23161 );
nor \U$29758 ( \30136 , \30134 , \30135 );
xnor \U$29759 ( \30137 , \30136 , \23007 );
and \U$29760 ( \30138 , \30132 , \30137 );
and \U$29761 ( \30139 , \30128 , \30137 );
or \U$29762 ( \30140 , \30133 , \30138 , \30139 );
and \U$29763 ( \30141 , \22716 , \25692 );
and \U$29764 ( \30142 , \22611 , \25690 );
nor \U$29765 ( \30143 , \30141 , \30142 );
xnor \U$29766 ( \30144 , \30143 , \25549 );
and \U$29767 ( \30145 , \22837 , \25369 );
and \U$29768 ( \30146 , \22721 , \25367 );
nor \U$29769 ( \30147 , \30145 , \30146 );
xnor \U$29770 ( \30148 , \30147 , \25123 );
and \U$29771 ( \30149 , \30144 , \30148 );
and \U$29772 ( \30150 , \23128 , \24974 );
and \U$29773 ( \30151 , \22952 , \24972 );
nor \U$29774 ( \30152 , \30150 , \30151 );
xnor \U$29775 ( \30153 , \30152 , \24787 );
and \U$29776 ( \30154 , \30148 , \30153 );
and \U$29777 ( \30155 , \30144 , \30153 );
or \U$29778 ( \30156 , \30149 , \30154 , \30155 );
and \U$29779 ( \30157 , \30140 , \30156 );
and \U$29780 ( \30158 , \23379 , \24661 );
and \U$29781 ( \30159 , \23136 , \24659 );
nor \U$29782 ( \30160 , \30158 , \30159 );
xnor \U$29783 ( \30161 , \30160 , \24456 );
and \U$29784 ( \30162 , \23570 , \24255 );
and \U$29785 ( \30163 , \23384 , \24253 );
nor \U$29786 ( \30164 , \30162 , \30163 );
xnor \U$29787 ( \30165 , \30164 , \24106 );
and \U$29788 ( \30166 , \30161 , \30165 );
and \U$29789 ( \30167 , \23978 , \23933 );
and \U$29790 ( \30168 , \23714 , \23931 );
nor \U$29791 ( \30169 , \30167 , \30168 );
xnor \U$29792 ( \30170 , \30169 , \23791 );
and \U$29793 ( \30171 , \30165 , \30170 );
and \U$29794 ( \30172 , \30161 , \30170 );
or \U$29795 ( \30173 , \30166 , \30171 , \30172 );
and \U$29796 ( \30174 , \30156 , \30173 );
and \U$29797 ( \30175 , \30140 , \30173 );
or \U$29798 ( \30176 , \30157 , \30174 , \30175 );
and \U$29799 ( \30177 , \27837 , \21916 );
and \U$29800 ( \30178 , \27494 , \21914 );
nor \U$29801 ( \30179 , \30177 , \30178 );
xnor \U$29802 ( \30180 , \30179 , \21867 );
and \U$29803 ( \30181 , \28342 , \21815 );
and \U$29804 ( \30182 , \28039 , \21813 );
nor \U$29805 ( \30183 , \30181 , \30182 );
xnor \U$29806 ( \30184 , \30183 , \21774 );
and \U$29807 ( \30185 , \30180 , \30184 );
and \U$29808 ( \30186 , \29040 , \21745 );
and \U$29809 ( \30187 , \28514 , \21743 );
nor \U$29810 ( \30188 , \30186 , \30187 );
xnor \U$29811 ( \30189 , \30188 , \21715 );
and \U$29812 ( \30190 , \30184 , \30189 );
and \U$29813 ( \30191 , \30180 , \30189 );
or \U$29814 ( \30192 , \30185 , \30190 , \30191 );
and \U$29815 ( \30193 , \26585 , \22333 );
and \U$29816 ( \30194 , \26116 , \22331 );
nor \U$29817 ( \30195 , \30193 , \30194 );
xnor \U$29818 ( \30196 , \30195 , \22239 );
and \U$29819 ( \30197 , \26854 , \22163 );
and \U$29820 ( \30198 , \26590 , \22161 );
nor \U$29821 ( \30199 , \30197 , \30198 );
xnor \U$29822 ( \30200 , \30199 , \22091 );
and \U$29823 ( \30201 , \30196 , \30200 );
and \U$29824 ( \30202 , \27485 , \22029 );
and \U$29825 ( \30203 , \27113 , \22027 );
nor \U$29826 ( \30204 , \30202 , \30203 );
xnor \U$29827 ( \30205 , \30204 , \21986 );
and \U$29828 ( \30206 , \30200 , \30205 );
and \U$29829 ( \30207 , \30196 , \30205 );
or \U$29830 ( \30208 , \30201 , \30206 , \30207 );
and \U$29831 ( \30209 , \30192 , \30208 );
and \U$29832 ( \30210 , \25348 , \22891 );
and \U$29833 ( \30211 , \25226 , \22889 );
nor \U$29834 ( \30212 , \30210 , \30211 );
xnor \U$29835 ( \30213 , \30212 , \22778 );
and \U$29836 ( \30214 , \25609 , \22697 );
and \U$29837 ( \30215 , \25353 , \22695 );
nor \U$29838 ( \30216 , \30214 , \30215 );
xnor \U$29839 ( \30217 , \30216 , \22561 );
and \U$29840 ( \30218 , \30213 , \30217 );
and \U$29841 ( \30219 , \26108 , \22497 );
and \U$29842 ( \30220 , \25806 , \22495 );
nor \U$29843 ( \30221 , \30219 , \30220 );
xnor \U$29844 ( \30222 , \30221 , \22419 );
and \U$29845 ( \30223 , \30217 , \30222 );
and \U$29846 ( \30224 , \30213 , \30222 );
or \U$29847 ( \30225 , \30218 , \30223 , \30224 );
and \U$29848 ( \30226 , \30208 , \30225 );
and \U$29849 ( \30227 , \30192 , \30225 );
or \U$29850 ( \30228 , \30209 , \30226 , \30227 );
and \U$29851 ( \30229 , \30176 , \30228 );
xor \U$29852 ( \30230 , \29350 , \29858 );
xor \U$29853 ( \30231 , \29858 , \29859 );
not \U$29854 ( \30232 , \30231 );
and \U$29855 ( \30233 , \30230 , \30232 );
and \U$29856 ( \30234 , \21653 , \30233 );
not \U$29857 ( \30235 , \30234 );
xnor \U$29858 ( \30236 , \30235 , \29862 );
and \U$29859 ( \30237 , \21685 , \29671 );
and \U$29860 ( \30238 , \21667 , \29669 );
nor \U$29861 ( \30239 , \30237 , \30238 );
xnor \U$29862 ( \30240 , \30239 , \29353 );
and \U$29863 ( \30241 , \30236 , \30240 );
and \U$29864 ( \30242 , \21754 , \29104 );
and \U$29865 ( \30243 , \21706 , \29102 );
nor \U$29866 ( \30244 , \30242 , \30243 );
xnor \U$29867 ( \30245 , \30244 , \28855 );
and \U$29868 ( \30246 , \30240 , \30245 );
and \U$29869 ( \30247 , \30236 , \30245 );
or \U$29870 ( \30248 , \30241 , \30246 , \30247 );
and \U$29871 ( \30249 , \22126 , \26983 );
and \U$29872 ( \30250 , \22046 , \26981 );
nor \U$29873 ( \30251 , \30249 , \30250 );
xnor \U$29874 ( \30252 , \30251 , \26742 );
and \U$29875 ( \30253 , \22262 , \26517 );
and \U$29876 ( \30254 , \22200 , \26515 );
nor \U$29877 ( \30255 , \30253 , \30254 );
xnor \U$29878 ( \30256 , \30255 , \26329 );
and \U$29879 ( \30257 , \30252 , \30256 );
and \U$29880 ( \30258 , \22523 , \26143 );
and \U$29881 ( \30259 , \22325 , \26141 );
nor \U$29882 ( \30260 , \30258 , \30259 );
xnor \U$29883 ( \30261 , \30260 , \25911 );
and \U$29884 ( \30262 , \30256 , \30261 );
and \U$29885 ( \30263 , \30252 , \30261 );
or \U$29886 ( \30264 , \30257 , \30262 , \30263 );
and \U$29887 ( \30265 , \30248 , \30264 );
and \U$29888 ( \30266 , \21831 , \28575 );
and \U$29889 ( \30267 , \21762 , \28573 );
nor \U$29890 ( \30268 , \30266 , \30267 );
xnor \U$29891 ( \30269 , \30268 , \28315 );
and \U$29892 ( \30270 , \21890 , \28081 );
and \U$29893 ( \30271 , \21836 , \28079 );
nor \U$29894 ( \30272 , \30270 , \30271 );
xnor \U$29895 ( \30273 , \30272 , \27766 );
and \U$29896 ( \30274 , \30269 , \30273 );
and \U$29897 ( \30275 , \22018 , \27572 );
and \U$29898 ( \30276 , \21941 , \27570 );
nor \U$29899 ( \30277 , \30275 , \30276 );
xnor \U$29900 ( \30278 , \30277 , \27232 );
and \U$29901 ( \30279 , \30273 , \30278 );
and \U$29902 ( \30280 , \30269 , \30278 );
or \U$29903 ( \30281 , \30274 , \30279 , \30280 );
and \U$29904 ( \30282 , \30264 , \30281 );
and \U$29905 ( \30283 , \30248 , \30281 );
or \U$29906 ( \30284 , \30265 , \30282 , \30283 );
and \U$29907 ( \30285 , \30228 , \30284 );
and \U$29908 ( \30286 , \30176 , \30284 );
or \U$29909 ( \30287 , \30229 , \30285 , \30286 );
xor \U$29910 ( \30288 , \29880 , \29884 );
xor \U$29911 ( \30289 , \30288 , \29889 );
xor \U$29912 ( \30290 , \29915 , \29919 );
xor \U$29913 ( \30291 , \30290 , \29924 );
and \U$29914 ( \30292 , \30289 , \30291 );
xor \U$29915 ( \30293 , \29932 , \29936 );
xor \U$29916 ( \30294 , \30293 , \29941 );
and \U$29917 ( \30295 , \30291 , \30294 );
and \U$29918 ( \30296 , \30289 , \30294 );
or \U$29919 ( \30297 , \30292 , \30295 , \30296 );
xor \U$29920 ( \30298 , \29899 , \29903 );
xor \U$29921 ( \30299 , \30298 , \29908 );
xor \U$29922 ( \30300 , \29952 , \29956 );
xor \U$29923 ( \30301 , \30300 , \29961 );
and \U$29924 ( \30302 , \30299 , \30301 );
xor \U$29925 ( \30303 , \29968 , \29972 );
xor \U$29926 ( \30304 , \30303 , \29977 );
and \U$29927 ( \30305 , \30301 , \30304 );
and \U$29928 ( \30306 , \30299 , \30304 );
or \U$29929 ( \30307 , \30302 , \30305 , \30306 );
and \U$29930 ( \30308 , \30297 , \30307 );
and \U$29931 ( \30309 , \29710 , \21697 );
and \U$29932 ( \30310 , \29464 , \21695 );
nor \U$29933 ( \30311 , \30309 , \30310 );
xnor \U$29934 ( \30312 , \30311 , \21678 );
and \U$29935 ( \30313 , \30034 , \21660 );
and \U$29936 ( \30314 , \29715 , \21658 );
nor \U$29937 ( \30315 , \30313 , \30314 );
xnor \U$29938 ( \30316 , \30315 , \21665 );
and \U$29939 ( \30317 , \30312 , \30316 );
buf \U$29940 ( \30318 , RIc22b048_186);
and \U$29941 ( \30319 , \30318 , \21654 );
and \U$29942 ( \30320 , \30316 , \30319 );
and \U$29943 ( \30321 , \30312 , \30319 );
or \U$29944 ( \30322 , \30317 , \30320 , \30321 );
xor \U$29945 ( \30323 , \30028 , \30032 );
xor \U$29946 ( \30324 , \30323 , \30035 );
and \U$29947 ( \30325 , \30322 , \30324 );
xor \U$29948 ( \30326 , \29985 , \29989 );
xor \U$29949 ( \30327 , \30326 , \29994 );
and \U$29950 ( \30328 , \30324 , \30327 );
and \U$29951 ( \30329 , \30322 , \30327 );
or \U$29952 ( \30330 , \30325 , \30328 , \30329 );
and \U$29953 ( \30331 , \30307 , \30330 );
and \U$29954 ( \30332 , \30297 , \30330 );
or \U$29955 ( \30333 , \30308 , \30331 , \30332 );
and \U$29956 ( \30334 , \30287 , \30333 );
xor \U$29957 ( \30335 , \29674 , \29678 );
xor \U$29958 ( \30336 , \30335 , \29683 );
xor \U$29959 ( \30337 , \29691 , \29695 );
xor \U$29960 ( \30338 , \30337 , \29700 );
and \U$29961 ( \30339 , \30336 , \30338 );
xor \U$29962 ( \30340 , \30005 , \30007 );
xor \U$29963 ( \30341 , \30340 , \30010 );
and \U$29964 ( \30342 , \30338 , \30341 );
and \U$29965 ( \30343 , \30336 , \30341 );
or \U$29966 ( \30344 , \30339 , \30342 , \30343 );
and \U$29967 ( \30345 , \30333 , \30344 );
and \U$29968 ( \30346 , \30287 , \30344 );
or \U$29969 ( \30347 , \30334 , \30345 , \30346 );
xor \U$29970 ( \30348 , \29964 , \29980 );
xor \U$29971 ( \30349 , \30348 , \29997 );
xor \U$29972 ( \30350 , \30015 , \30017 );
xor \U$29973 ( \30351 , \30350 , \30020 );
and \U$29974 ( \30352 , \30349 , \30351 );
xor \U$29975 ( \30353 , \30038 , \30040 );
xor \U$29976 ( \30354 , \30353 , \30042 );
and \U$29977 ( \30355 , \30351 , \30354 );
and \U$29978 ( \30356 , \30349 , \30354 );
or \U$29979 ( \30357 , \30352 , \30355 , \30356 );
xor \U$29980 ( \30358 , \29667 , \29686 );
xor \U$29981 ( \30359 , \30358 , \29703 );
and \U$29982 ( \30360 , \30357 , \30359 );
xor \U$29983 ( \30361 , \30075 , \30077 );
xor \U$29984 ( \30362 , \30361 , \30080 );
and \U$29985 ( \30363 , \30359 , \30362 );
and \U$29986 ( \30364 , \30357 , \30362 );
or \U$29987 ( \30365 , \30360 , \30363 , \30364 );
and \U$29988 ( \30366 , \30347 , \30365 );
xor \U$29989 ( \30367 , \29895 , \29947 );
xor \U$29990 ( \30368 , \30367 , \30000 );
xor \U$29991 ( \30369 , \30013 , \30023 );
xor \U$29992 ( \30370 , \30369 , \30045 );
and \U$29993 ( \30371 , \30368 , \30370 );
xor \U$29994 ( \30372 , \30051 , \30053 );
xor \U$29995 ( \30373 , \30372 , \30056 );
and \U$29996 ( \30374 , \30370 , \30373 );
and \U$29997 ( \30375 , \30368 , \30373 );
or \U$29998 ( \30376 , \30371 , \30374 , \30375 );
and \U$29999 ( \30377 , \30365 , \30376 );
and \U$30000 ( \30378 , \30347 , \30376 );
or \U$30001 ( \30379 , \30366 , \30377 , \30378 );
xor \U$30002 ( \30380 , \30003 , \30048 );
xor \U$30003 ( \30381 , \30380 , \30059 );
xor \U$30004 ( \30382 , \30064 , \30066 );
xor \U$30005 ( \30383 , \30382 , \30069 );
and \U$30006 ( \30384 , \30381 , \30383 );
xor \U$30007 ( \30385 , \30083 , \30085 );
xor \U$30008 ( \30386 , \30385 , \30088 );
and \U$30009 ( \30387 , \30383 , \30386 );
and \U$30010 ( \30388 , \30381 , \30386 );
or \U$30011 ( \30389 , \30384 , \30387 , \30388 );
and \U$30012 ( \30390 , \30379 , \30389 );
xor \U$30013 ( \30391 , \29709 , \29750 );
xor \U$30014 ( \30392 , \30391 , \29769 );
and \U$30015 ( \30393 , \30389 , \30392 );
and \U$30016 ( \30394 , \30379 , \30392 );
or \U$30017 ( \30395 , \30390 , \30393 , \30394 );
xor \U$30018 ( \30396 , \30062 , \30072 );
xor \U$30019 ( \30397 , \30396 , \30091 );
xor \U$30020 ( \30398 , \30096 , \30098 );
xor \U$30021 ( \30399 , \30398 , \30101 );
and \U$30022 ( \30400 , \30397 , \30399 );
and \U$30023 ( \30401 , \30395 , \30400 );
xor \U$30024 ( \30402 , \29772 , \29797 );
xor \U$30025 ( \30403 , \30402 , \29808 );
and \U$30026 ( \30404 , \30400 , \30403 );
and \U$30027 ( \30405 , \30395 , \30403 );
or \U$30028 ( \30406 , \30401 , \30404 , \30405 );
xor \U$30029 ( \30407 , \30110 , \30112 );
xor \U$30030 ( \30408 , \30407 , \30115 );
and \U$30031 ( \30409 , \30406 , \30408 );
and \U$30032 ( \30410 , \30124 , \30409 );
xor \U$30033 ( \30411 , \30124 , \30409 );
xor \U$30034 ( \30412 , \30406 , \30408 );
xor \U$30035 ( \30413 , \30180 , \30184 );
xor \U$30036 ( \30414 , \30413 , \30189 );
xor \U$30037 ( \30415 , \30196 , \30200 );
xor \U$30038 ( \30416 , \30415 , \30205 );
and \U$30039 ( \30417 , \30414 , \30416 );
xor \U$30040 ( \30418 , \30213 , \30217 );
xor \U$30041 ( \30419 , \30418 , \30222 );
and \U$30042 ( \30420 , \30416 , \30419 );
and \U$30043 ( \30421 , \30414 , \30419 );
or \U$30044 ( \30422 , \30417 , \30420 , \30421 );
xor \U$30045 ( \30423 , \30128 , \30132 );
xor \U$30046 ( \30424 , \30423 , \30137 );
xor \U$30047 ( \30425 , \30144 , \30148 );
xor \U$30048 ( \30426 , \30425 , \30153 );
and \U$30049 ( \30427 , \30424 , \30426 );
xor \U$30050 ( \30428 , \30161 , \30165 );
xor \U$30051 ( \30429 , \30428 , \30170 );
and \U$30052 ( \30430 , \30426 , \30429 );
and \U$30053 ( \30431 , \30424 , \30429 );
or \U$30054 ( \30432 , \30427 , \30430 , \30431 );
and \U$30055 ( \30433 , \30422 , \30432 );
and \U$30056 ( \30434 , \29464 , \21745 );
and \U$30057 ( \30435 , \29040 , \21743 );
nor \U$30058 ( \30436 , \30434 , \30435 );
xnor \U$30059 ( \30437 , \30436 , \21715 );
and \U$30060 ( \30438 , \29715 , \21697 );
and \U$30061 ( \30439 , \29710 , \21695 );
nor \U$30062 ( \30440 , \30438 , \30439 );
xnor \U$30063 ( \30441 , \30440 , \21678 );
and \U$30064 ( \30442 , \30437 , \30441 );
and \U$30065 ( \30443 , \30318 , \21660 );
and \U$30066 ( \30444 , \30034 , \21658 );
nor \U$30067 ( \30445 , \30443 , \30444 );
xnor \U$30068 ( \30446 , \30445 , \21665 );
and \U$30069 ( \30447 , \30441 , \30446 );
and \U$30070 ( \30448 , \30437 , \30446 );
or \U$30071 ( \30449 , \30442 , \30447 , \30448 );
xor \U$30072 ( \30450 , \30312 , \30316 );
xor \U$30073 ( \30451 , \30450 , \30319 );
or \U$30074 ( \30452 , \30449 , \30451 );
and \U$30075 ( \30453 , \30432 , \30452 );
and \U$30076 ( \30454 , \30422 , \30452 );
or \U$30077 ( \30455 , \30433 , \30453 , \30454 );
buf \U$30078 ( \30456 , RIc225a08_60);
buf \U$30079 ( \30457 , RIc225990_61);
and \U$30080 ( \30458 , \30456 , \30457 );
not \U$30081 ( \30459 , \30458 );
and \U$30082 ( \30460 , \29859 , \30459 );
not \U$30083 ( \30461 , \30460 );
and \U$30084 ( \30462 , \21667 , \30233 );
and \U$30085 ( \30463 , \21653 , \30231 );
nor \U$30086 ( \30464 , \30462 , \30463 );
xnor \U$30087 ( \30465 , \30464 , \29862 );
and \U$30088 ( \30466 , \30461 , \30465 );
and \U$30089 ( \30467 , \21706 , \29671 );
and \U$30090 ( \30468 , \21685 , \29669 );
nor \U$30091 ( \30469 , \30467 , \30468 );
xnor \U$30092 ( \30470 , \30469 , \29353 );
and \U$30093 ( \30471 , \30465 , \30470 );
and \U$30094 ( \30472 , \30461 , \30470 );
or \U$30095 ( \30473 , \30466 , \30471 , \30472 );
and \U$30096 ( \30474 , \22046 , \27572 );
and \U$30097 ( \30475 , \22018 , \27570 );
nor \U$30098 ( \30476 , \30474 , \30475 );
xnor \U$30099 ( \30477 , \30476 , \27232 );
and \U$30100 ( \30478 , \22200 , \26983 );
and \U$30101 ( \30479 , \22126 , \26981 );
nor \U$30102 ( \30480 , \30478 , \30479 );
xnor \U$30103 ( \30481 , \30480 , \26742 );
and \U$30104 ( \30482 , \30477 , \30481 );
and \U$30105 ( \30483 , \22325 , \26517 );
and \U$30106 ( \30484 , \22262 , \26515 );
nor \U$30107 ( \30485 , \30483 , \30484 );
xnor \U$30108 ( \30486 , \30485 , \26329 );
and \U$30109 ( \30487 , \30481 , \30486 );
and \U$30110 ( \30488 , \30477 , \30486 );
or \U$30111 ( \30489 , \30482 , \30487 , \30488 );
and \U$30112 ( \30490 , \30473 , \30489 );
and \U$30113 ( \30491 , \21762 , \29104 );
and \U$30114 ( \30492 , \21754 , \29102 );
nor \U$30115 ( \30493 , \30491 , \30492 );
xnor \U$30116 ( \30494 , \30493 , \28855 );
and \U$30117 ( \30495 , \21836 , \28575 );
and \U$30118 ( \30496 , \21831 , \28573 );
nor \U$30119 ( \30497 , \30495 , \30496 );
xnor \U$30120 ( \30498 , \30497 , \28315 );
and \U$30121 ( \30499 , \30494 , \30498 );
and \U$30122 ( \30500 , \21941 , \28081 );
and \U$30123 ( \30501 , \21890 , \28079 );
nor \U$30124 ( \30502 , \30500 , \30501 );
xnor \U$30125 ( \30503 , \30502 , \27766 );
and \U$30126 ( \30504 , \30498 , \30503 );
and \U$30127 ( \30505 , \30494 , \30503 );
or \U$30128 ( \30506 , \30499 , \30504 , \30505 );
and \U$30129 ( \30507 , \30489 , \30506 );
and \U$30130 ( \30508 , \30473 , \30506 );
or \U$30131 ( \30509 , \30490 , \30507 , \30508 );
and \U$30132 ( \30510 , \23136 , \24974 );
and \U$30133 ( \30511 , \23128 , \24972 );
nor \U$30134 ( \30512 , \30510 , \30511 );
xnor \U$30135 ( \30513 , \30512 , \24787 );
and \U$30136 ( \30514 , \23384 , \24661 );
and \U$30137 ( \30515 , \23379 , \24659 );
nor \U$30138 ( \30516 , \30514 , \30515 );
xnor \U$30139 ( \30517 , \30516 , \24456 );
and \U$30140 ( \30518 , \30513 , \30517 );
and \U$30141 ( \30519 , \23714 , \24255 );
and \U$30142 ( \30520 , \23570 , \24253 );
nor \U$30143 ( \30521 , \30519 , \30520 );
xnor \U$30144 ( \30522 , \30521 , \24106 );
and \U$30145 ( \30523 , \30517 , \30522 );
and \U$30146 ( \30524 , \30513 , \30522 );
or \U$30147 ( \30525 , \30518 , \30523 , \30524 );
and \U$30148 ( \30526 , \24003 , \23933 );
and \U$30149 ( \30527 , \23978 , \23931 );
nor \U$30150 ( \30528 , \30526 , \30527 );
xnor \U$30151 ( \30529 , \30528 , \23791 );
and \U$30152 ( \30530 , \24344 , \23637 );
and \U$30153 ( \30531 , \24177 , \23635 );
nor \U$30154 ( \30532 , \30530 , \30531 );
xnor \U$30155 ( \30533 , \30532 , \23500 );
and \U$30156 ( \30534 , \30529 , \30533 );
and \U$30157 ( \30535 , \24601 , \23431 );
and \U$30158 ( \30536 , \24482 , \23429 );
nor \U$30159 ( \30537 , \30535 , \30536 );
xnor \U$30160 ( \30538 , \30537 , \23279 );
and \U$30161 ( \30539 , \30533 , \30538 );
and \U$30162 ( \30540 , \30529 , \30538 );
or \U$30163 ( \30541 , \30534 , \30539 , \30540 );
and \U$30164 ( \30542 , \30525 , \30541 );
and \U$30165 ( \30543 , \22611 , \26143 );
and \U$30166 ( \30544 , \22523 , \26141 );
nor \U$30167 ( \30545 , \30543 , \30544 );
xnor \U$30168 ( \30546 , \30545 , \25911 );
and \U$30169 ( \30547 , \22721 , \25692 );
and \U$30170 ( \30548 , \22716 , \25690 );
nor \U$30171 ( \30549 , \30547 , \30548 );
xnor \U$30172 ( \30550 , \30549 , \25549 );
and \U$30173 ( \30551 , \30546 , \30550 );
and \U$30174 ( \30552 , \22952 , \25369 );
and \U$30175 ( \30553 , \22837 , \25367 );
nor \U$30176 ( \30554 , \30552 , \30553 );
xnor \U$30177 ( \30555 , \30554 , \25123 );
and \U$30178 ( \30556 , \30550 , \30555 );
and \U$30179 ( \30557 , \30546 , \30555 );
or \U$30180 ( \30558 , \30551 , \30556 , \30557 );
and \U$30181 ( \30559 , \30541 , \30558 );
and \U$30182 ( \30560 , \30525 , \30558 );
or \U$30183 ( \30561 , \30542 , \30559 , \30560 );
and \U$30184 ( \30562 , \30509 , \30561 );
and \U$30185 ( \30563 , \27494 , \22029 );
and \U$30186 ( \30564 , \27485 , \22027 );
nor \U$30187 ( \30565 , \30563 , \30564 );
xnor \U$30188 ( \30566 , \30565 , \21986 );
and \U$30189 ( \30567 , \28039 , \21916 );
and \U$30190 ( \30568 , \27837 , \21914 );
nor \U$30191 ( \30569 , \30567 , \30568 );
xnor \U$30192 ( \30570 , \30569 , \21867 );
and \U$30193 ( \30571 , \30566 , \30570 );
and \U$30194 ( \30572 , \28514 , \21815 );
and \U$30195 ( \30573 , \28342 , \21813 );
nor \U$30196 ( \30574 , \30572 , \30573 );
xnor \U$30197 ( \30575 , \30574 , \21774 );
and \U$30198 ( \30576 , \30570 , \30575 );
and \U$30199 ( \30577 , \30566 , \30575 );
or \U$30200 ( \30578 , \30571 , \30576 , \30577 );
and \U$30201 ( \30579 , \26116 , \22497 );
and \U$30202 ( \30580 , \26108 , \22495 );
nor \U$30203 ( \30581 , \30579 , \30580 );
xnor \U$30204 ( \30582 , \30581 , \22419 );
and \U$30205 ( \30583 , \26590 , \22333 );
and \U$30206 ( \30584 , \26585 , \22331 );
nor \U$30207 ( \30585 , \30583 , \30584 );
xnor \U$30208 ( \30586 , \30585 , \22239 );
and \U$30209 ( \30587 , \30582 , \30586 );
and \U$30210 ( \30588 , \27113 , \22163 );
and \U$30211 ( \30589 , \26854 , \22161 );
nor \U$30212 ( \30590 , \30588 , \30589 );
xnor \U$30213 ( \30591 , \30590 , \22091 );
and \U$30214 ( \30592 , \30586 , \30591 );
and \U$30215 ( \30593 , \30582 , \30591 );
or \U$30216 ( \30594 , \30587 , \30592 , \30593 );
and \U$30217 ( \30595 , \30578 , \30594 );
and \U$30218 ( \30596 , \25226 , \23163 );
and \U$30219 ( \30597 , \25018 , \23161 );
nor \U$30220 ( \30598 , \30596 , \30597 );
xnor \U$30221 ( \30599 , \30598 , \23007 );
and \U$30222 ( \30600 , \25353 , \22891 );
and \U$30223 ( \30601 , \25348 , \22889 );
nor \U$30224 ( \30602 , \30600 , \30601 );
xnor \U$30225 ( \30603 , \30602 , \22778 );
and \U$30226 ( \30604 , \30599 , \30603 );
and \U$30227 ( \30605 , \25806 , \22697 );
and \U$30228 ( \30606 , \25609 , \22695 );
nor \U$30229 ( \30607 , \30605 , \30606 );
xnor \U$30230 ( \30608 , \30607 , \22561 );
and \U$30231 ( \30609 , \30603 , \30608 );
and \U$30232 ( \30610 , \30599 , \30608 );
or \U$30233 ( \30611 , \30604 , \30609 , \30610 );
and \U$30234 ( \30612 , \30594 , \30611 );
and \U$30235 ( \30613 , \30578 , \30611 );
or \U$30236 ( \30614 , \30595 , \30612 , \30613 );
and \U$30237 ( \30615 , \30561 , \30614 );
and \U$30238 ( \30616 , \30509 , \30614 );
or \U$30239 ( \30617 , \30562 , \30615 , \30616 );
and \U$30240 ( \30618 , \30455 , \30617 );
xor \U$30241 ( \30619 , \30236 , \30240 );
xor \U$30242 ( \30620 , \30619 , \30245 );
xor \U$30243 ( \30621 , \30252 , \30256 );
xor \U$30244 ( \30622 , \30621 , \30261 );
and \U$30245 ( \30623 , \30620 , \30622 );
xor \U$30246 ( \30624 , \30269 , \30273 );
xor \U$30247 ( \30625 , \30624 , \30278 );
and \U$30248 ( \30626 , \30622 , \30625 );
and \U$30249 ( \30627 , \30620 , \30625 );
or \U$30250 ( \30628 , \30623 , \30626 , \30627 );
xor \U$30251 ( \30629 , \29845 , \29849 );
xor \U$30252 ( \30630 , \30629 , \29854 );
and \U$30253 ( \30631 , \30628 , \30630 );
xor \U$30254 ( \30632 , \29863 , \29867 );
xor \U$30255 ( \30633 , \30632 , \29872 );
and \U$30256 ( \30634 , \30630 , \30633 );
and \U$30257 ( \30635 , \30628 , \30633 );
or \U$30258 ( \30636 , \30631 , \30634 , \30635 );
and \U$30259 ( \30637 , \30617 , \30636 );
and \U$30260 ( \30638 , \30455 , \30636 );
or \U$30261 ( \30639 , \30618 , \30637 , \30638 );
xor \U$30262 ( \30640 , \30140 , \30156 );
xor \U$30263 ( \30641 , \30640 , \30173 );
xor \U$30264 ( \30642 , \30192 , \30208 );
xor \U$30265 ( \30643 , \30642 , \30225 );
and \U$30266 ( \30644 , \30641 , \30643 );
xor \U$30267 ( \30645 , \30248 , \30264 );
xor \U$30268 ( \30646 , \30645 , \30281 );
and \U$30269 ( \30647 , \30643 , \30646 );
and \U$30270 ( \30648 , \30641 , \30646 );
or \U$30271 ( \30649 , \30644 , \30647 , \30648 );
xor \U$30272 ( \30650 , \30289 , \30291 );
xor \U$30273 ( \30651 , \30650 , \30294 );
xor \U$30274 ( \30652 , \30299 , \30301 );
xor \U$30275 ( \30653 , \30652 , \30304 );
and \U$30276 ( \30654 , \30651 , \30653 );
xor \U$30277 ( \30655 , \30322 , \30324 );
xor \U$30278 ( \30656 , \30655 , \30327 );
and \U$30279 ( \30657 , \30653 , \30656 );
and \U$30280 ( \30658 , \30651 , \30656 );
or \U$30281 ( \30659 , \30654 , \30657 , \30658 );
and \U$30282 ( \30660 , \30649 , \30659 );
xor \U$30283 ( \30661 , \29911 , \29927 );
xor \U$30284 ( \30662 , \30661 , \29944 );
and \U$30285 ( \30663 , \30659 , \30662 );
and \U$30286 ( \30664 , \30649 , \30662 );
or \U$30287 ( \30665 , \30660 , \30663 , \30664 );
and \U$30288 ( \30666 , \30639 , \30665 );
xor \U$30289 ( \30667 , \29857 , \29875 );
xor \U$30290 ( \30668 , \30667 , \29892 );
xor \U$30291 ( \30669 , \30336 , \30338 );
xor \U$30292 ( \30670 , \30669 , \30341 );
and \U$30293 ( \30671 , \30668 , \30670 );
xor \U$30294 ( \30672 , \30349 , \30351 );
xor \U$30295 ( \30673 , \30672 , \30354 );
and \U$30296 ( \30674 , \30670 , \30673 );
and \U$30297 ( \30675 , \30668 , \30673 );
or \U$30298 ( \30676 , \30671 , \30674 , \30675 );
and \U$30299 ( \30677 , \30665 , \30676 );
and \U$30300 ( \30678 , \30639 , \30676 );
or \U$30301 ( \30679 , \30666 , \30677 , \30678 );
xor \U$30302 ( \30680 , \30287 , \30333 );
xor \U$30303 ( \30681 , \30680 , \30344 );
xor \U$30304 ( \30682 , \30357 , \30359 );
xor \U$30305 ( \30683 , \30682 , \30362 );
and \U$30306 ( \30684 , \30681 , \30683 );
xor \U$30307 ( \30685 , \30368 , \30370 );
xor \U$30308 ( \30686 , \30685 , \30373 );
and \U$30309 ( \30687 , \30683 , \30686 );
and \U$30310 ( \30688 , \30681 , \30686 );
or \U$30311 ( \30689 , \30684 , \30687 , \30688 );
and \U$30312 ( \30690 , \30679 , \30689 );
xor \U$30313 ( \30691 , \30381 , \30383 );
xor \U$30314 ( \30692 , \30691 , \30386 );
and \U$30315 ( \30693 , \30689 , \30692 );
and \U$30316 ( \30694 , \30679 , \30692 );
or \U$30317 ( \30695 , \30690 , \30693 , \30694 );
xor \U$30318 ( \30696 , \30379 , \30389 );
xor \U$30319 ( \30697 , \30696 , \30392 );
and \U$30320 ( \30698 , \30695 , \30697 );
xor \U$30321 ( \30699 , \30397 , \30399 );
and \U$30322 ( \30700 , \30697 , \30699 );
and \U$30323 ( \30701 , \30695 , \30699 );
or \U$30324 ( \30702 , \30698 , \30700 , \30701 );
xor \U$30325 ( \30703 , \30395 , \30400 );
xor \U$30326 ( \30704 , \30703 , \30403 );
and \U$30327 ( \30705 , \30702 , \30704 );
xor \U$30328 ( \30706 , \30094 , \30104 );
xor \U$30329 ( \30707 , \30706 , \30107 );
and \U$30330 ( \30708 , \30704 , \30707 );
and \U$30331 ( \30709 , \30702 , \30707 );
or \U$30332 ( \30710 , \30705 , \30708 , \30709 );
and \U$30333 ( \30711 , \30412 , \30710 );
xor \U$30334 ( \30712 , \30412 , \30710 );
xor \U$30335 ( \30713 , \30702 , \30704 );
xor \U$30336 ( \30714 , \30713 , \30707 );
and \U$30337 ( \30715 , \26585 , \22497 );
and \U$30338 ( \30716 , \26116 , \22495 );
nor \U$30339 ( \30717 , \30715 , \30716 );
xnor \U$30340 ( \30718 , \30717 , \22419 );
and \U$30341 ( \30719 , \26854 , \22333 );
and \U$30342 ( \30720 , \26590 , \22331 );
nor \U$30343 ( \30721 , \30719 , \30720 );
xnor \U$30344 ( \30722 , \30721 , \22239 );
and \U$30345 ( \30723 , \30718 , \30722 );
and \U$30346 ( \30724 , \27485 , \22163 );
and \U$30347 ( \30725 , \27113 , \22161 );
nor \U$30348 ( \30726 , \30724 , \30725 );
xnor \U$30349 ( \30727 , \30726 , \22091 );
and \U$30350 ( \30728 , \30722 , \30727 );
and \U$30351 ( \30729 , \30718 , \30727 );
or \U$30352 ( \30730 , \30723 , \30728 , \30729 );
and \U$30353 ( \30731 , \25348 , \23163 );
and \U$30354 ( \30732 , \25226 , \23161 );
nor \U$30355 ( \30733 , \30731 , \30732 );
xnor \U$30356 ( \30734 , \30733 , \23007 );
and \U$30357 ( \30735 , \25609 , \22891 );
and \U$30358 ( \30736 , \25353 , \22889 );
nor \U$30359 ( \30737 , \30735 , \30736 );
xnor \U$30360 ( \30738 , \30737 , \22778 );
and \U$30361 ( \30739 , \30734 , \30738 );
and \U$30362 ( \30740 , \26108 , \22697 );
and \U$30363 ( \30741 , \25806 , \22695 );
nor \U$30364 ( \30742 , \30740 , \30741 );
xnor \U$30365 ( \30743 , \30742 , \22561 );
and \U$30366 ( \30744 , \30738 , \30743 );
and \U$30367 ( \30745 , \30734 , \30743 );
or \U$30368 ( \30746 , \30739 , \30744 , \30745 );
and \U$30369 ( \30747 , \30730 , \30746 );
and \U$30370 ( \30748 , \27837 , \22029 );
and \U$30371 ( \30749 , \27494 , \22027 );
nor \U$30372 ( \30750 , \30748 , \30749 );
xnor \U$30373 ( \30751 , \30750 , \21986 );
and \U$30374 ( \30752 , \28342 , \21916 );
and \U$30375 ( \30753 , \28039 , \21914 );
nor \U$30376 ( \30754 , \30752 , \30753 );
xnor \U$30377 ( \30755 , \30754 , \21867 );
and \U$30378 ( \30756 , \30751 , \30755 );
and \U$30379 ( \30757 , \29040 , \21815 );
and \U$30380 ( \30758 , \28514 , \21813 );
nor \U$30381 ( \30759 , \30757 , \30758 );
xnor \U$30382 ( \30760 , \30759 , \21774 );
and \U$30383 ( \30761 , \30755 , \30760 );
and \U$30384 ( \30762 , \30751 , \30760 );
or \U$30385 ( \30763 , \30756 , \30761 , \30762 );
and \U$30386 ( \30764 , \30746 , \30763 );
and \U$30387 ( \30765 , \30730 , \30763 );
or \U$30388 ( \30766 , \30747 , \30764 , \30765 );
xor \U$30389 ( \30767 , \29859 , \30456 );
xor \U$30390 ( \30768 , \30456 , \30457 );
not \U$30391 ( \30769 , \30768 );
and \U$30392 ( \30770 , \30767 , \30769 );
and \U$30393 ( \30771 , \21653 , \30770 );
not \U$30394 ( \30772 , \30771 );
xnor \U$30395 ( \30773 , \30772 , \30460 );
and \U$30396 ( \30774 , \21685 , \30233 );
and \U$30397 ( \30775 , \21667 , \30231 );
nor \U$30398 ( \30776 , \30774 , \30775 );
xnor \U$30399 ( \30777 , \30776 , \29862 );
and \U$30400 ( \30778 , \30773 , \30777 );
and \U$30401 ( \30779 , \21754 , \29671 );
and \U$30402 ( \30780 , \21706 , \29669 );
nor \U$30403 ( \30781 , \30779 , \30780 );
xnor \U$30404 ( \30782 , \30781 , \29353 );
and \U$30405 ( \30783 , \30777 , \30782 );
and \U$30406 ( \30784 , \30773 , \30782 );
or \U$30407 ( \30785 , \30778 , \30783 , \30784 );
and \U$30408 ( \30786 , \22126 , \27572 );
and \U$30409 ( \30787 , \22046 , \27570 );
nor \U$30410 ( \30788 , \30786 , \30787 );
xnor \U$30411 ( \30789 , \30788 , \27232 );
and \U$30412 ( \30790 , \22262 , \26983 );
and \U$30413 ( \30791 , \22200 , \26981 );
nor \U$30414 ( \30792 , \30790 , \30791 );
xnor \U$30415 ( \30793 , \30792 , \26742 );
and \U$30416 ( \30794 , \30789 , \30793 );
and \U$30417 ( \30795 , \22523 , \26517 );
and \U$30418 ( \30796 , \22325 , \26515 );
nor \U$30419 ( \30797 , \30795 , \30796 );
xnor \U$30420 ( \30798 , \30797 , \26329 );
and \U$30421 ( \30799 , \30793 , \30798 );
and \U$30422 ( \30800 , \30789 , \30798 );
or \U$30423 ( \30801 , \30794 , \30799 , \30800 );
and \U$30424 ( \30802 , \30785 , \30801 );
and \U$30425 ( \30803 , \21831 , \29104 );
and \U$30426 ( \30804 , \21762 , \29102 );
nor \U$30427 ( \30805 , \30803 , \30804 );
xnor \U$30428 ( \30806 , \30805 , \28855 );
and \U$30429 ( \30807 , \21890 , \28575 );
and \U$30430 ( \30808 , \21836 , \28573 );
nor \U$30431 ( \30809 , \30807 , \30808 );
xnor \U$30432 ( \30810 , \30809 , \28315 );
and \U$30433 ( \30811 , \30806 , \30810 );
and \U$30434 ( \30812 , \22018 , \28081 );
and \U$30435 ( \30813 , \21941 , \28079 );
nor \U$30436 ( \30814 , \30812 , \30813 );
xnor \U$30437 ( \30815 , \30814 , \27766 );
and \U$30438 ( \30816 , \30810 , \30815 );
and \U$30439 ( \30817 , \30806 , \30815 );
or \U$30440 ( \30818 , \30811 , \30816 , \30817 );
and \U$30441 ( \30819 , \30801 , \30818 );
and \U$30442 ( \30820 , \30785 , \30818 );
or \U$30443 ( \30821 , \30802 , \30819 , \30820 );
and \U$30444 ( \30822 , \30766 , \30821 );
and \U$30445 ( \30823 , \22716 , \26143 );
and \U$30446 ( \30824 , \22611 , \26141 );
nor \U$30447 ( \30825 , \30823 , \30824 );
xnor \U$30448 ( \30826 , \30825 , \25911 );
and \U$30449 ( \30827 , \22837 , \25692 );
and \U$30450 ( \30828 , \22721 , \25690 );
nor \U$30451 ( \30829 , \30827 , \30828 );
xnor \U$30452 ( \30830 , \30829 , \25549 );
and \U$30453 ( \30831 , \30826 , \30830 );
and \U$30454 ( \30832 , \23128 , \25369 );
and \U$30455 ( \30833 , \22952 , \25367 );
nor \U$30456 ( \30834 , \30832 , \30833 );
xnor \U$30457 ( \30835 , \30834 , \25123 );
and \U$30458 ( \30836 , \30830 , \30835 );
and \U$30459 ( \30837 , \30826 , \30835 );
or \U$30460 ( \30838 , \30831 , \30836 , \30837 );
and \U$30461 ( \30839 , \24177 , \23933 );
and \U$30462 ( \30840 , \24003 , \23931 );
nor \U$30463 ( \30841 , \30839 , \30840 );
xnor \U$30464 ( \30842 , \30841 , \23791 );
and \U$30465 ( \30843 , \24482 , \23637 );
and \U$30466 ( \30844 , \24344 , \23635 );
nor \U$30467 ( \30845 , \30843 , \30844 );
xnor \U$30468 ( \30846 , \30845 , \23500 );
and \U$30469 ( \30847 , \30842 , \30846 );
and \U$30470 ( \30848 , \25018 , \23431 );
and \U$30471 ( \30849 , \24601 , \23429 );
nor \U$30472 ( \30850 , \30848 , \30849 );
xnor \U$30473 ( \30851 , \30850 , \23279 );
and \U$30474 ( \30852 , \30846 , \30851 );
and \U$30475 ( \30853 , \30842 , \30851 );
or \U$30476 ( \30854 , \30847 , \30852 , \30853 );
and \U$30477 ( \30855 , \30838 , \30854 );
and \U$30478 ( \30856 , \23379 , \24974 );
and \U$30479 ( \30857 , \23136 , \24972 );
nor \U$30480 ( \30858 , \30856 , \30857 );
xnor \U$30481 ( \30859 , \30858 , \24787 );
and \U$30482 ( \30860 , \23570 , \24661 );
and \U$30483 ( \30861 , \23384 , \24659 );
nor \U$30484 ( \30862 , \30860 , \30861 );
xnor \U$30485 ( \30863 , \30862 , \24456 );
and \U$30486 ( \30864 , \30859 , \30863 );
and \U$30487 ( \30865 , \23978 , \24255 );
and \U$30488 ( \30866 , \23714 , \24253 );
nor \U$30489 ( \30867 , \30865 , \30866 );
xnor \U$30490 ( \30868 , \30867 , \24106 );
and \U$30491 ( \30869 , \30863 , \30868 );
and \U$30492 ( \30870 , \30859 , \30868 );
or \U$30493 ( \30871 , \30864 , \30869 , \30870 );
and \U$30494 ( \30872 , \30854 , \30871 );
and \U$30495 ( \30873 , \30838 , \30871 );
or \U$30496 ( \30874 , \30855 , \30872 , \30873 );
and \U$30497 ( \30875 , \30821 , \30874 );
and \U$30498 ( \30876 , \30766 , \30874 );
or \U$30499 ( \30877 , \30822 , \30875 , \30876 );
and \U$30500 ( \30878 , \29710 , \21745 );
and \U$30501 ( \30879 , \29464 , \21743 );
nor \U$30502 ( \30880 , \30878 , \30879 );
xnor \U$30503 ( \30881 , \30880 , \21715 );
and \U$30504 ( \30882 , \30034 , \21697 );
and \U$30505 ( \30883 , \29715 , \21695 );
nor \U$30506 ( \30884 , \30882 , \30883 );
xnor \U$30507 ( \30885 , \30884 , \21678 );
and \U$30508 ( \30886 , \30881 , \30885 );
buf \U$30509 ( \30887 , RIc22b0c0_187);
and \U$30510 ( \30888 , \30887 , \21660 );
and \U$30511 ( \30889 , \30318 , \21658 );
nor \U$30512 ( \30890 , \30888 , \30889 );
xnor \U$30513 ( \30891 , \30890 , \21665 );
and \U$30514 ( \30892 , \30885 , \30891 );
and \U$30515 ( \30893 , \30881 , \30891 );
or \U$30516 ( \30894 , \30886 , \30892 , \30893 );
buf \U$30517 ( \30895 , RIc22b138_188);
and \U$30518 ( \30896 , \30895 , \21654 );
buf \U$30519 ( \30897 , \30896 );
and \U$30520 ( \30898 , \30894 , \30897 );
and \U$30521 ( \30899 , \30887 , \21654 );
and \U$30522 ( \30900 , \30897 , \30899 );
and \U$30523 ( \30901 , \30894 , \30899 );
or \U$30524 ( \30902 , \30898 , \30900 , \30901 );
xor \U$30525 ( \30903 , \30437 , \30441 );
xor \U$30526 ( \30904 , \30903 , \30446 );
xor \U$30527 ( \30905 , \30566 , \30570 );
xor \U$30528 ( \30906 , \30905 , \30575 );
and \U$30529 ( \30907 , \30904 , \30906 );
xor \U$30530 ( \30908 , \30582 , \30586 );
xor \U$30531 ( \30909 , \30908 , \30591 );
and \U$30532 ( \30910 , \30906 , \30909 );
and \U$30533 ( \30911 , \30904 , \30909 );
or \U$30534 ( \30912 , \30907 , \30910 , \30911 );
and \U$30535 ( \30913 , \30902 , \30912 );
xor \U$30536 ( \30914 , \30599 , \30603 );
xor \U$30537 ( \30915 , \30914 , \30608 );
xor \U$30538 ( \30916 , \30513 , \30517 );
xor \U$30539 ( \30917 , \30916 , \30522 );
and \U$30540 ( \30918 , \30915 , \30917 );
xor \U$30541 ( \30919 , \30529 , \30533 );
xor \U$30542 ( \30920 , \30919 , \30538 );
and \U$30543 ( \30921 , \30917 , \30920 );
and \U$30544 ( \30922 , \30915 , \30920 );
or \U$30545 ( \30923 , \30918 , \30921 , \30922 );
and \U$30546 ( \30924 , \30912 , \30923 );
and \U$30547 ( \30925 , \30902 , \30923 );
or \U$30548 ( \30926 , \30913 , \30924 , \30925 );
and \U$30549 ( \30927 , \30877 , \30926 );
xor \U$30550 ( \30928 , \30477 , \30481 );
xor \U$30551 ( \30929 , \30928 , \30486 );
xor \U$30552 ( \30930 , \30494 , \30498 );
xor \U$30553 ( \30931 , \30930 , \30503 );
and \U$30554 ( \30932 , \30929 , \30931 );
xor \U$30555 ( \30933 , \30546 , \30550 );
xor \U$30556 ( \30934 , \30933 , \30555 );
and \U$30557 ( \30935 , \30931 , \30934 );
and \U$30558 ( \30936 , \30929 , \30934 );
or \U$30559 ( \30937 , \30932 , \30935 , \30936 );
xor \U$30560 ( \30938 , \30620 , \30622 );
xor \U$30561 ( \30939 , \30938 , \30625 );
and \U$30562 ( \30940 , \30937 , \30939 );
xor \U$30563 ( \30941 , \30424 , \30426 );
xor \U$30564 ( \30942 , \30941 , \30429 );
and \U$30565 ( \30943 , \30939 , \30942 );
and \U$30566 ( \30944 , \30937 , \30942 );
or \U$30567 ( \30945 , \30940 , \30943 , \30944 );
and \U$30568 ( \30946 , \30926 , \30945 );
and \U$30569 ( \30947 , \30877 , \30945 );
or \U$30570 ( \30948 , \30927 , \30946 , \30947 );
xor \U$30571 ( \30949 , \30422 , \30432 );
xor \U$30572 ( \30950 , \30949 , \30452 );
xor \U$30573 ( \30951 , \30509 , \30561 );
xor \U$30574 ( \30952 , \30951 , \30614 );
and \U$30575 ( \30953 , \30950 , \30952 );
xor \U$30576 ( \30954 , \30628 , \30630 );
xor \U$30577 ( \30955 , \30954 , \30633 );
and \U$30578 ( \30956 , \30952 , \30955 );
and \U$30579 ( \30957 , \30950 , \30955 );
or \U$30580 ( \30958 , \30953 , \30956 , \30957 );
and \U$30581 ( \30959 , \30948 , \30958 );
xor \U$30582 ( \30960 , \30578 , \30594 );
xor \U$30583 ( \30961 , \30960 , \30611 );
xor \U$30584 ( \30962 , \30414 , \30416 );
xor \U$30585 ( \30963 , \30962 , \30419 );
and \U$30586 ( \30964 , \30961 , \30963 );
xnor \U$30587 ( \30965 , \30449 , \30451 );
and \U$30588 ( \30966 , \30963 , \30965 );
and \U$30589 ( \30967 , \30961 , \30965 );
or \U$30590 ( \30968 , \30964 , \30966 , \30967 );
xor \U$30591 ( \30969 , \30641 , \30643 );
xor \U$30592 ( \30970 , \30969 , \30646 );
and \U$30593 ( \30971 , \30968 , \30970 );
xor \U$30594 ( \30972 , \30651 , \30653 );
xor \U$30595 ( \30973 , \30972 , \30656 );
and \U$30596 ( \30974 , \30970 , \30973 );
and \U$30597 ( \30975 , \30968 , \30973 );
or \U$30598 ( \30976 , \30971 , \30974 , \30975 );
and \U$30599 ( \30977 , \30958 , \30976 );
and \U$30600 ( \30978 , \30948 , \30976 );
or \U$30601 ( \30979 , \30959 , \30977 , \30978 );
xor \U$30602 ( \30980 , \30176 , \30228 );
xor \U$30603 ( \30981 , \30980 , \30284 );
xor \U$30604 ( \30982 , \30297 , \30307 );
xor \U$30605 ( \30983 , \30982 , \30330 );
and \U$30606 ( \30984 , \30981 , \30983 );
xor \U$30607 ( \30985 , \30668 , \30670 );
xor \U$30608 ( \30986 , \30985 , \30673 );
and \U$30609 ( \30987 , \30983 , \30986 );
and \U$30610 ( \30988 , \30981 , \30986 );
or \U$30611 ( \30989 , \30984 , \30987 , \30988 );
and \U$30612 ( \30990 , \30979 , \30989 );
xor \U$30613 ( \30991 , \30681 , \30683 );
xor \U$30614 ( \30992 , \30991 , \30686 );
and \U$30615 ( \30993 , \30989 , \30992 );
and \U$30616 ( \30994 , \30979 , \30992 );
or \U$30617 ( \30995 , \30990 , \30993 , \30994 );
xor \U$30618 ( \30996 , \30347 , \30365 );
xor \U$30619 ( \30997 , \30996 , \30376 );
and \U$30620 ( \30998 , \30995 , \30997 );
xor \U$30621 ( \30999 , \30679 , \30689 );
xor \U$30622 ( \31000 , \30999 , \30692 );
and \U$30623 ( \31001 , \30997 , \31000 );
and \U$30624 ( \31002 , \30995 , \31000 );
or \U$30625 ( \31003 , \30998 , \31001 , \31002 );
xor \U$30626 ( \31004 , \30695 , \30697 );
xor \U$30627 ( \31005 , \31004 , \30699 );
and \U$30628 ( \31006 , \31003 , \31005 );
and \U$30629 ( \31007 , \30714 , \31006 );
xor \U$30630 ( \31008 , \30714 , \31006 );
xor \U$30631 ( \31009 , \31003 , \31005 );
and \U$30632 ( \31010 , \24003 , \24255 );
and \U$30633 ( \31011 , \23978 , \24253 );
nor \U$30634 ( \31012 , \31010 , \31011 );
xnor \U$30635 ( \31013 , \31012 , \24106 );
and \U$30636 ( \31014 , \24344 , \23933 );
and \U$30637 ( \31015 , \24177 , \23931 );
nor \U$30638 ( \31016 , \31014 , \31015 );
xnor \U$30639 ( \31017 , \31016 , \23791 );
and \U$30640 ( \31018 , \31013 , \31017 );
and \U$30641 ( \31019 , \24601 , \23637 );
and \U$30642 ( \31020 , \24482 , \23635 );
nor \U$30643 ( \31021 , \31019 , \31020 );
xnor \U$30644 ( \31022 , \31021 , \23500 );
and \U$30645 ( \31023 , \31017 , \31022 );
and \U$30646 ( \31024 , \31013 , \31022 );
or \U$30647 ( \31025 , \31018 , \31023 , \31024 );
and \U$30648 ( \31026 , \23136 , \25369 );
and \U$30649 ( \31027 , \23128 , \25367 );
nor \U$30650 ( \31028 , \31026 , \31027 );
xnor \U$30651 ( \31029 , \31028 , \25123 );
and \U$30652 ( \31030 , \23384 , \24974 );
and \U$30653 ( \31031 , \23379 , \24972 );
nor \U$30654 ( \31032 , \31030 , \31031 );
xnor \U$30655 ( \31033 , \31032 , \24787 );
and \U$30656 ( \31034 , \31029 , \31033 );
and \U$30657 ( \31035 , \23714 , \24661 );
and \U$30658 ( \31036 , \23570 , \24659 );
nor \U$30659 ( \31037 , \31035 , \31036 );
xnor \U$30660 ( \31038 , \31037 , \24456 );
and \U$30661 ( \31039 , \31033 , \31038 );
and \U$30662 ( \31040 , \31029 , \31038 );
or \U$30663 ( \31041 , \31034 , \31039 , \31040 );
and \U$30664 ( \31042 , \31025 , \31041 );
and \U$30665 ( \31043 , \22611 , \26517 );
and \U$30666 ( \31044 , \22523 , \26515 );
nor \U$30667 ( \31045 , \31043 , \31044 );
xnor \U$30668 ( \31046 , \31045 , \26329 );
and \U$30669 ( \31047 , \22721 , \26143 );
and \U$30670 ( \31048 , \22716 , \26141 );
nor \U$30671 ( \31049 , \31047 , \31048 );
xnor \U$30672 ( \31050 , \31049 , \25911 );
and \U$30673 ( \31051 , \31046 , \31050 );
and \U$30674 ( \31052 , \22952 , \25692 );
and \U$30675 ( \31053 , \22837 , \25690 );
nor \U$30676 ( \31054 , \31052 , \31053 );
xnor \U$30677 ( \31055 , \31054 , \25549 );
and \U$30678 ( \31056 , \31050 , \31055 );
and \U$30679 ( \31057 , \31046 , \31055 );
or \U$30680 ( \31058 , \31051 , \31056 , \31057 );
and \U$30681 ( \31059 , \31041 , \31058 );
and \U$30682 ( \31060 , \31025 , \31058 );
or \U$30683 ( \31061 , \31042 , \31059 , \31060 );
and \U$30684 ( \31062 , \22046 , \28081 );
and \U$30685 ( \31063 , \22018 , \28079 );
nor \U$30686 ( \31064 , \31062 , \31063 );
xnor \U$30687 ( \31065 , \31064 , \27766 );
and \U$30688 ( \31066 , \22200 , \27572 );
and \U$30689 ( \31067 , \22126 , \27570 );
nor \U$30690 ( \31068 , \31066 , \31067 );
xnor \U$30691 ( \31069 , \31068 , \27232 );
and \U$30692 ( \31070 , \31065 , \31069 );
and \U$30693 ( \31071 , \22325 , \26983 );
and \U$30694 ( \31072 , \22262 , \26981 );
nor \U$30695 ( \31073 , \31071 , \31072 );
xnor \U$30696 ( \31074 , \31073 , \26742 );
and \U$30697 ( \31075 , \31069 , \31074 );
and \U$30698 ( \31076 , \31065 , \31074 );
or \U$30699 ( \31077 , \31070 , \31075 , \31076 );
and \U$30700 ( \31078 , \21762 , \29671 );
and \U$30701 ( \31079 , \21754 , \29669 );
nor \U$30702 ( \31080 , \31078 , \31079 );
xnor \U$30703 ( \31081 , \31080 , \29353 );
and \U$30704 ( \31082 , \21836 , \29104 );
and \U$30705 ( \31083 , \21831 , \29102 );
nor \U$30706 ( \31084 , \31082 , \31083 );
xnor \U$30707 ( \31085 , \31084 , \28855 );
and \U$30708 ( \31086 , \31081 , \31085 );
and \U$30709 ( \31087 , \21941 , \28575 );
and \U$30710 ( \31088 , \21890 , \28573 );
nor \U$30711 ( \31089 , \31087 , \31088 );
xnor \U$30712 ( \31090 , \31089 , \28315 );
and \U$30713 ( \31091 , \31085 , \31090 );
and \U$30714 ( \31092 , \31081 , \31090 );
or \U$30715 ( \31093 , \31086 , \31091 , \31092 );
and \U$30716 ( \31094 , \31077 , \31093 );
buf \U$30717 ( \31095 , RIc225918_62);
buf \U$30718 ( \31096 , RIc2258a0_63);
and \U$30719 ( \31097 , \31095 , \31096 );
not \U$30720 ( \31098 , \31097 );
and \U$30721 ( \31099 , \30457 , \31098 );
not \U$30722 ( \31100 , \31099 );
and \U$30723 ( \31101 , \21667 , \30770 );
and \U$30724 ( \31102 , \21653 , \30768 );
nor \U$30725 ( \31103 , \31101 , \31102 );
xnor \U$30726 ( \31104 , \31103 , \30460 );
and \U$30727 ( \31105 , \31100 , \31104 );
and \U$30728 ( \31106 , \21706 , \30233 );
and \U$30729 ( \31107 , \21685 , \30231 );
nor \U$30730 ( \31108 , \31106 , \31107 );
xnor \U$30731 ( \31109 , \31108 , \29862 );
and \U$30732 ( \31110 , \31104 , \31109 );
and \U$30733 ( \31111 , \31100 , \31109 );
or \U$30734 ( \31112 , \31105 , \31110 , \31111 );
and \U$30735 ( \31113 , \31093 , \31112 );
and \U$30736 ( \31114 , \31077 , \31112 );
or \U$30737 ( \31115 , \31094 , \31113 , \31114 );
and \U$30738 ( \31116 , \31061 , \31115 );
and \U$30739 ( \31117 , \27494 , \22163 );
and \U$30740 ( \31118 , \27485 , \22161 );
nor \U$30741 ( \31119 , \31117 , \31118 );
xnor \U$30742 ( \31120 , \31119 , \22091 );
and \U$30743 ( \31121 , \28039 , \22029 );
and \U$30744 ( \31122 , \27837 , \22027 );
nor \U$30745 ( \31123 , \31121 , \31122 );
xnor \U$30746 ( \31124 , \31123 , \21986 );
and \U$30747 ( \31125 , \31120 , \31124 );
and \U$30748 ( \31126 , \28514 , \21916 );
and \U$30749 ( \31127 , \28342 , \21914 );
nor \U$30750 ( \31128 , \31126 , \31127 );
xnor \U$30751 ( \31129 , \31128 , \21867 );
and \U$30752 ( \31130 , \31124 , \31129 );
and \U$30753 ( \31131 , \31120 , \31129 );
or \U$30754 ( \31132 , \31125 , \31130 , \31131 );
and \U$30755 ( \31133 , \26116 , \22697 );
and \U$30756 ( \31134 , \26108 , \22695 );
nor \U$30757 ( \31135 , \31133 , \31134 );
xnor \U$30758 ( \31136 , \31135 , \22561 );
and \U$30759 ( \31137 , \26590 , \22497 );
and \U$30760 ( \31138 , \26585 , \22495 );
nor \U$30761 ( \31139 , \31137 , \31138 );
xnor \U$30762 ( \31140 , \31139 , \22419 );
and \U$30763 ( \31141 , \31136 , \31140 );
and \U$30764 ( \31142 , \27113 , \22333 );
and \U$30765 ( \31143 , \26854 , \22331 );
nor \U$30766 ( \31144 , \31142 , \31143 );
xnor \U$30767 ( \31145 , \31144 , \22239 );
and \U$30768 ( \31146 , \31140 , \31145 );
and \U$30769 ( \31147 , \31136 , \31145 );
or \U$30770 ( \31148 , \31141 , \31146 , \31147 );
and \U$30771 ( \31149 , \31132 , \31148 );
and \U$30772 ( \31150 , \25226 , \23431 );
and \U$30773 ( \31151 , \25018 , \23429 );
nor \U$30774 ( \31152 , \31150 , \31151 );
xnor \U$30775 ( \31153 , \31152 , \23279 );
and \U$30776 ( \31154 , \25353 , \23163 );
and \U$30777 ( \31155 , \25348 , \23161 );
nor \U$30778 ( \31156 , \31154 , \31155 );
xnor \U$30779 ( \31157 , \31156 , \23007 );
and \U$30780 ( \31158 , \31153 , \31157 );
and \U$30781 ( \31159 , \25806 , \22891 );
and \U$30782 ( \31160 , \25609 , \22889 );
nor \U$30783 ( \31161 , \31159 , \31160 );
xnor \U$30784 ( \31162 , \31161 , \22778 );
and \U$30785 ( \31163 , \31157 , \31162 );
and \U$30786 ( \31164 , \31153 , \31162 );
or \U$30787 ( \31165 , \31158 , \31163 , \31164 );
and \U$30788 ( \31166 , \31148 , \31165 );
and \U$30789 ( \31167 , \31132 , \31165 );
or \U$30790 ( \31168 , \31149 , \31166 , \31167 );
and \U$30791 ( \31169 , \31115 , \31168 );
and \U$30792 ( \31170 , \31061 , \31168 );
or \U$30793 ( \31171 , \31116 , \31169 , \31170 );
xor \U$30794 ( \31172 , \30826 , \30830 );
xor \U$30795 ( \31173 , \31172 , \30835 );
xor \U$30796 ( \31174 , \30842 , \30846 );
xor \U$30797 ( \31175 , \31174 , \30851 );
and \U$30798 ( \31176 , \31173 , \31175 );
xor \U$30799 ( \31177 , \30859 , \30863 );
xor \U$30800 ( \31178 , \31177 , \30868 );
and \U$30801 ( \31179 , \31175 , \31178 );
and \U$30802 ( \31180 , \31173 , \31178 );
or \U$30803 ( \31181 , \31176 , \31179 , \31180 );
xor \U$30804 ( \31182 , \30718 , \30722 );
xor \U$30805 ( \31183 , \31182 , \30727 );
xor \U$30806 ( \31184 , \30734 , \30738 );
xor \U$30807 ( \31185 , \31184 , \30743 );
and \U$30808 ( \31186 , \31183 , \31185 );
xor \U$30809 ( \31187 , \30751 , \30755 );
xor \U$30810 ( \31188 , \31187 , \30760 );
and \U$30811 ( \31189 , \31185 , \31188 );
and \U$30812 ( \31190 , \31183 , \31188 );
or \U$30813 ( \31191 , \31186 , \31189 , \31190 );
and \U$30814 ( \31192 , \31181 , \31191 );
and \U$30815 ( \31193 , \29464 , \21815 );
and \U$30816 ( \31194 , \29040 , \21813 );
nor \U$30817 ( \31195 , \31193 , \31194 );
xnor \U$30818 ( \31196 , \31195 , \21774 );
and \U$30819 ( \31197 , \29715 , \21745 );
and \U$30820 ( \31198 , \29710 , \21743 );
nor \U$30821 ( \31199 , \31197 , \31198 );
xnor \U$30822 ( \31200 , \31199 , \21715 );
and \U$30823 ( \31201 , \31196 , \31200 );
and \U$30824 ( \31202 , \30318 , \21697 );
and \U$30825 ( \31203 , \30034 , \21695 );
nor \U$30826 ( \31204 , \31202 , \31203 );
xnor \U$30827 ( \31205 , \31204 , \21678 );
and \U$30828 ( \31206 , \31200 , \31205 );
and \U$30829 ( \31207 , \31196 , \31205 );
or \U$30830 ( \31208 , \31201 , \31206 , \31207 );
xor \U$30831 ( \31209 , \30881 , \30885 );
xor \U$30832 ( \31210 , \31209 , \30891 );
and \U$30833 ( \31211 , \31208 , \31210 );
not \U$30834 ( \31212 , \30896 );
and \U$30835 ( \31213 , \31210 , \31212 );
and \U$30836 ( \31214 , \31208 , \31212 );
or \U$30837 ( \31215 , \31211 , \31213 , \31214 );
and \U$30838 ( \31216 , \31191 , \31215 );
and \U$30839 ( \31217 , \31181 , \31215 );
or \U$30840 ( \31218 , \31192 , \31216 , \31217 );
and \U$30841 ( \31219 , \31171 , \31218 );
xor \U$30842 ( \31220 , \30773 , \30777 );
xor \U$30843 ( \31221 , \31220 , \30782 );
xor \U$30844 ( \31222 , \30789 , \30793 );
xor \U$30845 ( \31223 , \31222 , \30798 );
and \U$30846 ( \31224 , \31221 , \31223 );
xor \U$30847 ( \31225 , \30806 , \30810 );
xor \U$30848 ( \31226 , \31225 , \30815 );
and \U$30849 ( \31227 , \31223 , \31226 );
and \U$30850 ( \31228 , \31221 , \31226 );
or \U$30851 ( \31229 , \31224 , \31227 , \31228 );
xor \U$30852 ( \31230 , \30461 , \30465 );
xor \U$30853 ( \31231 , \31230 , \30470 );
and \U$30854 ( \31232 , \31229 , \31231 );
xor \U$30855 ( \31233 , \30929 , \30931 );
xor \U$30856 ( \31234 , \31233 , \30934 );
and \U$30857 ( \31235 , \31231 , \31234 );
and \U$30858 ( \31236 , \31229 , \31234 );
or \U$30859 ( \31237 , \31232 , \31235 , \31236 );
and \U$30860 ( \31238 , \31218 , \31237 );
and \U$30861 ( \31239 , \31171 , \31237 );
or \U$30862 ( \31240 , \31219 , \31238 , \31239 );
xor \U$30863 ( \31241 , \30730 , \30746 );
xor \U$30864 ( \31242 , \31241 , \30763 );
xor \U$30865 ( \31243 , \30785 , \30801 );
xor \U$30866 ( \31244 , \31243 , \30818 );
and \U$30867 ( \31245 , \31242 , \31244 );
xor \U$30868 ( \31246 , \30838 , \30854 );
xor \U$30869 ( \31247 , \31246 , \30871 );
and \U$30870 ( \31248 , \31244 , \31247 );
and \U$30871 ( \31249 , \31242 , \31247 );
or \U$30872 ( \31250 , \31245 , \31248 , \31249 );
xor \U$30873 ( \31251 , \30894 , \30897 );
xor \U$30874 ( \31252 , \31251 , \30899 );
xor \U$30875 ( \31253 , \30904 , \30906 );
xor \U$30876 ( \31254 , \31253 , \30909 );
and \U$30877 ( \31255 , \31252 , \31254 );
xor \U$30878 ( \31256 , \30915 , \30917 );
xor \U$30879 ( \31257 , \31256 , \30920 );
and \U$30880 ( \31258 , \31254 , \31257 );
and \U$30881 ( \31259 , \31252 , \31257 );
or \U$30882 ( \31260 , \31255 , \31258 , \31259 );
and \U$30883 ( \31261 , \31250 , \31260 );
xor \U$30884 ( \31262 , \30525 , \30541 );
xor \U$30885 ( \31263 , \31262 , \30558 );
and \U$30886 ( \31264 , \31260 , \31263 );
and \U$30887 ( \31265 , \31250 , \31263 );
or \U$30888 ( \31266 , \31261 , \31264 , \31265 );
and \U$30889 ( \31267 , \31240 , \31266 );
xor \U$30890 ( \31268 , \30473 , \30489 );
xor \U$30891 ( \31269 , \31268 , \30506 );
xor \U$30892 ( \31270 , \30937 , \30939 );
xor \U$30893 ( \31271 , \31270 , \30942 );
and \U$30894 ( \31272 , \31269 , \31271 );
xor \U$30895 ( \31273 , \30961 , \30963 );
xor \U$30896 ( \31274 , \31273 , \30965 );
and \U$30897 ( \31275 , \31271 , \31274 );
and \U$30898 ( \31276 , \31269 , \31274 );
or \U$30899 ( \31277 , \31272 , \31275 , \31276 );
and \U$30900 ( \31278 , \31266 , \31277 );
and \U$30901 ( \31279 , \31240 , \31277 );
or \U$30902 ( \31280 , \31267 , \31278 , \31279 );
xor \U$30903 ( \31281 , \30877 , \30926 );
xor \U$30904 ( \31282 , \31281 , \30945 );
xor \U$30905 ( \31283 , \30950 , \30952 );
xor \U$30906 ( \31284 , \31283 , \30955 );
and \U$30907 ( \31285 , \31282 , \31284 );
xor \U$30908 ( \31286 , \30968 , \30970 );
xor \U$30909 ( \31287 , \31286 , \30973 );
and \U$30910 ( \31288 , \31284 , \31287 );
and \U$30911 ( \31289 , \31282 , \31287 );
or \U$30912 ( \31290 , \31285 , \31288 , \31289 );
and \U$30913 ( \31291 , \31280 , \31290 );
xor \U$30914 ( \31292 , \30649 , \30659 );
xor \U$30915 ( \31293 , \31292 , \30662 );
and \U$30916 ( \31294 , \31290 , \31293 );
and \U$30917 ( \31295 , \31280 , \31293 );
or \U$30918 ( \31296 , \31291 , \31294 , \31295 );
xor \U$30919 ( \31297 , \30455 , \30617 );
xor \U$30920 ( \31298 , \31297 , \30636 );
xor \U$30921 ( \31299 , \30948 , \30958 );
xor \U$30922 ( \31300 , \31299 , \30976 );
and \U$30923 ( \31301 , \31298 , \31300 );
xor \U$30924 ( \31302 , \30981 , \30983 );
xor \U$30925 ( \31303 , \31302 , \30986 );
and \U$30926 ( \31304 , \31300 , \31303 );
and \U$30927 ( \31305 , \31298 , \31303 );
or \U$30928 ( \31306 , \31301 , \31304 , \31305 );
and \U$30929 ( \31307 , \31296 , \31306 );
xor \U$30930 ( \31308 , \30639 , \30665 );
xor \U$30931 ( \31309 , \31308 , \30676 );
and \U$30932 ( \31310 , \31306 , \31309 );
and \U$30933 ( \31311 , \31296 , \31309 );
or \U$30934 ( \31312 , \31307 , \31310 , \31311 );
xor \U$30935 ( \31313 , \30995 , \30997 );
xor \U$30936 ( \31314 , \31313 , \31000 );
and \U$30937 ( \31315 , \31312 , \31314 );
and \U$30938 ( \31316 , \31009 , \31315 );
xor \U$30939 ( \31317 , \31009 , \31315 );
xor \U$30940 ( \31318 , \31312 , \31314 );
and \U$30941 ( \31319 , \22126 , \28081 );
and \U$30942 ( \31320 , \22046 , \28079 );
nor \U$30943 ( \31321 , \31319 , \31320 );
xnor \U$30944 ( \31322 , \31321 , \27766 );
and \U$30945 ( \31323 , \22262 , \27572 );
and \U$30946 ( \31324 , \22200 , \27570 );
nor \U$30947 ( \31325 , \31323 , \31324 );
xnor \U$30948 ( \31326 , \31325 , \27232 );
and \U$30949 ( \31327 , \31322 , \31326 );
and \U$30950 ( \31328 , \22523 , \26983 );
and \U$30951 ( \31329 , \22325 , \26981 );
nor \U$30952 ( \31330 , \31328 , \31329 );
xnor \U$30953 ( \31331 , \31330 , \26742 );
and \U$30954 ( \31332 , \31326 , \31331 );
and \U$30955 ( \31333 , \31322 , \31331 );
or \U$30956 ( \31334 , \31327 , \31332 , \31333 );
xor \U$30957 ( \31335 , \30457 , \31095 );
xor \U$30958 ( \31336 , \31095 , \31096 );
not \U$30959 ( \31337 , \31336 );
and \U$30960 ( \31338 , \31335 , \31337 );
and \U$30961 ( \31339 , \21653 , \31338 );
not \U$30962 ( \31340 , \31339 );
xnor \U$30963 ( \31341 , \31340 , \31099 );
and \U$30964 ( \31342 , \21685 , \30770 );
and \U$30965 ( \31343 , \21667 , \30768 );
nor \U$30966 ( \31344 , \31342 , \31343 );
xnor \U$30967 ( \31345 , \31344 , \30460 );
and \U$30968 ( \31346 , \31341 , \31345 );
and \U$30969 ( \31347 , \21754 , \30233 );
and \U$30970 ( \31348 , \21706 , \30231 );
nor \U$30971 ( \31349 , \31347 , \31348 );
xnor \U$30972 ( \31350 , \31349 , \29862 );
and \U$30973 ( \31351 , \31345 , \31350 );
and \U$30974 ( \31352 , \31341 , \31350 );
or \U$30975 ( \31353 , \31346 , \31351 , \31352 );
and \U$30976 ( \31354 , \31334 , \31353 );
and \U$30977 ( \31355 , \21831 , \29671 );
and \U$30978 ( \31356 , \21762 , \29669 );
nor \U$30979 ( \31357 , \31355 , \31356 );
xnor \U$30980 ( \31358 , \31357 , \29353 );
and \U$30981 ( \31359 , \21890 , \29104 );
and \U$30982 ( \31360 , \21836 , \29102 );
nor \U$30983 ( \31361 , \31359 , \31360 );
xnor \U$30984 ( \31362 , \31361 , \28855 );
and \U$30985 ( \31363 , \31358 , \31362 );
and \U$30986 ( \31364 , \22018 , \28575 );
and \U$30987 ( \31365 , \21941 , \28573 );
nor \U$30988 ( \31366 , \31364 , \31365 );
xnor \U$30989 ( \31367 , \31366 , \28315 );
and \U$30990 ( \31368 , \31362 , \31367 );
and \U$30991 ( \31369 , \31358 , \31367 );
or \U$30992 ( \31370 , \31363 , \31368 , \31369 );
and \U$30993 ( \31371 , \31353 , \31370 );
and \U$30994 ( \31372 , \31334 , \31370 );
or \U$30995 ( \31373 , \31354 , \31371 , \31372 );
and \U$30996 ( \31374 , \27837 , \22163 );
and \U$30997 ( \31375 , \27494 , \22161 );
nor \U$30998 ( \31376 , \31374 , \31375 );
xnor \U$30999 ( \31377 , \31376 , \22091 );
and \U$31000 ( \31378 , \28342 , \22029 );
and \U$31001 ( \31379 , \28039 , \22027 );
nor \U$31002 ( \31380 , \31378 , \31379 );
xnor \U$31003 ( \31381 , \31380 , \21986 );
and \U$31004 ( \31382 , \31377 , \31381 );
and \U$31005 ( \31383 , \29040 , \21916 );
and \U$31006 ( \31384 , \28514 , \21914 );
nor \U$31007 ( \31385 , \31383 , \31384 );
xnor \U$31008 ( \31386 , \31385 , \21867 );
and \U$31009 ( \31387 , \31381 , \31386 );
and \U$31010 ( \31388 , \31377 , \31386 );
or \U$31011 ( \31389 , \31382 , \31387 , \31388 );
and \U$31012 ( \31390 , \25348 , \23431 );
and \U$31013 ( \31391 , \25226 , \23429 );
nor \U$31014 ( \31392 , \31390 , \31391 );
xnor \U$31015 ( \31393 , \31392 , \23279 );
and \U$31016 ( \31394 , \25609 , \23163 );
and \U$31017 ( \31395 , \25353 , \23161 );
nor \U$31018 ( \31396 , \31394 , \31395 );
xnor \U$31019 ( \31397 , \31396 , \23007 );
and \U$31020 ( \31398 , \31393 , \31397 );
and \U$31021 ( \31399 , \26108 , \22891 );
and \U$31022 ( \31400 , \25806 , \22889 );
nor \U$31023 ( \31401 , \31399 , \31400 );
xnor \U$31024 ( \31402 , \31401 , \22778 );
and \U$31025 ( \31403 , \31397 , \31402 );
and \U$31026 ( \31404 , \31393 , \31402 );
or \U$31027 ( \31405 , \31398 , \31403 , \31404 );
and \U$31028 ( \31406 , \31389 , \31405 );
and \U$31029 ( \31407 , \26585 , \22697 );
and \U$31030 ( \31408 , \26116 , \22695 );
nor \U$31031 ( \31409 , \31407 , \31408 );
xnor \U$31032 ( \31410 , \31409 , \22561 );
and \U$31033 ( \31411 , \26854 , \22497 );
and \U$31034 ( \31412 , \26590 , \22495 );
nor \U$31035 ( \31413 , \31411 , \31412 );
xnor \U$31036 ( \31414 , \31413 , \22419 );
and \U$31037 ( \31415 , \31410 , \31414 );
and \U$31038 ( \31416 , \27485 , \22333 );
and \U$31039 ( \31417 , \27113 , \22331 );
nor \U$31040 ( \31418 , \31416 , \31417 );
xnor \U$31041 ( \31419 , \31418 , \22239 );
and \U$31042 ( \31420 , \31414 , \31419 );
and \U$31043 ( \31421 , \31410 , \31419 );
or \U$31044 ( \31422 , \31415 , \31420 , \31421 );
and \U$31045 ( \31423 , \31405 , \31422 );
and \U$31046 ( \31424 , \31389 , \31422 );
or \U$31047 ( \31425 , \31406 , \31423 , \31424 );
and \U$31048 ( \31426 , \31373 , \31425 );
and \U$31049 ( \31427 , \22716 , \26517 );
and \U$31050 ( \31428 , \22611 , \26515 );
nor \U$31051 ( \31429 , \31427 , \31428 );
xnor \U$31052 ( \31430 , \31429 , \26329 );
and \U$31053 ( \31431 , \22837 , \26143 );
and \U$31054 ( \31432 , \22721 , \26141 );
nor \U$31055 ( \31433 , \31431 , \31432 );
xnor \U$31056 ( \31434 , \31433 , \25911 );
and \U$31057 ( \31435 , \31430 , \31434 );
and \U$31058 ( \31436 , \23128 , \25692 );
and \U$31059 ( \31437 , \22952 , \25690 );
nor \U$31060 ( \31438 , \31436 , \31437 );
xnor \U$31061 ( \31439 , \31438 , \25549 );
and \U$31062 ( \31440 , \31434 , \31439 );
and \U$31063 ( \31441 , \31430 , \31439 );
or \U$31064 ( \31442 , \31435 , \31440 , \31441 );
and \U$31065 ( \31443 , \24177 , \24255 );
and \U$31066 ( \31444 , \24003 , \24253 );
nor \U$31067 ( \31445 , \31443 , \31444 );
xnor \U$31068 ( \31446 , \31445 , \24106 );
and \U$31069 ( \31447 , \24482 , \23933 );
and \U$31070 ( \31448 , \24344 , \23931 );
nor \U$31071 ( \31449 , \31447 , \31448 );
xnor \U$31072 ( \31450 , \31449 , \23791 );
and \U$31073 ( \31451 , \31446 , \31450 );
and \U$31074 ( \31452 , \25018 , \23637 );
and \U$31075 ( \31453 , \24601 , \23635 );
nor \U$31076 ( \31454 , \31452 , \31453 );
xnor \U$31077 ( \31455 , \31454 , \23500 );
and \U$31078 ( \31456 , \31450 , \31455 );
and \U$31079 ( \31457 , \31446 , \31455 );
or \U$31080 ( \31458 , \31451 , \31456 , \31457 );
and \U$31081 ( \31459 , \31442 , \31458 );
and \U$31082 ( \31460 , \23379 , \25369 );
and \U$31083 ( \31461 , \23136 , \25367 );
nor \U$31084 ( \31462 , \31460 , \31461 );
xnor \U$31085 ( \31463 , \31462 , \25123 );
and \U$31086 ( \31464 , \23570 , \24974 );
and \U$31087 ( \31465 , \23384 , \24972 );
nor \U$31088 ( \31466 , \31464 , \31465 );
xnor \U$31089 ( \31467 , \31466 , \24787 );
and \U$31090 ( \31468 , \31463 , \31467 );
and \U$31091 ( \31469 , \23978 , \24661 );
and \U$31092 ( \31470 , \23714 , \24659 );
nor \U$31093 ( \31471 , \31469 , \31470 );
xnor \U$31094 ( \31472 , \31471 , \24456 );
and \U$31095 ( \31473 , \31467 , \31472 );
and \U$31096 ( \31474 , \31463 , \31472 );
or \U$31097 ( \31475 , \31468 , \31473 , \31474 );
and \U$31098 ( \31476 , \31458 , \31475 );
and \U$31099 ( \31477 , \31442 , \31475 );
or \U$31100 ( \31478 , \31459 , \31476 , \31477 );
and \U$31101 ( \31479 , \31425 , \31478 );
and \U$31102 ( \31480 , \31373 , \31478 );
or \U$31103 ( \31481 , \31426 , \31479 , \31480 );
and \U$31104 ( \31482 , \29710 , \21815 );
and \U$31105 ( \31483 , \29464 , \21813 );
nor \U$31106 ( \31484 , \31482 , \31483 );
xnor \U$31107 ( \31485 , \31484 , \21774 );
and \U$31108 ( \31486 , \30034 , \21745 );
and \U$31109 ( \31487 , \29715 , \21743 );
nor \U$31110 ( \31488 , \31486 , \31487 );
xnor \U$31111 ( \31489 , \31488 , \21715 );
and \U$31112 ( \31490 , \31485 , \31489 );
and \U$31113 ( \31491 , \30887 , \21697 );
and \U$31114 ( \31492 , \30318 , \21695 );
nor \U$31115 ( \31493 , \31491 , \31492 );
xnor \U$31116 ( \31494 , \31493 , \21678 );
and \U$31117 ( \31495 , \31489 , \31494 );
and \U$31118 ( \31496 , \31485 , \31494 );
or \U$31119 ( \31497 , \31490 , \31495 , \31496 );
buf \U$31120 ( \31498 , RIc22b1b0_189);
and \U$31121 ( \31499 , \31498 , \21660 );
and \U$31122 ( \31500 , \30895 , \21658 );
nor \U$31123 ( \31501 , \31499 , \31500 );
xnor \U$31124 ( \31502 , \31501 , \21665 );
buf \U$31125 ( \31503 , RIc22b228_190);
and \U$31126 ( \31504 , \31503 , \21654 );
or \U$31127 ( \31505 , \31502 , \31504 );
and \U$31128 ( \31506 , \31497 , \31505 );
and \U$31129 ( \31507 , \30895 , \21660 );
and \U$31130 ( \31508 , \30887 , \21658 );
nor \U$31131 ( \31509 , \31507 , \31508 );
xnor \U$31132 ( \31510 , \31509 , \21665 );
and \U$31133 ( \31511 , \31505 , \31510 );
and \U$31134 ( \31512 , \31497 , \31510 );
or \U$31135 ( \31513 , \31506 , \31511 , \31512 );
and \U$31136 ( \31514 , \31498 , \21654 );
xor \U$31137 ( \31515 , \31120 , \31124 );
xor \U$31138 ( \31516 , \31515 , \31129 );
and \U$31139 ( \31517 , \31514 , \31516 );
xor \U$31140 ( \31518 , \31196 , \31200 );
xor \U$31141 ( \31519 , \31518 , \31205 );
and \U$31142 ( \31520 , \31516 , \31519 );
and \U$31143 ( \31521 , \31514 , \31519 );
or \U$31144 ( \31522 , \31517 , \31520 , \31521 );
and \U$31145 ( \31523 , \31513 , \31522 );
xor \U$31146 ( \31524 , \31013 , \31017 );
xor \U$31147 ( \31525 , \31524 , \31022 );
xor \U$31148 ( \31526 , \31136 , \31140 );
xor \U$31149 ( \31527 , \31526 , \31145 );
and \U$31150 ( \31528 , \31525 , \31527 );
xor \U$31151 ( \31529 , \31153 , \31157 );
xor \U$31152 ( \31530 , \31529 , \31162 );
and \U$31153 ( \31531 , \31527 , \31530 );
and \U$31154 ( \31532 , \31525 , \31530 );
or \U$31155 ( \31533 , \31528 , \31531 , \31532 );
and \U$31156 ( \31534 , \31522 , \31533 );
and \U$31157 ( \31535 , \31513 , \31533 );
or \U$31158 ( \31536 , \31523 , \31534 , \31535 );
and \U$31159 ( \31537 , \31481 , \31536 );
xor \U$31160 ( \31538 , \31065 , \31069 );
xor \U$31161 ( \31539 , \31538 , \31074 );
xor \U$31162 ( \31540 , \31029 , \31033 );
xor \U$31163 ( \31541 , \31540 , \31038 );
and \U$31164 ( \31542 , \31539 , \31541 );
xor \U$31165 ( \31543 , \31046 , \31050 );
xor \U$31166 ( \31544 , \31543 , \31055 );
and \U$31167 ( \31545 , \31541 , \31544 );
and \U$31168 ( \31546 , \31539 , \31544 );
or \U$31169 ( \31547 , \31542 , \31545 , \31546 );
xor \U$31170 ( \31548 , \31081 , \31085 );
xor \U$31171 ( \31549 , \31548 , \31090 );
xor \U$31172 ( \31550 , \31100 , \31104 );
xor \U$31173 ( \31551 , \31550 , \31109 );
and \U$31174 ( \31552 , \31549 , \31551 );
and \U$31175 ( \31553 , \31547 , \31552 );
xor \U$31176 ( \31554 , \31221 , \31223 );
xor \U$31177 ( \31555 , \31554 , \31226 );
and \U$31178 ( \31556 , \31552 , \31555 );
and \U$31179 ( \31557 , \31547 , \31555 );
or \U$31180 ( \31558 , \31553 , \31556 , \31557 );
and \U$31181 ( \31559 , \31536 , \31558 );
and \U$31182 ( \31560 , \31481 , \31558 );
or \U$31183 ( \31561 , \31537 , \31559 , \31560 );
xor \U$31184 ( \31562 , \31025 , \31041 );
xor \U$31185 ( \31563 , \31562 , \31058 );
xor \U$31186 ( \31564 , \31077 , \31093 );
xor \U$31187 ( \31565 , \31564 , \31112 );
and \U$31188 ( \31566 , \31563 , \31565 );
xor \U$31189 ( \31567 , \31132 , \31148 );
xor \U$31190 ( \31568 , \31567 , \31165 );
and \U$31191 ( \31569 , \31565 , \31568 );
and \U$31192 ( \31570 , \31563 , \31568 );
or \U$31193 ( \31571 , \31566 , \31569 , \31570 );
xor \U$31194 ( \31572 , \31173 , \31175 );
xor \U$31195 ( \31573 , \31572 , \31178 );
xor \U$31196 ( \31574 , \31183 , \31185 );
xor \U$31197 ( \31575 , \31574 , \31188 );
and \U$31198 ( \31576 , \31573 , \31575 );
xor \U$31199 ( \31577 , \31208 , \31210 );
xor \U$31200 ( \31578 , \31577 , \31212 );
and \U$31201 ( \31579 , \31575 , \31578 );
and \U$31202 ( \31580 , \31573 , \31578 );
or \U$31203 ( \31581 , \31576 , \31579 , \31580 );
and \U$31204 ( \31582 , \31571 , \31581 );
xor \U$31205 ( \31583 , \31242 , \31244 );
xor \U$31206 ( \31584 , \31583 , \31247 );
and \U$31207 ( \31585 , \31581 , \31584 );
and \U$31208 ( \31586 , \31571 , \31584 );
or \U$31209 ( \31587 , \31582 , \31585 , \31586 );
and \U$31210 ( \31588 , \31561 , \31587 );
xor \U$31211 ( \31589 , \31181 , \31191 );
xor \U$31212 ( \31590 , \31589 , \31215 );
xor \U$31213 ( \31591 , \31252 , \31254 );
xor \U$31214 ( \31592 , \31591 , \31257 );
and \U$31215 ( \31593 , \31590 , \31592 );
xor \U$31216 ( \31594 , \31229 , \31231 );
xor \U$31217 ( \31595 , \31594 , \31234 );
and \U$31218 ( \31596 , \31592 , \31595 );
and \U$31219 ( \31597 , \31590 , \31595 );
or \U$31220 ( \31598 , \31593 , \31596 , \31597 );
and \U$31221 ( \31599 , \31587 , \31598 );
and \U$31222 ( \31600 , \31561 , \31598 );
or \U$31223 ( \31601 , \31588 , \31599 , \31600 );
xor \U$31224 ( \31602 , \30766 , \30821 );
xor \U$31225 ( \31603 , \31602 , \30874 );
xor \U$31226 ( \31604 , \30902 , \30912 );
xor \U$31227 ( \31605 , \31604 , \30923 );
and \U$31228 ( \31606 , \31603 , \31605 );
xor \U$31229 ( \31607 , \31269 , \31271 );
xor \U$31230 ( \31608 , \31607 , \31274 );
and \U$31231 ( \31609 , \31605 , \31608 );
and \U$31232 ( \31610 , \31603 , \31608 );
or \U$31233 ( \31611 , \31606 , \31609 , \31610 );
and \U$31234 ( \31612 , \31601 , \31611 );
xor \U$31235 ( \31613 , \31282 , \31284 );
xor \U$31236 ( \31614 , \31613 , \31287 );
and \U$31237 ( \31615 , \31611 , \31614 );
and \U$31238 ( \31616 , \31601 , \31614 );
or \U$31239 ( \31617 , \31612 , \31615 , \31616 );
xor \U$31240 ( \31618 , \31280 , \31290 );
xor \U$31241 ( \31619 , \31618 , \31293 );
and \U$31242 ( \31620 , \31617 , \31619 );
xor \U$31243 ( \31621 , \31298 , \31300 );
xor \U$31244 ( \31622 , \31621 , \31303 );
and \U$31245 ( \31623 , \31619 , \31622 );
and \U$31246 ( \31624 , \31617 , \31622 );
or \U$31247 ( \31625 , \31620 , \31623 , \31624 );
xor \U$31248 ( \31626 , \31296 , \31306 );
xor \U$31249 ( \31627 , \31626 , \31309 );
and \U$31250 ( \31628 , \31625 , \31627 );
xor \U$31251 ( \31629 , \30979 , \30989 );
xor \U$31252 ( \31630 , \31629 , \30992 );
and \U$31253 ( \31631 , \31627 , \31630 );
and \U$31254 ( \31632 , \31625 , \31630 );
or \U$31255 ( \31633 , \31628 , \31631 , \31632 );
and \U$31256 ( \31634 , \31318 , \31633 );
xor \U$31257 ( \31635 , \31318 , \31633 );
xor \U$31258 ( \31636 , \31625 , \31627 );
xor \U$31259 ( \31637 , \31636 , \31630 );
xor \U$31260 ( \31638 , \31446 , \31450 );
xor \U$31261 ( \31639 , \31638 , \31455 );
xor \U$31262 ( \31640 , \31463 , \31467 );
xor \U$31263 ( \31641 , \31640 , \31472 );
and \U$31264 ( \31642 , \31639 , \31641 );
xor \U$31265 ( \31643 , \31393 , \31397 );
xor \U$31266 ( \31644 , \31643 , \31402 );
and \U$31267 ( \31645 , \31641 , \31644 );
and \U$31268 ( \31646 , \31639 , \31644 );
or \U$31269 ( \31647 , \31642 , \31645 , \31646 );
xor \U$31270 ( \31648 , \31377 , \31381 );
xor \U$31271 ( \31649 , \31648 , \31386 );
xor \U$31272 ( \31650 , \31485 , \31489 );
xor \U$31273 ( \31651 , \31650 , \31494 );
and \U$31274 ( \31652 , \31649 , \31651 );
xor \U$31275 ( \31653 , \31410 , \31414 );
xor \U$31276 ( \31654 , \31653 , \31419 );
and \U$31277 ( \31655 , \31651 , \31654 );
and \U$31278 ( \31656 , \31649 , \31654 );
or \U$31279 ( \31657 , \31652 , \31655 , \31656 );
and \U$31280 ( \31658 , \31647 , \31657 );
and \U$31281 ( \31659 , \29464 , \21916 );
and \U$31282 ( \31660 , \29040 , \21914 );
nor \U$31283 ( \31661 , \31659 , \31660 );
xnor \U$31284 ( \31662 , \31661 , \21867 );
and \U$31285 ( \31663 , \29715 , \21815 );
and \U$31286 ( \31664 , \29710 , \21813 );
nor \U$31287 ( \31665 , \31663 , \31664 );
xnor \U$31288 ( \31666 , \31665 , \21774 );
and \U$31289 ( \31667 , \31662 , \31666 );
and \U$31290 ( \31668 , \30318 , \21745 );
and \U$31291 ( \31669 , \30034 , \21743 );
nor \U$31292 ( \31670 , \31668 , \31669 );
xnor \U$31293 ( \31671 , \31670 , \21715 );
and \U$31294 ( \31672 , \31666 , \31671 );
and \U$31295 ( \31673 , \31662 , \31671 );
or \U$31296 ( \31674 , \31667 , \31672 , \31673 );
and \U$31297 ( \31675 , \30895 , \21697 );
and \U$31298 ( \31676 , \30887 , \21695 );
nor \U$31299 ( \31677 , \31675 , \31676 );
xnor \U$31300 ( \31678 , \31677 , \21678 );
and \U$31301 ( \31679 , \31503 , \21660 );
and \U$31302 ( \31680 , \31498 , \21658 );
nor \U$31303 ( \31681 , \31679 , \31680 );
xnor \U$31304 ( \31682 , \31681 , \21665 );
and \U$31305 ( \31683 , \31678 , \31682 );
buf \U$31306 ( \31684 , RIc22b2a0_191);
and \U$31307 ( \31685 , \31684 , \21654 );
and \U$31308 ( \31686 , \31682 , \31685 );
and \U$31309 ( \31687 , \31678 , \31685 );
or \U$31310 ( \31688 , \31683 , \31686 , \31687 );
and \U$31311 ( \31689 , \31674 , \31688 );
xnor \U$31312 ( \31690 , \31502 , \31504 );
and \U$31313 ( \31691 , \31688 , \31690 );
and \U$31314 ( \31692 , \31674 , \31690 );
or \U$31315 ( \31693 , \31689 , \31691 , \31692 );
and \U$31316 ( \31694 , \31657 , \31693 );
and \U$31317 ( \31695 , \31647 , \31693 );
or \U$31318 ( \31696 , \31658 , \31694 , \31695 );
not \U$31319 ( \31697 , \31096 );
and \U$31320 ( \31698 , \21667 , \31338 );
and \U$31321 ( \31699 , \21653 , \31336 );
nor \U$31322 ( \31700 , \31698 , \31699 );
xnor \U$31323 ( \31701 , \31700 , \31099 );
and \U$31324 ( \31702 , \31697 , \31701 );
and \U$31325 ( \31703 , \21706 , \30770 );
and \U$31326 ( \31704 , \21685 , \30768 );
nor \U$31327 ( \31705 , \31703 , \31704 );
xnor \U$31328 ( \31706 , \31705 , \30460 );
and \U$31329 ( \31707 , \31701 , \31706 );
and \U$31330 ( \31708 , \31697 , \31706 );
or \U$31331 ( \31709 , \31702 , \31707 , \31708 );
and \U$31332 ( \31710 , \21762 , \30233 );
and \U$31333 ( \31711 , \21754 , \30231 );
nor \U$31334 ( \31712 , \31710 , \31711 );
xnor \U$31335 ( \31713 , \31712 , \29862 );
and \U$31336 ( \31714 , \21836 , \29671 );
and \U$31337 ( \31715 , \21831 , \29669 );
nor \U$31338 ( \31716 , \31714 , \31715 );
xnor \U$31339 ( \31717 , \31716 , \29353 );
and \U$31340 ( \31718 , \31713 , \31717 );
and \U$31341 ( \31719 , \21941 , \29104 );
and \U$31342 ( \31720 , \21890 , \29102 );
nor \U$31343 ( \31721 , \31719 , \31720 );
xnor \U$31344 ( \31722 , \31721 , \28855 );
and \U$31345 ( \31723 , \31717 , \31722 );
and \U$31346 ( \31724 , \31713 , \31722 );
or \U$31347 ( \31725 , \31718 , \31723 , \31724 );
and \U$31348 ( \31726 , \31709 , \31725 );
and \U$31349 ( \31727 , \22046 , \28575 );
and \U$31350 ( \31728 , \22018 , \28573 );
nor \U$31351 ( \31729 , \31727 , \31728 );
xnor \U$31352 ( \31730 , \31729 , \28315 );
and \U$31353 ( \31731 , \22200 , \28081 );
and \U$31354 ( \31732 , \22126 , \28079 );
nor \U$31355 ( \31733 , \31731 , \31732 );
xnor \U$31356 ( \31734 , \31733 , \27766 );
and \U$31357 ( \31735 , \31730 , \31734 );
and \U$31358 ( \31736 , \22325 , \27572 );
and \U$31359 ( \31737 , \22262 , \27570 );
nor \U$31360 ( \31738 , \31736 , \31737 );
xnor \U$31361 ( \31739 , \31738 , \27232 );
and \U$31362 ( \31740 , \31734 , \31739 );
and \U$31363 ( \31741 , \31730 , \31739 );
or \U$31364 ( \31742 , \31735 , \31740 , \31741 );
and \U$31365 ( \31743 , \31725 , \31742 );
and \U$31366 ( \31744 , \31709 , \31742 );
or \U$31367 ( \31745 , \31726 , \31743 , \31744 );
and \U$31368 ( \31746 , \26116 , \22891 );
and \U$31369 ( \31747 , \26108 , \22889 );
nor \U$31370 ( \31748 , \31746 , \31747 );
xnor \U$31371 ( \31749 , \31748 , \22778 );
and \U$31372 ( \31750 , \26590 , \22697 );
and \U$31373 ( \31751 , \26585 , \22695 );
nor \U$31374 ( \31752 , \31750 , \31751 );
xnor \U$31375 ( \31753 , \31752 , \22561 );
and \U$31376 ( \31754 , \31749 , \31753 );
and \U$31377 ( \31755 , \27113 , \22497 );
and \U$31378 ( \31756 , \26854 , \22495 );
nor \U$31379 ( \31757 , \31755 , \31756 );
xnor \U$31380 ( \31758 , \31757 , \22419 );
and \U$31381 ( \31759 , \31753 , \31758 );
and \U$31382 ( \31760 , \31749 , \31758 );
or \U$31383 ( \31761 , \31754 , \31759 , \31760 );
and \U$31384 ( \31762 , \25226 , \23637 );
and \U$31385 ( \31763 , \25018 , \23635 );
nor \U$31386 ( \31764 , \31762 , \31763 );
xnor \U$31387 ( \31765 , \31764 , \23500 );
and \U$31388 ( \31766 , \25353 , \23431 );
and \U$31389 ( \31767 , \25348 , \23429 );
nor \U$31390 ( \31768 , \31766 , \31767 );
xnor \U$31391 ( \31769 , \31768 , \23279 );
and \U$31392 ( \31770 , \31765 , \31769 );
and \U$31393 ( \31771 , \25806 , \23163 );
and \U$31394 ( \31772 , \25609 , \23161 );
nor \U$31395 ( \31773 , \31771 , \31772 );
xnor \U$31396 ( \31774 , \31773 , \23007 );
and \U$31397 ( \31775 , \31769 , \31774 );
and \U$31398 ( \31776 , \31765 , \31774 );
or \U$31399 ( \31777 , \31770 , \31775 , \31776 );
and \U$31400 ( \31778 , \31761 , \31777 );
and \U$31401 ( \31779 , \27494 , \22333 );
and \U$31402 ( \31780 , \27485 , \22331 );
nor \U$31403 ( \31781 , \31779 , \31780 );
xnor \U$31404 ( \31782 , \31781 , \22239 );
and \U$31405 ( \31783 , \28039 , \22163 );
and \U$31406 ( \31784 , \27837 , \22161 );
nor \U$31407 ( \31785 , \31783 , \31784 );
xnor \U$31408 ( \31786 , \31785 , \22091 );
and \U$31409 ( \31787 , \31782 , \31786 );
and \U$31410 ( \31788 , \28514 , \22029 );
and \U$31411 ( \31789 , \28342 , \22027 );
nor \U$31412 ( \31790 , \31788 , \31789 );
xnor \U$31413 ( \31791 , \31790 , \21986 );
and \U$31414 ( \31792 , \31786 , \31791 );
and \U$31415 ( \31793 , \31782 , \31791 );
or \U$31416 ( \31794 , \31787 , \31792 , \31793 );
and \U$31417 ( \31795 , \31777 , \31794 );
and \U$31418 ( \31796 , \31761 , \31794 );
or \U$31419 ( \31797 , \31778 , \31795 , \31796 );
and \U$31420 ( \31798 , \31745 , \31797 );
and \U$31421 ( \31799 , \23136 , \25692 );
and \U$31422 ( \31800 , \23128 , \25690 );
nor \U$31423 ( \31801 , \31799 , \31800 );
xnor \U$31424 ( \31802 , \31801 , \25549 );
and \U$31425 ( \31803 , \23384 , \25369 );
and \U$31426 ( \31804 , \23379 , \25367 );
nor \U$31427 ( \31805 , \31803 , \31804 );
xnor \U$31428 ( \31806 , \31805 , \25123 );
and \U$31429 ( \31807 , \31802 , \31806 );
and \U$31430 ( \31808 , \23714 , \24974 );
and \U$31431 ( \31809 , \23570 , \24972 );
nor \U$31432 ( \31810 , \31808 , \31809 );
xnor \U$31433 ( \31811 , \31810 , \24787 );
and \U$31434 ( \31812 , \31806 , \31811 );
and \U$31435 ( \31813 , \31802 , \31811 );
or \U$31436 ( \31814 , \31807 , \31812 , \31813 );
and \U$31437 ( \31815 , \24003 , \24661 );
and \U$31438 ( \31816 , \23978 , \24659 );
nor \U$31439 ( \31817 , \31815 , \31816 );
xnor \U$31440 ( \31818 , \31817 , \24456 );
and \U$31441 ( \31819 , \24344 , \24255 );
and \U$31442 ( \31820 , \24177 , \24253 );
nor \U$31443 ( \31821 , \31819 , \31820 );
xnor \U$31444 ( \31822 , \31821 , \24106 );
and \U$31445 ( \31823 , \31818 , \31822 );
and \U$31446 ( \31824 , \24601 , \23933 );
and \U$31447 ( \31825 , \24482 , \23931 );
nor \U$31448 ( \31826 , \31824 , \31825 );
xnor \U$31449 ( \31827 , \31826 , \23791 );
and \U$31450 ( \31828 , \31822 , \31827 );
and \U$31451 ( \31829 , \31818 , \31827 );
or \U$31452 ( \31830 , \31823 , \31828 , \31829 );
and \U$31453 ( \31831 , \31814 , \31830 );
and \U$31454 ( \31832 , \22611 , \26983 );
and \U$31455 ( \31833 , \22523 , \26981 );
nor \U$31456 ( \31834 , \31832 , \31833 );
xnor \U$31457 ( \31835 , \31834 , \26742 );
and \U$31458 ( \31836 , \22721 , \26517 );
and \U$31459 ( \31837 , \22716 , \26515 );
nor \U$31460 ( \31838 , \31836 , \31837 );
xnor \U$31461 ( \31839 , \31838 , \26329 );
and \U$31462 ( \31840 , \31835 , \31839 );
and \U$31463 ( \31841 , \22952 , \26143 );
and \U$31464 ( \31842 , \22837 , \26141 );
nor \U$31465 ( \31843 , \31841 , \31842 );
xnor \U$31466 ( \31844 , \31843 , \25911 );
and \U$31467 ( \31845 , \31839 , \31844 );
and \U$31468 ( \31846 , \31835 , \31844 );
or \U$31469 ( \31847 , \31840 , \31845 , \31846 );
and \U$31470 ( \31848 , \31830 , \31847 );
and \U$31471 ( \31849 , \31814 , \31847 );
or \U$31472 ( \31850 , \31831 , \31848 , \31849 );
and \U$31473 ( \31851 , \31797 , \31850 );
and \U$31474 ( \31852 , \31745 , \31850 );
or \U$31475 ( \31853 , \31798 , \31851 , \31852 );
and \U$31476 ( \31854 , \31696 , \31853 );
xor \U$31477 ( \31855 , \31430 , \31434 );
xor \U$31478 ( \31856 , \31855 , \31439 );
xor \U$31479 ( \31857 , \31322 , \31326 );
xor \U$31480 ( \31858 , \31857 , \31331 );
and \U$31481 ( \31859 , \31856 , \31858 );
xor \U$31482 ( \31860 , \31358 , \31362 );
xor \U$31483 ( \31861 , \31860 , \31367 );
and \U$31484 ( \31862 , \31858 , \31861 );
and \U$31485 ( \31863 , \31856 , \31861 );
or \U$31486 ( \31864 , \31859 , \31862 , \31863 );
xor \U$31487 ( \31865 , \31539 , \31541 );
xor \U$31488 ( \31866 , \31865 , \31544 );
and \U$31489 ( \31867 , \31864 , \31866 );
xor \U$31490 ( \31868 , \31549 , \31551 );
and \U$31491 ( \31869 , \31866 , \31868 );
and \U$31492 ( \31870 , \31864 , \31868 );
or \U$31493 ( \31871 , \31867 , \31869 , \31870 );
and \U$31494 ( \31872 , \31853 , \31871 );
and \U$31495 ( \31873 , \31696 , \31871 );
or \U$31496 ( \31874 , \31854 , \31872 , \31873 );
xor \U$31497 ( \31875 , \31334 , \31353 );
xor \U$31498 ( \31876 , \31875 , \31370 );
xor \U$31499 ( \31877 , \31389 , \31405 );
xor \U$31500 ( \31878 , \31877 , \31422 );
and \U$31501 ( \31879 , \31876 , \31878 );
xor \U$31502 ( \31880 , \31442 , \31458 );
xor \U$31503 ( \31881 , \31880 , \31475 );
and \U$31504 ( \31882 , \31878 , \31881 );
and \U$31505 ( \31883 , \31876 , \31881 );
or \U$31506 ( \31884 , \31879 , \31882 , \31883 );
xor \U$31507 ( \31885 , \31497 , \31505 );
xor \U$31508 ( \31886 , \31885 , \31510 );
xor \U$31509 ( \31887 , \31514 , \31516 );
xor \U$31510 ( \31888 , \31887 , \31519 );
and \U$31511 ( \31889 , \31886 , \31888 );
xor \U$31512 ( \31890 , \31525 , \31527 );
xor \U$31513 ( \31891 , \31890 , \31530 );
and \U$31514 ( \31892 , \31888 , \31891 );
and \U$31515 ( \31893 , \31886 , \31891 );
or \U$31516 ( \31894 , \31889 , \31892 , \31893 );
and \U$31517 ( \31895 , \31884 , \31894 );
xor \U$31518 ( \31896 , \31563 , \31565 );
xor \U$31519 ( \31897 , \31896 , \31568 );
and \U$31520 ( \31898 , \31894 , \31897 );
and \U$31521 ( \31899 , \31884 , \31897 );
or \U$31522 ( \31900 , \31895 , \31898 , \31899 );
and \U$31523 ( \31901 , \31874 , \31900 );
xor \U$31524 ( \31902 , \31513 , \31522 );
xor \U$31525 ( \31903 , \31902 , \31533 );
xor \U$31526 ( \31904 , \31547 , \31552 );
xor \U$31527 ( \31905 , \31904 , \31555 );
and \U$31528 ( \31906 , \31903 , \31905 );
xor \U$31529 ( \31907 , \31573 , \31575 );
xor \U$31530 ( \31908 , \31907 , \31578 );
and \U$31531 ( \31909 , \31905 , \31908 );
and \U$31532 ( \31910 , \31903 , \31908 );
or \U$31533 ( \31911 , \31906 , \31909 , \31910 );
and \U$31534 ( \31912 , \31900 , \31911 );
and \U$31535 ( \31913 , \31874 , \31911 );
or \U$31536 ( \31914 , \31901 , \31912 , \31913 );
xor \U$31537 ( \31915 , \31061 , \31115 );
xor \U$31538 ( \31916 , \31915 , \31168 );
xor \U$31539 ( \31917 , \31571 , \31581 );
xor \U$31540 ( \31918 , \31917 , \31584 );
and \U$31541 ( \31919 , \31916 , \31918 );
xor \U$31542 ( \31920 , \31590 , \31592 );
xor \U$31543 ( \31921 , \31920 , \31595 );
and \U$31544 ( \31922 , \31918 , \31921 );
and \U$31545 ( \31923 , \31916 , \31921 );
or \U$31546 ( \31924 , \31919 , \31922 , \31923 );
and \U$31547 ( \31925 , \31914 , \31924 );
xor \U$31548 ( \31926 , \31250 , \31260 );
xor \U$31549 ( \31927 , \31926 , \31263 );
and \U$31550 ( \31928 , \31924 , \31927 );
and \U$31551 ( \31929 , \31914 , \31927 );
or \U$31552 ( \31930 , \31925 , \31928 , \31929 );
xor \U$31553 ( \31931 , \31171 , \31218 );
xor \U$31554 ( \31932 , \31931 , \31237 );
xor \U$31555 ( \31933 , \31561 , \31587 );
xor \U$31556 ( \31934 , \31933 , \31598 );
and \U$31557 ( \31935 , \31932 , \31934 );
xor \U$31558 ( \31936 , \31603 , \31605 );
xor \U$31559 ( \31937 , \31936 , \31608 );
and \U$31560 ( \31938 , \31934 , \31937 );
and \U$31561 ( \31939 , \31932 , \31937 );
or \U$31562 ( \31940 , \31935 , \31938 , \31939 );
and \U$31563 ( \31941 , \31930 , \31940 );
xor \U$31564 ( \31942 , \31240 , \31266 );
xor \U$31565 ( \31943 , \31942 , \31277 );
and \U$31566 ( \31944 , \31940 , \31943 );
and \U$31567 ( \31945 , \31930 , \31943 );
or \U$31568 ( \31946 , \31941 , \31944 , \31945 );
xor \U$31569 ( \31947 , \31617 , \31619 );
xor \U$31570 ( \31948 , \31947 , \31622 );
and \U$31571 ( \31949 , \31946 , \31948 );
and \U$31572 ( \31950 , \31637 , \31949 );
xor \U$31573 ( \31951 , \31637 , \31949 );
xor \U$31574 ( \31952 , \31946 , \31948 );
xor \U$31575 ( \31953 , \31749 , \31753 );
xor \U$31576 ( \31954 , \31953 , \31758 );
xor \U$31577 ( \31955 , \31765 , \31769 );
xor \U$31578 ( \31956 , \31955 , \31774 );
and \U$31579 ( \31957 , \31954 , \31956 );
xor \U$31580 ( \31958 , \31818 , \31822 );
xor \U$31581 ( \31959 , \31958 , \31827 );
and \U$31582 ( \31960 , \31956 , \31959 );
and \U$31583 ( \31961 , \31954 , \31959 );
or \U$31584 ( \31962 , \31957 , \31960 , \31961 );
xor \U$31585 ( \31963 , \31662 , \31666 );
xor \U$31586 ( \31964 , \31963 , \31671 );
xor \U$31587 ( \31965 , \31678 , \31682 );
xor \U$31588 ( \31966 , \31965 , \31685 );
and \U$31589 ( \31967 , \31964 , \31966 );
xor \U$31590 ( \31968 , \31782 , \31786 );
xor \U$31591 ( \31969 , \31968 , \31791 );
and \U$31592 ( \31970 , \31966 , \31969 );
and \U$31593 ( \31971 , \31964 , \31969 );
or \U$31594 ( \31972 , \31967 , \31970 , \31971 );
and \U$31595 ( \31973 , \31962 , \31972 );
and \U$31596 ( \31974 , \29040 , \22029 );
and \U$31597 ( \31975 , \28514 , \22027 );
nor \U$31598 ( \31976 , \31974 , \31975 );
xnor \U$31599 ( \31977 , \31976 , \21986 );
and \U$31600 ( \31978 , \29710 , \21916 );
and \U$31601 ( \31979 , \29464 , \21914 );
nor \U$31602 ( \31980 , \31978 , \31979 );
xnor \U$31603 ( \31981 , \31980 , \21867 );
and \U$31604 ( \31982 , \31977 , \31981 );
and \U$31605 ( \31983 , \30034 , \21815 );
and \U$31606 ( \31984 , \29715 , \21813 );
nor \U$31607 ( \31985 , \31983 , \31984 );
xnor \U$31608 ( \31986 , \31985 , \21774 );
and \U$31609 ( \31987 , \31981 , \31986 );
and \U$31610 ( \31988 , \31977 , \31986 );
or \U$31611 ( \31989 , \31982 , \31987 , \31988 );
and \U$31612 ( \31990 , \30887 , \21745 );
and \U$31613 ( \31991 , \30318 , \21743 );
nor \U$31614 ( \31992 , \31990 , \31991 );
xnor \U$31615 ( \31993 , \31992 , \21715 );
and \U$31616 ( \31994 , \31498 , \21697 );
and \U$31617 ( \31995 , \30895 , \21695 );
nor \U$31618 ( \31996 , \31994 , \31995 );
xnor \U$31619 ( \31997 , \31996 , \21678 );
and \U$31620 ( \31998 , \31993 , \31997 );
and \U$31621 ( \31999 , \31684 , \21660 );
and \U$31622 ( \32000 , \31503 , \21658 );
nor \U$31623 ( \32001 , \31999 , \32000 );
xnor \U$31624 ( \32002 , \32001 , \21665 );
and \U$31625 ( \32003 , \31997 , \32002 );
and \U$31626 ( \32004 , \31993 , \32002 );
or \U$31627 ( \32005 , \31998 , \32003 , \32004 );
or \U$31628 ( \32006 , \31989 , \32005 );
and \U$31629 ( \32007 , \31972 , \32006 );
and \U$31630 ( \32008 , \31962 , \32006 );
or \U$31631 ( \32009 , \31973 , \32007 , \32008 );
and \U$31632 ( \32010 , \26108 , \23163 );
and \U$31633 ( \32011 , \25806 , \23161 );
nor \U$31634 ( \32012 , \32010 , \32011 );
xnor \U$31635 ( \32013 , \32012 , \23007 );
and \U$31636 ( \32014 , \26585 , \22891 );
and \U$31637 ( \32015 , \26116 , \22889 );
nor \U$31638 ( \32016 , \32014 , \32015 );
xnor \U$31639 ( \32017 , \32016 , \22778 );
and \U$31640 ( \32018 , \32013 , \32017 );
and \U$31641 ( \32019 , \26854 , \22697 );
and \U$31642 ( \32020 , \26590 , \22695 );
nor \U$31643 ( \32021 , \32019 , \32020 );
xnor \U$31644 ( \32022 , \32021 , \22561 );
and \U$31645 ( \32023 , \32017 , \32022 );
and \U$31646 ( \32024 , \32013 , \32022 );
or \U$31647 ( \32025 , \32018 , \32023 , \32024 );
and \U$31648 ( \32026 , \27485 , \22497 );
and \U$31649 ( \32027 , \27113 , \22495 );
nor \U$31650 ( \32028 , \32026 , \32027 );
xnor \U$31651 ( \32029 , \32028 , \22419 );
and \U$31652 ( \32030 , \27837 , \22333 );
and \U$31653 ( \32031 , \27494 , \22331 );
nor \U$31654 ( \32032 , \32030 , \32031 );
xnor \U$31655 ( \32033 , \32032 , \22239 );
and \U$31656 ( \32034 , \32029 , \32033 );
and \U$31657 ( \32035 , \28342 , \22163 );
and \U$31658 ( \32036 , \28039 , \22161 );
nor \U$31659 ( \32037 , \32035 , \32036 );
xnor \U$31660 ( \32038 , \32037 , \22091 );
and \U$31661 ( \32039 , \32033 , \32038 );
and \U$31662 ( \32040 , \32029 , \32038 );
or \U$31663 ( \32041 , \32034 , \32039 , \32040 );
and \U$31664 ( \32042 , \32025 , \32041 );
and \U$31665 ( \32043 , \25018 , \23933 );
and \U$31666 ( \32044 , \24601 , \23931 );
nor \U$31667 ( \32045 , \32043 , \32044 );
xnor \U$31668 ( \32046 , \32045 , \23791 );
and \U$31669 ( \32047 , \25348 , \23637 );
and \U$31670 ( \32048 , \25226 , \23635 );
nor \U$31671 ( \32049 , \32047 , \32048 );
xnor \U$31672 ( \32050 , \32049 , \23500 );
and \U$31673 ( \32051 , \32046 , \32050 );
and \U$31674 ( \32052 , \25609 , \23431 );
and \U$31675 ( \32053 , \25353 , \23429 );
nor \U$31676 ( \32054 , \32052 , \32053 );
xnor \U$31677 ( \32055 , \32054 , \23279 );
and \U$31678 ( \32056 , \32050 , \32055 );
and \U$31679 ( \32057 , \32046 , \32055 );
or \U$31680 ( \32058 , \32051 , \32056 , \32057 );
and \U$31681 ( \32059 , \32041 , \32058 );
and \U$31682 ( \32060 , \32025 , \32058 );
or \U$31683 ( \32061 , \32042 , \32059 , \32060 );
and \U$31684 ( \32062 , \23128 , \26143 );
and \U$31685 ( \32063 , \22952 , \26141 );
nor \U$31686 ( \32064 , \32062 , \32063 );
xnor \U$31687 ( \32065 , \32064 , \25911 );
and \U$31688 ( \32066 , \23379 , \25692 );
and \U$31689 ( \32067 , \23136 , \25690 );
nor \U$31690 ( \32068 , \32066 , \32067 );
xnor \U$31691 ( \32069 , \32068 , \25549 );
and \U$31692 ( \32070 , \32065 , \32069 );
and \U$31693 ( \32071 , \23570 , \25369 );
and \U$31694 ( \32072 , \23384 , \25367 );
nor \U$31695 ( \32073 , \32071 , \32072 );
xnor \U$31696 ( \32074 , \32073 , \25123 );
and \U$31697 ( \32075 , \32069 , \32074 );
and \U$31698 ( \32076 , \32065 , \32074 );
or \U$31699 ( \32077 , \32070 , \32075 , \32076 );
and \U$31700 ( \32078 , \23978 , \24974 );
and \U$31701 ( \32079 , \23714 , \24972 );
nor \U$31702 ( \32080 , \32078 , \32079 );
xnor \U$31703 ( \32081 , \32080 , \24787 );
and \U$31704 ( \32082 , \24177 , \24661 );
and \U$31705 ( \32083 , \24003 , \24659 );
nor \U$31706 ( \32084 , \32082 , \32083 );
xnor \U$31707 ( \32085 , \32084 , \24456 );
and \U$31708 ( \32086 , \32081 , \32085 );
and \U$31709 ( \32087 , \24482 , \24255 );
and \U$31710 ( \32088 , \24344 , \24253 );
nor \U$31711 ( \32089 , \32087 , \32088 );
xnor \U$31712 ( \32090 , \32089 , \24106 );
and \U$31713 ( \32091 , \32085 , \32090 );
and \U$31714 ( \32092 , \32081 , \32090 );
or \U$31715 ( \32093 , \32086 , \32091 , \32092 );
and \U$31716 ( \32094 , \32077 , \32093 );
and \U$31717 ( \32095 , \22523 , \27572 );
and \U$31718 ( \32096 , \22325 , \27570 );
nor \U$31719 ( \32097 , \32095 , \32096 );
xnor \U$31720 ( \32098 , \32097 , \27232 );
and \U$31721 ( \32099 , \22716 , \26983 );
and \U$31722 ( \32100 , \22611 , \26981 );
nor \U$31723 ( \32101 , \32099 , \32100 );
xnor \U$31724 ( \32102 , \32101 , \26742 );
and \U$31725 ( \32103 , \32098 , \32102 );
and \U$31726 ( \32104 , \22837 , \26517 );
and \U$31727 ( \32105 , \22721 , \26515 );
nor \U$31728 ( \32106 , \32104 , \32105 );
xnor \U$31729 ( \32107 , \32106 , \26329 );
and \U$31730 ( \32108 , \32102 , \32107 );
and \U$31731 ( \32109 , \32098 , \32107 );
or \U$31732 ( \32110 , \32103 , \32108 , \32109 );
and \U$31733 ( \32111 , \32093 , \32110 );
and \U$31734 ( \32112 , \32077 , \32110 );
or \U$31735 ( \32113 , \32094 , \32111 , \32112 );
and \U$31736 ( \32114 , \32061 , \32113 );
and \U$31737 ( \32115 , \21754 , \30770 );
and \U$31738 ( \32116 , \21706 , \30768 );
nor \U$31739 ( \32117 , \32115 , \32116 );
xnor \U$31740 ( \32118 , \32117 , \30460 );
and \U$31741 ( \32119 , \21831 , \30233 );
and \U$31742 ( \32120 , \21762 , \30231 );
nor \U$31743 ( \32121 , \32119 , \32120 );
xnor \U$31744 ( \32122 , \32121 , \29862 );
and \U$31745 ( \32123 , \32118 , \32122 );
and \U$31746 ( \32124 , \21890 , \29671 );
and \U$31747 ( \32125 , \21836 , \29669 );
nor \U$31748 ( \32126 , \32124 , \32125 );
xnor \U$31749 ( \32127 , \32126 , \29353 );
and \U$31750 ( \32128 , \32122 , \32127 );
and \U$31751 ( \32129 , \32118 , \32127 );
or \U$31752 ( \32130 , \32123 , \32128 , \32129 );
and \U$31753 ( \32131 , \22018 , \29104 );
and \U$31754 ( \32132 , \21941 , \29102 );
nor \U$31755 ( \32133 , \32131 , \32132 );
xnor \U$31756 ( \32134 , \32133 , \28855 );
and \U$31757 ( \32135 , \22126 , \28575 );
and \U$31758 ( \32136 , \22046 , \28573 );
nor \U$31759 ( \32137 , \32135 , \32136 );
xnor \U$31760 ( \32138 , \32137 , \28315 );
and \U$31761 ( \32139 , \32134 , \32138 );
and \U$31762 ( \32140 , \22262 , \28081 );
and \U$31763 ( \32141 , \22200 , \28079 );
nor \U$31764 ( \32142 , \32140 , \32141 );
xnor \U$31765 ( \32143 , \32142 , \27766 );
and \U$31766 ( \32144 , \32138 , \32143 );
and \U$31767 ( \32145 , \32134 , \32143 );
or \U$31768 ( \32146 , \32139 , \32144 , \32145 );
and \U$31769 ( \32147 , \32130 , \32146 );
buf \U$31770 ( \32148 , RIc225828_64);
xor \U$31771 ( \32149 , \31096 , \32148 );
not \U$31772 ( \32150 , \32148 );
and \U$31773 ( \32151 , \32149 , \32150 );
and \U$31774 ( \32152 , \21653 , \32151 );
not \U$31775 ( \32153 , \32152 );
xnor \U$31776 ( \32154 , \32153 , \31096 );
and \U$31777 ( \32155 , \21685 , \31338 );
and \U$31778 ( \32156 , \21667 , \31336 );
nor \U$31779 ( \32157 , \32155 , \32156 );
xnor \U$31780 ( \32158 , \32157 , \31099 );
and \U$31781 ( \32159 , \32154 , \32158 );
and \U$31782 ( \32160 , \32146 , \32159 );
and \U$31783 ( \32161 , \32130 , \32159 );
or \U$31784 ( \32162 , \32147 , \32160 , \32161 );
and \U$31785 ( \32163 , \32113 , \32162 );
and \U$31786 ( \32164 , \32061 , \32162 );
or \U$31787 ( \32165 , \32114 , \32163 , \32164 );
and \U$31788 ( \32166 , \32009 , \32165 );
xor \U$31789 ( \32167 , \31802 , \31806 );
xor \U$31790 ( \32168 , \32167 , \31811 );
xor \U$31791 ( \32169 , \31730 , \31734 );
xor \U$31792 ( \32170 , \32169 , \31739 );
and \U$31793 ( \32171 , \32168 , \32170 );
xor \U$31794 ( \32172 , \31835 , \31839 );
xor \U$31795 ( \32173 , \32172 , \31844 );
and \U$31796 ( \32174 , \32170 , \32173 );
and \U$31797 ( \32175 , \32168 , \32173 );
or \U$31798 ( \32176 , \32171 , \32174 , \32175 );
xor \U$31799 ( \32177 , \31697 , \31701 );
xor \U$31800 ( \32178 , \32177 , \31706 );
xor \U$31801 ( \32179 , \31713 , \31717 );
xor \U$31802 ( \32180 , \32179 , \31722 );
and \U$31803 ( \32181 , \32178 , \32180 );
and \U$31804 ( \32182 , \32176 , \32181 );
xor \U$31805 ( \32183 , \31341 , \31345 );
xor \U$31806 ( \32184 , \32183 , \31350 );
and \U$31807 ( \32185 , \32181 , \32184 );
and \U$31808 ( \32186 , \32176 , \32184 );
or \U$31809 ( \32187 , \32182 , \32185 , \32186 );
and \U$31810 ( \32188 , \32165 , \32187 );
and \U$31811 ( \32189 , \32009 , \32187 );
or \U$31812 ( \32190 , \32166 , \32188 , \32189 );
xor \U$31813 ( \32191 , \31856 , \31858 );
xor \U$31814 ( \32192 , \32191 , \31861 );
xor \U$31815 ( \32193 , \31639 , \31641 );
xor \U$31816 ( \32194 , \32193 , \31644 );
and \U$31817 ( \32195 , \32192 , \32194 );
xor \U$31818 ( \32196 , \31649 , \31651 );
xor \U$31819 ( \32197 , \32196 , \31654 );
and \U$31820 ( \32198 , \32194 , \32197 );
and \U$31821 ( \32199 , \32192 , \32197 );
or \U$31822 ( \32200 , \32195 , \32198 , \32199 );
xor \U$31823 ( \32201 , \31761 , \31777 );
xor \U$31824 ( \32202 , \32201 , \31794 );
xor \U$31825 ( \32203 , \31814 , \31830 );
xor \U$31826 ( \32204 , \32203 , \31847 );
and \U$31827 ( \32205 , \32202 , \32204 );
xor \U$31828 ( \32206 , \31674 , \31688 );
xor \U$31829 ( \32207 , \32206 , \31690 );
and \U$31830 ( \32208 , \32204 , \32207 );
and \U$31831 ( \32209 , \32202 , \32207 );
or \U$31832 ( \32210 , \32205 , \32208 , \32209 );
and \U$31833 ( \32211 , \32200 , \32210 );
xor \U$31834 ( \32212 , \31876 , \31878 );
xor \U$31835 ( \32213 , \32212 , \31881 );
and \U$31836 ( \32214 , \32210 , \32213 );
and \U$31837 ( \32215 , \32200 , \32213 );
or \U$31838 ( \32216 , \32211 , \32214 , \32215 );
and \U$31839 ( \32217 , \32190 , \32216 );
xor \U$31840 ( \32218 , \31647 , \31657 );
xor \U$31841 ( \32219 , \32218 , \31693 );
xor \U$31842 ( \32220 , \31886 , \31888 );
xor \U$31843 ( \32221 , \32220 , \31891 );
and \U$31844 ( \32222 , \32219 , \32221 );
xor \U$31845 ( \32223 , \31864 , \31866 );
xor \U$31846 ( \32224 , \32223 , \31868 );
and \U$31847 ( \32225 , \32221 , \32224 );
and \U$31848 ( \32226 , \32219 , \32224 );
or \U$31849 ( \32227 , \32222 , \32225 , \32226 );
and \U$31850 ( \32228 , \32216 , \32227 );
and \U$31851 ( \32229 , \32190 , \32227 );
or \U$31852 ( \32230 , \32217 , \32228 , \32229 );
xor \U$31853 ( \32231 , \31373 , \31425 );
xor \U$31854 ( \32232 , \32231 , \31478 );
xor \U$31855 ( \32233 , \31884 , \31894 );
xor \U$31856 ( \32234 , \32233 , \31897 );
and \U$31857 ( \32235 , \32232 , \32234 );
xor \U$31858 ( \32236 , \31903 , \31905 );
xor \U$31859 ( \32237 , \32236 , \31908 );
and \U$31860 ( \32238 , \32234 , \32237 );
and \U$31861 ( \32239 , \32232 , \32237 );
or \U$31862 ( \32240 , \32235 , \32238 , \32239 );
and \U$31863 ( \32241 , \32230 , \32240 );
xor \U$31864 ( \32242 , \31481 , \31536 );
xor \U$31865 ( \32243 , \32242 , \31558 );
and \U$31866 ( \32244 , \32240 , \32243 );
and \U$31867 ( \32245 , \32230 , \32243 );
or \U$31868 ( \32246 , \32241 , \32244 , \32245 );
xor \U$31869 ( \32247 , \31914 , \31924 );
xor \U$31870 ( \32248 , \32247 , \31927 );
and \U$31871 ( \32249 , \32246 , \32248 );
xor \U$31872 ( \32250 , \31932 , \31934 );
xor \U$31873 ( \32251 , \32250 , \31937 );
and \U$31874 ( \32252 , \32248 , \32251 );
and \U$31875 ( \32253 , \32246 , \32251 );
or \U$31876 ( \32254 , \32249 , \32252 , \32253 );
xor \U$31877 ( \32255 , \31930 , \31940 );
xor \U$31878 ( \32256 , \32255 , \31943 );
and \U$31879 ( \32257 , \32254 , \32256 );
xor \U$31880 ( \32258 , \31601 , \31611 );
xor \U$31881 ( \32259 , \32258 , \31614 );
and \U$31882 ( \32260 , \32256 , \32259 );
and \U$31883 ( \32261 , \32254 , \32259 );
or \U$31884 ( \32262 , \32257 , \32260 , \32261 );
and \U$31885 ( \32263 , \31952 , \32262 );
xor \U$31886 ( \32264 , \31952 , \32262 );
xor \U$31887 ( \32265 , \32254 , \32256 );
xor \U$31888 ( \32266 , \32265 , \32259 );
xor \U$31889 ( \32267 , \32013 , \32017 );
xor \U$31890 ( \32268 , \32267 , \32022 );
xor \U$31891 ( \32269 , \31977 , \31981 );
xor \U$31892 ( \32270 , \32269 , \31986 );
and \U$31893 ( \32271 , \32268 , \32270 );
xor \U$31894 ( \32272 , \32029 , \32033 );
xor \U$31895 ( \32273 , \32272 , \32038 );
and \U$31896 ( \32274 , \32270 , \32273 );
and \U$31897 ( \32275 , \32268 , \32273 );
or \U$31898 ( \32276 , \32271 , \32274 , \32275 );
xor \U$31899 ( \32277 , \32065 , \32069 );
xor \U$31900 ( \32278 , \32277 , \32074 );
xor \U$31901 ( \32279 , \32081 , \32085 );
xor \U$31902 ( \32280 , \32279 , \32090 );
and \U$31903 ( \32281 , \32278 , \32280 );
xor \U$31904 ( \32282 , \32046 , \32050 );
xor \U$31905 ( \32283 , \32282 , \32055 );
and \U$31906 ( \32284 , \32280 , \32283 );
and \U$31907 ( \32285 , \32278 , \32283 );
or \U$31908 ( \32286 , \32281 , \32284 , \32285 );
and \U$31909 ( \32287 , \32276 , \32286 );
and \U$31910 ( \32288 , \29715 , \21916 );
and \U$31911 ( \32289 , \29710 , \21914 );
nor \U$31912 ( \32290 , \32288 , \32289 );
xnor \U$31913 ( \32291 , \32290 , \21867 );
and \U$31914 ( \32292 , \30318 , \21815 );
and \U$31915 ( \32293 , \30034 , \21813 );
nor \U$31916 ( \32294 , \32292 , \32293 );
xnor \U$31917 ( \32295 , \32294 , \21774 );
and \U$31918 ( \32296 , \32291 , \32295 );
and \U$31919 ( \32297 , \30895 , \21745 );
and \U$31920 ( \32298 , \30887 , \21743 );
nor \U$31921 ( \32299 , \32297 , \32298 );
xnor \U$31922 ( \32300 , \32299 , \21715 );
and \U$31923 ( \32301 , \32295 , \32300 );
and \U$31924 ( \32302 , \32291 , \32300 );
or \U$31925 ( \32303 , \32296 , \32301 , \32302 );
buf \U$31926 ( \32304 , RIc22b318_192);
nand \U$31927 ( \32305 , \32304 , \21654 );
not \U$31928 ( \32306 , \32305 );
and \U$31929 ( \32307 , \32303 , \32306 );
xor \U$31930 ( \32308 , \31993 , \31997 );
xor \U$31931 ( \32309 , \32308 , \32002 );
and \U$31932 ( \32310 , \32306 , \32309 );
and \U$31933 ( \32311 , \32303 , \32309 );
or \U$31934 ( \32312 , \32307 , \32310 , \32311 );
and \U$31935 ( \32313 , \32286 , \32312 );
and \U$31936 ( \32314 , \32276 , \32312 );
or \U$31937 ( \32315 , \32287 , \32313 , \32314 );
and \U$31938 ( \32316 , \23384 , \25692 );
and \U$31939 ( \32317 , \23379 , \25690 );
nor \U$31940 ( \32318 , \32316 , \32317 );
xnor \U$31941 ( \32319 , \32318 , \25549 );
and \U$31942 ( \32320 , \23714 , \25369 );
and \U$31943 ( \32321 , \23570 , \25367 );
nor \U$31944 ( \32322 , \32320 , \32321 );
xnor \U$31945 ( \32323 , \32322 , \25123 );
and \U$31946 ( \32324 , \32319 , \32323 );
and \U$31947 ( \32325 , \24003 , \24974 );
and \U$31948 ( \32326 , \23978 , \24972 );
nor \U$31949 ( \32327 , \32325 , \32326 );
xnor \U$31950 ( \32328 , \32327 , \24787 );
and \U$31951 ( \32329 , \32323 , \32328 );
and \U$31952 ( \32330 , \32319 , \32328 );
or \U$31953 ( \32331 , \32324 , \32329 , \32330 );
and \U$31954 ( \32332 , \22721 , \26983 );
and \U$31955 ( \32333 , \22716 , \26981 );
nor \U$31956 ( \32334 , \32332 , \32333 );
xnor \U$31957 ( \32335 , \32334 , \26742 );
and \U$31958 ( \32336 , \22952 , \26517 );
and \U$31959 ( \32337 , \22837 , \26515 );
nor \U$31960 ( \32338 , \32336 , \32337 );
xnor \U$31961 ( \32339 , \32338 , \26329 );
and \U$31962 ( \32340 , \32335 , \32339 );
and \U$31963 ( \32341 , \23136 , \26143 );
and \U$31964 ( \32342 , \23128 , \26141 );
nor \U$31965 ( \32343 , \32341 , \32342 );
xnor \U$31966 ( \32344 , \32343 , \25911 );
and \U$31967 ( \32345 , \32339 , \32344 );
and \U$31968 ( \32346 , \32335 , \32344 );
or \U$31969 ( \32347 , \32340 , \32345 , \32346 );
and \U$31970 ( \32348 , \32331 , \32347 );
and \U$31971 ( \32349 , \24344 , \24661 );
and \U$31972 ( \32350 , \24177 , \24659 );
nor \U$31973 ( \32351 , \32349 , \32350 );
xnor \U$31974 ( \32352 , \32351 , \24456 );
and \U$31975 ( \32353 , \24601 , \24255 );
and \U$31976 ( \32354 , \24482 , \24253 );
nor \U$31977 ( \32355 , \32353 , \32354 );
xnor \U$31978 ( \32356 , \32355 , \24106 );
and \U$31979 ( \32357 , \32352 , \32356 );
and \U$31980 ( \32358 , \25226 , \23933 );
and \U$31981 ( \32359 , \25018 , \23931 );
nor \U$31982 ( \32360 , \32358 , \32359 );
xnor \U$31983 ( \32361 , \32360 , \23791 );
and \U$31984 ( \32362 , \32356 , \32361 );
and \U$31985 ( \32363 , \32352 , \32361 );
or \U$31986 ( \32364 , \32357 , \32362 , \32363 );
and \U$31987 ( \32365 , \32347 , \32364 );
and \U$31988 ( \32366 , \32331 , \32364 );
or \U$31989 ( \32367 , \32348 , \32365 , \32366 );
and \U$31990 ( \32368 , \22200 , \28575 );
and \U$31991 ( \32369 , \22126 , \28573 );
nor \U$31992 ( \32370 , \32368 , \32369 );
xnor \U$31993 ( \32371 , \32370 , \28315 );
and \U$31994 ( \32372 , \22325 , \28081 );
and \U$31995 ( \32373 , \22262 , \28079 );
nor \U$31996 ( \32374 , \32372 , \32373 );
xnor \U$31997 ( \32375 , \32374 , \27766 );
and \U$31998 ( \32376 , \32371 , \32375 );
and \U$31999 ( \32377 , \22611 , \27572 );
and \U$32000 ( \32378 , \22523 , \27570 );
nor \U$32001 ( \32379 , \32377 , \32378 );
xnor \U$32002 ( \32380 , \32379 , \27232 );
and \U$32003 ( \32381 , \32375 , \32380 );
and \U$32004 ( \32382 , \32371 , \32380 );
or \U$32005 ( \32383 , \32376 , \32381 , \32382 );
and \U$32006 ( \32384 , \21836 , \30233 );
and \U$32007 ( \32385 , \21831 , \30231 );
nor \U$32008 ( \32386 , \32384 , \32385 );
xnor \U$32009 ( \32387 , \32386 , \29862 );
and \U$32010 ( \32388 , \21941 , \29671 );
and \U$32011 ( \32389 , \21890 , \29669 );
nor \U$32012 ( \32390 , \32388 , \32389 );
xnor \U$32013 ( \32391 , \32390 , \29353 );
and \U$32014 ( \32392 , \32387 , \32391 );
and \U$32015 ( \32393 , \22046 , \29104 );
and \U$32016 ( \32394 , \22018 , \29102 );
nor \U$32017 ( \32395 , \32393 , \32394 );
xnor \U$32018 ( \32396 , \32395 , \28855 );
and \U$32019 ( \32397 , \32391 , \32396 );
and \U$32020 ( \32398 , \32387 , \32396 );
or \U$32021 ( \32399 , \32392 , \32397 , \32398 );
and \U$32022 ( \32400 , \32383 , \32399 );
and \U$32023 ( \32401 , \21667 , \32151 );
and \U$32024 ( \32402 , \21653 , \32148 );
nor \U$32025 ( \32403 , \32401 , \32402 );
xnor \U$32026 ( \32404 , \32403 , \31096 );
and \U$32027 ( \32405 , \21706 , \31338 );
and \U$32028 ( \32406 , \21685 , \31336 );
nor \U$32029 ( \32407 , \32405 , \32406 );
xnor \U$32030 ( \32408 , \32407 , \31099 );
and \U$32031 ( \32409 , \32404 , \32408 );
and \U$32032 ( \32410 , \21762 , \30770 );
and \U$32033 ( \32411 , \21754 , \30768 );
nor \U$32034 ( \32412 , \32410 , \32411 );
xnor \U$32035 ( \32413 , \32412 , \30460 );
and \U$32036 ( \32414 , \32408 , \32413 );
and \U$32037 ( \32415 , \32404 , \32413 );
or \U$32038 ( \32416 , \32409 , \32414 , \32415 );
and \U$32039 ( \32417 , \32399 , \32416 );
and \U$32040 ( \32418 , \32383 , \32416 );
or \U$32041 ( \32419 , \32400 , \32417 , \32418 );
and \U$32042 ( \32420 , \32367 , \32419 );
and \U$32043 ( \32421 , \26590 , \22891 );
and \U$32044 ( \32422 , \26585 , \22889 );
nor \U$32045 ( \32423 , \32421 , \32422 );
xnor \U$32046 ( \32424 , \32423 , \22778 );
and \U$32047 ( \32425 , \27113 , \22697 );
and \U$32048 ( \32426 , \26854 , \22695 );
nor \U$32049 ( \32427 , \32425 , \32426 );
xnor \U$32050 ( \32428 , \32427 , \22561 );
and \U$32051 ( \32429 , \32424 , \32428 );
and \U$32052 ( \32430 , \27494 , \22497 );
and \U$32053 ( \32431 , \27485 , \22495 );
nor \U$32054 ( \32432 , \32430 , \32431 );
xnor \U$32055 ( \32433 , \32432 , \22419 );
and \U$32056 ( \32434 , \32428 , \32433 );
and \U$32057 ( \32435 , \32424 , \32433 );
or \U$32058 ( \32436 , \32429 , \32434 , \32435 );
and \U$32059 ( \32437 , \25353 , \23637 );
and \U$32060 ( \32438 , \25348 , \23635 );
nor \U$32061 ( \32439 , \32437 , \32438 );
xnor \U$32062 ( \32440 , \32439 , \23500 );
and \U$32063 ( \32441 , \25806 , \23431 );
and \U$32064 ( \32442 , \25609 , \23429 );
nor \U$32065 ( \32443 , \32441 , \32442 );
xnor \U$32066 ( \32444 , \32443 , \23279 );
and \U$32067 ( \32445 , \32440 , \32444 );
and \U$32068 ( \32446 , \26116 , \23163 );
and \U$32069 ( \32447 , \26108 , \23161 );
nor \U$32070 ( \32448 , \32446 , \32447 );
xnor \U$32071 ( \32449 , \32448 , \23007 );
and \U$32072 ( \32450 , \32444 , \32449 );
and \U$32073 ( \32451 , \32440 , \32449 );
or \U$32074 ( \32452 , \32445 , \32450 , \32451 );
and \U$32075 ( \32453 , \32436 , \32452 );
and \U$32076 ( \32454 , \28039 , \22333 );
and \U$32077 ( \32455 , \27837 , \22331 );
nor \U$32078 ( \32456 , \32454 , \32455 );
xnor \U$32079 ( \32457 , \32456 , \22239 );
and \U$32080 ( \32458 , \28514 , \22163 );
and \U$32081 ( \32459 , \28342 , \22161 );
nor \U$32082 ( \32460 , \32458 , \32459 );
xnor \U$32083 ( \32461 , \32460 , \22091 );
and \U$32084 ( \32462 , \32457 , \32461 );
and \U$32085 ( \32463 , \29464 , \22029 );
and \U$32086 ( \32464 , \29040 , \22027 );
nor \U$32087 ( \32465 , \32463 , \32464 );
xnor \U$32088 ( \32466 , \32465 , \21986 );
and \U$32089 ( \32467 , \32461 , \32466 );
and \U$32090 ( \32468 , \32457 , \32466 );
or \U$32091 ( \32469 , \32462 , \32467 , \32468 );
and \U$32092 ( \32470 , \32452 , \32469 );
and \U$32093 ( \32471 , \32436 , \32469 );
or \U$32094 ( \32472 , \32453 , \32470 , \32471 );
and \U$32095 ( \32473 , \32419 , \32472 );
and \U$32096 ( \32474 , \32367 , \32472 );
or \U$32097 ( \32475 , \32420 , \32473 , \32474 );
and \U$32098 ( \32476 , \32315 , \32475 );
xor \U$32099 ( \32477 , \32118 , \32122 );
xor \U$32100 ( \32478 , \32477 , \32127 );
xor \U$32101 ( \32479 , \32134 , \32138 );
xor \U$32102 ( \32480 , \32479 , \32143 );
and \U$32103 ( \32481 , \32478 , \32480 );
xor \U$32104 ( \32482 , \32098 , \32102 );
xor \U$32105 ( \32483 , \32482 , \32107 );
and \U$32106 ( \32484 , \32480 , \32483 );
and \U$32107 ( \32485 , \32478 , \32483 );
or \U$32108 ( \32486 , \32481 , \32484 , \32485 );
xor \U$32109 ( \32487 , \32168 , \32170 );
xor \U$32110 ( \32488 , \32487 , \32173 );
and \U$32111 ( \32489 , \32486 , \32488 );
xor \U$32112 ( \32490 , \32178 , \32180 );
and \U$32113 ( \32491 , \32488 , \32490 );
and \U$32114 ( \32492 , \32486 , \32490 );
or \U$32115 ( \32493 , \32489 , \32491 , \32492 );
and \U$32116 ( \32494 , \32475 , \32493 );
and \U$32117 ( \32495 , \32315 , \32493 );
or \U$32118 ( \32496 , \32476 , \32494 , \32495 );
xor \U$32119 ( \32497 , \32025 , \32041 );
xor \U$32120 ( \32498 , \32497 , \32058 );
xor \U$32121 ( \32499 , \32077 , \32093 );
xor \U$32122 ( \32500 , \32499 , \32110 );
and \U$32123 ( \32501 , \32498 , \32500 );
xor \U$32124 ( \32502 , \32130 , \32146 );
xor \U$32125 ( \32503 , \32502 , \32159 );
and \U$32126 ( \32504 , \32500 , \32503 );
and \U$32127 ( \32505 , \32498 , \32503 );
or \U$32128 ( \32506 , \32501 , \32504 , \32505 );
xor \U$32129 ( \32507 , \31954 , \31956 );
xor \U$32130 ( \32508 , \32507 , \31959 );
xor \U$32131 ( \32509 , \31964 , \31966 );
xor \U$32132 ( \32510 , \32509 , \31969 );
and \U$32133 ( \32511 , \32508 , \32510 );
xnor \U$32134 ( \32512 , \31989 , \32005 );
and \U$32135 ( \32513 , \32510 , \32512 );
and \U$32136 ( \32514 , \32508 , \32512 );
or \U$32137 ( \32515 , \32511 , \32513 , \32514 );
and \U$32138 ( \32516 , \32506 , \32515 );
xor \U$32139 ( \32517 , \31709 , \31725 );
xor \U$32140 ( \32518 , \32517 , \31742 );
and \U$32141 ( \32519 , \32515 , \32518 );
and \U$32142 ( \32520 , \32506 , \32518 );
or \U$32143 ( \32521 , \32516 , \32519 , \32520 );
and \U$32144 ( \32522 , \32496 , \32521 );
xor \U$32145 ( \32523 , \32176 , \32181 );
xor \U$32146 ( \32524 , \32523 , \32184 );
xor \U$32147 ( \32525 , \32192 , \32194 );
xor \U$32148 ( \32526 , \32525 , \32197 );
and \U$32149 ( \32527 , \32524 , \32526 );
xor \U$32150 ( \32528 , \32202 , \32204 );
xor \U$32151 ( \32529 , \32528 , \32207 );
and \U$32152 ( \32530 , \32526 , \32529 );
and \U$32153 ( \32531 , \32524 , \32529 );
or \U$32154 ( \32532 , \32527 , \32530 , \32531 );
and \U$32155 ( \32533 , \32521 , \32532 );
and \U$32156 ( \32534 , \32496 , \32532 );
or \U$32157 ( \32535 , \32522 , \32533 , \32534 );
xor \U$32158 ( \32536 , \31745 , \31797 );
xor \U$32159 ( \32537 , \32536 , \31850 );
xor \U$32160 ( \32538 , \32200 , \32210 );
xor \U$32161 ( \32539 , \32538 , \32213 );
and \U$32162 ( \32540 , \32537 , \32539 );
xor \U$32163 ( \32541 , \32219 , \32221 );
xor \U$32164 ( \32542 , \32541 , \32224 );
and \U$32165 ( \32543 , \32539 , \32542 );
and \U$32166 ( \32544 , \32537 , \32542 );
or \U$32167 ( \32545 , \32540 , \32543 , \32544 );
and \U$32168 ( \32546 , \32535 , \32545 );
xor \U$32169 ( \32547 , \31696 , \31853 );
xor \U$32170 ( \32548 , \32547 , \31871 );
and \U$32171 ( \32549 , \32545 , \32548 );
and \U$32172 ( \32550 , \32535 , \32548 );
or \U$32173 ( \32551 , \32546 , \32549 , \32550 );
xor \U$32174 ( \32552 , \32190 , \32216 );
xor \U$32175 ( \32553 , \32552 , \32227 );
xor \U$32176 ( \32554 , \32232 , \32234 );
xor \U$32177 ( \32555 , \32554 , \32237 );
and \U$32178 ( \32556 , \32553 , \32555 );
and \U$32179 ( \32557 , \32551 , \32556 );
xor \U$32180 ( \32558 , \31916 , \31918 );
xor \U$32181 ( \32559 , \32558 , \31921 );
and \U$32182 ( \32560 , \32556 , \32559 );
and \U$32183 ( \32561 , \32551 , \32559 );
or \U$32184 ( \32562 , \32557 , \32560 , \32561 );
xor \U$32185 ( \32563 , \31874 , \31900 );
xor \U$32186 ( \32564 , \32563 , \31911 );
xor \U$32187 ( \32565 , \32230 , \32240 );
xor \U$32188 ( \32566 , \32565 , \32243 );
and \U$32189 ( \32567 , \32564 , \32566 );
and \U$32190 ( \32568 , \32562 , \32567 );
xor \U$32191 ( \32569 , \32246 , \32248 );
xor \U$32192 ( \32570 , \32569 , \32251 );
and \U$32193 ( \32571 , \32567 , \32570 );
and \U$32194 ( \32572 , \32562 , \32570 );
or \U$32195 ( \32573 , \32568 , \32571 , \32572 );
and \U$32196 ( \32574 , \32266 , \32573 );
xor \U$32197 ( \32575 , \32266 , \32573 );
xor \U$32198 ( \32576 , \32562 , \32567 );
xor \U$32199 ( \32577 , \32576 , \32570 );
and \U$32200 ( \32578 , \31498 , \21745 );
and \U$32201 ( \32579 , \30895 , \21743 );
nor \U$32202 ( \32580 , \32578 , \32579 );
xnor \U$32203 ( \32581 , \32580 , \21715 );
and \U$32204 ( \32582 , \31684 , \21697 );
and \U$32205 ( \32583 , \31503 , \21695 );
nor \U$32206 ( \32584 , \32582 , \32583 );
xnor \U$32207 ( \32585 , \32584 , \21678 );
and \U$32208 ( \32586 , \32581 , \32585 );
nand \U$32209 ( \32587 , \32304 , \21658 );
xnor \U$32210 ( \32588 , \32587 , \21665 );
and \U$32211 ( \32589 , \32585 , \32588 );
and \U$32212 ( \32590 , \32581 , \32588 );
or \U$32213 ( \32591 , \32586 , \32589 , \32590 );
and \U$32214 ( \32592 , \29710 , \22029 );
and \U$32215 ( \32593 , \29464 , \22027 );
nor \U$32216 ( \32594 , \32592 , \32593 );
xnor \U$32217 ( \32595 , \32594 , \21986 );
and \U$32218 ( \32596 , \30034 , \21916 );
and \U$32219 ( \32597 , \29715 , \21914 );
nor \U$32220 ( \32598 , \32596 , \32597 );
xnor \U$32221 ( \32599 , \32598 , \21867 );
and \U$32222 ( \32600 , \32595 , \32599 );
and \U$32223 ( \32601 , \30887 , \21815 );
and \U$32224 ( \32602 , \30318 , \21813 );
nor \U$32225 ( \32603 , \32601 , \32602 );
xnor \U$32226 ( \32604 , \32603 , \21774 );
and \U$32227 ( \32605 , \32599 , \32604 );
and \U$32228 ( \32606 , \32595 , \32604 );
or \U$32229 ( \32607 , \32600 , \32605 , \32606 );
and \U$32230 ( \32608 , \32591 , \32607 );
and \U$32231 ( \32609 , \31503 , \21697 );
and \U$32232 ( \32610 , \31498 , \21695 );
nor \U$32233 ( \32611 , \32609 , \32610 );
xnor \U$32234 ( \32612 , \32611 , \21678 );
and \U$32235 ( \32613 , \32607 , \32612 );
and \U$32236 ( \32614 , \32591 , \32612 );
or \U$32237 ( \32615 , \32608 , \32613 , \32614 );
and \U$32238 ( \32616 , \32304 , \21660 );
and \U$32239 ( \32617 , \31684 , \21658 );
nor \U$32240 ( \32618 , \32616 , \32617 );
xnor \U$32241 ( \32619 , \32618 , \21665 );
xor \U$32242 ( \32620 , \32457 , \32461 );
xor \U$32243 ( \32621 , \32620 , \32466 );
and \U$32244 ( \32622 , \32619 , \32621 );
xor \U$32245 ( \32623 , \32291 , \32295 );
xor \U$32246 ( \32624 , \32623 , \32300 );
and \U$32247 ( \32625 , \32621 , \32624 );
and \U$32248 ( \32626 , \32619 , \32624 );
or \U$32249 ( \32627 , \32622 , \32625 , \32626 );
and \U$32250 ( \32628 , \32615 , \32627 );
xor \U$32251 ( \32629 , \32424 , \32428 );
xor \U$32252 ( \32630 , \32629 , \32433 );
xor \U$32253 ( \32631 , \32440 , \32444 );
xor \U$32254 ( \32632 , \32631 , \32449 );
and \U$32255 ( \32633 , \32630 , \32632 );
xor \U$32256 ( \32634 , \32352 , \32356 );
xor \U$32257 ( \32635 , \32634 , \32361 );
and \U$32258 ( \32636 , \32632 , \32635 );
and \U$32259 ( \32637 , \32630 , \32635 );
or \U$32260 ( \32638 , \32633 , \32636 , \32637 );
and \U$32261 ( \32639 , \32627 , \32638 );
and \U$32262 ( \32640 , \32615 , \32638 );
or \U$32263 ( \32641 , \32628 , \32639 , \32640 );
and \U$32264 ( \32642 , \26585 , \23163 );
and \U$32265 ( \32643 , \26116 , \23161 );
nor \U$32266 ( \32644 , \32642 , \32643 );
xnor \U$32267 ( \32645 , \32644 , \23007 );
and \U$32268 ( \32646 , \26854 , \22891 );
and \U$32269 ( \32647 , \26590 , \22889 );
nor \U$32270 ( \32648 , \32646 , \32647 );
xnor \U$32271 ( \32649 , \32648 , \22778 );
and \U$32272 ( \32650 , \32645 , \32649 );
and \U$32273 ( \32651 , \27485 , \22697 );
and \U$32274 ( \32652 , \27113 , \22695 );
nor \U$32275 ( \32653 , \32651 , \32652 );
xnor \U$32276 ( \32654 , \32653 , \22561 );
and \U$32277 ( \32655 , \32649 , \32654 );
and \U$32278 ( \32656 , \32645 , \32654 );
or \U$32279 ( \32657 , \32650 , \32655 , \32656 );
and \U$32280 ( \32658 , \25348 , \23933 );
and \U$32281 ( \32659 , \25226 , \23931 );
nor \U$32282 ( \32660 , \32658 , \32659 );
xnor \U$32283 ( \32661 , \32660 , \23791 );
and \U$32284 ( \32662 , \25609 , \23637 );
and \U$32285 ( \32663 , \25353 , \23635 );
nor \U$32286 ( \32664 , \32662 , \32663 );
xnor \U$32287 ( \32665 , \32664 , \23500 );
and \U$32288 ( \32666 , \32661 , \32665 );
and \U$32289 ( \32667 , \26108 , \23431 );
and \U$32290 ( \32668 , \25806 , \23429 );
nor \U$32291 ( \32669 , \32667 , \32668 );
xnor \U$32292 ( \32670 , \32669 , \23279 );
and \U$32293 ( \32671 , \32665 , \32670 );
and \U$32294 ( \32672 , \32661 , \32670 );
or \U$32295 ( \32673 , \32666 , \32671 , \32672 );
and \U$32296 ( \32674 , \32657 , \32673 );
and \U$32297 ( \32675 , \27837 , \22497 );
and \U$32298 ( \32676 , \27494 , \22495 );
nor \U$32299 ( \32677 , \32675 , \32676 );
xnor \U$32300 ( \32678 , \32677 , \22419 );
and \U$32301 ( \32679 , \28342 , \22333 );
and \U$32302 ( \32680 , \28039 , \22331 );
nor \U$32303 ( \32681 , \32679 , \32680 );
xnor \U$32304 ( \32682 , \32681 , \22239 );
and \U$32305 ( \32683 , \32678 , \32682 );
and \U$32306 ( \32684 , \29040 , \22163 );
and \U$32307 ( \32685 , \28514 , \22161 );
nor \U$32308 ( \32686 , \32684 , \32685 );
xnor \U$32309 ( \32687 , \32686 , \22091 );
and \U$32310 ( \32688 , \32682 , \32687 );
and \U$32311 ( \32689 , \32678 , \32687 );
or \U$32312 ( \32690 , \32683 , \32688 , \32689 );
and \U$32313 ( \32691 , \32673 , \32690 );
and \U$32314 ( \32692 , \32657 , \32690 );
or \U$32315 ( \32693 , \32674 , \32691 , \32692 );
and \U$32316 ( \32694 , \22126 , \29104 );
and \U$32317 ( \32695 , \22046 , \29102 );
nor \U$32318 ( \32696 , \32694 , \32695 );
xnor \U$32319 ( \32697 , \32696 , \28855 );
and \U$32320 ( \32698 , \22262 , \28575 );
and \U$32321 ( \32699 , \22200 , \28573 );
nor \U$32322 ( \32700 , \32698 , \32699 );
xnor \U$32323 ( \32701 , \32700 , \28315 );
and \U$32324 ( \32702 , \32697 , \32701 );
and \U$32325 ( \32703 , \22523 , \28081 );
and \U$32326 ( \32704 , \22325 , \28079 );
nor \U$32327 ( \32705 , \32703 , \32704 );
xnor \U$32328 ( \32706 , \32705 , \27766 );
and \U$32329 ( \32707 , \32701 , \32706 );
and \U$32330 ( \32708 , \32697 , \32706 );
or \U$32331 ( \32709 , \32702 , \32707 , \32708 );
and \U$32332 ( \32710 , \21685 , \32151 );
and \U$32333 ( \32711 , \21667 , \32148 );
nor \U$32334 ( \32712 , \32710 , \32711 );
xnor \U$32335 ( \32713 , \32712 , \31096 );
and \U$32336 ( \32714 , \21754 , \31338 );
and \U$32337 ( \32715 , \21706 , \31336 );
nor \U$32338 ( \32716 , \32714 , \32715 );
xnor \U$32339 ( \32717 , \32716 , \31099 );
and \U$32340 ( \32718 , \32713 , \32717 );
and \U$32341 ( \32719 , \32717 , \21665 );
and \U$32342 ( \32720 , \32713 , \21665 );
or \U$32343 ( \32721 , \32718 , \32719 , \32720 );
and \U$32344 ( \32722 , \32709 , \32721 );
and \U$32345 ( \32723 , \21831 , \30770 );
and \U$32346 ( \32724 , \21762 , \30768 );
nor \U$32347 ( \32725 , \32723 , \32724 );
xnor \U$32348 ( \32726 , \32725 , \30460 );
and \U$32349 ( \32727 , \21890 , \30233 );
and \U$32350 ( \32728 , \21836 , \30231 );
nor \U$32351 ( \32729 , \32727 , \32728 );
xnor \U$32352 ( \32730 , \32729 , \29862 );
and \U$32353 ( \32731 , \32726 , \32730 );
and \U$32354 ( \32732 , \22018 , \29671 );
and \U$32355 ( \32733 , \21941 , \29669 );
nor \U$32356 ( \32734 , \32732 , \32733 );
xnor \U$32357 ( \32735 , \32734 , \29353 );
and \U$32358 ( \32736 , \32730 , \32735 );
and \U$32359 ( \32737 , \32726 , \32735 );
or \U$32360 ( \32738 , \32731 , \32736 , \32737 );
and \U$32361 ( \32739 , \32721 , \32738 );
and \U$32362 ( \32740 , \32709 , \32738 );
or \U$32363 ( \32741 , \32722 , \32739 , \32740 );
and \U$32364 ( \32742 , \32693 , \32741 );
and \U$32365 ( \32743 , \23379 , \26143 );
and \U$32366 ( \32744 , \23136 , \26141 );
nor \U$32367 ( \32745 , \32743 , \32744 );
xnor \U$32368 ( \32746 , \32745 , \25911 );
and \U$32369 ( \32747 , \23570 , \25692 );
and \U$32370 ( \32748 , \23384 , \25690 );
nor \U$32371 ( \32749 , \32747 , \32748 );
xnor \U$32372 ( \32750 , \32749 , \25549 );
and \U$32373 ( \32751 , \32746 , \32750 );
and \U$32374 ( \32752 , \23978 , \25369 );
and \U$32375 ( \32753 , \23714 , \25367 );
nor \U$32376 ( \32754 , \32752 , \32753 );
xnor \U$32377 ( \32755 , \32754 , \25123 );
and \U$32378 ( \32756 , \32750 , \32755 );
and \U$32379 ( \32757 , \32746 , \32755 );
or \U$32380 ( \32758 , \32751 , \32756 , \32757 );
and \U$32381 ( \32759 , \22716 , \27572 );
and \U$32382 ( \32760 , \22611 , \27570 );
nor \U$32383 ( \32761 , \32759 , \32760 );
xnor \U$32384 ( \32762 , \32761 , \27232 );
and \U$32385 ( \32763 , \22837 , \26983 );
and \U$32386 ( \32764 , \22721 , \26981 );
nor \U$32387 ( \32765 , \32763 , \32764 );
xnor \U$32388 ( \32766 , \32765 , \26742 );
and \U$32389 ( \32767 , \32762 , \32766 );
and \U$32390 ( \32768 , \23128 , \26517 );
and \U$32391 ( \32769 , \22952 , \26515 );
nor \U$32392 ( \32770 , \32768 , \32769 );
xnor \U$32393 ( \32771 , \32770 , \26329 );
and \U$32394 ( \32772 , \32766 , \32771 );
and \U$32395 ( \32773 , \32762 , \32771 );
or \U$32396 ( \32774 , \32767 , \32772 , \32773 );
and \U$32397 ( \32775 , \32758 , \32774 );
and \U$32398 ( \32776 , \24177 , \24974 );
and \U$32399 ( \32777 , \24003 , \24972 );
nor \U$32400 ( \32778 , \32776 , \32777 );
xnor \U$32401 ( \32779 , \32778 , \24787 );
and \U$32402 ( \32780 , \24482 , \24661 );
and \U$32403 ( \32781 , \24344 , \24659 );
nor \U$32404 ( \32782 , \32780 , \32781 );
xnor \U$32405 ( \32783 , \32782 , \24456 );
and \U$32406 ( \32784 , \32779 , \32783 );
and \U$32407 ( \32785 , \25018 , \24255 );
and \U$32408 ( \32786 , \24601 , \24253 );
nor \U$32409 ( \32787 , \32785 , \32786 );
xnor \U$32410 ( \32788 , \32787 , \24106 );
and \U$32411 ( \32789 , \32783 , \32788 );
and \U$32412 ( \32790 , \32779 , \32788 );
or \U$32413 ( \32791 , \32784 , \32789 , \32790 );
and \U$32414 ( \32792 , \32774 , \32791 );
and \U$32415 ( \32793 , \32758 , \32791 );
or \U$32416 ( \32794 , \32775 , \32792 , \32793 );
and \U$32417 ( \32795 , \32741 , \32794 );
and \U$32418 ( \32796 , \32693 , \32794 );
or \U$32419 ( \32797 , \32742 , \32795 , \32796 );
and \U$32420 ( \32798 , \32641 , \32797 );
xor \U$32421 ( \32799 , \32319 , \32323 );
xor \U$32422 ( \32800 , \32799 , \32328 );
xor \U$32423 ( \32801 , \32335 , \32339 );
xor \U$32424 ( \32802 , \32801 , \32344 );
and \U$32425 ( \32803 , \32800 , \32802 );
xor \U$32426 ( \32804 , \32371 , \32375 );
xor \U$32427 ( \32805 , \32804 , \32380 );
and \U$32428 ( \32806 , \32802 , \32805 );
and \U$32429 ( \32807 , \32800 , \32805 );
or \U$32430 ( \32808 , \32803 , \32806 , \32807 );
xor \U$32431 ( \32809 , \32387 , \32391 );
xor \U$32432 ( \32810 , \32809 , \32396 );
xor \U$32433 ( \32811 , \32404 , \32408 );
xor \U$32434 ( \32812 , \32811 , \32413 );
and \U$32435 ( \32813 , \32810 , \32812 );
and \U$32436 ( \32814 , \32808 , \32813 );
xor \U$32437 ( \32815 , \32154 , \32158 );
and \U$32438 ( \32816 , \32813 , \32815 );
and \U$32439 ( \32817 , \32808 , \32815 );
or \U$32440 ( \32818 , \32814 , \32816 , \32817 );
and \U$32441 ( \32819 , \32797 , \32818 );
and \U$32442 ( \32820 , \32641 , \32818 );
or \U$32443 ( \32821 , \32798 , \32819 , \32820 );
xor \U$32444 ( \32822 , \32331 , \32347 );
xor \U$32445 ( \32823 , \32822 , \32364 );
xor \U$32446 ( \32824 , \32436 , \32452 );
xor \U$32447 ( \32825 , \32824 , \32469 );
and \U$32448 ( \32826 , \32823 , \32825 );
xor \U$32449 ( \32827 , \32303 , \32306 );
xor \U$32450 ( \32828 , \32827 , \32309 );
and \U$32451 ( \32829 , \32825 , \32828 );
and \U$32452 ( \32830 , \32823 , \32828 );
or \U$32453 ( \32831 , \32826 , \32829 , \32830 );
xor \U$32454 ( \32832 , \32478 , \32480 );
xor \U$32455 ( \32833 , \32832 , \32483 );
xor \U$32456 ( \32834 , \32268 , \32270 );
xor \U$32457 ( \32835 , \32834 , \32273 );
and \U$32458 ( \32836 , \32833 , \32835 );
xor \U$32459 ( \32837 , \32278 , \32280 );
xor \U$32460 ( \32838 , \32837 , \32283 );
and \U$32461 ( \32839 , \32835 , \32838 );
and \U$32462 ( \32840 , \32833 , \32838 );
or \U$32463 ( \32841 , \32836 , \32839 , \32840 );
and \U$32464 ( \32842 , \32831 , \32841 );
xor \U$32465 ( \32843 , \32498 , \32500 );
xor \U$32466 ( \32844 , \32843 , \32503 );
and \U$32467 ( \32845 , \32841 , \32844 );
and \U$32468 ( \32846 , \32831 , \32844 );
or \U$32469 ( \32847 , \32842 , \32845 , \32846 );
and \U$32470 ( \32848 , \32821 , \32847 );
xor \U$32471 ( \32849 , \32276 , \32286 );
xor \U$32472 ( \32850 , \32849 , \32312 );
xor \U$32473 ( \32851 , \32508 , \32510 );
xor \U$32474 ( \32852 , \32851 , \32512 );
and \U$32475 ( \32853 , \32850 , \32852 );
xor \U$32476 ( \32854 , \32486 , \32488 );
xor \U$32477 ( \32855 , \32854 , \32490 );
and \U$32478 ( \32856 , \32852 , \32855 );
and \U$32479 ( \32857 , \32850 , \32855 );
or \U$32480 ( \32858 , \32853 , \32856 , \32857 );
and \U$32481 ( \32859 , \32847 , \32858 );
and \U$32482 ( \32860 , \32821 , \32858 );
or \U$32483 ( \32861 , \32848 , \32859 , \32860 );
xor \U$32484 ( \32862 , \31962 , \31972 );
xor \U$32485 ( \32863 , \32862 , \32006 );
xor \U$32486 ( \32864 , \32061 , \32113 );
xor \U$32487 ( \32865 , \32864 , \32162 );
and \U$32488 ( \32866 , \32863 , \32865 );
xor \U$32489 ( \32867 , \32524 , \32526 );
xor \U$32490 ( \32868 , \32867 , \32529 );
and \U$32491 ( \32869 , \32865 , \32868 );
and \U$32492 ( \32870 , \32863 , \32868 );
or \U$32493 ( \32871 , \32866 , \32869 , \32870 );
and \U$32494 ( \32872 , \32861 , \32871 );
xor \U$32495 ( \32873 , \32009 , \32165 );
xor \U$32496 ( \32874 , \32873 , \32187 );
and \U$32497 ( \32875 , \32871 , \32874 );
and \U$32498 ( \32876 , \32861 , \32874 );
or \U$32499 ( \32877 , \32872 , \32875 , \32876 );
xor \U$32500 ( \32878 , \32535 , \32545 );
xor \U$32501 ( \32879 , \32878 , \32548 );
and \U$32502 ( \32880 , \32877 , \32879 );
xor \U$32503 ( \32881 , \32553 , \32555 );
and \U$32504 ( \32882 , \32879 , \32881 );
and \U$32505 ( \32883 , \32877 , \32881 );
or \U$32506 ( \32884 , \32880 , \32882 , \32883 );
xor \U$32507 ( \32885 , \32551 , \32556 );
xor \U$32508 ( \32886 , \32885 , \32559 );
and \U$32509 ( \32887 , \32884 , \32886 );
xor \U$32510 ( \32888 , \32564 , \32566 );
and \U$32511 ( \32889 , \32886 , \32888 );
and \U$32512 ( \32890 , \32884 , \32888 );
or \U$32513 ( \32891 , \32887 , \32889 , \32890 );
and \U$32514 ( \32892 , \32577 , \32891 );
xor \U$32515 ( \32893 , \32577 , \32891 );
xor \U$32516 ( \32894 , \32884 , \32886 );
xor \U$32517 ( \32895 , \32894 , \32888 );
and \U$32518 ( \32896 , \21941 , \30233 );
and \U$32519 ( \32897 , \21890 , \30231 );
nor \U$32520 ( \32898 , \32896 , \32897 );
xnor \U$32521 ( \32899 , \32898 , \29862 );
and \U$32522 ( \32900 , \22046 , \29671 );
and \U$32523 ( \32901 , \22018 , \29669 );
nor \U$32524 ( \32902 , \32900 , \32901 );
xnor \U$32525 ( \32903 , \32902 , \29353 );
and \U$32526 ( \32904 , \32899 , \32903 );
and \U$32527 ( \32905 , \22200 , \29104 );
and \U$32528 ( \32906 , \22126 , \29102 );
nor \U$32529 ( \32907 , \32905 , \32906 );
xnor \U$32530 ( \32908 , \32907 , \28855 );
and \U$32531 ( \32909 , \32903 , \32908 );
and \U$32532 ( \32910 , \32899 , \32908 );
or \U$32533 ( \32911 , \32904 , \32909 , \32910 );
and \U$32534 ( \32912 , \21706 , \32151 );
and \U$32535 ( \32913 , \21685 , \32148 );
nor \U$32536 ( \32914 , \32912 , \32913 );
xnor \U$32537 ( \32915 , \32914 , \31096 );
and \U$32538 ( \32916 , \21762 , \31338 );
and \U$32539 ( \32917 , \21754 , \31336 );
nor \U$32540 ( \32918 , \32916 , \32917 );
xnor \U$32541 ( \32919 , \32918 , \31099 );
and \U$32542 ( \32920 , \32915 , \32919 );
and \U$32543 ( \32921 , \21836 , \30770 );
and \U$32544 ( \32922 , \21831 , \30768 );
nor \U$32545 ( \32923 , \32921 , \32922 );
xnor \U$32546 ( \32924 , \32923 , \30460 );
and \U$32547 ( \32925 , \32919 , \32924 );
and \U$32548 ( \32926 , \32915 , \32924 );
or \U$32549 ( \32927 , \32920 , \32925 , \32926 );
and \U$32550 ( \32928 , \32911 , \32927 );
and \U$32551 ( \32929 , \22325 , \28575 );
and \U$32552 ( \32930 , \22262 , \28573 );
nor \U$32553 ( \32931 , \32929 , \32930 );
xnor \U$32554 ( \32932 , \32931 , \28315 );
and \U$32555 ( \32933 , \22611 , \28081 );
and \U$32556 ( \32934 , \22523 , \28079 );
nor \U$32557 ( \32935 , \32933 , \32934 );
xnor \U$32558 ( \32936 , \32935 , \27766 );
and \U$32559 ( \32937 , \32932 , \32936 );
and \U$32560 ( \32938 , \22721 , \27572 );
and \U$32561 ( \32939 , \22716 , \27570 );
nor \U$32562 ( \32940 , \32938 , \32939 );
xnor \U$32563 ( \32941 , \32940 , \27232 );
and \U$32564 ( \32942 , \32936 , \32941 );
and \U$32565 ( \32943 , \32932 , \32941 );
or \U$32566 ( \32944 , \32937 , \32942 , \32943 );
and \U$32567 ( \32945 , \32927 , \32944 );
and \U$32568 ( \32946 , \32911 , \32944 );
or \U$32569 ( \32947 , \32928 , \32945 , \32946 );
and \U$32570 ( \32948 , \27113 , \22891 );
and \U$32571 ( \32949 , \26854 , \22889 );
nor \U$32572 ( \32950 , \32948 , \32949 );
xnor \U$32573 ( \32951 , \32950 , \22778 );
and \U$32574 ( \32952 , \27494 , \22697 );
and \U$32575 ( \32953 , \27485 , \22695 );
nor \U$32576 ( \32954 , \32952 , \32953 );
xnor \U$32577 ( \32955 , \32954 , \22561 );
and \U$32578 ( \32956 , \32951 , \32955 );
and \U$32579 ( \32957 , \28039 , \22497 );
and \U$32580 ( \32958 , \27837 , \22495 );
nor \U$32581 ( \32959 , \32957 , \32958 );
xnor \U$32582 ( \32960 , \32959 , \22419 );
and \U$32583 ( \32961 , \32955 , \32960 );
and \U$32584 ( \32962 , \32951 , \32960 );
or \U$32585 ( \32963 , \32956 , \32961 , \32962 );
and \U$32586 ( \32964 , \28514 , \22333 );
and \U$32587 ( \32965 , \28342 , \22331 );
nor \U$32588 ( \32966 , \32964 , \32965 );
xnor \U$32589 ( \32967 , \32966 , \22239 );
and \U$32590 ( \32968 , \29464 , \22163 );
and \U$32591 ( \32969 , \29040 , \22161 );
nor \U$32592 ( \32970 , \32968 , \32969 );
xnor \U$32593 ( \32971 , \32970 , \22091 );
and \U$32594 ( \32972 , \32967 , \32971 );
and \U$32595 ( \32973 , \29715 , \22029 );
and \U$32596 ( \32974 , \29710 , \22027 );
nor \U$32597 ( \32975 , \32973 , \32974 );
xnor \U$32598 ( \32976 , \32975 , \21986 );
and \U$32599 ( \32977 , \32971 , \32976 );
and \U$32600 ( \32978 , \32967 , \32976 );
or \U$32601 ( \32979 , \32972 , \32977 , \32978 );
and \U$32602 ( \32980 , \32963 , \32979 );
and \U$32603 ( \32981 , \25806 , \23637 );
and \U$32604 ( \32982 , \25609 , \23635 );
nor \U$32605 ( \32983 , \32981 , \32982 );
xnor \U$32606 ( \32984 , \32983 , \23500 );
and \U$32607 ( \32985 , \26116 , \23431 );
and \U$32608 ( \32986 , \26108 , \23429 );
nor \U$32609 ( \32987 , \32985 , \32986 );
xnor \U$32610 ( \32988 , \32987 , \23279 );
and \U$32611 ( \32989 , \32984 , \32988 );
and \U$32612 ( \32990 , \26590 , \23163 );
and \U$32613 ( \32991 , \26585 , \23161 );
nor \U$32614 ( \32992 , \32990 , \32991 );
xnor \U$32615 ( \32993 , \32992 , \23007 );
and \U$32616 ( \32994 , \32988 , \32993 );
and \U$32617 ( \32995 , \32984 , \32993 );
or \U$32618 ( \32996 , \32989 , \32994 , \32995 );
and \U$32619 ( \32997 , \32979 , \32996 );
and \U$32620 ( \32998 , \32963 , \32996 );
or \U$32621 ( \32999 , \32980 , \32997 , \32998 );
and \U$32622 ( \33000 , \32947 , \32999 );
and \U$32623 ( \33001 , \22952 , \26983 );
and \U$32624 ( \33002 , \22837 , \26981 );
nor \U$32625 ( \33003 , \33001 , \33002 );
xnor \U$32626 ( \33004 , \33003 , \26742 );
and \U$32627 ( \33005 , \23136 , \26517 );
and \U$32628 ( \33006 , \23128 , \26515 );
nor \U$32629 ( \33007 , \33005 , \33006 );
xnor \U$32630 ( \33008 , \33007 , \26329 );
and \U$32631 ( \33009 , \33004 , \33008 );
and \U$32632 ( \33010 , \23384 , \26143 );
and \U$32633 ( \33011 , \23379 , \26141 );
nor \U$32634 ( \33012 , \33010 , \33011 );
xnor \U$32635 ( \33013 , \33012 , \25911 );
and \U$32636 ( \33014 , \33008 , \33013 );
and \U$32637 ( \33015 , \33004 , \33013 );
or \U$32638 ( \33016 , \33009 , \33014 , \33015 );
and \U$32639 ( \33017 , \24601 , \24661 );
and \U$32640 ( \33018 , \24482 , \24659 );
nor \U$32641 ( \33019 , \33017 , \33018 );
xnor \U$32642 ( \33020 , \33019 , \24456 );
and \U$32643 ( \33021 , \25226 , \24255 );
and \U$32644 ( \33022 , \25018 , \24253 );
nor \U$32645 ( \33023 , \33021 , \33022 );
xnor \U$32646 ( \33024 , \33023 , \24106 );
and \U$32647 ( \33025 , \33020 , \33024 );
and \U$32648 ( \33026 , \25353 , \23933 );
and \U$32649 ( \33027 , \25348 , \23931 );
nor \U$32650 ( \33028 , \33026 , \33027 );
xnor \U$32651 ( \33029 , \33028 , \23791 );
and \U$32652 ( \33030 , \33024 , \33029 );
and \U$32653 ( \33031 , \33020 , \33029 );
or \U$32654 ( \33032 , \33025 , \33030 , \33031 );
and \U$32655 ( \33033 , \33016 , \33032 );
and \U$32656 ( \33034 , \23714 , \25692 );
and \U$32657 ( \33035 , \23570 , \25690 );
nor \U$32658 ( \33036 , \33034 , \33035 );
xnor \U$32659 ( \33037 , \33036 , \25549 );
and \U$32660 ( \33038 , \24003 , \25369 );
and \U$32661 ( \33039 , \23978 , \25367 );
nor \U$32662 ( \33040 , \33038 , \33039 );
xnor \U$32663 ( \33041 , \33040 , \25123 );
and \U$32664 ( \33042 , \33037 , \33041 );
and \U$32665 ( \33043 , \24344 , \24974 );
and \U$32666 ( \33044 , \24177 , \24972 );
nor \U$32667 ( \33045 , \33043 , \33044 );
xnor \U$32668 ( \33046 , \33045 , \24787 );
and \U$32669 ( \33047 , \33041 , \33046 );
and \U$32670 ( \33048 , \33037 , \33046 );
or \U$32671 ( \33049 , \33042 , \33047 , \33048 );
and \U$32672 ( \33050 , \33032 , \33049 );
and \U$32673 ( \33051 , \33016 , \33049 );
or \U$32674 ( \33052 , \33033 , \33050 , \33051 );
and \U$32675 ( \33053 , \32999 , \33052 );
and \U$32676 ( \33054 , \32947 , \33052 );
or \U$32677 ( \33055 , \33000 , \33053 , \33054 );
xor \U$32678 ( \33056 , \32746 , \32750 );
xor \U$32679 ( \33057 , \33056 , \32755 );
xor \U$32680 ( \33058 , \32762 , \32766 );
xor \U$32681 ( \33059 , \33058 , \32771 );
and \U$32682 ( \33060 , \33057 , \33059 );
xor \U$32683 ( \33061 , \32779 , \32783 );
xor \U$32684 ( \33062 , \33061 , \32788 );
and \U$32685 ( \33063 , \33059 , \33062 );
and \U$32686 ( \33064 , \33057 , \33062 );
or \U$32687 ( \33065 , \33060 , \33063 , \33064 );
and \U$32688 ( \33066 , \30318 , \21916 );
and \U$32689 ( \33067 , \30034 , \21914 );
nor \U$32690 ( \33068 , \33066 , \33067 );
xnor \U$32691 ( \33069 , \33068 , \21867 );
and \U$32692 ( \33070 , \30895 , \21815 );
and \U$32693 ( \33071 , \30887 , \21813 );
nor \U$32694 ( \33072 , \33070 , \33071 );
xnor \U$32695 ( \33073 , \33072 , \21774 );
and \U$32696 ( \33074 , \33069 , \33073 );
and \U$32697 ( \33075 , \31503 , \21745 );
and \U$32698 ( \33076 , \31498 , \21743 );
nor \U$32699 ( \33077 , \33075 , \33076 );
xnor \U$32700 ( \33078 , \33077 , \21715 );
and \U$32701 ( \33079 , \33073 , \33078 );
and \U$32702 ( \33080 , \33069 , \33078 );
or \U$32703 ( \33081 , \33074 , \33079 , \33080 );
xor \U$32704 ( \33082 , \32581 , \32585 );
xor \U$32705 ( \33083 , \33082 , \32588 );
and \U$32706 ( \33084 , \33081 , \33083 );
xor \U$32707 ( \33085 , \32595 , \32599 );
xor \U$32708 ( \33086 , \33085 , \32604 );
and \U$32709 ( \33087 , \33083 , \33086 );
and \U$32710 ( \33088 , \33081 , \33086 );
or \U$32711 ( \33089 , \33084 , \33087 , \33088 );
and \U$32712 ( \33090 , \33065 , \33089 );
xor \U$32713 ( \33091 , \32645 , \32649 );
xor \U$32714 ( \33092 , \33091 , \32654 );
xor \U$32715 ( \33093 , \32661 , \32665 );
xor \U$32716 ( \33094 , \33093 , \32670 );
and \U$32717 ( \33095 , \33092 , \33094 );
xor \U$32718 ( \33096 , \32678 , \32682 );
xor \U$32719 ( \33097 , \33096 , \32687 );
and \U$32720 ( \33098 , \33094 , \33097 );
and \U$32721 ( \33099 , \33092 , \33097 );
or \U$32722 ( \33100 , \33095 , \33098 , \33099 );
and \U$32723 ( \33101 , \33089 , \33100 );
and \U$32724 ( \33102 , \33065 , \33100 );
or \U$32725 ( \33103 , \33090 , \33101 , \33102 );
and \U$32726 ( \33104 , \33055 , \33103 );
xor \U$32727 ( \33105 , \32697 , \32701 );
xor \U$32728 ( \33106 , \33105 , \32706 );
xor \U$32729 ( \33107 , \32713 , \32717 );
xor \U$32730 ( \33108 , \33107 , \21665 );
and \U$32731 ( \33109 , \33106 , \33108 );
xor \U$32732 ( \33110 , \32726 , \32730 );
xor \U$32733 ( \33111 , \33110 , \32735 );
and \U$32734 ( \33112 , \33108 , \33111 );
and \U$32735 ( \33113 , \33106 , \33111 );
or \U$32736 ( \33114 , \33109 , \33112 , \33113 );
xor \U$32737 ( \33115 , \32800 , \32802 );
xor \U$32738 ( \33116 , \33115 , \32805 );
and \U$32739 ( \33117 , \33114 , \33116 );
xor \U$32740 ( \33118 , \32810 , \32812 );
and \U$32741 ( \33119 , \33116 , \33118 );
and \U$32742 ( \33120 , \33114 , \33118 );
or \U$32743 ( \33121 , \33117 , \33119 , \33120 );
and \U$32744 ( \33122 , \33103 , \33121 );
and \U$32745 ( \33123 , \33055 , \33121 );
or \U$32746 ( \33124 , \33104 , \33122 , \33123 );
xor \U$32747 ( \33125 , \32657 , \32673 );
xor \U$32748 ( \33126 , \33125 , \32690 );
xor \U$32749 ( \33127 , \32709 , \32721 );
xor \U$32750 ( \33128 , \33127 , \32738 );
and \U$32751 ( \33129 , \33126 , \33128 );
xor \U$32752 ( \33130 , \32758 , \32774 );
xor \U$32753 ( \33131 , \33130 , \32791 );
and \U$32754 ( \33132 , \33128 , \33131 );
and \U$32755 ( \33133 , \33126 , \33131 );
or \U$32756 ( \33134 , \33129 , \33132 , \33133 );
xor \U$32757 ( \33135 , \32591 , \32607 );
xor \U$32758 ( \33136 , \33135 , \32612 );
xor \U$32759 ( \33137 , \32619 , \32621 );
xor \U$32760 ( \33138 , \33137 , \32624 );
and \U$32761 ( \33139 , \33136 , \33138 );
xor \U$32762 ( \33140 , \32630 , \32632 );
xor \U$32763 ( \33141 , \33140 , \32635 );
and \U$32764 ( \33142 , \33138 , \33141 );
and \U$32765 ( \33143 , \33136 , \33141 );
or \U$32766 ( \33144 , \33139 , \33142 , \33143 );
and \U$32767 ( \33145 , \33134 , \33144 );
xor \U$32768 ( \33146 , \32383 , \32399 );
xor \U$32769 ( \33147 , \33146 , \32416 );
and \U$32770 ( \33148 , \33144 , \33147 );
and \U$32771 ( \33149 , \33134 , \33147 );
or \U$32772 ( \33150 , \33145 , \33148 , \33149 );
and \U$32773 ( \33151 , \33124 , \33150 );
xor \U$32774 ( \33152 , \32823 , \32825 );
xor \U$32775 ( \33153 , \33152 , \32828 );
xor \U$32776 ( \33154 , \32833 , \32835 );
xor \U$32777 ( \33155 , \33154 , \32838 );
and \U$32778 ( \33156 , \33153 , \33155 );
xor \U$32779 ( \33157 , \32808 , \32813 );
xor \U$32780 ( \33158 , \33157 , \32815 );
and \U$32781 ( \33159 , \33155 , \33158 );
and \U$32782 ( \33160 , \33153 , \33158 );
or \U$32783 ( \33161 , \33156 , \33159 , \33160 );
and \U$32784 ( \33162 , \33150 , \33161 );
and \U$32785 ( \33163 , \33124 , \33161 );
or \U$32786 ( \33164 , \33151 , \33162 , \33163 );
xor \U$32787 ( \33165 , \32367 , \32419 );
xor \U$32788 ( \33166 , \33165 , \32472 );
xor \U$32789 ( \33167 , \32831 , \32841 );
xor \U$32790 ( \33168 , \33167 , \32844 );
and \U$32791 ( \33169 , \33166 , \33168 );
xor \U$32792 ( \33170 , \32850 , \32852 );
xor \U$32793 ( \33171 , \33170 , \32855 );
and \U$32794 ( \33172 , \33168 , \33171 );
and \U$32795 ( \33173 , \33166 , \33171 );
or \U$32796 ( \33174 , \33169 , \33172 , \33173 );
and \U$32797 ( \33175 , \33164 , \33174 );
xor \U$32798 ( \33176 , \32506 , \32515 );
xor \U$32799 ( \33177 , \33176 , \32518 );
and \U$32800 ( \33178 , \33174 , \33177 );
and \U$32801 ( \33179 , \33164 , \33177 );
or \U$32802 ( \33180 , \33175 , \33178 , \33179 );
xor \U$32803 ( \33181 , \32315 , \32475 );
xor \U$32804 ( \33182 , \33181 , \32493 );
xor \U$32805 ( \33183 , \32821 , \32847 );
xor \U$32806 ( \33184 , \33183 , \32858 );
and \U$32807 ( \33185 , \33182 , \33184 );
xor \U$32808 ( \33186 , \32863 , \32865 );
xor \U$32809 ( \33187 , \33186 , \32868 );
and \U$32810 ( \33188 , \33184 , \33187 );
and \U$32811 ( \33189 , \33182 , \33187 );
or \U$32812 ( \33190 , \33185 , \33188 , \33189 );
and \U$32813 ( \33191 , \33180 , \33190 );
xor \U$32814 ( \33192 , \32537 , \32539 );
xor \U$32815 ( \33193 , \33192 , \32542 );
and \U$32816 ( \33194 , \33190 , \33193 );
and \U$32817 ( \33195 , \33180 , \33193 );
or \U$32818 ( \33196 , \33191 , \33194 , \33195 );
xor \U$32819 ( \33197 , \32496 , \32521 );
xor \U$32820 ( \33198 , \33197 , \32532 );
xor \U$32821 ( \33199 , \32861 , \32871 );
xor \U$32822 ( \33200 , \33199 , \32874 );
and \U$32823 ( \33201 , \33198 , \33200 );
and \U$32824 ( \33202 , \33196 , \33201 );
xor \U$32825 ( \33203 , \32877 , \32879 );
xor \U$32826 ( \33204 , \33203 , \32881 );
and \U$32827 ( \33205 , \33201 , \33204 );
and \U$32828 ( \33206 , \33196 , \33204 );
or \U$32829 ( \33207 , \33202 , \33205 , \33206 );
and \U$32830 ( \33208 , \32895 , \33207 );
xor \U$32831 ( \33209 , \32895 , \33207 );
xor \U$32832 ( \33210 , \33196 , \33201 );
xor \U$32833 ( \33211 , \33210 , \33204 );
and \U$32834 ( \33212 , \28342 , \22497 );
and \U$32835 ( \33213 , \28039 , \22495 );
nor \U$32836 ( \33214 , \33212 , \33213 );
xnor \U$32837 ( \33215 , \33214 , \22419 );
and \U$32838 ( \33216 , \29040 , \22333 );
and \U$32839 ( \33217 , \28514 , \22331 );
nor \U$32840 ( \33218 , \33216 , \33217 );
xnor \U$32841 ( \33219 , \33218 , \22239 );
and \U$32842 ( \33220 , \33215 , \33219 );
and \U$32843 ( \33221 , \29710 , \22163 );
and \U$32844 ( \33222 , \29464 , \22161 );
nor \U$32845 ( \33223 , \33221 , \33222 );
xnor \U$32846 ( \33224 , \33223 , \22091 );
and \U$32847 ( \33225 , \33219 , \33224 );
and \U$32848 ( \33226 , \33215 , \33224 );
or \U$32849 ( \33227 , \33220 , \33225 , \33226 );
and \U$32850 ( \33228 , \25609 , \23933 );
and \U$32851 ( \33229 , \25353 , \23931 );
nor \U$32852 ( \33230 , \33228 , \33229 );
xnor \U$32853 ( \33231 , \33230 , \23791 );
and \U$32854 ( \33232 , \26108 , \23637 );
and \U$32855 ( \33233 , \25806 , \23635 );
nor \U$32856 ( \33234 , \33232 , \33233 );
xnor \U$32857 ( \33235 , \33234 , \23500 );
and \U$32858 ( \33236 , \33231 , \33235 );
and \U$32859 ( \33237 , \26585 , \23431 );
and \U$32860 ( \33238 , \26116 , \23429 );
nor \U$32861 ( \33239 , \33237 , \33238 );
xnor \U$32862 ( \33240 , \33239 , \23279 );
and \U$32863 ( \33241 , \33235 , \33240 );
and \U$32864 ( \33242 , \33231 , \33240 );
or \U$32865 ( \33243 , \33236 , \33241 , \33242 );
and \U$32866 ( \33244 , \33227 , \33243 );
and \U$32867 ( \33245 , \26854 , \23163 );
and \U$32868 ( \33246 , \26590 , \23161 );
nor \U$32869 ( \33247 , \33245 , \33246 );
xnor \U$32870 ( \33248 , \33247 , \23007 );
and \U$32871 ( \33249 , \27485 , \22891 );
and \U$32872 ( \33250 , \27113 , \22889 );
nor \U$32873 ( \33251 , \33249 , \33250 );
xnor \U$32874 ( \33252 , \33251 , \22778 );
and \U$32875 ( \33253 , \33248 , \33252 );
and \U$32876 ( \33254 , \27837 , \22697 );
and \U$32877 ( \33255 , \27494 , \22695 );
nor \U$32878 ( \33256 , \33254 , \33255 );
xnor \U$32879 ( \33257 , \33256 , \22561 );
and \U$32880 ( \33258 , \33252 , \33257 );
and \U$32881 ( \33259 , \33248 , \33257 );
or \U$32882 ( \33260 , \33253 , \33258 , \33259 );
and \U$32883 ( \33261 , \33243 , \33260 );
and \U$32884 ( \33262 , \33227 , \33260 );
or \U$32885 ( \33263 , \33244 , \33261 , \33262 );
and \U$32886 ( \33264 , \22262 , \29104 );
and \U$32887 ( \33265 , \22200 , \29102 );
nor \U$32888 ( \33266 , \33264 , \33265 );
xnor \U$32889 ( \33267 , \33266 , \28855 );
and \U$32890 ( \33268 , \22523 , \28575 );
and \U$32891 ( \33269 , \22325 , \28573 );
nor \U$32892 ( \33270 , \33268 , \33269 );
xnor \U$32893 ( \33271 , \33270 , \28315 );
and \U$32894 ( \33272 , \33267 , \33271 );
and \U$32895 ( \33273 , \22716 , \28081 );
and \U$32896 ( \33274 , \22611 , \28079 );
nor \U$32897 ( \33275 , \33273 , \33274 );
xnor \U$32898 ( \33276 , \33275 , \27766 );
and \U$32899 ( \33277 , \33271 , \33276 );
and \U$32900 ( \33278 , \33267 , \33276 );
or \U$32901 ( \33279 , \33272 , \33277 , \33278 );
and \U$32902 ( \33280 , \21890 , \30770 );
and \U$32903 ( \33281 , \21836 , \30768 );
nor \U$32904 ( \33282 , \33280 , \33281 );
xnor \U$32905 ( \33283 , \33282 , \30460 );
and \U$32906 ( \33284 , \22018 , \30233 );
and \U$32907 ( \33285 , \21941 , \30231 );
nor \U$32908 ( \33286 , \33284 , \33285 );
xnor \U$32909 ( \33287 , \33286 , \29862 );
and \U$32910 ( \33288 , \33283 , \33287 );
and \U$32911 ( \33289 , \22126 , \29671 );
and \U$32912 ( \33290 , \22046 , \29669 );
nor \U$32913 ( \33291 , \33289 , \33290 );
xnor \U$32914 ( \33292 , \33291 , \29353 );
and \U$32915 ( \33293 , \33287 , \33292 );
and \U$32916 ( \33294 , \33283 , \33292 );
or \U$32917 ( \33295 , \33288 , \33293 , \33294 );
and \U$32918 ( \33296 , \33279 , \33295 );
and \U$32919 ( \33297 , \21754 , \32151 );
and \U$32920 ( \33298 , \21706 , \32148 );
nor \U$32921 ( \33299 , \33297 , \33298 );
xnor \U$32922 ( \33300 , \33299 , \31096 );
and \U$32923 ( \33301 , \21831 , \31338 );
and \U$32924 ( \33302 , \21762 , \31336 );
nor \U$32925 ( \33303 , \33301 , \33302 );
xnor \U$32926 ( \33304 , \33303 , \31099 );
and \U$32927 ( \33305 , \33300 , \33304 );
and \U$32928 ( \33306 , \33304 , \21678 );
and \U$32929 ( \33307 , \33300 , \21678 );
or \U$32930 ( \33308 , \33305 , \33306 , \33307 );
and \U$32931 ( \33309 , \33295 , \33308 );
and \U$32932 ( \33310 , \33279 , \33308 );
or \U$32933 ( \33311 , \33296 , \33309 , \33310 );
and \U$32934 ( \33312 , \33263 , \33311 );
and \U$32935 ( \33313 , \22837 , \27572 );
and \U$32936 ( \33314 , \22721 , \27570 );
nor \U$32937 ( \33315 , \33313 , \33314 );
xnor \U$32938 ( \33316 , \33315 , \27232 );
and \U$32939 ( \33317 , \23128 , \26983 );
and \U$32940 ( \33318 , \22952 , \26981 );
nor \U$32941 ( \33319 , \33317 , \33318 );
xnor \U$32942 ( \33320 , \33319 , \26742 );
and \U$32943 ( \33321 , \33316 , \33320 );
and \U$32944 ( \33322 , \23379 , \26517 );
and \U$32945 ( \33323 , \23136 , \26515 );
nor \U$32946 ( \33324 , \33322 , \33323 );
xnor \U$32947 ( \33325 , \33324 , \26329 );
and \U$32948 ( \33326 , \33320 , \33325 );
and \U$32949 ( \33327 , \33316 , \33325 );
or \U$32950 ( \33328 , \33321 , \33326 , \33327 );
and \U$32951 ( \33329 , \23570 , \26143 );
and \U$32952 ( \33330 , \23384 , \26141 );
nor \U$32953 ( \33331 , \33329 , \33330 );
xnor \U$32954 ( \33332 , \33331 , \25911 );
and \U$32955 ( \33333 , \23978 , \25692 );
and \U$32956 ( \33334 , \23714 , \25690 );
nor \U$32957 ( \33335 , \33333 , \33334 );
xnor \U$32958 ( \33336 , \33335 , \25549 );
and \U$32959 ( \33337 , \33332 , \33336 );
and \U$32960 ( \33338 , \24177 , \25369 );
and \U$32961 ( \33339 , \24003 , \25367 );
nor \U$32962 ( \33340 , \33338 , \33339 );
xnor \U$32963 ( \33341 , \33340 , \25123 );
and \U$32964 ( \33342 , \33336 , \33341 );
and \U$32965 ( \33343 , \33332 , \33341 );
or \U$32966 ( \33344 , \33337 , \33342 , \33343 );
and \U$32967 ( \33345 , \33328 , \33344 );
and \U$32968 ( \33346 , \24482 , \24974 );
and \U$32969 ( \33347 , \24344 , \24972 );
nor \U$32970 ( \33348 , \33346 , \33347 );
xnor \U$32971 ( \33349 , \33348 , \24787 );
and \U$32972 ( \33350 , \25018 , \24661 );
and \U$32973 ( \33351 , \24601 , \24659 );
nor \U$32974 ( \33352 , \33350 , \33351 );
xnor \U$32975 ( \33353 , \33352 , \24456 );
and \U$32976 ( \33354 , \33349 , \33353 );
and \U$32977 ( \33355 , \25348 , \24255 );
and \U$32978 ( \33356 , \25226 , \24253 );
nor \U$32979 ( \33357 , \33355 , \33356 );
xnor \U$32980 ( \33358 , \33357 , \24106 );
and \U$32981 ( \33359 , \33353 , \33358 );
and \U$32982 ( \33360 , \33349 , \33358 );
or \U$32983 ( \33361 , \33354 , \33359 , \33360 );
and \U$32984 ( \33362 , \33344 , \33361 );
and \U$32985 ( \33363 , \33328 , \33361 );
or \U$32986 ( \33364 , \33345 , \33362 , \33363 );
and \U$32987 ( \33365 , \33311 , \33364 );
and \U$32988 ( \33366 , \33263 , \33364 );
or \U$32989 ( \33367 , \33312 , \33365 , \33366 );
and \U$32990 ( \33368 , \30034 , \22029 );
and \U$32991 ( \33369 , \29715 , \22027 );
nor \U$32992 ( \33370 , \33368 , \33369 );
xnor \U$32993 ( \33371 , \33370 , \21986 );
and \U$32994 ( \33372 , \30887 , \21916 );
and \U$32995 ( \33373 , \30318 , \21914 );
nor \U$32996 ( \33374 , \33372 , \33373 );
xnor \U$32997 ( \33375 , \33374 , \21867 );
and \U$32998 ( \33376 , \33371 , \33375 );
and \U$32999 ( \33377 , \31498 , \21815 );
and \U$33000 ( \33378 , \30895 , \21813 );
nor \U$33001 ( \33379 , \33377 , \33378 );
xnor \U$33002 ( \33380 , \33379 , \21774 );
and \U$33003 ( \33381 , \33375 , \33380 );
and \U$33004 ( \33382 , \33371 , \33380 );
or \U$33005 ( \33383 , \33376 , \33381 , \33382 );
and \U$33006 ( \33384 , \31684 , \21745 );
and \U$33007 ( \33385 , \31503 , \21743 );
nor \U$33008 ( \33386 , \33384 , \33385 );
xnor \U$33009 ( \33387 , \33386 , \21715 );
nand \U$33010 ( \33388 , \32304 , \21695 );
xnor \U$33011 ( \33389 , \33388 , \21678 );
and \U$33012 ( \33390 , \33387 , \33389 );
and \U$33013 ( \33391 , \33383 , \33390 );
and \U$33014 ( \33392 , \32304 , \21697 );
and \U$33015 ( \33393 , \31684 , \21695 );
nor \U$33016 ( \33394 , \33392 , \33393 );
xnor \U$33017 ( \33395 , \33394 , \21678 );
and \U$33018 ( \33396 , \33390 , \33395 );
and \U$33019 ( \33397 , \33383 , \33395 );
or \U$33020 ( \33398 , \33391 , \33396 , \33397 );
xor \U$33021 ( \33399 , \32984 , \32988 );
xor \U$33022 ( \33400 , \33399 , \32993 );
xor \U$33023 ( \33401 , \33020 , \33024 );
xor \U$33024 ( \33402 , \33401 , \33029 );
and \U$33025 ( \33403 , \33400 , \33402 );
xor \U$33026 ( \33404 , \33037 , \33041 );
xor \U$33027 ( \33405 , \33404 , \33046 );
and \U$33028 ( \33406 , \33402 , \33405 );
and \U$33029 ( \33407 , \33400 , \33405 );
or \U$33030 ( \33408 , \33403 , \33406 , \33407 );
and \U$33031 ( \33409 , \33398 , \33408 );
xor \U$33032 ( \33410 , \32951 , \32955 );
xor \U$33033 ( \33411 , \33410 , \32960 );
xor \U$33034 ( \33412 , \32967 , \32971 );
xor \U$33035 ( \33413 , \33412 , \32976 );
and \U$33036 ( \33414 , \33411 , \33413 );
xor \U$33037 ( \33415 , \33069 , \33073 );
xor \U$33038 ( \33416 , \33415 , \33078 );
and \U$33039 ( \33417 , \33413 , \33416 );
and \U$33040 ( \33418 , \33411 , \33416 );
or \U$33041 ( \33419 , \33414 , \33417 , \33418 );
and \U$33042 ( \33420 , \33408 , \33419 );
and \U$33043 ( \33421 , \33398 , \33419 );
or \U$33044 ( \33422 , \33409 , \33420 , \33421 );
and \U$33045 ( \33423 , \33367 , \33422 );
xor \U$33046 ( \33424 , \32899 , \32903 );
xor \U$33047 ( \33425 , \33424 , \32908 );
xor \U$33048 ( \33426 , \33004 , \33008 );
xor \U$33049 ( \33427 , \33426 , \33013 );
and \U$33050 ( \33428 , \33425 , \33427 );
xor \U$33051 ( \33429 , \32932 , \32936 );
xor \U$33052 ( \33430 , \33429 , \32941 );
and \U$33053 ( \33431 , \33427 , \33430 );
and \U$33054 ( \33432 , \33425 , \33430 );
or \U$33055 ( \33433 , \33428 , \33431 , \33432 );
xor \U$33056 ( \33434 , \33106 , \33108 );
xor \U$33057 ( \33435 , \33434 , \33111 );
and \U$33058 ( \33436 , \33433 , \33435 );
xor \U$33059 ( \33437 , \33057 , \33059 );
xor \U$33060 ( \33438 , \33437 , \33062 );
and \U$33061 ( \33439 , \33435 , \33438 );
and \U$33062 ( \33440 , \33433 , \33438 );
or \U$33063 ( \33441 , \33436 , \33439 , \33440 );
and \U$33064 ( \33442 , \33422 , \33441 );
and \U$33065 ( \33443 , \33367 , \33441 );
or \U$33066 ( \33444 , \33423 , \33442 , \33443 );
xor \U$33067 ( \33445 , \32963 , \32979 );
xor \U$33068 ( \33446 , \33445 , \32996 );
xor \U$33069 ( \33447 , \33081 , \33083 );
xor \U$33070 ( \33448 , \33447 , \33086 );
and \U$33071 ( \33449 , \33446 , \33448 );
xor \U$33072 ( \33450 , \33092 , \33094 );
xor \U$33073 ( \33451 , \33450 , \33097 );
and \U$33074 ( \33452 , \33448 , \33451 );
and \U$33075 ( \33453 , \33446 , \33451 );
or \U$33076 ( \33454 , \33449 , \33452 , \33453 );
xor \U$33077 ( \33455 , \33126 , \33128 );
xor \U$33078 ( \33456 , \33455 , \33131 );
and \U$33079 ( \33457 , \33454 , \33456 );
xor \U$33080 ( \33458 , \33136 , \33138 );
xor \U$33081 ( \33459 , \33458 , \33141 );
and \U$33082 ( \33460 , \33456 , \33459 );
and \U$33083 ( \33461 , \33454 , \33459 );
or \U$33084 ( \33462 , \33457 , \33460 , \33461 );
and \U$33085 ( \33463 , \33444 , \33462 );
xor \U$33086 ( \33464 , \32947 , \32999 );
xor \U$33087 ( \33465 , \33464 , \33052 );
xor \U$33088 ( \33466 , \33065 , \33089 );
xor \U$33089 ( \33467 , \33466 , \33100 );
and \U$33090 ( \33468 , \33465 , \33467 );
xor \U$33091 ( \33469 , \33114 , \33116 );
xor \U$33092 ( \33470 , \33469 , \33118 );
and \U$33093 ( \33471 , \33467 , \33470 );
and \U$33094 ( \33472 , \33465 , \33470 );
or \U$33095 ( \33473 , \33468 , \33471 , \33472 );
and \U$33096 ( \33474 , \33462 , \33473 );
and \U$33097 ( \33475 , \33444 , \33473 );
or \U$33098 ( \33476 , \33463 , \33474 , \33475 );
xor \U$33099 ( \33477 , \32615 , \32627 );
xor \U$33100 ( \33478 , \33477 , \32638 );
xor \U$33101 ( \33479 , \32693 , \32741 );
xor \U$33102 ( \33480 , \33479 , \32794 );
and \U$33103 ( \33481 , \33478 , \33480 );
xor \U$33104 ( \33482 , \33153 , \33155 );
xor \U$33105 ( \33483 , \33482 , \33158 );
and \U$33106 ( \33484 , \33480 , \33483 );
and \U$33107 ( \33485 , \33478 , \33483 );
or \U$33108 ( \33486 , \33481 , \33484 , \33485 );
and \U$33109 ( \33487 , \33476 , \33486 );
xor \U$33110 ( \33488 , \32641 , \32797 );
xor \U$33111 ( \33489 , \33488 , \32818 );
and \U$33112 ( \33490 , \33486 , \33489 );
and \U$33113 ( \33491 , \33476 , \33489 );
or \U$33114 ( \33492 , \33487 , \33490 , \33491 );
xor \U$33115 ( \33493 , \33164 , \33174 );
xor \U$33116 ( \33494 , \33493 , \33177 );
and \U$33117 ( \33495 , \33492 , \33494 );
xor \U$33118 ( \33496 , \33182 , \33184 );
xor \U$33119 ( \33497 , \33496 , \33187 );
and \U$33120 ( \33498 , \33494 , \33497 );
and \U$33121 ( \33499 , \33492 , \33497 );
or \U$33122 ( \33500 , \33495 , \33498 , \33499 );
xor \U$33123 ( \33501 , \33180 , \33190 );
xor \U$33124 ( \33502 , \33501 , \33193 );
and \U$33125 ( \33503 , \33500 , \33502 );
xor \U$33126 ( \33504 , \33198 , \33200 );
and \U$33127 ( \33505 , \33502 , \33504 );
and \U$33128 ( \33506 , \33500 , \33504 );
or \U$33129 ( \33507 , \33503 , \33505 , \33506 );
and \U$33130 ( \33508 , \33211 , \33507 );
xor \U$33131 ( \33509 , \33211 , \33507 );
xor \U$33132 ( \33510 , \33500 , \33502 );
xor \U$33133 ( \33511 , \33510 , \33504 );
xor \U$33134 ( \33512 , \33215 , \33219 );
xor \U$33135 ( \33513 , \33512 , \33224 );
xor \U$33136 ( \33514 , \33231 , \33235 );
xor \U$33137 ( \33515 , \33514 , \33240 );
and \U$33138 ( \33516 , \33513 , \33515 );
xor \U$33139 ( \33517 , \33248 , \33252 );
xor \U$33140 ( \33518 , \33517 , \33257 );
and \U$33141 ( \33519 , \33515 , \33518 );
and \U$33142 ( \33520 , \33513 , \33518 );
or \U$33143 ( \33521 , \33516 , \33519 , \33520 );
xor \U$33144 ( \33522 , \33316 , \33320 );
xor \U$33145 ( \33523 , \33522 , \33325 );
xor \U$33146 ( \33524 , \33332 , \33336 );
xor \U$33147 ( \33525 , \33524 , \33341 );
and \U$33148 ( \33526 , \33523 , \33525 );
xor \U$33149 ( \33527 , \33349 , \33353 );
xor \U$33150 ( \33528 , \33527 , \33358 );
and \U$33151 ( \33529 , \33525 , \33528 );
and \U$33152 ( \33530 , \33523 , \33528 );
or \U$33153 ( \33531 , \33526 , \33529 , \33530 );
and \U$33154 ( \33532 , \33521 , \33531 );
and \U$33155 ( \33533 , \30895 , \21916 );
and \U$33156 ( \33534 , \30887 , \21914 );
nor \U$33157 ( \33535 , \33533 , \33534 );
xnor \U$33158 ( \33536 , \33535 , \21867 );
and \U$33159 ( \33537 , \31503 , \21815 );
and \U$33160 ( \33538 , \31498 , \21813 );
nor \U$33161 ( \33539 , \33537 , \33538 );
xnor \U$33162 ( \33540 , \33539 , \21774 );
and \U$33163 ( \33541 , \33536 , \33540 );
and \U$33164 ( \33542 , \32304 , \21745 );
and \U$33165 ( \33543 , \31684 , \21743 );
nor \U$33166 ( \33544 , \33542 , \33543 );
xnor \U$33167 ( \33545 , \33544 , \21715 );
and \U$33168 ( \33546 , \33540 , \33545 );
and \U$33169 ( \33547 , \33536 , \33545 );
or \U$33170 ( \33548 , \33541 , \33546 , \33547 );
xor \U$33171 ( \33549 , \33371 , \33375 );
xor \U$33172 ( \33550 , \33549 , \33380 );
and \U$33173 ( \33551 , \33548 , \33550 );
xor \U$33174 ( \33552 , \33387 , \33389 );
and \U$33175 ( \33553 , \33550 , \33552 );
and \U$33176 ( \33554 , \33548 , \33552 );
or \U$33177 ( \33555 , \33551 , \33553 , \33554 );
and \U$33178 ( \33556 , \33531 , \33555 );
and \U$33179 ( \33557 , \33521 , \33555 );
or \U$33180 ( \33558 , \33532 , \33556 , \33557 );
and \U$33181 ( \33559 , \25226 , \24661 );
and \U$33182 ( \33560 , \25018 , \24659 );
nor \U$33183 ( \33561 , \33559 , \33560 );
xnor \U$33184 ( \33562 , \33561 , \24456 );
and \U$33185 ( \33563 , \25353 , \24255 );
and \U$33186 ( \33564 , \25348 , \24253 );
nor \U$33187 ( \33565 , \33563 , \33564 );
xnor \U$33188 ( \33566 , \33565 , \24106 );
and \U$33189 ( \33567 , \33562 , \33566 );
and \U$33190 ( \33568 , \25806 , \23933 );
and \U$33191 ( \33569 , \25609 , \23931 );
nor \U$33192 ( \33570 , \33568 , \33569 );
xnor \U$33193 ( \33571 , \33570 , \23791 );
and \U$33194 ( \33572 , \33566 , \33571 );
and \U$33195 ( \33573 , \33562 , \33571 );
or \U$33196 ( \33574 , \33567 , \33572 , \33573 );
and \U$33197 ( \33575 , \23136 , \26983 );
and \U$33198 ( \33576 , \23128 , \26981 );
nor \U$33199 ( \33577 , \33575 , \33576 );
xnor \U$33200 ( \33578 , \33577 , \26742 );
and \U$33201 ( \33579 , \23384 , \26517 );
and \U$33202 ( \33580 , \23379 , \26515 );
nor \U$33203 ( \33581 , \33579 , \33580 );
xnor \U$33204 ( \33582 , \33581 , \26329 );
and \U$33205 ( \33583 , \33578 , \33582 );
and \U$33206 ( \33584 , \23714 , \26143 );
and \U$33207 ( \33585 , \23570 , \26141 );
nor \U$33208 ( \33586 , \33584 , \33585 );
xnor \U$33209 ( \33587 , \33586 , \25911 );
and \U$33210 ( \33588 , \33582 , \33587 );
and \U$33211 ( \33589 , \33578 , \33587 );
or \U$33212 ( \33590 , \33583 , \33588 , \33589 );
and \U$33213 ( \33591 , \33574 , \33590 );
and \U$33214 ( \33592 , \24003 , \25692 );
and \U$33215 ( \33593 , \23978 , \25690 );
nor \U$33216 ( \33594 , \33592 , \33593 );
xnor \U$33217 ( \33595 , \33594 , \25549 );
and \U$33218 ( \33596 , \24344 , \25369 );
and \U$33219 ( \33597 , \24177 , \25367 );
nor \U$33220 ( \33598 , \33596 , \33597 );
xnor \U$33221 ( \33599 , \33598 , \25123 );
and \U$33222 ( \33600 , \33595 , \33599 );
and \U$33223 ( \33601 , \24601 , \24974 );
and \U$33224 ( \33602 , \24482 , \24972 );
nor \U$33225 ( \33603 , \33601 , \33602 );
xnor \U$33226 ( \33604 , \33603 , \24787 );
and \U$33227 ( \33605 , \33599 , \33604 );
and \U$33228 ( \33606 , \33595 , \33604 );
or \U$33229 ( \33607 , \33600 , \33605 , \33606 );
and \U$33230 ( \33608 , \33590 , \33607 );
and \U$33231 ( \33609 , \33574 , \33607 );
or \U$33232 ( \33610 , \33591 , \33608 , \33609 );
and \U$33233 ( \33611 , \22611 , \28575 );
and \U$33234 ( \33612 , \22523 , \28573 );
nor \U$33235 ( \33613 , \33611 , \33612 );
xnor \U$33236 ( \33614 , \33613 , \28315 );
and \U$33237 ( \33615 , \22721 , \28081 );
and \U$33238 ( \33616 , \22716 , \28079 );
nor \U$33239 ( \33617 , \33615 , \33616 );
xnor \U$33240 ( \33618 , \33617 , \27766 );
and \U$33241 ( \33619 , \33614 , \33618 );
and \U$33242 ( \33620 , \22952 , \27572 );
and \U$33243 ( \33621 , \22837 , \27570 );
nor \U$33244 ( \33622 , \33620 , \33621 );
xnor \U$33245 ( \33623 , \33622 , \27232 );
and \U$33246 ( \33624 , \33618 , \33623 );
and \U$33247 ( \33625 , \33614 , \33623 );
or \U$33248 ( \33626 , \33619 , \33624 , \33625 );
and \U$33249 ( \33627 , \21762 , \32151 );
and \U$33250 ( \33628 , \21754 , \32148 );
nor \U$33251 ( \33629 , \33627 , \33628 );
xnor \U$33252 ( \33630 , \33629 , \31096 );
and \U$33253 ( \33631 , \21836 , \31338 );
and \U$33254 ( \33632 , \21831 , \31336 );
nor \U$33255 ( \33633 , \33631 , \33632 );
xnor \U$33256 ( \33634 , \33633 , \31099 );
and \U$33257 ( \33635 , \33630 , \33634 );
and \U$33258 ( \33636 , \21941 , \30770 );
and \U$33259 ( \33637 , \21890 , \30768 );
nor \U$33260 ( \33638 , \33636 , \33637 );
xnor \U$33261 ( \33639 , \33638 , \30460 );
and \U$33262 ( \33640 , \33634 , \33639 );
and \U$33263 ( \33641 , \33630 , \33639 );
or \U$33264 ( \33642 , \33635 , \33640 , \33641 );
and \U$33265 ( \33643 , \33626 , \33642 );
and \U$33266 ( \33644 , \22046 , \30233 );
and \U$33267 ( \33645 , \22018 , \30231 );
nor \U$33268 ( \33646 , \33644 , \33645 );
xnor \U$33269 ( \33647 , \33646 , \29862 );
and \U$33270 ( \33648 , \22200 , \29671 );
and \U$33271 ( \33649 , \22126 , \29669 );
nor \U$33272 ( \33650 , \33648 , \33649 );
xnor \U$33273 ( \33651 , \33650 , \29353 );
and \U$33274 ( \33652 , \33647 , \33651 );
and \U$33275 ( \33653 , \22325 , \29104 );
and \U$33276 ( \33654 , \22262 , \29102 );
nor \U$33277 ( \33655 , \33653 , \33654 );
xnor \U$33278 ( \33656 , \33655 , \28855 );
and \U$33279 ( \33657 , \33651 , \33656 );
and \U$33280 ( \33658 , \33647 , \33656 );
or \U$33281 ( \33659 , \33652 , \33657 , \33658 );
and \U$33282 ( \33660 , \33642 , \33659 );
and \U$33283 ( \33661 , \33626 , \33659 );
or \U$33284 ( \33662 , \33643 , \33660 , \33661 );
and \U$33285 ( \33663 , \33610 , \33662 );
and \U$33286 ( \33664 , \26116 , \23637 );
and \U$33287 ( \33665 , \26108 , \23635 );
nor \U$33288 ( \33666 , \33664 , \33665 );
xnor \U$33289 ( \33667 , \33666 , \23500 );
and \U$33290 ( \33668 , \26590 , \23431 );
and \U$33291 ( \33669 , \26585 , \23429 );
nor \U$33292 ( \33670 , \33668 , \33669 );
xnor \U$33293 ( \33671 , \33670 , \23279 );
and \U$33294 ( \33672 , \33667 , \33671 );
and \U$33295 ( \33673 , \27113 , \23163 );
and \U$33296 ( \33674 , \26854 , \23161 );
nor \U$33297 ( \33675 , \33673 , \33674 );
xnor \U$33298 ( \33676 , \33675 , \23007 );
and \U$33299 ( \33677 , \33671 , \33676 );
and \U$33300 ( \33678 , \33667 , \33676 );
or \U$33301 ( \33679 , \33672 , \33677 , \33678 );
and \U$33302 ( \33680 , \29464 , \22333 );
and \U$33303 ( \33681 , \29040 , \22331 );
nor \U$33304 ( \33682 , \33680 , \33681 );
xnor \U$33305 ( \33683 , \33682 , \22239 );
and \U$33306 ( \33684 , \29715 , \22163 );
and \U$33307 ( \33685 , \29710 , \22161 );
nor \U$33308 ( \33686 , \33684 , \33685 );
xnor \U$33309 ( \33687 , \33686 , \22091 );
and \U$33310 ( \33688 , \33683 , \33687 );
and \U$33311 ( \33689 , \30318 , \22029 );
and \U$33312 ( \33690 , \30034 , \22027 );
nor \U$33313 ( \33691 , \33689 , \33690 );
xnor \U$33314 ( \33692 , \33691 , \21986 );
and \U$33315 ( \33693 , \33687 , \33692 );
and \U$33316 ( \33694 , \33683 , \33692 );
or \U$33317 ( \33695 , \33688 , \33693 , \33694 );
and \U$33318 ( \33696 , \33679 , \33695 );
and \U$33319 ( \33697 , \27494 , \22891 );
and \U$33320 ( \33698 , \27485 , \22889 );
nor \U$33321 ( \33699 , \33697 , \33698 );
xnor \U$33322 ( \33700 , \33699 , \22778 );
and \U$33323 ( \33701 , \28039 , \22697 );
and \U$33324 ( \33702 , \27837 , \22695 );
nor \U$33325 ( \33703 , \33701 , \33702 );
xnor \U$33326 ( \33704 , \33703 , \22561 );
and \U$33327 ( \33705 , \33700 , \33704 );
and \U$33328 ( \33706 , \28514 , \22497 );
and \U$33329 ( \33707 , \28342 , \22495 );
nor \U$33330 ( \33708 , \33706 , \33707 );
xnor \U$33331 ( \33709 , \33708 , \22419 );
and \U$33332 ( \33710 , \33704 , \33709 );
and \U$33333 ( \33711 , \33700 , \33709 );
or \U$33334 ( \33712 , \33705 , \33710 , \33711 );
and \U$33335 ( \33713 , \33695 , \33712 );
and \U$33336 ( \33714 , \33679 , \33712 );
or \U$33337 ( \33715 , \33696 , \33713 , \33714 );
and \U$33338 ( \33716 , \33662 , \33715 );
and \U$33339 ( \33717 , \33610 , \33715 );
or \U$33340 ( \33718 , \33663 , \33716 , \33717 );
and \U$33341 ( \33719 , \33558 , \33718 );
xor \U$33342 ( \33720 , \33267 , \33271 );
xor \U$33343 ( \33721 , \33720 , \33276 );
xor \U$33344 ( \33722 , \33283 , \33287 );
xor \U$33345 ( \33723 , \33722 , \33292 );
and \U$33346 ( \33724 , \33721 , \33723 );
xor \U$33347 ( \33725 , \33300 , \33304 );
xor \U$33348 ( \33726 , \33725 , \21678 );
and \U$33349 ( \33727 , \33723 , \33726 );
and \U$33350 ( \33728 , \33721 , \33726 );
or \U$33351 ( \33729 , \33724 , \33727 , \33728 );
xor \U$33352 ( \33730 , \32915 , \32919 );
xor \U$33353 ( \33731 , \33730 , \32924 );
and \U$33354 ( \33732 , \33729 , \33731 );
xor \U$33355 ( \33733 , \33425 , \33427 );
xor \U$33356 ( \33734 , \33733 , \33430 );
and \U$33357 ( \33735 , \33731 , \33734 );
and \U$33358 ( \33736 , \33729 , \33734 );
or \U$33359 ( \33737 , \33732 , \33735 , \33736 );
and \U$33360 ( \33738 , \33718 , \33737 );
and \U$33361 ( \33739 , \33558 , \33737 );
or \U$33362 ( \33740 , \33719 , \33738 , \33739 );
xor \U$33363 ( \33741 , \33227 , \33243 );
xor \U$33364 ( \33742 , \33741 , \33260 );
xor \U$33365 ( \33743 , \33279 , \33295 );
xor \U$33366 ( \33744 , \33743 , \33308 );
and \U$33367 ( \33745 , \33742 , \33744 );
xor \U$33368 ( \33746 , \33328 , \33344 );
xor \U$33369 ( \33747 , \33746 , \33361 );
and \U$33370 ( \33748 , \33744 , \33747 );
and \U$33371 ( \33749 , \33742 , \33747 );
or \U$33372 ( \33750 , \33745 , \33748 , \33749 );
xor \U$33373 ( \33751 , \33383 , \33390 );
xor \U$33374 ( \33752 , \33751 , \33395 );
xor \U$33375 ( \33753 , \33400 , \33402 );
xor \U$33376 ( \33754 , \33753 , \33405 );
and \U$33377 ( \33755 , \33752 , \33754 );
xor \U$33378 ( \33756 , \33411 , \33413 );
xor \U$33379 ( \33757 , \33756 , \33416 );
and \U$33380 ( \33758 , \33754 , \33757 );
and \U$33381 ( \33759 , \33752 , \33757 );
or \U$33382 ( \33760 , \33755 , \33758 , \33759 );
and \U$33383 ( \33761 , \33750 , \33760 );
xor \U$33384 ( \33762 , \33016 , \33032 );
xor \U$33385 ( \33763 , \33762 , \33049 );
and \U$33386 ( \33764 , \33760 , \33763 );
and \U$33387 ( \33765 , \33750 , \33763 );
or \U$33388 ( \33766 , \33761 , \33764 , \33765 );
and \U$33389 ( \33767 , \33740 , \33766 );
xor \U$33390 ( \33768 , \32911 , \32927 );
xor \U$33391 ( \33769 , \33768 , \32944 );
xor \U$33392 ( \33770 , \33446 , \33448 );
xor \U$33393 ( \33771 , \33770 , \33451 );
and \U$33394 ( \33772 , \33769 , \33771 );
xor \U$33395 ( \33773 , \33433 , \33435 );
xor \U$33396 ( \33774 , \33773 , \33438 );
and \U$33397 ( \33775 , \33771 , \33774 );
and \U$33398 ( \33776 , \33769 , \33774 );
or \U$33399 ( \33777 , \33772 , \33775 , \33776 );
and \U$33400 ( \33778 , \33766 , \33777 );
and \U$33401 ( \33779 , \33740 , \33777 );
or \U$33402 ( \33780 , \33767 , \33778 , \33779 );
xor \U$33403 ( \33781 , \33367 , \33422 );
xor \U$33404 ( \33782 , \33781 , \33441 );
xor \U$33405 ( \33783 , \33454 , \33456 );
xor \U$33406 ( \33784 , \33783 , \33459 );
and \U$33407 ( \33785 , \33782 , \33784 );
xor \U$33408 ( \33786 , \33465 , \33467 );
xor \U$33409 ( \33787 , \33786 , \33470 );
and \U$33410 ( \33788 , \33784 , \33787 );
and \U$33411 ( \33789 , \33782 , \33787 );
or \U$33412 ( \33790 , \33785 , \33788 , \33789 );
and \U$33413 ( \33791 , \33780 , \33790 );
xor \U$33414 ( \33792 , \33134 , \33144 );
xor \U$33415 ( \33793 , \33792 , \33147 );
and \U$33416 ( \33794 , \33790 , \33793 );
and \U$33417 ( \33795 , \33780 , \33793 );
or \U$33418 ( \33796 , \33791 , \33794 , \33795 );
xor \U$33419 ( \33797 , \33055 , \33103 );
xor \U$33420 ( \33798 , \33797 , \33121 );
xor \U$33421 ( \33799 , \33444 , \33462 );
xor \U$33422 ( \33800 , \33799 , \33473 );
and \U$33423 ( \33801 , \33798 , \33800 );
xor \U$33424 ( \33802 , \33478 , \33480 );
xor \U$33425 ( \33803 , \33802 , \33483 );
and \U$33426 ( \33804 , \33800 , \33803 );
and \U$33427 ( \33805 , \33798 , \33803 );
or \U$33428 ( \33806 , \33801 , \33804 , \33805 );
and \U$33429 ( \33807 , \33796 , \33806 );
xor \U$33430 ( \33808 , \33166 , \33168 );
xor \U$33431 ( \33809 , \33808 , \33171 );
and \U$33432 ( \33810 , \33806 , \33809 );
and \U$33433 ( \33811 , \33796 , \33809 );
or \U$33434 ( \33812 , \33807 , \33810 , \33811 );
xor \U$33435 ( \33813 , \33124 , \33150 );
xor \U$33436 ( \33814 , \33813 , \33161 );
xor \U$33437 ( \33815 , \33476 , \33486 );
xor \U$33438 ( \33816 , \33815 , \33489 );
and \U$33439 ( \33817 , \33814 , \33816 );
and \U$33440 ( \33818 , \33812 , \33817 );
xor \U$33441 ( \33819 , \33492 , \33494 );
xor \U$33442 ( \33820 , \33819 , \33497 );
and \U$33443 ( \33821 , \33817 , \33820 );
and \U$33444 ( \33822 , \33812 , \33820 );
or \U$33445 ( \33823 , \33818 , \33821 , \33822 );
and \U$33446 ( \33824 , \33511 , \33823 );
xor \U$33447 ( \33825 , \33511 , \33823 );
xor \U$33448 ( \33826 , \33812 , \33817 );
xor \U$33449 ( \33827 , \33826 , \33820 );
xor \U$33450 ( \33828 , \33562 , \33566 );
xor \U$33451 ( \33829 , \33828 , \33571 );
xor \U$33452 ( \33830 , \33667 , \33671 );
xor \U$33453 ( \33831 , \33830 , \33676 );
and \U$33454 ( \33832 , \33829 , \33831 );
xor \U$33455 ( \33833 , \33700 , \33704 );
xor \U$33456 ( \33834 , \33833 , \33709 );
and \U$33457 ( \33835 , \33831 , \33834 );
and \U$33458 ( \33836 , \33829 , \33834 );
or \U$33459 ( \33837 , \33832 , \33835 , \33836 );
and \U$33460 ( \33838 , \30887 , \22029 );
and \U$33461 ( \33839 , \30318 , \22027 );
nor \U$33462 ( \33840 , \33838 , \33839 );
xnor \U$33463 ( \33841 , \33840 , \21986 );
and \U$33464 ( \33842 , \31498 , \21916 );
and \U$33465 ( \33843 , \30895 , \21914 );
nor \U$33466 ( \33844 , \33842 , \33843 );
xnor \U$33467 ( \33845 , \33844 , \21867 );
and \U$33468 ( \33846 , \33841 , \33845 );
and \U$33469 ( \33847 , \31684 , \21815 );
and \U$33470 ( \33848 , \31503 , \21813 );
nor \U$33471 ( \33849 , \33847 , \33848 );
xnor \U$33472 ( \33850 , \33849 , \21774 );
and \U$33473 ( \33851 , \33845 , \33850 );
and \U$33474 ( \33852 , \33841 , \33850 );
or \U$33475 ( \33853 , \33846 , \33851 , \33852 );
xor \U$33476 ( \33854 , \33683 , \33687 );
xor \U$33477 ( \33855 , \33854 , \33692 );
and \U$33478 ( \33856 , \33853 , \33855 );
xor \U$33479 ( \33857 , \33536 , \33540 );
xor \U$33480 ( \33858 , \33857 , \33545 );
and \U$33481 ( \33859 , \33855 , \33858 );
and \U$33482 ( \33860 , \33853 , \33858 );
or \U$33483 ( \33861 , \33856 , \33859 , \33860 );
and \U$33484 ( \33862 , \33837 , \33861 );
xor \U$33485 ( \33863 , \33614 , \33618 );
xor \U$33486 ( \33864 , \33863 , \33623 );
xor \U$33487 ( \33865 , \33578 , \33582 );
xor \U$33488 ( \33866 , \33865 , \33587 );
and \U$33489 ( \33867 , \33864 , \33866 );
xor \U$33490 ( \33868 , \33595 , \33599 );
xor \U$33491 ( \33869 , \33868 , \33604 );
and \U$33492 ( \33870 , \33866 , \33869 );
and \U$33493 ( \33871 , \33864 , \33869 );
or \U$33494 ( \33872 , \33867 , \33870 , \33871 );
and \U$33495 ( \33873 , \33861 , \33872 );
and \U$33496 ( \33874 , \33837 , \33872 );
or \U$33497 ( \33875 , \33862 , \33873 , \33874 );
and \U$33498 ( \33876 , \22523 , \29104 );
and \U$33499 ( \33877 , \22325 , \29102 );
nor \U$33500 ( \33878 , \33876 , \33877 );
xnor \U$33501 ( \33879 , \33878 , \28855 );
and \U$33502 ( \33880 , \22716 , \28575 );
and \U$33503 ( \33881 , \22611 , \28573 );
nor \U$33504 ( \33882 , \33880 , \33881 );
xnor \U$33505 ( \33883 , \33882 , \28315 );
and \U$33506 ( \33884 , \33879 , \33883 );
and \U$33507 ( \33885 , \22837 , \28081 );
and \U$33508 ( \33886 , \22721 , \28079 );
nor \U$33509 ( \33887 , \33885 , \33886 );
xnor \U$33510 ( \33888 , \33887 , \27766 );
and \U$33511 ( \33889 , \33883 , \33888 );
and \U$33512 ( \33890 , \33879 , \33888 );
or \U$33513 ( \33891 , \33884 , \33889 , \33890 );
and \U$33514 ( \33892 , \21831 , \32151 );
and \U$33515 ( \33893 , \21762 , \32148 );
nor \U$33516 ( \33894 , \33892 , \33893 );
xnor \U$33517 ( \33895 , \33894 , \31096 );
and \U$33518 ( \33896 , \21890 , \31338 );
and \U$33519 ( \33897 , \21836 , \31336 );
nor \U$33520 ( \33898 , \33896 , \33897 );
xnor \U$33521 ( \33899 , \33898 , \31099 );
and \U$33522 ( \33900 , \33895 , \33899 );
and \U$33523 ( \33901 , \33899 , \21715 );
and \U$33524 ( \33902 , \33895 , \21715 );
or \U$33525 ( \33903 , \33900 , \33901 , \33902 );
and \U$33526 ( \33904 , \33891 , \33903 );
and \U$33527 ( \33905 , \22018 , \30770 );
and \U$33528 ( \33906 , \21941 , \30768 );
nor \U$33529 ( \33907 , \33905 , \33906 );
xnor \U$33530 ( \33908 , \33907 , \30460 );
and \U$33531 ( \33909 , \22126 , \30233 );
and \U$33532 ( \33910 , \22046 , \30231 );
nor \U$33533 ( \33911 , \33909 , \33910 );
xnor \U$33534 ( \33912 , \33911 , \29862 );
and \U$33535 ( \33913 , \33908 , \33912 );
and \U$33536 ( \33914 , \22262 , \29671 );
and \U$33537 ( \33915 , \22200 , \29669 );
nor \U$33538 ( \33916 , \33914 , \33915 );
xnor \U$33539 ( \33917 , \33916 , \29353 );
and \U$33540 ( \33918 , \33912 , \33917 );
and \U$33541 ( \33919 , \33908 , \33917 );
or \U$33542 ( \33920 , \33913 , \33918 , \33919 );
and \U$33543 ( \33921 , \33903 , \33920 );
and \U$33544 ( \33922 , \33891 , \33920 );
or \U$33545 ( \33923 , \33904 , \33921 , \33922 );
and \U$33546 ( \33924 , \25018 , \24974 );
and \U$33547 ( \33925 , \24601 , \24972 );
nor \U$33548 ( \33926 , \33924 , \33925 );
xnor \U$33549 ( \33927 , \33926 , \24787 );
and \U$33550 ( \33928 , \25348 , \24661 );
and \U$33551 ( \33929 , \25226 , \24659 );
nor \U$33552 ( \33930 , \33928 , \33929 );
xnor \U$33553 ( \33931 , \33930 , \24456 );
and \U$33554 ( \33932 , \33927 , \33931 );
and \U$33555 ( \33933 , \25609 , \24255 );
and \U$33556 ( \33934 , \25353 , \24253 );
nor \U$33557 ( \33935 , \33933 , \33934 );
xnor \U$33558 ( \33936 , \33935 , \24106 );
and \U$33559 ( \33937 , \33931 , \33936 );
and \U$33560 ( \33938 , \33927 , \33936 );
or \U$33561 ( \33939 , \33932 , \33937 , \33938 );
and \U$33562 ( \33940 , \23978 , \26143 );
and \U$33563 ( \33941 , \23714 , \26141 );
nor \U$33564 ( \33942 , \33940 , \33941 );
xnor \U$33565 ( \33943 , \33942 , \25911 );
and \U$33566 ( \33944 , \24177 , \25692 );
and \U$33567 ( \33945 , \24003 , \25690 );
nor \U$33568 ( \33946 , \33944 , \33945 );
xnor \U$33569 ( \33947 , \33946 , \25549 );
and \U$33570 ( \33948 , \33943 , \33947 );
and \U$33571 ( \33949 , \24482 , \25369 );
and \U$33572 ( \33950 , \24344 , \25367 );
nor \U$33573 ( \33951 , \33949 , \33950 );
xnor \U$33574 ( \33952 , \33951 , \25123 );
and \U$33575 ( \33953 , \33947 , \33952 );
and \U$33576 ( \33954 , \33943 , \33952 );
or \U$33577 ( \33955 , \33948 , \33953 , \33954 );
and \U$33578 ( \33956 , \33939 , \33955 );
and \U$33579 ( \33957 , \23128 , \27572 );
and \U$33580 ( \33958 , \22952 , \27570 );
nor \U$33581 ( \33959 , \33957 , \33958 );
xnor \U$33582 ( \33960 , \33959 , \27232 );
and \U$33583 ( \33961 , \23379 , \26983 );
and \U$33584 ( \33962 , \23136 , \26981 );
nor \U$33585 ( \33963 , \33961 , \33962 );
xnor \U$33586 ( \33964 , \33963 , \26742 );
and \U$33587 ( \33965 , \33960 , \33964 );
and \U$33588 ( \33966 , \23570 , \26517 );
and \U$33589 ( \33967 , \23384 , \26515 );
nor \U$33590 ( \33968 , \33966 , \33967 );
xnor \U$33591 ( \33969 , \33968 , \26329 );
and \U$33592 ( \33970 , \33964 , \33969 );
and \U$33593 ( \33971 , \33960 , \33969 );
or \U$33594 ( \33972 , \33965 , \33970 , \33971 );
and \U$33595 ( \33973 , \33955 , \33972 );
and \U$33596 ( \33974 , \33939 , \33972 );
or \U$33597 ( \33975 , \33956 , \33973 , \33974 );
and \U$33598 ( \33976 , \33923 , \33975 );
and \U$33599 ( \33977 , \26108 , \23933 );
and \U$33600 ( \33978 , \25806 , \23931 );
nor \U$33601 ( \33979 , \33977 , \33978 );
xnor \U$33602 ( \33980 , \33979 , \23791 );
and \U$33603 ( \33981 , \26585 , \23637 );
and \U$33604 ( \33982 , \26116 , \23635 );
nor \U$33605 ( \33983 , \33981 , \33982 );
xnor \U$33606 ( \33984 , \33983 , \23500 );
and \U$33607 ( \33985 , \33980 , \33984 );
and \U$33608 ( \33986 , \26854 , \23431 );
and \U$33609 ( \33987 , \26590 , \23429 );
nor \U$33610 ( \33988 , \33986 , \33987 );
xnor \U$33611 ( \33989 , \33988 , \23279 );
and \U$33612 ( \33990 , \33984 , \33989 );
and \U$33613 ( \33991 , \33980 , \33989 );
or \U$33614 ( \33992 , \33985 , \33990 , \33991 );
and \U$33615 ( \33993 , \27485 , \23163 );
and \U$33616 ( \33994 , \27113 , \23161 );
nor \U$33617 ( \33995 , \33993 , \33994 );
xnor \U$33618 ( \33996 , \33995 , \23007 );
and \U$33619 ( \33997 , \27837 , \22891 );
and \U$33620 ( \33998 , \27494 , \22889 );
nor \U$33621 ( \33999 , \33997 , \33998 );
xnor \U$33622 ( \34000 , \33999 , \22778 );
and \U$33623 ( \34001 , \33996 , \34000 );
and \U$33624 ( \34002 , \28342 , \22697 );
and \U$33625 ( \34003 , \28039 , \22695 );
nor \U$33626 ( \34004 , \34002 , \34003 );
xnor \U$33627 ( \34005 , \34004 , \22561 );
and \U$33628 ( \34006 , \34000 , \34005 );
and \U$33629 ( \34007 , \33996 , \34005 );
or \U$33630 ( \34008 , \34001 , \34006 , \34007 );
and \U$33631 ( \34009 , \33992 , \34008 );
and \U$33632 ( \34010 , \29040 , \22497 );
and \U$33633 ( \34011 , \28514 , \22495 );
nor \U$33634 ( \34012 , \34010 , \34011 );
xnor \U$33635 ( \34013 , \34012 , \22419 );
and \U$33636 ( \34014 , \29710 , \22333 );
and \U$33637 ( \34015 , \29464 , \22331 );
nor \U$33638 ( \34016 , \34014 , \34015 );
xnor \U$33639 ( \34017 , \34016 , \22239 );
and \U$33640 ( \34018 , \34013 , \34017 );
and \U$33641 ( \34019 , \30034 , \22163 );
and \U$33642 ( \34020 , \29715 , \22161 );
nor \U$33643 ( \34021 , \34019 , \34020 );
xnor \U$33644 ( \34022 , \34021 , \22091 );
and \U$33645 ( \34023 , \34017 , \34022 );
and \U$33646 ( \34024 , \34013 , \34022 );
or \U$33647 ( \34025 , \34018 , \34023 , \34024 );
and \U$33648 ( \34026 , \34008 , \34025 );
and \U$33649 ( \34027 , \33992 , \34025 );
or \U$33650 ( \34028 , \34009 , \34026 , \34027 );
and \U$33651 ( \34029 , \33975 , \34028 );
and \U$33652 ( \34030 , \33923 , \34028 );
or \U$33653 ( \34031 , \33976 , \34029 , \34030 );
and \U$33654 ( \34032 , \33875 , \34031 );
xor \U$33655 ( \34033 , \33721 , \33723 );
xor \U$33656 ( \34034 , \34033 , \33726 );
xor \U$33657 ( \34035 , \33513 , \33515 );
xor \U$33658 ( \34036 , \34035 , \33518 );
and \U$33659 ( \34037 , \34034 , \34036 );
xor \U$33660 ( \34038 , \33523 , \33525 );
xor \U$33661 ( \34039 , \34038 , \33528 );
and \U$33662 ( \34040 , \34036 , \34039 );
and \U$33663 ( \34041 , \34034 , \34039 );
or \U$33664 ( \34042 , \34037 , \34040 , \34041 );
and \U$33665 ( \34043 , \34031 , \34042 );
and \U$33666 ( \34044 , \33875 , \34042 );
or \U$33667 ( \34045 , \34032 , \34043 , \34044 );
xor \U$33668 ( \34046 , \33574 , \33590 );
xor \U$33669 ( \34047 , \34046 , \33607 );
xor \U$33670 ( \34048 , \33679 , \33695 );
xor \U$33671 ( \34049 , \34048 , \33712 );
and \U$33672 ( \34050 , \34047 , \34049 );
xor \U$33673 ( \34051 , \33548 , \33550 );
xor \U$33674 ( \34052 , \34051 , \33552 );
and \U$33675 ( \34053 , \34049 , \34052 );
and \U$33676 ( \34054 , \34047 , \34052 );
or \U$33677 ( \34055 , \34050 , \34053 , \34054 );
xor \U$33678 ( \34056 , \33742 , \33744 );
xor \U$33679 ( \34057 , \34056 , \33747 );
and \U$33680 ( \34058 , \34055 , \34057 );
xor \U$33681 ( \34059 , \33752 , \33754 );
xor \U$33682 ( \34060 , \34059 , \33757 );
and \U$33683 ( \34061 , \34057 , \34060 );
and \U$33684 ( \34062 , \34055 , \34060 );
or \U$33685 ( \34063 , \34058 , \34061 , \34062 );
and \U$33686 ( \34064 , \34045 , \34063 );
xor \U$33687 ( \34065 , \33521 , \33531 );
xor \U$33688 ( \34066 , \34065 , \33555 );
xor \U$33689 ( \34067 , \33610 , \33662 );
xor \U$33690 ( \34068 , \34067 , \33715 );
and \U$33691 ( \34069 , \34066 , \34068 );
xor \U$33692 ( \34070 , \33729 , \33731 );
xor \U$33693 ( \34071 , \34070 , \33734 );
and \U$33694 ( \34072 , \34068 , \34071 );
and \U$33695 ( \34073 , \34066 , \34071 );
or \U$33696 ( \34074 , \34069 , \34072 , \34073 );
and \U$33697 ( \34075 , \34063 , \34074 );
and \U$33698 ( \34076 , \34045 , \34074 );
or \U$33699 ( \34077 , \34064 , \34075 , \34076 );
xor \U$33700 ( \34078 , \33263 , \33311 );
xor \U$33701 ( \34079 , \34078 , \33364 );
xor \U$33702 ( \34080 , \33398 , \33408 );
xor \U$33703 ( \34081 , \34080 , \33419 );
and \U$33704 ( \34082 , \34079 , \34081 );
xor \U$33705 ( \34083 , \33769 , \33771 );
xor \U$33706 ( \34084 , \34083 , \33774 );
and \U$33707 ( \34085 , \34081 , \34084 );
and \U$33708 ( \34086 , \34079 , \34084 );
or \U$33709 ( \34087 , \34082 , \34085 , \34086 );
and \U$33710 ( \34088 , \34077 , \34087 );
xor \U$33711 ( \34089 , \33782 , \33784 );
xor \U$33712 ( \34090 , \34089 , \33787 );
and \U$33713 ( \34091 , \34087 , \34090 );
and \U$33714 ( \34092 , \34077 , \34090 );
or \U$33715 ( \34093 , \34088 , \34091 , \34092 );
xor \U$33716 ( \34094 , \33780 , \33790 );
xor \U$33717 ( \34095 , \34094 , \33793 );
and \U$33718 ( \34096 , \34093 , \34095 );
xor \U$33719 ( \34097 , \33798 , \33800 );
xor \U$33720 ( \34098 , \34097 , \33803 );
and \U$33721 ( \34099 , \34095 , \34098 );
and \U$33722 ( \34100 , \34093 , \34098 );
or \U$33723 ( \34101 , \34096 , \34099 , \34100 );
xor \U$33724 ( \34102 , \33796 , \33806 );
xor \U$33725 ( \34103 , \34102 , \33809 );
and \U$33726 ( \34104 , \34101 , \34103 );
xor \U$33727 ( \34105 , \33814 , \33816 );
and \U$33728 ( \34106 , \34103 , \34105 );
and \U$33729 ( \34107 , \34101 , \34105 );
or \U$33730 ( \34108 , \34104 , \34106 , \34107 );
and \U$33731 ( \34109 , \33827 , \34108 );
xor \U$33732 ( \34110 , \33827 , \34108 );
xor \U$33733 ( \34111 , \34101 , \34103 );
xor \U$33734 ( \34112 , \34111 , \34105 );
and \U$33735 ( \34113 , \24344 , \25692 );
and \U$33736 ( \34114 , \24177 , \25690 );
nor \U$33737 ( \34115 , \34113 , \34114 );
xnor \U$33738 ( \34116 , \34115 , \25549 );
and \U$33739 ( \34117 , \24601 , \25369 );
and \U$33740 ( \34118 , \24482 , \25367 );
nor \U$33741 ( \34119 , \34117 , \34118 );
xnor \U$33742 ( \34120 , \34119 , \25123 );
and \U$33743 ( \34121 , \34116 , \34120 );
and \U$33744 ( \34122 , \25226 , \24974 );
and \U$33745 ( \34123 , \25018 , \24972 );
nor \U$33746 ( \34124 , \34122 , \34123 );
xnor \U$33747 ( \34125 , \34124 , \24787 );
and \U$33748 ( \34126 , \34120 , \34125 );
and \U$33749 ( \34127 , \34116 , \34125 );
or \U$33750 ( \34128 , \34121 , \34126 , \34127 );
and \U$33751 ( \34129 , \25353 , \24661 );
and \U$33752 ( \34130 , \25348 , \24659 );
nor \U$33753 ( \34131 , \34129 , \34130 );
xnor \U$33754 ( \34132 , \34131 , \24456 );
and \U$33755 ( \34133 , \25806 , \24255 );
and \U$33756 ( \34134 , \25609 , \24253 );
nor \U$33757 ( \34135 , \34133 , \34134 );
xnor \U$33758 ( \34136 , \34135 , \24106 );
and \U$33759 ( \34137 , \34132 , \34136 );
and \U$33760 ( \34138 , \26116 , \23933 );
and \U$33761 ( \34139 , \26108 , \23931 );
nor \U$33762 ( \34140 , \34138 , \34139 );
xnor \U$33763 ( \34141 , \34140 , \23791 );
and \U$33764 ( \34142 , \34136 , \34141 );
and \U$33765 ( \34143 , \34132 , \34141 );
or \U$33766 ( \34144 , \34137 , \34142 , \34143 );
and \U$33767 ( \34145 , \34128 , \34144 );
and \U$33768 ( \34146 , \23384 , \26983 );
and \U$33769 ( \34147 , \23379 , \26981 );
nor \U$33770 ( \34148 , \34146 , \34147 );
xnor \U$33771 ( \34149 , \34148 , \26742 );
and \U$33772 ( \34150 , \23714 , \26517 );
and \U$33773 ( \34151 , \23570 , \26515 );
nor \U$33774 ( \34152 , \34150 , \34151 );
xnor \U$33775 ( \34153 , \34152 , \26329 );
and \U$33776 ( \34154 , \34149 , \34153 );
and \U$33777 ( \34155 , \24003 , \26143 );
and \U$33778 ( \34156 , \23978 , \26141 );
nor \U$33779 ( \34157 , \34155 , \34156 );
xnor \U$33780 ( \34158 , \34157 , \25911 );
and \U$33781 ( \34159 , \34153 , \34158 );
and \U$33782 ( \34160 , \34149 , \34158 );
or \U$33783 ( \34161 , \34154 , \34159 , \34160 );
and \U$33784 ( \34162 , \34144 , \34161 );
and \U$33785 ( \34163 , \34128 , \34161 );
or \U$33786 ( \34164 , \34145 , \34162 , \34163 );
and \U$33787 ( \34165 , \28039 , \22891 );
and \U$33788 ( \34166 , \27837 , \22889 );
nor \U$33789 ( \34167 , \34165 , \34166 );
xnor \U$33790 ( \34168 , \34167 , \22778 );
and \U$33791 ( \34169 , \28514 , \22697 );
and \U$33792 ( \34170 , \28342 , \22695 );
nor \U$33793 ( \34171 , \34169 , \34170 );
xnor \U$33794 ( \34172 , \34171 , \22561 );
and \U$33795 ( \34173 , \34168 , \34172 );
and \U$33796 ( \34174 , \29464 , \22497 );
and \U$33797 ( \34175 , \29040 , \22495 );
nor \U$33798 ( \34176 , \34174 , \34175 );
xnor \U$33799 ( \34177 , \34176 , \22419 );
and \U$33800 ( \34178 , \34172 , \34177 );
and \U$33801 ( \34179 , \34168 , \34177 );
or \U$33802 ( \34180 , \34173 , \34178 , \34179 );
and \U$33803 ( \34181 , \29715 , \22333 );
and \U$33804 ( \34182 , \29710 , \22331 );
nor \U$33805 ( \34183 , \34181 , \34182 );
xnor \U$33806 ( \34184 , \34183 , \22239 );
and \U$33807 ( \34185 , \30318 , \22163 );
and \U$33808 ( \34186 , \30034 , \22161 );
nor \U$33809 ( \34187 , \34185 , \34186 );
xnor \U$33810 ( \34188 , \34187 , \22091 );
and \U$33811 ( \34189 , \34184 , \34188 );
and \U$33812 ( \34190 , \30895 , \22029 );
and \U$33813 ( \34191 , \30887 , \22027 );
nor \U$33814 ( \34192 , \34190 , \34191 );
xnor \U$33815 ( \34193 , \34192 , \21986 );
and \U$33816 ( \34194 , \34188 , \34193 );
and \U$33817 ( \34195 , \34184 , \34193 );
or \U$33818 ( \34196 , \34189 , \34194 , \34195 );
and \U$33819 ( \34197 , \34180 , \34196 );
and \U$33820 ( \34198 , \26590 , \23637 );
and \U$33821 ( \34199 , \26585 , \23635 );
nor \U$33822 ( \34200 , \34198 , \34199 );
xnor \U$33823 ( \34201 , \34200 , \23500 );
and \U$33824 ( \34202 , \27113 , \23431 );
and \U$33825 ( \34203 , \26854 , \23429 );
nor \U$33826 ( \34204 , \34202 , \34203 );
xnor \U$33827 ( \34205 , \34204 , \23279 );
and \U$33828 ( \34206 , \34201 , \34205 );
and \U$33829 ( \34207 , \27494 , \23163 );
and \U$33830 ( \34208 , \27485 , \23161 );
nor \U$33831 ( \34209 , \34207 , \34208 );
xnor \U$33832 ( \34210 , \34209 , \23007 );
and \U$33833 ( \34211 , \34205 , \34210 );
and \U$33834 ( \34212 , \34201 , \34210 );
or \U$33835 ( \34213 , \34206 , \34211 , \34212 );
and \U$33836 ( \34214 , \34196 , \34213 );
and \U$33837 ( \34215 , \34180 , \34213 );
or \U$33838 ( \34216 , \34197 , \34214 , \34215 );
and \U$33839 ( \34217 , \34164 , \34216 );
and \U$33840 ( \34218 , \21836 , \32151 );
and \U$33841 ( \34219 , \21831 , \32148 );
nor \U$33842 ( \34220 , \34218 , \34219 );
xnor \U$33843 ( \34221 , \34220 , \31096 );
and \U$33844 ( \34222 , \21941 , \31338 );
and \U$33845 ( \34223 , \21890 , \31336 );
nor \U$33846 ( \34224 , \34222 , \34223 );
xnor \U$33847 ( \34225 , \34224 , \31099 );
and \U$33848 ( \34226 , \34221 , \34225 );
and \U$33849 ( \34227 , \22046 , \30770 );
and \U$33850 ( \34228 , \22018 , \30768 );
nor \U$33851 ( \34229 , \34227 , \34228 );
xnor \U$33852 ( \34230 , \34229 , \30460 );
and \U$33853 ( \34231 , \34225 , \34230 );
and \U$33854 ( \34232 , \34221 , \34230 );
or \U$33855 ( \34233 , \34226 , \34231 , \34232 );
and \U$33856 ( \34234 , \22200 , \30233 );
and \U$33857 ( \34235 , \22126 , \30231 );
nor \U$33858 ( \34236 , \34234 , \34235 );
xnor \U$33859 ( \34237 , \34236 , \29862 );
and \U$33860 ( \34238 , \22325 , \29671 );
and \U$33861 ( \34239 , \22262 , \29669 );
nor \U$33862 ( \34240 , \34238 , \34239 );
xnor \U$33863 ( \34241 , \34240 , \29353 );
and \U$33864 ( \34242 , \34237 , \34241 );
and \U$33865 ( \34243 , \22611 , \29104 );
and \U$33866 ( \34244 , \22523 , \29102 );
nor \U$33867 ( \34245 , \34243 , \34244 );
xnor \U$33868 ( \34246 , \34245 , \28855 );
and \U$33869 ( \34247 , \34241 , \34246 );
and \U$33870 ( \34248 , \34237 , \34246 );
or \U$33871 ( \34249 , \34242 , \34247 , \34248 );
and \U$33872 ( \34250 , \34233 , \34249 );
and \U$33873 ( \34251 , \22721 , \28575 );
and \U$33874 ( \34252 , \22716 , \28573 );
nor \U$33875 ( \34253 , \34251 , \34252 );
xnor \U$33876 ( \34254 , \34253 , \28315 );
and \U$33877 ( \34255 , \22952 , \28081 );
and \U$33878 ( \34256 , \22837 , \28079 );
nor \U$33879 ( \34257 , \34255 , \34256 );
xnor \U$33880 ( \34258 , \34257 , \27766 );
and \U$33881 ( \34259 , \34254 , \34258 );
and \U$33882 ( \34260 , \23136 , \27572 );
and \U$33883 ( \34261 , \23128 , \27570 );
nor \U$33884 ( \34262 , \34260 , \34261 );
xnor \U$33885 ( \34263 , \34262 , \27232 );
and \U$33886 ( \34264 , \34258 , \34263 );
and \U$33887 ( \34265 , \34254 , \34263 );
or \U$33888 ( \34266 , \34259 , \34264 , \34265 );
and \U$33889 ( \34267 , \34249 , \34266 );
and \U$33890 ( \34268 , \34233 , \34266 );
or \U$33891 ( \34269 , \34250 , \34267 , \34268 );
and \U$33892 ( \34270 , \34216 , \34269 );
and \U$33893 ( \34271 , \34164 , \34269 );
or \U$33894 ( \34272 , \34217 , \34270 , \34271 );
xor \U$33895 ( \34273 , \33879 , \33883 );
xor \U$33896 ( \34274 , \34273 , \33888 );
xor \U$33897 ( \34275 , \33943 , \33947 );
xor \U$33898 ( \34276 , \34275 , \33952 );
and \U$33899 ( \34277 , \34274 , \34276 );
xor \U$33900 ( \34278 , \33960 , \33964 );
xor \U$33901 ( \34279 , \34278 , \33969 );
and \U$33902 ( \34280 , \34276 , \34279 );
and \U$33903 ( \34281 , \34274 , \34279 );
or \U$33904 ( \34282 , \34277 , \34280 , \34281 );
xor \U$33905 ( \34283 , \33927 , \33931 );
xor \U$33906 ( \34284 , \34283 , \33936 );
xor \U$33907 ( \34285 , \33980 , \33984 );
xor \U$33908 ( \34286 , \34285 , \33989 );
and \U$33909 ( \34287 , \34284 , \34286 );
xor \U$33910 ( \34288 , \33996 , \34000 );
xor \U$33911 ( \34289 , \34288 , \34005 );
and \U$33912 ( \34290 , \34286 , \34289 );
and \U$33913 ( \34291 , \34284 , \34289 );
or \U$33914 ( \34292 , \34287 , \34290 , \34291 );
and \U$33915 ( \34293 , \34282 , \34292 );
nand \U$33916 ( \34294 , \32304 , \21743 );
xnor \U$33917 ( \34295 , \34294 , \21715 );
xor \U$33918 ( \34296 , \34013 , \34017 );
xor \U$33919 ( \34297 , \34296 , \34022 );
and \U$33920 ( \34298 , \34295 , \34297 );
xor \U$33921 ( \34299 , \33841 , \33845 );
xor \U$33922 ( \34300 , \34299 , \33850 );
and \U$33923 ( \34301 , \34297 , \34300 );
and \U$33924 ( \34302 , \34295 , \34300 );
or \U$33925 ( \34303 , \34298 , \34301 , \34302 );
and \U$33926 ( \34304 , \34292 , \34303 );
and \U$33927 ( \34305 , \34282 , \34303 );
or \U$33928 ( \34306 , \34293 , \34304 , \34305 );
and \U$33929 ( \34307 , \34272 , \34306 );
xor \U$33930 ( \34308 , \33630 , \33634 );
xor \U$33931 ( \34309 , \34308 , \33639 );
xor \U$33932 ( \34310 , \33647 , \33651 );
xor \U$33933 ( \34311 , \34310 , \33656 );
and \U$33934 ( \34312 , \34309 , \34311 );
xor \U$33935 ( \34313 , \33864 , \33866 );
xor \U$33936 ( \34314 , \34313 , \33869 );
and \U$33937 ( \34315 , \34311 , \34314 );
and \U$33938 ( \34316 , \34309 , \34314 );
or \U$33939 ( \34317 , \34312 , \34315 , \34316 );
and \U$33940 ( \34318 , \34306 , \34317 );
and \U$33941 ( \34319 , \34272 , \34317 );
or \U$33942 ( \34320 , \34307 , \34318 , \34319 );
xor \U$33943 ( \34321 , \33837 , \33861 );
xor \U$33944 ( \34322 , \34321 , \33872 );
xor \U$33945 ( \34323 , \33923 , \33975 );
xor \U$33946 ( \34324 , \34323 , \34028 );
and \U$33947 ( \34325 , \34322 , \34324 );
xor \U$33948 ( \34326 , \34034 , \34036 );
xor \U$33949 ( \34327 , \34326 , \34039 );
and \U$33950 ( \34328 , \34324 , \34327 );
and \U$33951 ( \34329 , \34322 , \34327 );
or \U$33952 ( \34330 , \34325 , \34328 , \34329 );
and \U$33953 ( \34331 , \34320 , \34330 );
xor \U$33954 ( \34332 , \33992 , \34008 );
xor \U$33955 ( \34333 , \34332 , \34025 );
xor \U$33956 ( \34334 , \33829 , \33831 );
xor \U$33957 ( \34335 , \34334 , \33834 );
and \U$33958 ( \34336 , \34333 , \34335 );
xor \U$33959 ( \34337 , \33853 , \33855 );
xor \U$33960 ( \34338 , \34337 , \33858 );
and \U$33961 ( \34339 , \34335 , \34338 );
and \U$33962 ( \34340 , \34333 , \34338 );
or \U$33963 ( \34341 , \34336 , \34339 , \34340 );
xor \U$33964 ( \34342 , \33626 , \33642 );
xor \U$33965 ( \34343 , \34342 , \33659 );
and \U$33966 ( \34344 , \34341 , \34343 );
xor \U$33967 ( \34345 , \34047 , \34049 );
xor \U$33968 ( \34346 , \34345 , \34052 );
and \U$33969 ( \34347 , \34343 , \34346 );
and \U$33970 ( \34348 , \34341 , \34346 );
or \U$33971 ( \34349 , \34344 , \34347 , \34348 );
and \U$33972 ( \34350 , \34330 , \34349 );
and \U$33973 ( \34351 , \34320 , \34349 );
or \U$33974 ( \34352 , \34331 , \34350 , \34351 );
xor \U$33975 ( \34353 , \33875 , \34031 );
xor \U$33976 ( \34354 , \34353 , \34042 );
xor \U$33977 ( \34355 , \34055 , \34057 );
xor \U$33978 ( \34356 , \34355 , \34060 );
and \U$33979 ( \34357 , \34354 , \34356 );
xor \U$33980 ( \34358 , \34066 , \34068 );
xor \U$33981 ( \34359 , \34358 , \34071 );
and \U$33982 ( \34360 , \34356 , \34359 );
and \U$33983 ( \34361 , \34354 , \34359 );
or \U$33984 ( \34362 , \34357 , \34360 , \34361 );
and \U$33985 ( \34363 , \34352 , \34362 );
xor \U$33986 ( \34364 , \33750 , \33760 );
xor \U$33987 ( \34365 , \34364 , \33763 );
and \U$33988 ( \34366 , \34362 , \34365 );
and \U$33989 ( \34367 , \34352 , \34365 );
or \U$33990 ( \34368 , \34363 , \34366 , \34367 );
xor \U$33991 ( \34369 , \33558 , \33718 );
xor \U$33992 ( \34370 , \34369 , \33737 );
xor \U$33993 ( \34371 , \34045 , \34063 );
xor \U$33994 ( \34372 , \34371 , \34074 );
and \U$33995 ( \34373 , \34370 , \34372 );
xor \U$33996 ( \34374 , \34079 , \34081 );
xor \U$33997 ( \34375 , \34374 , \34084 );
and \U$33998 ( \34376 , \34372 , \34375 );
and \U$33999 ( \34377 , \34370 , \34375 );
or \U$34000 ( \34378 , \34373 , \34376 , \34377 );
and \U$34001 ( \34379 , \34368 , \34378 );
xor \U$34002 ( \34380 , \33740 , \33766 );
xor \U$34003 ( \34381 , \34380 , \33777 );
and \U$34004 ( \34382 , \34378 , \34381 );
and \U$34005 ( \34383 , \34368 , \34381 );
or \U$34006 ( \34384 , \34379 , \34382 , \34383 );
xor \U$34007 ( \34385 , \34093 , \34095 );
xor \U$34008 ( \34386 , \34385 , \34098 );
and \U$34009 ( \34387 , \34384 , \34386 );
and \U$34010 ( \34388 , \34112 , \34387 );
xor \U$34011 ( \34389 , \34112 , \34387 );
xor \U$34012 ( \34390 , \34384 , \34386 );
and \U$34013 ( \34391 , \31498 , \22029 );
and \U$34014 ( \34392 , \30895 , \22027 );
nor \U$34015 ( \34393 , \34391 , \34392 );
xnor \U$34016 ( \34394 , \34393 , \21986 );
and \U$34017 ( \34395 , \31684 , \21916 );
and \U$34018 ( \34396 , \31503 , \21914 );
nor \U$34019 ( \34397 , \34395 , \34396 );
xnor \U$34020 ( \34398 , \34397 , \21867 );
and \U$34021 ( \34399 , \34394 , \34398 );
nand \U$34022 ( \34400 , \32304 , \21813 );
xnor \U$34023 ( \34401 , \34400 , \21774 );
and \U$34024 ( \34402 , \34398 , \34401 );
and \U$34025 ( \34403 , \34394 , \34401 );
or \U$34026 ( \34404 , \34399 , \34402 , \34403 );
and \U$34027 ( \34405 , \31503 , \21916 );
and \U$34028 ( \34406 , \31498 , \21914 );
nor \U$34029 ( \34407 , \34405 , \34406 );
xnor \U$34030 ( \34408 , \34407 , \21867 );
and \U$34031 ( \34409 , \34404 , \34408 );
and \U$34032 ( \34410 , \32304 , \21815 );
and \U$34033 ( \34411 , \31684 , \21813 );
nor \U$34034 ( \34412 , \34410 , \34411 );
xnor \U$34035 ( \34413 , \34412 , \21774 );
and \U$34036 ( \34414 , \34408 , \34413 );
and \U$34037 ( \34415 , \34404 , \34413 );
or \U$34038 ( \34416 , \34409 , \34414 , \34415 );
xor \U$34039 ( \34417 , \34168 , \34172 );
xor \U$34040 ( \34418 , \34417 , \34177 );
xor \U$34041 ( \34419 , \34184 , \34188 );
xor \U$34042 ( \34420 , \34419 , \34193 );
and \U$34043 ( \34421 , \34418 , \34420 );
xor \U$34044 ( \34422 , \34201 , \34205 );
xor \U$34045 ( \34423 , \34422 , \34210 );
and \U$34046 ( \34424 , \34420 , \34423 );
and \U$34047 ( \34425 , \34418 , \34423 );
or \U$34048 ( \34426 , \34421 , \34424 , \34425 );
and \U$34049 ( \34427 , \34416 , \34426 );
xor \U$34050 ( \34428 , \34116 , \34120 );
xor \U$34051 ( \34429 , \34428 , \34125 );
xor \U$34052 ( \34430 , \34132 , \34136 );
xor \U$34053 ( \34431 , \34430 , \34141 );
and \U$34054 ( \34432 , \34429 , \34431 );
xor \U$34055 ( \34433 , \34149 , \34153 );
xor \U$34056 ( \34434 , \34433 , \34158 );
and \U$34057 ( \34435 , \34431 , \34434 );
and \U$34058 ( \34436 , \34429 , \34434 );
or \U$34059 ( \34437 , \34432 , \34435 , \34436 );
and \U$34060 ( \34438 , \34426 , \34437 );
and \U$34061 ( \34439 , \34416 , \34437 );
or \U$34062 ( \34440 , \34427 , \34438 , \34439 );
and \U$34063 ( \34441 , \22126 , \30770 );
and \U$34064 ( \34442 , \22046 , \30768 );
nor \U$34065 ( \34443 , \34441 , \34442 );
xnor \U$34066 ( \34444 , \34443 , \30460 );
and \U$34067 ( \34445 , \22262 , \30233 );
and \U$34068 ( \34446 , \22200 , \30231 );
nor \U$34069 ( \34447 , \34445 , \34446 );
xnor \U$34070 ( \34448 , \34447 , \29862 );
and \U$34071 ( \34449 , \34444 , \34448 );
and \U$34072 ( \34450 , \22523 , \29671 );
and \U$34073 ( \34451 , \22325 , \29669 );
nor \U$34074 ( \34452 , \34450 , \34451 );
xnor \U$34075 ( \34453 , \34452 , \29353 );
and \U$34076 ( \34454 , \34448 , \34453 );
and \U$34077 ( \34455 , \34444 , \34453 );
or \U$34078 ( \34456 , \34449 , \34454 , \34455 );
and \U$34079 ( \34457 , \22716 , \29104 );
and \U$34080 ( \34458 , \22611 , \29102 );
nor \U$34081 ( \34459 , \34457 , \34458 );
xnor \U$34082 ( \34460 , \34459 , \28855 );
and \U$34083 ( \34461 , \22837 , \28575 );
and \U$34084 ( \34462 , \22721 , \28573 );
nor \U$34085 ( \34463 , \34461 , \34462 );
xnor \U$34086 ( \34464 , \34463 , \28315 );
and \U$34087 ( \34465 , \34460 , \34464 );
and \U$34088 ( \34466 , \23128 , \28081 );
and \U$34089 ( \34467 , \22952 , \28079 );
nor \U$34090 ( \34468 , \34466 , \34467 );
xnor \U$34091 ( \34469 , \34468 , \27766 );
and \U$34092 ( \34470 , \34464 , \34469 );
and \U$34093 ( \34471 , \34460 , \34469 );
or \U$34094 ( \34472 , \34465 , \34470 , \34471 );
and \U$34095 ( \34473 , \34456 , \34472 );
and \U$34096 ( \34474 , \21890 , \32151 );
and \U$34097 ( \34475 , \21836 , \32148 );
nor \U$34098 ( \34476 , \34474 , \34475 );
xnor \U$34099 ( \34477 , \34476 , \31096 );
and \U$34100 ( \34478 , \22018 , \31338 );
and \U$34101 ( \34479 , \21941 , \31336 );
nor \U$34102 ( \34480 , \34478 , \34479 );
xnor \U$34103 ( \34481 , \34480 , \31099 );
and \U$34104 ( \34482 , \34477 , \34481 );
and \U$34105 ( \34483 , \34481 , \21774 );
and \U$34106 ( \34484 , \34477 , \21774 );
or \U$34107 ( \34485 , \34482 , \34483 , \34484 );
and \U$34108 ( \34486 , \34472 , \34485 );
and \U$34109 ( \34487 , \34456 , \34485 );
or \U$34110 ( \34488 , \34473 , \34486 , \34487 );
and \U$34111 ( \34489 , \25348 , \24974 );
and \U$34112 ( \34490 , \25226 , \24972 );
nor \U$34113 ( \34491 , \34489 , \34490 );
xnor \U$34114 ( \34492 , \34491 , \24787 );
and \U$34115 ( \34493 , \25609 , \24661 );
and \U$34116 ( \34494 , \25353 , \24659 );
nor \U$34117 ( \34495 , \34493 , \34494 );
xnor \U$34118 ( \34496 , \34495 , \24456 );
and \U$34119 ( \34497 , \34492 , \34496 );
and \U$34120 ( \34498 , \26108 , \24255 );
and \U$34121 ( \34499 , \25806 , \24253 );
nor \U$34122 ( \34500 , \34498 , \34499 );
xnor \U$34123 ( \34501 , \34500 , \24106 );
and \U$34124 ( \34502 , \34496 , \34501 );
and \U$34125 ( \34503 , \34492 , \34501 );
or \U$34126 ( \34504 , \34497 , \34502 , \34503 );
and \U$34127 ( \34505 , \23379 , \27572 );
and \U$34128 ( \34506 , \23136 , \27570 );
nor \U$34129 ( \34507 , \34505 , \34506 );
xnor \U$34130 ( \34508 , \34507 , \27232 );
and \U$34131 ( \34509 , \23570 , \26983 );
and \U$34132 ( \34510 , \23384 , \26981 );
nor \U$34133 ( \34511 , \34509 , \34510 );
xnor \U$34134 ( \34512 , \34511 , \26742 );
and \U$34135 ( \34513 , \34508 , \34512 );
and \U$34136 ( \34514 , \23978 , \26517 );
and \U$34137 ( \34515 , \23714 , \26515 );
nor \U$34138 ( \34516 , \34514 , \34515 );
xnor \U$34139 ( \34517 , \34516 , \26329 );
and \U$34140 ( \34518 , \34512 , \34517 );
and \U$34141 ( \34519 , \34508 , \34517 );
or \U$34142 ( \34520 , \34513 , \34518 , \34519 );
and \U$34143 ( \34521 , \34504 , \34520 );
and \U$34144 ( \34522 , \24177 , \26143 );
and \U$34145 ( \34523 , \24003 , \26141 );
nor \U$34146 ( \34524 , \34522 , \34523 );
xnor \U$34147 ( \34525 , \34524 , \25911 );
and \U$34148 ( \34526 , \24482 , \25692 );
and \U$34149 ( \34527 , \24344 , \25690 );
nor \U$34150 ( \34528 , \34526 , \34527 );
xnor \U$34151 ( \34529 , \34528 , \25549 );
and \U$34152 ( \34530 , \34525 , \34529 );
and \U$34153 ( \34531 , \25018 , \25369 );
and \U$34154 ( \34532 , \24601 , \25367 );
nor \U$34155 ( \34533 , \34531 , \34532 );
xnor \U$34156 ( \34534 , \34533 , \25123 );
and \U$34157 ( \34535 , \34529 , \34534 );
and \U$34158 ( \34536 , \34525 , \34534 );
or \U$34159 ( \34537 , \34530 , \34535 , \34536 );
and \U$34160 ( \34538 , \34520 , \34537 );
and \U$34161 ( \34539 , \34504 , \34537 );
or \U$34162 ( \34540 , \34521 , \34538 , \34539 );
and \U$34163 ( \34541 , \34488 , \34540 );
and \U$34164 ( \34542 , \27837 , \23163 );
and \U$34165 ( \34543 , \27494 , \23161 );
nor \U$34166 ( \34544 , \34542 , \34543 );
xnor \U$34167 ( \34545 , \34544 , \23007 );
and \U$34168 ( \34546 , \28342 , \22891 );
and \U$34169 ( \34547 , \28039 , \22889 );
nor \U$34170 ( \34548 , \34546 , \34547 );
xnor \U$34171 ( \34549 , \34548 , \22778 );
and \U$34172 ( \34550 , \34545 , \34549 );
and \U$34173 ( \34551 , \29040 , \22697 );
and \U$34174 ( \34552 , \28514 , \22695 );
nor \U$34175 ( \34553 , \34551 , \34552 );
xnor \U$34176 ( \34554 , \34553 , \22561 );
and \U$34177 ( \34555 , \34549 , \34554 );
and \U$34178 ( \34556 , \34545 , \34554 );
or \U$34179 ( \34557 , \34550 , \34555 , \34556 );
and \U$34180 ( \34558 , \29710 , \22497 );
and \U$34181 ( \34559 , \29464 , \22495 );
nor \U$34182 ( \34560 , \34558 , \34559 );
xnor \U$34183 ( \34561 , \34560 , \22419 );
and \U$34184 ( \34562 , \30034 , \22333 );
and \U$34185 ( \34563 , \29715 , \22331 );
nor \U$34186 ( \34564 , \34562 , \34563 );
xnor \U$34187 ( \34565 , \34564 , \22239 );
and \U$34188 ( \34566 , \34561 , \34565 );
and \U$34189 ( \34567 , \30887 , \22163 );
and \U$34190 ( \34568 , \30318 , \22161 );
nor \U$34191 ( \34569 , \34567 , \34568 );
xnor \U$34192 ( \34570 , \34569 , \22091 );
and \U$34193 ( \34571 , \34565 , \34570 );
and \U$34194 ( \34572 , \34561 , \34570 );
or \U$34195 ( \34573 , \34566 , \34571 , \34572 );
and \U$34196 ( \34574 , \34557 , \34573 );
and \U$34197 ( \34575 , \26585 , \23933 );
and \U$34198 ( \34576 , \26116 , \23931 );
nor \U$34199 ( \34577 , \34575 , \34576 );
xnor \U$34200 ( \34578 , \34577 , \23791 );
and \U$34201 ( \34579 , \26854 , \23637 );
and \U$34202 ( \34580 , \26590 , \23635 );
nor \U$34203 ( \34581 , \34579 , \34580 );
xnor \U$34204 ( \34582 , \34581 , \23500 );
and \U$34205 ( \34583 , \34578 , \34582 );
and \U$34206 ( \34584 , \27485 , \23431 );
and \U$34207 ( \34585 , \27113 , \23429 );
nor \U$34208 ( \34586 , \34584 , \34585 );
xnor \U$34209 ( \34587 , \34586 , \23279 );
and \U$34210 ( \34588 , \34582 , \34587 );
and \U$34211 ( \34589 , \34578 , \34587 );
or \U$34212 ( \34590 , \34583 , \34588 , \34589 );
and \U$34213 ( \34591 , \34573 , \34590 );
and \U$34214 ( \34592 , \34557 , \34590 );
or \U$34215 ( \34593 , \34574 , \34591 , \34592 );
and \U$34216 ( \34594 , \34540 , \34593 );
and \U$34217 ( \34595 , \34488 , \34593 );
or \U$34218 ( \34596 , \34541 , \34594 , \34595 );
and \U$34219 ( \34597 , \34440 , \34596 );
xor \U$34220 ( \34598 , \34221 , \34225 );
xor \U$34221 ( \34599 , \34598 , \34230 );
xor \U$34222 ( \34600 , \34237 , \34241 );
xor \U$34223 ( \34601 , \34600 , \34246 );
and \U$34224 ( \34602 , \34599 , \34601 );
xor \U$34225 ( \34603 , \34254 , \34258 );
xor \U$34226 ( \34604 , \34603 , \34263 );
and \U$34227 ( \34605 , \34601 , \34604 );
and \U$34228 ( \34606 , \34599 , \34604 );
or \U$34229 ( \34607 , \34602 , \34605 , \34606 );
xor \U$34230 ( \34608 , \33895 , \33899 );
xor \U$34231 ( \34609 , \34608 , \21715 );
and \U$34232 ( \34610 , \34607 , \34609 );
xor \U$34233 ( \34611 , \33908 , \33912 );
xor \U$34234 ( \34612 , \34611 , \33917 );
and \U$34235 ( \34613 , \34609 , \34612 );
and \U$34236 ( \34614 , \34607 , \34612 );
or \U$34237 ( \34615 , \34610 , \34613 , \34614 );
and \U$34238 ( \34616 , \34596 , \34615 );
and \U$34239 ( \34617 , \34440 , \34615 );
or \U$34240 ( \34618 , \34597 , \34616 , \34617 );
xor \U$34241 ( \34619 , \34128 , \34144 );
xor \U$34242 ( \34620 , \34619 , \34161 );
xor \U$34243 ( \34621 , \34180 , \34196 );
xor \U$34244 ( \34622 , \34621 , \34213 );
and \U$34245 ( \34623 , \34620 , \34622 );
xor \U$34246 ( \34624 , \34233 , \34249 );
xor \U$34247 ( \34625 , \34624 , \34266 );
and \U$34248 ( \34626 , \34622 , \34625 );
and \U$34249 ( \34627 , \34620 , \34625 );
or \U$34250 ( \34628 , \34623 , \34626 , \34627 );
xor \U$34251 ( \34629 , \34274 , \34276 );
xor \U$34252 ( \34630 , \34629 , \34279 );
xor \U$34253 ( \34631 , \34284 , \34286 );
xor \U$34254 ( \34632 , \34631 , \34289 );
and \U$34255 ( \34633 , \34630 , \34632 );
xor \U$34256 ( \34634 , \34295 , \34297 );
xor \U$34257 ( \34635 , \34634 , \34300 );
and \U$34258 ( \34636 , \34632 , \34635 );
and \U$34259 ( \34637 , \34630 , \34635 );
or \U$34260 ( \34638 , \34633 , \34636 , \34637 );
and \U$34261 ( \34639 , \34628 , \34638 );
xor \U$34262 ( \34640 , \33939 , \33955 );
xor \U$34263 ( \34641 , \34640 , \33972 );
and \U$34264 ( \34642 , \34638 , \34641 );
and \U$34265 ( \34643 , \34628 , \34641 );
or \U$34266 ( \34644 , \34639 , \34642 , \34643 );
and \U$34267 ( \34645 , \34618 , \34644 );
xor \U$34268 ( \34646 , \33891 , \33903 );
xor \U$34269 ( \34647 , \34646 , \33920 );
xor \U$34270 ( \34648 , \34309 , \34311 );
xor \U$34271 ( \34649 , \34648 , \34314 );
and \U$34272 ( \34650 , \34647 , \34649 );
xor \U$34273 ( \34651 , \34333 , \34335 );
xor \U$34274 ( \34652 , \34651 , \34338 );
and \U$34275 ( \34653 , \34649 , \34652 );
and \U$34276 ( \34654 , \34647 , \34652 );
or \U$34277 ( \34655 , \34650 , \34653 , \34654 );
and \U$34278 ( \34656 , \34644 , \34655 );
and \U$34279 ( \34657 , \34618 , \34655 );
or \U$34280 ( \34658 , \34645 , \34656 , \34657 );
xor \U$34281 ( \34659 , \34272 , \34306 );
xor \U$34282 ( \34660 , \34659 , \34317 );
xor \U$34283 ( \34661 , \34322 , \34324 );
xor \U$34284 ( \34662 , \34661 , \34327 );
and \U$34285 ( \34663 , \34660 , \34662 );
xor \U$34286 ( \34664 , \34341 , \34343 );
xor \U$34287 ( \34665 , \34664 , \34346 );
and \U$34288 ( \34666 , \34662 , \34665 );
and \U$34289 ( \34667 , \34660 , \34665 );
or \U$34290 ( \34668 , \34663 , \34666 , \34667 );
and \U$34291 ( \34669 , \34658 , \34668 );
xor \U$34292 ( \34670 , \34354 , \34356 );
xor \U$34293 ( \34671 , \34670 , \34359 );
and \U$34294 ( \34672 , \34668 , \34671 );
and \U$34295 ( \34673 , \34658 , \34671 );
or \U$34296 ( \34674 , \34669 , \34672 , \34673 );
xor \U$34297 ( \34675 , \34352 , \34362 );
xor \U$34298 ( \34676 , \34675 , \34365 );
and \U$34299 ( \34677 , \34674 , \34676 );
xor \U$34300 ( \34678 , \34370 , \34372 );
xor \U$34301 ( \34679 , \34678 , \34375 );
and \U$34302 ( \34680 , \34676 , \34679 );
and \U$34303 ( \34681 , \34674 , \34679 );
or \U$34304 ( \34682 , \34677 , \34680 , \34681 );
xor \U$34305 ( \34683 , \34368 , \34378 );
xor \U$34306 ( \34684 , \34683 , \34381 );
and \U$34307 ( \34685 , \34682 , \34684 );
xor \U$34308 ( \34686 , \34077 , \34087 );
xor \U$34309 ( \34687 , \34686 , \34090 );
and \U$34310 ( \34688 , \34684 , \34687 );
and \U$34311 ( \34689 , \34682 , \34687 );
or \U$34312 ( \34690 , \34685 , \34688 , \34689 );
and \U$34313 ( \34691 , \34390 , \34690 );
xor \U$34314 ( \34692 , \34390 , \34690 );
xor \U$34315 ( \34693 , \34682 , \34684 );
xor \U$34316 ( \34694 , \34693 , \34687 );
xor \U$34317 ( \34695 , \34444 , \34448 );
xor \U$34318 ( \34696 , \34695 , \34453 );
xor \U$34319 ( \34697 , \34460 , \34464 );
xor \U$34320 ( \34698 , \34697 , \34469 );
and \U$34321 ( \34699 , \34696 , \34698 );
xor \U$34322 ( \34700 , \34508 , \34512 );
xor \U$34323 ( \34701 , \34700 , \34517 );
and \U$34324 ( \34702 , \34698 , \34701 );
and \U$34325 ( \34703 , \34696 , \34701 );
or \U$34326 ( \34704 , \34699 , \34702 , \34703 );
xor \U$34327 ( \34705 , \34492 , \34496 );
xor \U$34328 ( \34706 , \34705 , \34501 );
xor \U$34329 ( \34707 , \34525 , \34529 );
xor \U$34330 ( \34708 , \34707 , \34534 );
and \U$34331 ( \34709 , \34706 , \34708 );
xor \U$34332 ( \34710 , \34578 , \34582 );
xor \U$34333 ( \34711 , \34710 , \34587 );
and \U$34334 ( \34712 , \34708 , \34711 );
and \U$34335 ( \34713 , \34706 , \34711 );
or \U$34336 ( \34714 , \34709 , \34712 , \34713 );
and \U$34337 ( \34715 , \34704 , \34714 );
xor \U$34338 ( \34716 , \34545 , \34549 );
xor \U$34339 ( \34717 , \34716 , \34554 );
xor \U$34340 ( \34718 , \34394 , \34398 );
xor \U$34341 ( \34719 , \34718 , \34401 );
and \U$34342 ( \34720 , \34717 , \34719 );
xor \U$34343 ( \34721 , \34561 , \34565 );
xor \U$34344 ( \34722 , \34721 , \34570 );
and \U$34345 ( \34723 , \34719 , \34722 );
and \U$34346 ( \34724 , \34717 , \34722 );
or \U$34347 ( \34725 , \34720 , \34723 , \34724 );
and \U$34348 ( \34726 , \34714 , \34725 );
and \U$34349 ( \34727 , \34704 , \34725 );
or \U$34350 ( \34728 , \34715 , \34726 , \34727 );
and \U$34351 ( \34729 , \23714 , \26983 );
and \U$34352 ( \34730 , \23570 , \26981 );
nor \U$34353 ( \34731 , \34729 , \34730 );
xnor \U$34354 ( \34732 , \34731 , \26742 );
and \U$34355 ( \34733 , \24003 , \26517 );
and \U$34356 ( \34734 , \23978 , \26515 );
nor \U$34357 ( \34735 , \34733 , \34734 );
xnor \U$34358 ( \34736 , \34735 , \26329 );
and \U$34359 ( \34737 , \34732 , \34736 );
and \U$34360 ( \34738 , \24344 , \26143 );
and \U$34361 ( \34739 , \24177 , \26141 );
nor \U$34362 ( \34740 , \34738 , \34739 );
xnor \U$34363 ( \34741 , \34740 , \25911 );
and \U$34364 ( \34742 , \34736 , \34741 );
and \U$34365 ( \34743 , \34732 , \34741 );
or \U$34366 ( \34744 , \34737 , \34742 , \34743 );
and \U$34367 ( \34745 , \25806 , \24661 );
and \U$34368 ( \34746 , \25609 , \24659 );
nor \U$34369 ( \34747 , \34745 , \34746 );
xnor \U$34370 ( \34748 , \34747 , \24456 );
and \U$34371 ( \34749 , \26116 , \24255 );
and \U$34372 ( \34750 , \26108 , \24253 );
nor \U$34373 ( \34751 , \34749 , \34750 );
xnor \U$34374 ( \34752 , \34751 , \24106 );
and \U$34375 ( \34753 , \34748 , \34752 );
and \U$34376 ( \34754 , \26590 , \23933 );
and \U$34377 ( \34755 , \26585 , \23931 );
nor \U$34378 ( \34756 , \34754 , \34755 );
xnor \U$34379 ( \34757 , \34756 , \23791 );
and \U$34380 ( \34758 , \34752 , \34757 );
and \U$34381 ( \34759 , \34748 , \34757 );
or \U$34382 ( \34760 , \34753 , \34758 , \34759 );
and \U$34383 ( \34761 , \34744 , \34760 );
and \U$34384 ( \34762 , \24601 , \25692 );
and \U$34385 ( \34763 , \24482 , \25690 );
nor \U$34386 ( \34764 , \34762 , \34763 );
xnor \U$34387 ( \34765 , \34764 , \25549 );
and \U$34388 ( \34766 , \25226 , \25369 );
and \U$34389 ( \34767 , \25018 , \25367 );
nor \U$34390 ( \34768 , \34766 , \34767 );
xnor \U$34391 ( \34769 , \34768 , \25123 );
and \U$34392 ( \34770 , \34765 , \34769 );
and \U$34393 ( \34771 , \25353 , \24974 );
and \U$34394 ( \34772 , \25348 , \24972 );
nor \U$34395 ( \34773 , \34771 , \34772 );
xnor \U$34396 ( \34774 , \34773 , \24787 );
and \U$34397 ( \34775 , \34769 , \34774 );
and \U$34398 ( \34776 , \34765 , \34774 );
or \U$34399 ( \34777 , \34770 , \34775 , \34776 );
and \U$34400 ( \34778 , \34760 , \34777 );
and \U$34401 ( \34779 , \34744 , \34777 );
or \U$34402 ( \34780 , \34761 , \34778 , \34779 );
and \U$34403 ( \34781 , \30318 , \22333 );
and \U$34404 ( \34782 , \30034 , \22331 );
nor \U$34405 ( \34783 , \34781 , \34782 );
xnor \U$34406 ( \34784 , \34783 , \22239 );
and \U$34407 ( \34785 , \30895 , \22163 );
and \U$34408 ( \34786 , \30887 , \22161 );
nor \U$34409 ( \34787 , \34785 , \34786 );
xnor \U$34410 ( \34788 , \34787 , \22091 );
and \U$34411 ( \34789 , \34784 , \34788 );
and \U$34412 ( \34790 , \31503 , \22029 );
and \U$34413 ( \34791 , \31498 , \22027 );
nor \U$34414 ( \34792 , \34790 , \34791 );
xnor \U$34415 ( \34793 , \34792 , \21986 );
and \U$34416 ( \34794 , \34788 , \34793 );
and \U$34417 ( \34795 , \34784 , \34793 );
or \U$34418 ( \34796 , \34789 , \34794 , \34795 );
and \U$34419 ( \34797 , \28514 , \22891 );
and \U$34420 ( \34798 , \28342 , \22889 );
nor \U$34421 ( \34799 , \34797 , \34798 );
xnor \U$34422 ( \34800 , \34799 , \22778 );
and \U$34423 ( \34801 , \29464 , \22697 );
and \U$34424 ( \34802 , \29040 , \22695 );
nor \U$34425 ( \34803 , \34801 , \34802 );
xnor \U$34426 ( \34804 , \34803 , \22561 );
and \U$34427 ( \34805 , \34800 , \34804 );
and \U$34428 ( \34806 , \29715 , \22497 );
and \U$34429 ( \34807 , \29710 , \22495 );
nor \U$34430 ( \34808 , \34806 , \34807 );
xnor \U$34431 ( \34809 , \34808 , \22419 );
and \U$34432 ( \34810 , \34804 , \34809 );
and \U$34433 ( \34811 , \34800 , \34809 );
or \U$34434 ( \34812 , \34805 , \34810 , \34811 );
and \U$34435 ( \34813 , \34796 , \34812 );
and \U$34436 ( \34814 , \27113 , \23637 );
and \U$34437 ( \34815 , \26854 , \23635 );
nor \U$34438 ( \34816 , \34814 , \34815 );
xnor \U$34439 ( \34817 , \34816 , \23500 );
and \U$34440 ( \34818 , \27494 , \23431 );
and \U$34441 ( \34819 , \27485 , \23429 );
nor \U$34442 ( \34820 , \34818 , \34819 );
xnor \U$34443 ( \34821 , \34820 , \23279 );
and \U$34444 ( \34822 , \34817 , \34821 );
and \U$34445 ( \34823 , \28039 , \23163 );
and \U$34446 ( \34824 , \27837 , \23161 );
nor \U$34447 ( \34825 , \34823 , \34824 );
xnor \U$34448 ( \34826 , \34825 , \23007 );
and \U$34449 ( \34827 , \34821 , \34826 );
and \U$34450 ( \34828 , \34817 , \34826 );
or \U$34451 ( \34829 , \34822 , \34827 , \34828 );
and \U$34452 ( \34830 , \34812 , \34829 );
and \U$34453 ( \34831 , \34796 , \34829 );
or \U$34454 ( \34832 , \34813 , \34830 , \34831 );
and \U$34455 ( \34833 , \34780 , \34832 );
and \U$34456 ( \34834 , \22952 , \28575 );
and \U$34457 ( \34835 , \22837 , \28573 );
nor \U$34458 ( \34836 , \34834 , \34835 );
xnor \U$34459 ( \34837 , \34836 , \28315 );
and \U$34460 ( \34838 , \23136 , \28081 );
and \U$34461 ( \34839 , \23128 , \28079 );
nor \U$34462 ( \34840 , \34838 , \34839 );
xnor \U$34463 ( \34841 , \34840 , \27766 );
and \U$34464 ( \34842 , \34837 , \34841 );
and \U$34465 ( \34843 , \23384 , \27572 );
and \U$34466 ( \34844 , \23379 , \27570 );
nor \U$34467 ( \34845 , \34843 , \34844 );
xnor \U$34468 ( \34846 , \34845 , \27232 );
and \U$34469 ( \34847 , \34841 , \34846 );
and \U$34470 ( \34848 , \34837 , \34846 );
or \U$34471 ( \34849 , \34842 , \34847 , \34848 );
and \U$34472 ( \34850 , \21941 , \32151 );
and \U$34473 ( \34851 , \21890 , \32148 );
nor \U$34474 ( \34852 , \34850 , \34851 );
xnor \U$34475 ( \34853 , \34852 , \31096 );
and \U$34476 ( \34854 , \22046 , \31338 );
and \U$34477 ( \34855 , \22018 , \31336 );
nor \U$34478 ( \34856 , \34854 , \34855 );
xnor \U$34479 ( \34857 , \34856 , \31099 );
and \U$34480 ( \34858 , \34853 , \34857 );
and \U$34481 ( \34859 , \22200 , \30770 );
and \U$34482 ( \34860 , \22126 , \30768 );
nor \U$34483 ( \34861 , \34859 , \34860 );
xnor \U$34484 ( \34862 , \34861 , \30460 );
and \U$34485 ( \34863 , \34857 , \34862 );
and \U$34486 ( \34864 , \34853 , \34862 );
or \U$34487 ( \34865 , \34858 , \34863 , \34864 );
and \U$34488 ( \34866 , \34849 , \34865 );
and \U$34489 ( \34867 , \22325 , \30233 );
and \U$34490 ( \34868 , \22262 , \30231 );
nor \U$34491 ( \34869 , \34867 , \34868 );
xnor \U$34492 ( \34870 , \34869 , \29862 );
and \U$34493 ( \34871 , \22611 , \29671 );
and \U$34494 ( \34872 , \22523 , \29669 );
nor \U$34495 ( \34873 , \34871 , \34872 );
xnor \U$34496 ( \34874 , \34873 , \29353 );
and \U$34497 ( \34875 , \34870 , \34874 );
and \U$34498 ( \34876 , \22721 , \29104 );
and \U$34499 ( \34877 , \22716 , \29102 );
nor \U$34500 ( \34878 , \34876 , \34877 );
xnor \U$34501 ( \34879 , \34878 , \28855 );
and \U$34502 ( \34880 , \34874 , \34879 );
and \U$34503 ( \34881 , \34870 , \34879 );
or \U$34504 ( \34882 , \34875 , \34880 , \34881 );
and \U$34505 ( \34883 , \34865 , \34882 );
and \U$34506 ( \34884 , \34849 , \34882 );
or \U$34507 ( \34885 , \34866 , \34883 , \34884 );
and \U$34508 ( \34886 , \34832 , \34885 );
and \U$34509 ( \34887 , \34780 , \34885 );
or \U$34510 ( \34888 , \34833 , \34886 , \34887 );
and \U$34511 ( \34889 , \34728 , \34888 );
xor \U$34512 ( \34890 , \34418 , \34420 );
xor \U$34513 ( \34891 , \34890 , \34423 );
xor \U$34514 ( \34892 , \34599 , \34601 );
xor \U$34515 ( \34893 , \34892 , \34604 );
and \U$34516 ( \34894 , \34891 , \34893 );
xor \U$34517 ( \34895 , \34429 , \34431 );
xor \U$34518 ( \34896 , \34895 , \34434 );
and \U$34519 ( \34897 , \34893 , \34896 );
and \U$34520 ( \34898 , \34891 , \34896 );
or \U$34521 ( \34899 , \34894 , \34897 , \34898 );
and \U$34522 ( \34900 , \34888 , \34899 );
and \U$34523 ( \34901 , \34728 , \34899 );
or \U$34524 ( \34902 , \34889 , \34900 , \34901 );
xor \U$34525 ( \34903 , \34416 , \34426 );
xor \U$34526 ( \34904 , \34903 , \34437 );
xor \U$34527 ( \34905 , \34488 , \34540 );
xor \U$34528 ( \34906 , \34905 , \34593 );
and \U$34529 ( \34907 , \34904 , \34906 );
xor \U$34530 ( \34908 , \34607 , \34609 );
xor \U$34531 ( \34909 , \34908 , \34612 );
and \U$34532 ( \34910 , \34906 , \34909 );
and \U$34533 ( \34911 , \34904 , \34909 );
or \U$34534 ( \34912 , \34907 , \34910 , \34911 );
and \U$34535 ( \34913 , \34902 , \34912 );
xor \U$34536 ( \34914 , \34404 , \34408 );
xor \U$34537 ( \34915 , \34914 , \34413 );
xor \U$34538 ( \34916 , \34504 , \34520 );
xor \U$34539 ( \34917 , \34916 , \34537 );
and \U$34540 ( \34918 , \34915 , \34917 );
xor \U$34541 ( \34919 , \34557 , \34573 );
xor \U$34542 ( \34920 , \34919 , \34590 );
and \U$34543 ( \34921 , \34917 , \34920 );
and \U$34544 ( \34922 , \34915 , \34920 );
or \U$34545 ( \34923 , \34918 , \34921 , \34922 );
xor \U$34546 ( \34924 , \34620 , \34622 );
xor \U$34547 ( \34925 , \34924 , \34625 );
and \U$34548 ( \34926 , \34923 , \34925 );
xor \U$34549 ( \34927 , \34630 , \34632 );
xor \U$34550 ( \34928 , \34927 , \34635 );
and \U$34551 ( \34929 , \34925 , \34928 );
and \U$34552 ( \34930 , \34923 , \34928 );
or \U$34553 ( \34931 , \34926 , \34929 , \34930 );
and \U$34554 ( \34932 , \34912 , \34931 );
and \U$34555 ( \34933 , \34902 , \34931 );
or \U$34556 ( \34934 , \34913 , \34932 , \34933 );
xor \U$34557 ( \34935 , \34164 , \34216 );
xor \U$34558 ( \34936 , \34935 , \34269 );
xor \U$34559 ( \34937 , \34282 , \34292 );
xor \U$34560 ( \34938 , \34937 , \34303 );
and \U$34561 ( \34939 , \34936 , \34938 );
xor \U$34562 ( \34940 , \34647 , \34649 );
xor \U$34563 ( \34941 , \34940 , \34652 );
and \U$34564 ( \34942 , \34938 , \34941 );
and \U$34565 ( \34943 , \34936 , \34941 );
or \U$34566 ( \34944 , \34939 , \34942 , \34943 );
and \U$34567 ( \34945 , \34934 , \34944 );
xor \U$34568 ( \34946 , \34660 , \34662 );
xor \U$34569 ( \34947 , \34946 , \34665 );
and \U$34570 ( \34948 , \34944 , \34947 );
and \U$34571 ( \34949 , \34934 , \34947 );
or \U$34572 ( \34950 , \34945 , \34948 , \34949 );
xor \U$34573 ( \34951 , \34320 , \34330 );
xor \U$34574 ( \34952 , \34951 , \34349 );
and \U$34575 ( \34953 , \34950 , \34952 );
xor \U$34576 ( \34954 , \34658 , \34668 );
xor \U$34577 ( \34955 , \34954 , \34671 );
and \U$34578 ( \34956 , \34952 , \34955 );
and \U$34579 ( \34957 , \34950 , \34955 );
or \U$34580 ( \34958 , \34953 , \34956 , \34957 );
xor \U$34581 ( \34959 , \34674 , \34676 );
xor \U$34582 ( \34960 , \34959 , \34679 );
and \U$34583 ( \34961 , \34958 , \34960 );
and \U$34584 ( \34962 , \34694 , \34961 );
xor \U$34585 ( \34963 , \34694 , \34961 );
xor \U$34586 ( \34964 , \34958 , \34960 );
xor \U$34587 ( \34965 , \34748 , \34752 );
xor \U$34588 ( \34966 , \34965 , \34757 );
xor \U$34589 ( \34967 , \34765 , \34769 );
xor \U$34590 ( \34968 , \34967 , \34774 );
and \U$34591 ( \34969 , \34966 , \34968 );
xor \U$34592 ( \34970 , \34817 , \34821 );
xor \U$34593 ( \34971 , \34970 , \34826 );
and \U$34594 ( \34972 , \34968 , \34971 );
and \U$34595 ( \34973 , \34966 , \34971 );
or \U$34596 ( \34974 , \34969 , \34972 , \34973 );
xor \U$34597 ( \34975 , \34732 , \34736 );
xor \U$34598 ( \34976 , \34975 , \34741 );
xor \U$34599 ( \34977 , \34837 , \34841 );
xor \U$34600 ( \34978 , \34977 , \34846 );
and \U$34601 ( \34979 , \34976 , \34978 );
xor \U$34602 ( \34980 , \34870 , \34874 );
xor \U$34603 ( \34981 , \34980 , \34879 );
and \U$34604 ( \34982 , \34978 , \34981 );
and \U$34605 ( \34983 , \34976 , \34981 );
or \U$34606 ( \34984 , \34979 , \34982 , \34983 );
and \U$34607 ( \34985 , \34974 , \34984 );
and \U$34608 ( \34986 , \32304 , \21916 );
and \U$34609 ( \34987 , \31684 , \21914 );
nor \U$34610 ( \34988 , \34986 , \34987 );
xnor \U$34611 ( \34989 , \34988 , \21867 );
xor \U$34612 ( \34990 , \34784 , \34788 );
xor \U$34613 ( \34991 , \34990 , \34793 );
and \U$34614 ( \34992 , \34989 , \34991 );
xor \U$34615 ( \34993 , \34800 , \34804 );
xor \U$34616 ( \34994 , \34993 , \34809 );
and \U$34617 ( \34995 , \34991 , \34994 );
and \U$34618 ( \34996 , \34989 , \34994 );
or \U$34619 ( \34997 , \34992 , \34995 , \34996 );
and \U$34620 ( \34998 , \34984 , \34997 );
and \U$34621 ( \34999 , \34974 , \34997 );
or \U$34622 ( \35000 , \34985 , \34998 , \34999 );
and \U$34623 ( \35001 , \22837 , \29104 );
and \U$34624 ( \35002 , \22721 , \29102 );
nor \U$34625 ( \35003 , \35001 , \35002 );
xnor \U$34626 ( \35004 , \35003 , \28855 );
and \U$34627 ( \35005 , \23128 , \28575 );
and \U$34628 ( \35006 , \22952 , \28573 );
nor \U$34629 ( \35007 , \35005 , \35006 );
xnor \U$34630 ( \35008 , \35007 , \28315 );
and \U$34631 ( \35009 , \35004 , \35008 );
and \U$34632 ( \35010 , \23379 , \28081 );
and \U$34633 ( \35011 , \23136 , \28079 );
nor \U$34634 ( \35012 , \35010 , \35011 );
xnor \U$34635 ( \35013 , \35012 , \27766 );
and \U$34636 ( \35014 , \35008 , \35013 );
and \U$34637 ( \35015 , \35004 , \35013 );
or \U$34638 ( \35016 , \35009 , \35014 , \35015 );
and \U$34639 ( \35017 , \22262 , \30770 );
and \U$34640 ( \35018 , \22200 , \30768 );
nor \U$34641 ( \35019 , \35017 , \35018 );
xnor \U$34642 ( \35020 , \35019 , \30460 );
and \U$34643 ( \35021 , \22523 , \30233 );
and \U$34644 ( \35022 , \22325 , \30231 );
nor \U$34645 ( \35023 , \35021 , \35022 );
xnor \U$34646 ( \35024 , \35023 , \29862 );
and \U$34647 ( \35025 , \35020 , \35024 );
and \U$34648 ( \35026 , \22716 , \29671 );
and \U$34649 ( \35027 , \22611 , \29669 );
nor \U$34650 ( \35028 , \35026 , \35027 );
xnor \U$34651 ( \35029 , \35028 , \29353 );
and \U$34652 ( \35030 , \35024 , \35029 );
and \U$34653 ( \35031 , \35020 , \35029 );
or \U$34654 ( \35032 , \35025 , \35030 , \35031 );
and \U$34655 ( \35033 , \35016 , \35032 );
and \U$34656 ( \35034 , \22018 , \32151 );
and \U$34657 ( \35035 , \21941 , \32148 );
nor \U$34658 ( \35036 , \35034 , \35035 );
xnor \U$34659 ( \35037 , \35036 , \31096 );
and \U$34660 ( \35038 , \22126 , \31338 );
and \U$34661 ( \35039 , \22046 , \31336 );
nor \U$34662 ( \35040 , \35038 , \35039 );
xnor \U$34663 ( \35041 , \35040 , \31099 );
and \U$34664 ( \35042 , \35037 , \35041 );
and \U$34665 ( \35043 , \35041 , \21867 );
and \U$34666 ( \35044 , \35037 , \21867 );
or \U$34667 ( \35045 , \35042 , \35043 , \35044 );
and \U$34668 ( \35046 , \35032 , \35045 );
and \U$34669 ( \35047 , \35016 , \35045 );
or \U$34670 ( \35048 , \35033 , \35046 , \35047 );
and \U$34671 ( \35049 , \30034 , \22497 );
and \U$34672 ( \35050 , \29715 , \22495 );
nor \U$34673 ( \35051 , \35049 , \35050 );
xnor \U$34674 ( \35052 , \35051 , \22419 );
and \U$34675 ( \35053 , \30887 , \22333 );
and \U$34676 ( \35054 , \30318 , \22331 );
nor \U$34677 ( \35055 , \35053 , \35054 );
xnor \U$34678 ( \35056 , \35055 , \22239 );
and \U$34679 ( \35057 , \35052 , \35056 );
and \U$34680 ( \35058 , \31498 , \22163 );
and \U$34681 ( \35059 , \30895 , \22161 );
nor \U$34682 ( \35060 , \35058 , \35059 );
xnor \U$34683 ( \35061 , \35060 , \22091 );
and \U$34684 ( \35062 , \35056 , \35061 );
and \U$34685 ( \35063 , \35052 , \35061 );
or \U$34686 ( \35064 , \35057 , \35062 , \35063 );
and \U$34687 ( \35065 , \26854 , \23933 );
and \U$34688 ( \35066 , \26590 , \23931 );
nor \U$34689 ( \35067 , \35065 , \35066 );
xnor \U$34690 ( \35068 , \35067 , \23791 );
and \U$34691 ( \35069 , \27485 , \23637 );
and \U$34692 ( \35070 , \27113 , \23635 );
nor \U$34693 ( \35071 , \35069 , \35070 );
xnor \U$34694 ( \35072 , \35071 , \23500 );
and \U$34695 ( \35073 , \35068 , \35072 );
and \U$34696 ( \35074 , \27837 , \23431 );
and \U$34697 ( \35075 , \27494 , \23429 );
nor \U$34698 ( \35076 , \35074 , \35075 );
xnor \U$34699 ( \35077 , \35076 , \23279 );
and \U$34700 ( \35078 , \35072 , \35077 );
and \U$34701 ( \35079 , \35068 , \35077 );
or \U$34702 ( \35080 , \35073 , \35078 , \35079 );
and \U$34703 ( \35081 , \35064 , \35080 );
and \U$34704 ( \35082 , \28342 , \23163 );
and \U$34705 ( \35083 , \28039 , \23161 );
nor \U$34706 ( \35084 , \35082 , \35083 );
xnor \U$34707 ( \35085 , \35084 , \23007 );
and \U$34708 ( \35086 , \29040 , \22891 );
and \U$34709 ( \35087 , \28514 , \22889 );
nor \U$34710 ( \35088 , \35086 , \35087 );
xnor \U$34711 ( \35089 , \35088 , \22778 );
and \U$34712 ( \35090 , \35085 , \35089 );
and \U$34713 ( \35091 , \29710 , \22697 );
and \U$34714 ( \35092 , \29464 , \22695 );
nor \U$34715 ( \35093 , \35091 , \35092 );
xnor \U$34716 ( \35094 , \35093 , \22561 );
and \U$34717 ( \35095 , \35089 , \35094 );
and \U$34718 ( \35096 , \35085 , \35094 );
or \U$34719 ( \35097 , \35090 , \35095 , \35096 );
and \U$34720 ( \35098 , \35080 , \35097 );
and \U$34721 ( \35099 , \35064 , \35097 );
or \U$34722 ( \35100 , \35081 , \35098 , \35099 );
and \U$34723 ( \35101 , \35048 , \35100 );
and \U$34724 ( \35102 , \25609 , \24974 );
and \U$34725 ( \35103 , \25353 , \24972 );
nor \U$34726 ( \35104 , \35102 , \35103 );
xnor \U$34727 ( \35105 , \35104 , \24787 );
and \U$34728 ( \35106 , \26108 , \24661 );
and \U$34729 ( \35107 , \25806 , \24659 );
nor \U$34730 ( \35108 , \35106 , \35107 );
xnor \U$34731 ( \35109 , \35108 , \24456 );
and \U$34732 ( \35110 , \35105 , \35109 );
and \U$34733 ( \35111 , \26585 , \24255 );
and \U$34734 ( \35112 , \26116 , \24253 );
nor \U$34735 ( \35113 , \35111 , \35112 );
xnor \U$34736 ( \35114 , \35113 , \24106 );
and \U$34737 ( \35115 , \35109 , \35114 );
and \U$34738 ( \35116 , \35105 , \35114 );
or \U$34739 ( \35117 , \35110 , \35115 , \35116 );
and \U$34740 ( \35118 , \24482 , \26143 );
and \U$34741 ( \35119 , \24344 , \26141 );
nor \U$34742 ( \35120 , \35118 , \35119 );
xnor \U$34743 ( \35121 , \35120 , \25911 );
and \U$34744 ( \35122 , \25018 , \25692 );
and \U$34745 ( \35123 , \24601 , \25690 );
nor \U$34746 ( \35124 , \35122 , \35123 );
xnor \U$34747 ( \35125 , \35124 , \25549 );
and \U$34748 ( \35126 , \35121 , \35125 );
and \U$34749 ( \35127 , \25348 , \25369 );
and \U$34750 ( \35128 , \25226 , \25367 );
nor \U$34751 ( \35129 , \35127 , \35128 );
xnor \U$34752 ( \35130 , \35129 , \25123 );
and \U$34753 ( \35131 , \35125 , \35130 );
and \U$34754 ( \35132 , \35121 , \35130 );
or \U$34755 ( \35133 , \35126 , \35131 , \35132 );
and \U$34756 ( \35134 , \35117 , \35133 );
and \U$34757 ( \35135 , \23570 , \27572 );
and \U$34758 ( \35136 , \23384 , \27570 );
nor \U$34759 ( \35137 , \35135 , \35136 );
xnor \U$34760 ( \35138 , \35137 , \27232 );
and \U$34761 ( \35139 , \23978 , \26983 );
and \U$34762 ( \35140 , \23714 , \26981 );
nor \U$34763 ( \35141 , \35139 , \35140 );
xnor \U$34764 ( \35142 , \35141 , \26742 );
and \U$34765 ( \35143 , \35138 , \35142 );
and \U$34766 ( \35144 , \24177 , \26517 );
and \U$34767 ( \35145 , \24003 , \26515 );
nor \U$34768 ( \35146 , \35144 , \35145 );
xnor \U$34769 ( \35147 , \35146 , \26329 );
and \U$34770 ( \35148 , \35142 , \35147 );
and \U$34771 ( \35149 , \35138 , \35147 );
or \U$34772 ( \35150 , \35143 , \35148 , \35149 );
and \U$34773 ( \35151 , \35133 , \35150 );
and \U$34774 ( \35152 , \35117 , \35150 );
or \U$34775 ( \35153 , \35134 , \35151 , \35152 );
and \U$34776 ( \35154 , \35100 , \35153 );
and \U$34777 ( \35155 , \35048 , \35153 );
or \U$34778 ( \35156 , \35101 , \35154 , \35155 );
and \U$34779 ( \35157 , \35000 , \35156 );
xor \U$34780 ( \35158 , \34477 , \34481 );
xor \U$34781 ( \35159 , \35158 , \21774 );
xor \U$34782 ( \35160 , \34696 , \34698 );
xor \U$34783 ( \35161 , \35160 , \34701 );
and \U$34784 ( \35162 , \35159 , \35161 );
xor \U$34785 ( \35163 , \34706 , \34708 );
xor \U$34786 ( \35164 , \35163 , \34711 );
and \U$34787 ( \35165 , \35161 , \35164 );
and \U$34788 ( \35166 , \35159 , \35164 );
or \U$34789 ( \35167 , \35162 , \35165 , \35166 );
and \U$34790 ( \35168 , \35156 , \35167 );
and \U$34791 ( \35169 , \35000 , \35167 );
or \U$34792 ( \35170 , \35157 , \35168 , \35169 );
xor \U$34793 ( \35171 , \34744 , \34760 );
xor \U$34794 ( \35172 , \35171 , \34777 );
xor \U$34795 ( \35173 , \34796 , \34812 );
xor \U$34796 ( \35174 , \35173 , \34829 );
and \U$34797 ( \35175 , \35172 , \35174 );
xor \U$34798 ( \35176 , \34717 , \34719 );
xor \U$34799 ( \35177 , \35176 , \34722 );
and \U$34800 ( \35178 , \35174 , \35177 );
and \U$34801 ( \35179 , \35172 , \35177 );
or \U$34802 ( \35180 , \35175 , \35178 , \35179 );
xor \U$34803 ( \35181 , \34456 , \34472 );
xor \U$34804 ( \35182 , \35181 , \34485 );
and \U$34805 ( \35183 , \35180 , \35182 );
xor \U$34806 ( \35184 , \34915 , \34917 );
xor \U$34807 ( \35185 , \35184 , \34920 );
and \U$34808 ( \35186 , \35182 , \35185 );
and \U$34809 ( \35187 , \35180 , \35185 );
or \U$34810 ( \35188 , \35183 , \35186 , \35187 );
and \U$34811 ( \35189 , \35170 , \35188 );
xor \U$34812 ( \35190 , \34704 , \34714 );
xor \U$34813 ( \35191 , \35190 , \34725 );
xor \U$34814 ( \35192 , \34780 , \34832 );
xor \U$34815 ( \35193 , \35192 , \34885 );
and \U$34816 ( \35194 , \35191 , \35193 );
xor \U$34817 ( \35195 , \34891 , \34893 );
xor \U$34818 ( \35196 , \35195 , \34896 );
and \U$34819 ( \35197 , \35193 , \35196 );
and \U$34820 ( \35198 , \35191 , \35196 );
or \U$34821 ( \35199 , \35194 , \35197 , \35198 );
and \U$34822 ( \35200 , \35188 , \35199 );
and \U$34823 ( \35201 , \35170 , \35199 );
or \U$34824 ( \35202 , \35189 , \35200 , \35201 );
xor \U$34825 ( \35203 , \34728 , \34888 );
xor \U$34826 ( \35204 , \35203 , \34899 );
xor \U$34827 ( \35205 , \34904 , \34906 );
xor \U$34828 ( \35206 , \35205 , \34909 );
and \U$34829 ( \35207 , \35204 , \35206 );
xor \U$34830 ( \35208 , \34923 , \34925 );
xor \U$34831 ( \35209 , \35208 , \34928 );
and \U$34832 ( \35210 , \35206 , \35209 );
and \U$34833 ( \35211 , \35204 , \35209 );
or \U$34834 ( \35212 , \35207 , \35210 , \35211 );
and \U$34835 ( \35213 , \35202 , \35212 );
xor \U$34836 ( \35214 , \34628 , \34638 );
xor \U$34837 ( \35215 , \35214 , \34641 );
and \U$34838 ( \35216 , \35212 , \35215 );
and \U$34839 ( \35217 , \35202 , \35215 );
or \U$34840 ( \35218 , \35213 , \35216 , \35217 );
xor \U$34841 ( \35219 , \34440 , \34596 );
xor \U$34842 ( \35220 , \35219 , \34615 );
xor \U$34843 ( \35221 , \34902 , \34912 );
xor \U$34844 ( \35222 , \35221 , \34931 );
and \U$34845 ( \35223 , \35220 , \35222 );
xor \U$34846 ( \35224 , \34936 , \34938 );
xor \U$34847 ( \35225 , \35224 , \34941 );
and \U$34848 ( \35226 , \35222 , \35225 );
and \U$34849 ( \35227 , \35220 , \35225 );
or \U$34850 ( \35228 , \35223 , \35226 , \35227 );
and \U$34851 ( \35229 , \35218 , \35228 );
xor \U$34852 ( \35230 , \34618 , \34644 );
xor \U$34853 ( \35231 , \35230 , \34655 );
and \U$34854 ( \35232 , \35228 , \35231 );
and \U$34855 ( \35233 , \35218 , \35231 );
or \U$34856 ( \35234 , \35229 , \35232 , \35233 );
xor \U$34857 ( \35235 , \34950 , \34952 );
xor \U$34858 ( \35236 , \35235 , \34955 );
and \U$34859 ( \35237 , \35234 , \35236 );
and \U$34860 ( \35238 , \34964 , \35237 );
xor \U$34861 ( \35239 , \34964 , \35237 );
xor \U$34862 ( \35240 , \35234 , \35236 );
xor \U$34863 ( \35241 , \35105 , \35109 );
xor \U$34864 ( \35242 , \35241 , \35114 );
xor \U$34865 ( \35243 , \35068 , \35072 );
xor \U$34866 ( \35244 , \35243 , \35077 );
and \U$34867 ( \35245 , \35242 , \35244 );
xor \U$34868 ( \35246 , \35085 , \35089 );
xor \U$34869 ( \35247 , \35246 , \35094 );
and \U$34870 ( \35248 , \35244 , \35247 );
and \U$34871 ( \35249 , \35242 , \35247 );
or \U$34872 ( \35250 , \35245 , \35248 , \35249 );
and \U$34873 ( \35251 , \31684 , \22029 );
and \U$34874 ( \35252 , \31503 , \22027 );
nor \U$34875 ( \35253 , \35251 , \35252 );
xnor \U$34876 ( \35254 , \35253 , \21986 );
nand \U$34877 ( \35255 , \32304 , \21914 );
xnor \U$34878 ( \35256 , \35255 , \21867 );
and \U$34879 ( \35257 , \35254 , \35256 );
xor \U$34880 ( \35258 , \35052 , \35056 );
xor \U$34881 ( \35259 , \35258 , \35061 );
and \U$34882 ( \35260 , \35256 , \35259 );
and \U$34883 ( \35261 , \35254 , \35259 );
or \U$34884 ( \35262 , \35257 , \35260 , \35261 );
and \U$34885 ( \35263 , \35250 , \35262 );
xor \U$34886 ( \35264 , \35004 , \35008 );
xor \U$34887 ( \35265 , \35264 , \35013 );
xor \U$34888 ( \35266 , \35121 , \35125 );
xor \U$34889 ( \35267 , \35266 , \35130 );
and \U$34890 ( \35268 , \35265 , \35267 );
xor \U$34891 ( \35269 , \35138 , \35142 );
xor \U$34892 ( \35270 , \35269 , \35147 );
and \U$34893 ( \35271 , \35267 , \35270 );
and \U$34894 ( \35272 , \35265 , \35270 );
or \U$34895 ( \35273 , \35268 , \35271 , \35272 );
and \U$34896 ( \35274 , \35262 , \35273 );
and \U$34897 ( \35275 , \35250 , \35273 );
or \U$34898 ( \35276 , \35263 , \35274 , \35275 );
and \U$34899 ( \35277 , \30895 , \22333 );
and \U$34900 ( \35278 , \30887 , \22331 );
nor \U$34901 ( \35279 , \35277 , \35278 );
xnor \U$34902 ( \35280 , \35279 , \22239 );
and \U$34903 ( \35281 , \31503 , \22163 );
and \U$34904 ( \35282 , \31498 , \22161 );
nor \U$34905 ( \35283 , \35281 , \35282 );
xnor \U$34906 ( \35284 , \35283 , \22091 );
and \U$34907 ( \35285 , \35280 , \35284 );
and \U$34908 ( \35286 , \32304 , \22029 );
and \U$34909 ( \35287 , \31684 , \22027 );
nor \U$34910 ( \35288 , \35286 , \35287 );
xnor \U$34911 ( \35289 , \35288 , \21986 );
and \U$34912 ( \35290 , \35284 , \35289 );
and \U$34913 ( \35291 , \35280 , \35289 );
or \U$34914 ( \35292 , \35285 , \35290 , \35291 );
and \U$34915 ( \35293 , \27494 , \23637 );
and \U$34916 ( \35294 , \27485 , \23635 );
nor \U$34917 ( \35295 , \35293 , \35294 );
xnor \U$34918 ( \35296 , \35295 , \23500 );
and \U$34919 ( \35297 , \28039 , \23431 );
and \U$34920 ( \35298 , \27837 , \23429 );
nor \U$34921 ( \35299 , \35297 , \35298 );
xnor \U$34922 ( \35300 , \35299 , \23279 );
and \U$34923 ( \35301 , \35296 , \35300 );
and \U$34924 ( \35302 , \28514 , \23163 );
and \U$34925 ( \35303 , \28342 , \23161 );
nor \U$34926 ( \35304 , \35302 , \35303 );
xnor \U$34927 ( \35305 , \35304 , \23007 );
and \U$34928 ( \35306 , \35300 , \35305 );
and \U$34929 ( \35307 , \35296 , \35305 );
or \U$34930 ( \35308 , \35301 , \35306 , \35307 );
and \U$34931 ( \35309 , \35292 , \35308 );
and \U$34932 ( \35310 , \29464 , \22891 );
and \U$34933 ( \35311 , \29040 , \22889 );
nor \U$34934 ( \35312 , \35310 , \35311 );
xnor \U$34935 ( \35313 , \35312 , \22778 );
and \U$34936 ( \35314 , \29715 , \22697 );
and \U$34937 ( \35315 , \29710 , \22695 );
nor \U$34938 ( \35316 , \35314 , \35315 );
xnor \U$34939 ( \35317 , \35316 , \22561 );
and \U$34940 ( \35318 , \35313 , \35317 );
and \U$34941 ( \35319 , \30318 , \22497 );
and \U$34942 ( \35320 , \30034 , \22495 );
nor \U$34943 ( \35321 , \35319 , \35320 );
xnor \U$34944 ( \35322 , \35321 , \22419 );
and \U$34945 ( \35323 , \35317 , \35322 );
and \U$34946 ( \35324 , \35313 , \35322 );
or \U$34947 ( \35325 , \35318 , \35323 , \35324 );
and \U$34948 ( \35326 , \35308 , \35325 );
and \U$34949 ( \35327 , \35292 , \35325 );
or \U$34950 ( \35328 , \35309 , \35326 , \35327 );
and \U$34951 ( \35329 , \22611 , \30233 );
and \U$34952 ( \35330 , \22523 , \30231 );
nor \U$34953 ( \35331 , \35329 , \35330 );
xnor \U$34954 ( \35332 , \35331 , \29862 );
and \U$34955 ( \35333 , \22721 , \29671 );
and \U$34956 ( \35334 , \22716 , \29669 );
nor \U$34957 ( \35335 , \35333 , \35334 );
xnor \U$34958 ( \35336 , \35335 , \29353 );
and \U$34959 ( \35337 , \35332 , \35336 );
and \U$34960 ( \35338 , \22952 , \29104 );
and \U$34961 ( \35339 , \22837 , \29102 );
nor \U$34962 ( \35340 , \35338 , \35339 );
xnor \U$34963 ( \35341 , \35340 , \28855 );
and \U$34964 ( \35342 , \35336 , \35341 );
and \U$34965 ( \35343 , \35332 , \35341 );
or \U$34966 ( \35344 , \35337 , \35342 , \35343 );
and \U$34967 ( \35345 , \23136 , \28575 );
and \U$34968 ( \35346 , \23128 , \28573 );
nor \U$34969 ( \35347 , \35345 , \35346 );
xnor \U$34970 ( \35348 , \35347 , \28315 );
and \U$34971 ( \35349 , \23384 , \28081 );
and \U$34972 ( \35350 , \23379 , \28079 );
nor \U$34973 ( \35351 , \35349 , \35350 );
xnor \U$34974 ( \35352 , \35351 , \27766 );
and \U$34975 ( \35353 , \35348 , \35352 );
and \U$34976 ( \35354 , \23714 , \27572 );
and \U$34977 ( \35355 , \23570 , \27570 );
nor \U$34978 ( \35356 , \35354 , \35355 );
xnor \U$34979 ( \35357 , \35356 , \27232 );
and \U$34980 ( \35358 , \35352 , \35357 );
and \U$34981 ( \35359 , \35348 , \35357 );
or \U$34982 ( \35360 , \35353 , \35358 , \35359 );
and \U$34983 ( \35361 , \35344 , \35360 );
and \U$34984 ( \35362 , \22046 , \32151 );
and \U$34985 ( \35363 , \22018 , \32148 );
nor \U$34986 ( \35364 , \35362 , \35363 );
xnor \U$34987 ( \35365 , \35364 , \31096 );
and \U$34988 ( \35366 , \22200 , \31338 );
and \U$34989 ( \35367 , \22126 , \31336 );
nor \U$34990 ( \35368 , \35366 , \35367 );
xnor \U$34991 ( \35369 , \35368 , \31099 );
and \U$34992 ( \35370 , \35365 , \35369 );
and \U$34993 ( \35371 , \22325 , \30770 );
and \U$34994 ( \35372 , \22262 , \30768 );
nor \U$34995 ( \35373 , \35371 , \35372 );
xnor \U$34996 ( \35374 , \35373 , \30460 );
and \U$34997 ( \35375 , \35369 , \35374 );
and \U$34998 ( \35376 , \35365 , \35374 );
or \U$34999 ( \35377 , \35370 , \35375 , \35376 );
and \U$35000 ( \35378 , \35360 , \35377 );
and \U$35001 ( \35379 , \35344 , \35377 );
or \U$35002 ( \35380 , \35361 , \35378 , \35379 );
and \U$35003 ( \35381 , \35328 , \35380 );
and \U$35004 ( \35382 , \26116 , \24661 );
and \U$35005 ( \35383 , \26108 , \24659 );
nor \U$35006 ( \35384 , \35382 , \35383 );
xnor \U$35007 ( \35385 , \35384 , \24456 );
and \U$35008 ( \35386 , \26590 , \24255 );
and \U$35009 ( \35387 , \26585 , \24253 );
nor \U$35010 ( \35388 , \35386 , \35387 );
xnor \U$35011 ( \35389 , \35388 , \24106 );
and \U$35012 ( \35390 , \35385 , \35389 );
and \U$35013 ( \35391 , \27113 , \23933 );
and \U$35014 ( \35392 , \26854 , \23931 );
nor \U$35015 ( \35393 , \35391 , \35392 );
xnor \U$35016 ( \35394 , \35393 , \23791 );
and \U$35017 ( \35395 , \35389 , \35394 );
and \U$35018 ( \35396 , \35385 , \35394 );
or \U$35019 ( \35397 , \35390 , \35395 , \35396 );
and \U$35020 ( \35398 , \25226 , \25692 );
and \U$35021 ( \35399 , \25018 , \25690 );
nor \U$35022 ( \35400 , \35398 , \35399 );
xnor \U$35023 ( \35401 , \35400 , \25549 );
and \U$35024 ( \35402 , \25353 , \25369 );
and \U$35025 ( \35403 , \25348 , \25367 );
nor \U$35026 ( \35404 , \35402 , \35403 );
xnor \U$35027 ( \35405 , \35404 , \25123 );
and \U$35028 ( \35406 , \35401 , \35405 );
and \U$35029 ( \35407 , \25806 , \24974 );
and \U$35030 ( \35408 , \25609 , \24972 );
nor \U$35031 ( \35409 , \35407 , \35408 );
xnor \U$35032 ( \35410 , \35409 , \24787 );
and \U$35033 ( \35411 , \35405 , \35410 );
and \U$35034 ( \35412 , \35401 , \35410 );
or \U$35035 ( \35413 , \35406 , \35411 , \35412 );
and \U$35036 ( \35414 , \35397 , \35413 );
and \U$35037 ( \35415 , \24003 , \26983 );
and \U$35038 ( \35416 , \23978 , \26981 );
nor \U$35039 ( \35417 , \35415 , \35416 );
xnor \U$35040 ( \35418 , \35417 , \26742 );
and \U$35041 ( \35419 , \24344 , \26517 );
and \U$35042 ( \35420 , \24177 , \26515 );
nor \U$35043 ( \35421 , \35419 , \35420 );
xnor \U$35044 ( \35422 , \35421 , \26329 );
and \U$35045 ( \35423 , \35418 , \35422 );
and \U$35046 ( \35424 , \24601 , \26143 );
and \U$35047 ( \35425 , \24482 , \26141 );
nor \U$35048 ( \35426 , \35424 , \35425 );
xnor \U$35049 ( \35427 , \35426 , \25911 );
and \U$35050 ( \35428 , \35422 , \35427 );
and \U$35051 ( \35429 , \35418 , \35427 );
or \U$35052 ( \35430 , \35423 , \35428 , \35429 );
and \U$35053 ( \35431 , \35413 , \35430 );
and \U$35054 ( \35432 , \35397 , \35430 );
or \U$35055 ( \35433 , \35414 , \35431 , \35432 );
and \U$35056 ( \35434 , \35380 , \35433 );
and \U$35057 ( \35435 , \35328 , \35433 );
or \U$35058 ( \35436 , \35381 , \35434 , \35435 );
and \U$35059 ( \35437 , \35276 , \35436 );
xor \U$35060 ( \35438 , \34853 , \34857 );
xor \U$35061 ( \35439 , \35438 , \34862 );
xor \U$35062 ( \35440 , \34966 , \34968 );
xor \U$35063 ( \35441 , \35440 , \34971 );
and \U$35064 ( \35442 , \35439 , \35441 );
xor \U$35065 ( \35443 , \34976 , \34978 );
xor \U$35066 ( \35444 , \35443 , \34981 );
and \U$35067 ( \35445 , \35441 , \35444 );
and \U$35068 ( \35446 , \35439 , \35444 );
or \U$35069 ( \35447 , \35442 , \35445 , \35446 );
and \U$35070 ( \35448 , \35436 , \35447 );
and \U$35071 ( \35449 , \35276 , \35447 );
or \U$35072 ( \35450 , \35437 , \35448 , \35449 );
xor \U$35073 ( \35451 , \35064 , \35080 );
xor \U$35074 ( \35452 , \35451 , \35097 );
xor \U$35075 ( \35453 , \35117 , \35133 );
xor \U$35076 ( \35454 , \35453 , \35150 );
and \U$35077 ( \35455 , \35452 , \35454 );
xor \U$35078 ( \35456 , \34989 , \34991 );
xor \U$35079 ( \35457 , \35456 , \34994 );
and \U$35080 ( \35458 , \35454 , \35457 );
and \U$35081 ( \35459 , \35452 , \35457 );
or \U$35082 ( \35460 , \35455 , \35458 , \35459 );
xor \U$35083 ( \35461 , \34849 , \34865 );
xor \U$35084 ( \35462 , \35461 , \34882 );
and \U$35085 ( \35463 , \35460 , \35462 );
xor \U$35086 ( \35464 , \35172 , \35174 );
xor \U$35087 ( \35465 , \35464 , \35177 );
and \U$35088 ( \35466 , \35462 , \35465 );
and \U$35089 ( \35467 , \35460 , \35465 );
or \U$35090 ( \35468 , \35463 , \35466 , \35467 );
and \U$35091 ( \35469 , \35450 , \35468 );
xor \U$35092 ( \35470 , \34974 , \34984 );
xor \U$35093 ( \35471 , \35470 , \34997 );
xor \U$35094 ( \35472 , \35048 , \35100 );
xor \U$35095 ( \35473 , \35472 , \35153 );
and \U$35096 ( \35474 , \35471 , \35473 );
xor \U$35097 ( \35475 , \35159 , \35161 );
xor \U$35098 ( \35476 , \35475 , \35164 );
and \U$35099 ( \35477 , \35473 , \35476 );
and \U$35100 ( \35478 , \35471 , \35476 );
or \U$35101 ( \35479 , \35474 , \35477 , \35478 );
and \U$35102 ( \35480 , \35468 , \35479 );
and \U$35103 ( \35481 , \35450 , \35479 );
or \U$35104 ( \35482 , \35469 , \35480 , \35481 );
xor \U$35105 ( \35483 , \35000 , \35156 );
xor \U$35106 ( \35484 , \35483 , \35167 );
xor \U$35107 ( \35485 , \35180 , \35182 );
xor \U$35108 ( \35486 , \35485 , \35185 );
and \U$35109 ( \35487 , \35484 , \35486 );
xor \U$35110 ( \35488 , \35191 , \35193 );
xor \U$35111 ( \35489 , \35488 , \35196 );
and \U$35112 ( \35490 , \35486 , \35489 );
and \U$35113 ( \35491 , \35484 , \35489 );
or \U$35114 ( \35492 , \35487 , \35490 , \35491 );
and \U$35115 ( \35493 , \35482 , \35492 );
xor \U$35116 ( \35494 , \35204 , \35206 );
xor \U$35117 ( \35495 , \35494 , \35209 );
and \U$35118 ( \35496 , \35492 , \35495 );
and \U$35119 ( \35497 , \35482 , \35495 );
or \U$35120 ( \35498 , \35493 , \35496 , \35497 );
xor \U$35121 ( \35499 , \35202 , \35212 );
xor \U$35122 ( \35500 , \35499 , \35215 );
and \U$35123 ( \35501 , \35498 , \35500 );
xor \U$35124 ( \35502 , \35220 , \35222 );
xor \U$35125 ( \35503 , \35502 , \35225 );
and \U$35126 ( \35504 , \35500 , \35503 );
and \U$35127 ( \35505 , \35498 , \35503 );
or \U$35128 ( \35506 , \35501 , \35504 , \35505 );
xor \U$35129 ( \35507 , \35218 , \35228 );
xor \U$35130 ( \35508 , \35507 , \35231 );
and \U$35131 ( \35509 , \35506 , \35508 );
xor \U$35132 ( \35510 , \34934 , \34944 );
xor \U$35133 ( \35511 , \35510 , \34947 );
and \U$35134 ( \35512 , \35508 , \35511 );
and \U$35135 ( \35513 , \35506 , \35511 );
or \U$35136 ( \35514 , \35509 , \35512 , \35513 );
and \U$35137 ( \35515 , \35240 , \35514 );
xor \U$35138 ( \35516 , \35240 , \35514 );
xor \U$35139 ( \35517 , \35506 , \35508 );
xor \U$35140 ( \35518 , \35517 , \35511 );
xor \U$35141 ( \35519 , \35385 , \35389 );
xor \U$35142 ( \35520 , \35519 , \35394 );
xor \U$35143 ( \35521 , \35401 , \35405 );
xor \U$35144 ( \35522 , \35521 , \35410 );
and \U$35145 ( \35523 , \35520 , \35522 );
xor \U$35146 ( \35524 , \35418 , \35422 );
xor \U$35147 ( \35525 , \35524 , \35427 );
and \U$35148 ( \35526 , \35522 , \35525 );
and \U$35149 ( \35527 , \35520 , \35525 );
or \U$35150 ( \35528 , \35523 , \35526 , \35527 );
xor \U$35151 ( \35529 , \35280 , \35284 );
xor \U$35152 ( \35530 , \35529 , \35289 );
xor \U$35153 ( \35531 , \35296 , \35300 );
xor \U$35154 ( \35532 , \35531 , \35305 );
and \U$35155 ( \35533 , \35530 , \35532 );
xor \U$35156 ( \35534 , \35313 , \35317 );
xor \U$35157 ( \35535 , \35534 , \35322 );
and \U$35158 ( \35536 , \35532 , \35535 );
and \U$35159 ( \35537 , \35530 , \35535 );
or \U$35160 ( \35538 , \35533 , \35536 , \35537 );
and \U$35161 ( \35539 , \35528 , \35538 );
xor \U$35162 ( \35540 , \35332 , \35336 );
xor \U$35163 ( \35541 , \35540 , \35341 );
xor \U$35164 ( \35542 , \35348 , \35352 );
xor \U$35165 ( \35543 , \35542 , \35357 );
and \U$35166 ( \35544 , \35541 , \35543 );
xor \U$35167 ( \35545 , \35365 , \35369 );
xor \U$35168 ( \35546 , \35545 , \35374 );
and \U$35169 ( \35547 , \35543 , \35546 );
and \U$35170 ( \35548 , \35541 , \35546 );
or \U$35171 ( \35549 , \35544 , \35547 , \35548 );
and \U$35172 ( \35550 , \35538 , \35549 );
and \U$35173 ( \35551 , \35528 , \35549 );
or \U$35174 ( \35552 , \35539 , \35550 , \35551 );
and \U$35175 ( \35553 , \26108 , \24974 );
and \U$35176 ( \35554 , \25806 , \24972 );
nor \U$35177 ( \35555 , \35553 , \35554 );
xnor \U$35178 ( \35556 , \35555 , \24787 );
and \U$35179 ( \35557 , \26585 , \24661 );
and \U$35180 ( \35558 , \26116 , \24659 );
nor \U$35181 ( \35559 , \35557 , \35558 );
xnor \U$35182 ( \35560 , \35559 , \24456 );
and \U$35183 ( \35561 , \35556 , \35560 );
and \U$35184 ( \35562 , \26854 , \24255 );
and \U$35185 ( \35563 , \26590 , \24253 );
nor \U$35186 ( \35564 , \35562 , \35563 );
xnor \U$35187 ( \35565 , \35564 , \24106 );
and \U$35188 ( \35566 , \35560 , \35565 );
and \U$35189 ( \35567 , \35556 , \35565 );
or \U$35190 ( \35568 , \35561 , \35566 , \35567 );
and \U$35191 ( \35569 , \23978 , \27572 );
and \U$35192 ( \35570 , \23714 , \27570 );
nor \U$35193 ( \35571 , \35569 , \35570 );
xnor \U$35194 ( \35572 , \35571 , \27232 );
and \U$35195 ( \35573 , \24177 , \26983 );
and \U$35196 ( \35574 , \24003 , \26981 );
nor \U$35197 ( \35575 , \35573 , \35574 );
xnor \U$35198 ( \35576 , \35575 , \26742 );
and \U$35199 ( \35577 , \35572 , \35576 );
and \U$35200 ( \35578 , \24482 , \26517 );
and \U$35201 ( \35579 , \24344 , \26515 );
nor \U$35202 ( \35580 , \35578 , \35579 );
xnor \U$35203 ( \35581 , \35580 , \26329 );
and \U$35204 ( \35582 , \35576 , \35581 );
and \U$35205 ( \35583 , \35572 , \35581 );
or \U$35206 ( \35584 , \35577 , \35582 , \35583 );
and \U$35207 ( \35585 , \35568 , \35584 );
and \U$35208 ( \35586 , \25018 , \26143 );
and \U$35209 ( \35587 , \24601 , \26141 );
nor \U$35210 ( \35588 , \35586 , \35587 );
xnor \U$35211 ( \35589 , \35588 , \25911 );
and \U$35212 ( \35590 , \25348 , \25692 );
and \U$35213 ( \35591 , \25226 , \25690 );
nor \U$35214 ( \35592 , \35590 , \35591 );
xnor \U$35215 ( \35593 , \35592 , \25549 );
and \U$35216 ( \35594 , \35589 , \35593 );
and \U$35217 ( \35595 , \25609 , \25369 );
and \U$35218 ( \35596 , \25353 , \25367 );
nor \U$35219 ( \35597 , \35595 , \35596 );
xnor \U$35220 ( \35598 , \35597 , \25123 );
and \U$35221 ( \35599 , \35593 , \35598 );
and \U$35222 ( \35600 , \35589 , \35598 );
or \U$35223 ( \35601 , \35594 , \35599 , \35600 );
and \U$35224 ( \35602 , \35584 , \35601 );
and \U$35225 ( \35603 , \35568 , \35601 );
or \U$35226 ( \35604 , \35585 , \35602 , \35603 );
and \U$35227 ( \35605 , \22523 , \30770 );
and \U$35228 ( \35606 , \22325 , \30768 );
nor \U$35229 ( \35607 , \35605 , \35606 );
xnor \U$35230 ( \35608 , \35607 , \30460 );
and \U$35231 ( \35609 , \22716 , \30233 );
and \U$35232 ( \35610 , \22611 , \30231 );
nor \U$35233 ( \35611 , \35609 , \35610 );
xnor \U$35234 ( \35612 , \35611 , \29862 );
and \U$35235 ( \35613 , \35608 , \35612 );
and \U$35236 ( \35614 , \22837 , \29671 );
and \U$35237 ( \35615 , \22721 , \29669 );
nor \U$35238 ( \35616 , \35614 , \35615 );
xnor \U$35239 ( \35617 , \35616 , \29353 );
and \U$35240 ( \35618 , \35612 , \35617 );
and \U$35241 ( \35619 , \35608 , \35617 );
or \U$35242 ( \35620 , \35613 , \35618 , \35619 );
and \U$35243 ( \35621 , \22126 , \32151 );
and \U$35244 ( \35622 , \22046 , \32148 );
nor \U$35245 ( \35623 , \35621 , \35622 );
xnor \U$35246 ( \35624 , \35623 , \31096 );
and \U$35247 ( \35625 , \22262 , \31338 );
and \U$35248 ( \35626 , \22200 , \31336 );
nor \U$35249 ( \35627 , \35625 , \35626 );
xnor \U$35250 ( \35628 , \35627 , \31099 );
and \U$35251 ( \35629 , \35624 , \35628 );
and \U$35252 ( \35630 , \35628 , \21986 );
and \U$35253 ( \35631 , \35624 , \21986 );
or \U$35254 ( \35632 , \35629 , \35630 , \35631 );
and \U$35255 ( \35633 , \35620 , \35632 );
and \U$35256 ( \35634 , \23128 , \29104 );
and \U$35257 ( \35635 , \22952 , \29102 );
nor \U$35258 ( \35636 , \35634 , \35635 );
xnor \U$35259 ( \35637 , \35636 , \28855 );
and \U$35260 ( \35638 , \23379 , \28575 );
and \U$35261 ( \35639 , \23136 , \28573 );
nor \U$35262 ( \35640 , \35638 , \35639 );
xnor \U$35263 ( \35641 , \35640 , \28315 );
and \U$35264 ( \35642 , \35637 , \35641 );
and \U$35265 ( \35643 , \23570 , \28081 );
and \U$35266 ( \35644 , \23384 , \28079 );
nor \U$35267 ( \35645 , \35643 , \35644 );
xnor \U$35268 ( \35646 , \35645 , \27766 );
and \U$35269 ( \35647 , \35641 , \35646 );
and \U$35270 ( \35648 , \35637 , \35646 );
or \U$35271 ( \35649 , \35642 , \35647 , \35648 );
and \U$35272 ( \35650 , \35632 , \35649 );
and \U$35273 ( \35651 , \35620 , \35649 );
or \U$35274 ( \35652 , \35633 , \35650 , \35651 );
and \U$35275 ( \35653 , \35604 , \35652 );
and \U$35276 ( \35654 , \30887 , \22497 );
and \U$35277 ( \35655 , \30318 , \22495 );
nor \U$35278 ( \35656 , \35654 , \35655 );
xnor \U$35279 ( \35657 , \35656 , \22419 );
and \U$35280 ( \35658 , \31498 , \22333 );
and \U$35281 ( \35659 , \30895 , \22331 );
nor \U$35282 ( \35660 , \35658 , \35659 );
xnor \U$35283 ( \35661 , \35660 , \22239 );
and \U$35284 ( \35662 , \35657 , \35661 );
and \U$35285 ( \35663 , \31684 , \22163 );
and \U$35286 ( \35664 , \31503 , \22161 );
nor \U$35287 ( \35665 , \35663 , \35664 );
xnor \U$35288 ( \35666 , \35665 , \22091 );
and \U$35289 ( \35667 , \35661 , \35666 );
and \U$35290 ( \35668 , \35657 , \35666 );
or \U$35291 ( \35669 , \35662 , \35667 , \35668 );
and \U$35292 ( \35670 , \27485 , \23933 );
and \U$35293 ( \35671 , \27113 , \23931 );
nor \U$35294 ( \35672 , \35670 , \35671 );
xnor \U$35295 ( \35673 , \35672 , \23791 );
and \U$35296 ( \35674 , \27837 , \23637 );
and \U$35297 ( \35675 , \27494 , \23635 );
nor \U$35298 ( \35676 , \35674 , \35675 );
xnor \U$35299 ( \35677 , \35676 , \23500 );
and \U$35300 ( \35678 , \35673 , \35677 );
and \U$35301 ( \35679 , \28342 , \23431 );
and \U$35302 ( \35680 , \28039 , \23429 );
nor \U$35303 ( \35681 , \35679 , \35680 );
xnor \U$35304 ( \35682 , \35681 , \23279 );
and \U$35305 ( \35683 , \35677 , \35682 );
and \U$35306 ( \35684 , \35673 , \35682 );
or \U$35307 ( \35685 , \35678 , \35683 , \35684 );
and \U$35308 ( \35686 , \35669 , \35685 );
and \U$35309 ( \35687 , \29040 , \23163 );
and \U$35310 ( \35688 , \28514 , \23161 );
nor \U$35311 ( \35689 , \35687 , \35688 );
xnor \U$35312 ( \35690 , \35689 , \23007 );
and \U$35313 ( \35691 , \29710 , \22891 );
and \U$35314 ( \35692 , \29464 , \22889 );
nor \U$35315 ( \35693 , \35691 , \35692 );
xnor \U$35316 ( \35694 , \35693 , \22778 );
and \U$35317 ( \35695 , \35690 , \35694 );
and \U$35318 ( \35696 , \30034 , \22697 );
and \U$35319 ( \35697 , \29715 , \22695 );
nor \U$35320 ( \35698 , \35696 , \35697 );
xnor \U$35321 ( \35699 , \35698 , \22561 );
and \U$35322 ( \35700 , \35694 , \35699 );
and \U$35323 ( \35701 , \35690 , \35699 );
or \U$35324 ( \35702 , \35695 , \35700 , \35701 );
and \U$35325 ( \35703 , \35685 , \35702 );
and \U$35326 ( \35704 , \35669 , \35702 );
or \U$35327 ( \35705 , \35686 , \35703 , \35704 );
and \U$35328 ( \35706 , \35652 , \35705 );
and \U$35329 ( \35707 , \35604 , \35705 );
or \U$35330 ( \35708 , \35653 , \35706 , \35707 );
and \U$35331 ( \35709 , \35552 , \35708 );
xor \U$35332 ( \35710 , \35020 , \35024 );
xor \U$35333 ( \35711 , \35710 , \35029 );
xor \U$35334 ( \35712 , \35037 , \35041 );
xor \U$35335 ( \35713 , \35712 , \21867 );
and \U$35336 ( \35714 , \35711 , \35713 );
xor \U$35337 ( \35715 , \35265 , \35267 );
xor \U$35338 ( \35716 , \35715 , \35270 );
and \U$35339 ( \35717 , \35713 , \35716 );
and \U$35340 ( \35718 , \35711 , \35716 );
or \U$35341 ( \35719 , \35714 , \35717 , \35718 );
and \U$35342 ( \35720 , \35708 , \35719 );
and \U$35343 ( \35721 , \35552 , \35719 );
or \U$35344 ( \35722 , \35709 , \35720 , \35721 );
xor \U$35345 ( \35723 , \35292 , \35308 );
xor \U$35346 ( \35724 , \35723 , \35325 );
xor \U$35347 ( \35725 , \35242 , \35244 );
xor \U$35348 ( \35726 , \35725 , \35247 );
and \U$35349 ( \35727 , \35724 , \35726 );
xor \U$35350 ( \35728 , \35254 , \35256 );
xor \U$35351 ( \35729 , \35728 , \35259 );
and \U$35352 ( \35730 , \35726 , \35729 );
and \U$35353 ( \35731 , \35724 , \35729 );
or \U$35354 ( \35732 , \35727 , \35730 , \35731 );
xor \U$35355 ( \35733 , \35344 , \35360 );
xor \U$35356 ( \35734 , \35733 , \35377 );
xor \U$35357 ( \35735 , \35397 , \35413 );
xor \U$35358 ( \35736 , \35735 , \35430 );
and \U$35359 ( \35737 , \35734 , \35736 );
and \U$35360 ( \35738 , \35732 , \35737 );
xor \U$35361 ( \35739 , \35016 , \35032 );
xor \U$35362 ( \35740 , \35739 , \35045 );
and \U$35363 ( \35741 , \35737 , \35740 );
and \U$35364 ( \35742 , \35732 , \35740 );
or \U$35365 ( \35743 , \35738 , \35741 , \35742 );
and \U$35366 ( \35744 , \35722 , \35743 );
xor \U$35367 ( \35745 , \35250 , \35262 );
xor \U$35368 ( \35746 , \35745 , \35273 );
xor \U$35369 ( \35747 , \35452 , \35454 );
xor \U$35370 ( \35748 , \35747 , \35457 );
and \U$35371 ( \35749 , \35746 , \35748 );
xor \U$35372 ( \35750 , \35439 , \35441 );
xor \U$35373 ( \35751 , \35750 , \35444 );
and \U$35374 ( \35752 , \35748 , \35751 );
and \U$35375 ( \35753 , \35746 , \35751 );
or \U$35376 ( \35754 , \35749 , \35752 , \35753 );
and \U$35377 ( \35755 , \35743 , \35754 );
and \U$35378 ( \35756 , \35722 , \35754 );
or \U$35379 ( \35757 , \35744 , \35755 , \35756 );
xor \U$35380 ( \35758 , \35276 , \35436 );
xor \U$35381 ( \35759 , \35758 , \35447 );
xor \U$35382 ( \35760 , \35460 , \35462 );
xor \U$35383 ( \35761 , \35760 , \35465 );
and \U$35384 ( \35762 , \35759 , \35761 );
xor \U$35385 ( \35763 , \35471 , \35473 );
xor \U$35386 ( \35764 , \35763 , \35476 );
and \U$35387 ( \35765 , \35761 , \35764 );
and \U$35388 ( \35766 , \35759 , \35764 );
or \U$35389 ( \35767 , \35762 , \35765 , \35766 );
and \U$35390 ( \35768 , \35757 , \35767 );
xor \U$35391 ( \35769 , \35484 , \35486 );
xor \U$35392 ( \35770 , \35769 , \35489 );
and \U$35393 ( \35771 , \35767 , \35770 );
and \U$35394 ( \35772 , \35757 , \35770 );
or \U$35395 ( \35773 , \35768 , \35771 , \35772 );
xor \U$35396 ( \35774 , \35170 , \35188 );
xor \U$35397 ( \35775 , \35774 , \35199 );
and \U$35398 ( \35776 , \35773 , \35775 );
xor \U$35399 ( \35777 , \35482 , \35492 );
xor \U$35400 ( \35778 , \35777 , \35495 );
and \U$35401 ( \35779 , \35775 , \35778 );
and \U$35402 ( \35780 , \35773 , \35778 );
or \U$35403 ( \35781 , \35776 , \35779 , \35780 );
xor \U$35404 ( \35782 , \35498 , \35500 );
xor \U$35405 ( \35783 , \35782 , \35503 );
and \U$35406 ( \35784 , \35781 , \35783 );
and \U$35407 ( \35785 , \35518 , \35784 );
xor \U$35408 ( \35786 , \35518 , \35784 );
xor \U$35409 ( \35787 , \35781 , \35783 );
and \U$35410 ( \35788 , \25353 , \25692 );
and \U$35411 ( \35789 , \25348 , \25690 );
nor \U$35412 ( \35790 , \35788 , \35789 );
xnor \U$35413 ( \35791 , \35790 , \25549 );
and \U$35414 ( \35792 , \25806 , \25369 );
and \U$35415 ( \35793 , \25609 , \25367 );
nor \U$35416 ( \35794 , \35792 , \35793 );
xnor \U$35417 ( \35795 , \35794 , \25123 );
and \U$35418 ( \35796 , \35791 , \35795 );
and \U$35419 ( \35797 , \26116 , \24974 );
and \U$35420 ( \35798 , \26108 , \24972 );
nor \U$35421 ( \35799 , \35797 , \35798 );
xnor \U$35422 ( \35800 , \35799 , \24787 );
and \U$35423 ( \35801 , \35795 , \35800 );
and \U$35424 ( \35802 , \35791 , \35800 );
or \U$35425 ( \35803 , \35796 , \35801 , \35802 );
and \U$35426 ( \35804 , \24344 , \26983 );
and \U$35427 ( \35805 , \24177 , \26981 );
nor \U$35428 ( \35806 , \35804 , \35805 );
xnor \U$35429 ( \35807 , \35806 , \26742 );
and \U$35430 ( \35808 , \24601 , \26517 );
and \U$35431 ( \35809 , \24482 , \26515 );
nor \U$35432 ( \35810 , \35808 , \35809 );
xnor \U$35433 ( \35811 , \35810 , \26329 );
and \U$35434 ( \35812 , \35807 , \35811 );
and \U$35435 ( \35813 , \25226 , \26143 );
and \U$35436 ( \35814 , \25018 , \26141 );
nor \U$35437 ( \35815 , \35813 , \35814 );
xnor \U$35438 ( \35816 , \35815 , \25911 );
and \U$35439 ( \35817 , \35811 , \35816 );
and \U$35440 ( \35818 , \35807 , \35816 );
or \U$35441 ( \35819 , \35812 , \35817 , \35818 );
and \U$35442 ( \35820 , \35803 , \35819 );
and \U$35443 ( \35821 , \26590 , \24661 );
and \U$35444 ( \35822 , \26585 , \24659 );
nor \U$35445 ( \35823 , \35821 , \35822 );
xnor \U$35446 ( \35824 , \35823 , \24456 );
and \U$35447 ( \35825 , \27113 , \24255 );
and \U$35448 ( \35826 , \26854 , \24253 );
nor \U$35449 ( \35827 , \35825 , \35826 );
xnor \U$35450 ( \35828 , \35827 , \24106 );
and \U$35451 ( \35829 , \35824 , \35828 );
and \U$35452 ( \35830 , \27494 , \23933 );
and \U$35453 ( \35831 , \27485 , \23931 );
nor \U$35454 ( \35832 , \35830 , \35831 );
xnor \U$35455 ( \35833 , \35832 , \23791 );
and \U$35456 ( \35834 , \35828 , \35833 );
and \U$35457 ( \35835 , \35824 , \35833 );
or \U$35458 ( \35836 , \35829 , \35834 , \35835 );
and \U$35459 ( \35837 , \35819 , \35836 );
and \U$35460 ( \35838 , \35803 , \35836 );
or \U$35461 ( \35839 , \35820 , \35837 , \35838 );
and \U$35462 ( \35840 , \29715 , \22891 );
and \U$35463 ( \35841 , \29710 , \22889 );
nor \U$35464 ( \35842 , \35840 , \35841 );
xnor \U$35465 ( \35843 , \35842 , \22778 );
and \U$35466 ( \35844 , \30318 , \22697 );
and \U$35467 ( \35845 , \30034 , \22695 );
nor \U$35468 ( \35846 , \35844 , \35845 );
xnor \U$35469 ( \35847 , \35846 , \22561 );
and \U$35470 ( \35848 , \35843 , \35847 );
and \U$35471 ( \35849 , \30895 , \22497 );
and \U$35472 ( \35850 , \30887 , \22495 );
nor \U$35473 ( \35851 , \35849 , \35850 );
xnor \U$35474 ( \35852 , \35851 , \22419 );
and \U$35475 ( \35853 , \35847 , \35852 );
and \U$35476 ( \35854 , \35843 , \35852 );
or \U$35477 ( \35855 , \35848 , \35853 , \35854 );
and \U$35478 ( \35856 , \28039 , \23637 );
and \U$35479 ( \35857 , \27837 , \23635 );
nor \U$35480 ( \35858 , \35856 , \35857 );
xnor \U$35481 ( \35859 , \35858 , \23500 );
and \U$35482 ( \35860 , \28514 , \23431 );
and \U$35483 ( \35861 , \28342 , \23429 );
nor \U$35484 ( \35862 , \35860 , \35861 );
xnor \U$35485 ( \35863 , \35862 , \23279 );
and \U$35486 ( \35864 , \35859 , \35863 );
and \U$35487 ( \35865 , \29464 , \23163 );
and \U$35488 ( \35866 , \29040 , \23161 );
nor \U$35489 ( \35867 , \35865 , \35866 );
xnor \U$35490 ( \35868 , \35867 , \23007 );
and \U$35491 ( \35869 , \35863 , \35868 );
and \U$35492 ( \35870 , \35859 , \35868 );
or \U$35493 ( \35871 , \35864 , \35869 , \35870 );
and \U$35494 ( \35872 , \35855 , \35871 );
and \U$35495 ( \35873 , \31503 , \22333 );
and \U$35496 ( \35874 , \31498 , \22331 );
nor \U$35497 ( \35875 , \35873 , \35874 );
xnor \U$35498 ( \35876 , \35875 , \22239 );
and \U$35499 ( \35877 , \32304 , \22163 );
and \U$35500 ( \35878 , \31684 , \22161 );
nor \U$35501 ( \35879 , \35877 , \35878 );
xnor \U$35502 ( \35880 , \35879 , \22091 );
and \U$35503 ( \35881 , \35876 , \35880 );
and \U$35504 ( \35882 , \35871 , \35881 );
and \U$35505 ( \35883 , \35855 , \35881 );
or \U$35506 ( \35884 , \35872 , \35882 , \35883 );
and \U$35507 ( \35885 , \35839 , \35884 );
and \U$35508 ( \35886 , \23384 , \28575 );
and \U$35509 ( \35887 , \23379 , \28573 );
nor \U$35510 ( \35888 , \35886 , \35887 );
xnor \U$35511 ( \35889 , \35888 , \28315 );
and \U$35512 ( \35890 , \23714 , \28081 );
and \U$35513 ( \35891 , \23570 , \28079 );
nor \U$35514 ( \35892 , \35890 , \35891 );
xnor \U$35515 ( \35893 , \35892 , \27766 );
and \U$35516 ( \35894 , \35889 , \35893 );
and \U$35517 ( \35895 , \24003 , \27572 );
and \U$35518 ( \35896 , \23978 , \27570 );
nor \U$35519 ( \35897 , \35895 , \35896 );
xnor \U$35520 ( \35898 , \35897 , \27232 );
and \U$35521 ( \35899 , \35893 , \35898 );
and \U$35522 ( \35900 , \35889 , \35898 );
or \U$35523 ( \35901 , \35894 , \35899 , \35900 );
and \U$35524 ( \35902 , \22200 , \32151 );
and \U$35525 ( \35903 , \22126 , \32148 );
nor \U$35526 ( \35904 , \35902 , \35903 );
xnor \U$35527 ( \35905 , \35904 , \31096 );
and \U$35528 ( \35906 , \22325 , \31338 );
and \U$35529 ( \35907 , \22262 , \31336 );
nor \U$35530 ( \35908 , \35906 , \35907 );
xnor \U$35531 ( \35909 , \35908 , \31099 );
and \U$35532 ( \35910 , \35905 , \35909 );
and \U$35533 ( \35911 , \22611 , \30770 );
and \U$35534 ( \35912 , \22523 , \30768 );
nor \U$35535 ( \35913 , \35911 , \35912 );
xnor \U$35536 ( \35914 , \35913 , \30460 );
and \U$35537 ( \35915 , \35909 , \35914 );
and \U$35538 ( \35916 , \35905 , \35914 );
or \U$35539 ( \35917 , \35910 , \35915 , \35916 );
and \U$35540 ( \35918 , \35901 , \35917 );
and \U$35541 ( \35919 , \22721 , \30233 );
and \U$35542 ( \35920 , \22716 , \30231 );
nor \U$35543 ( \35921 , \35919 , \35920 );
xnor \U$35544 ( \35922 , \35921 , \29862 );
and \U$35545 ( \35923 , \22952 , \29671 );
and \U$35546 ( \35924 , \22837 , \29669 );
nor \U$35547 ( \35925 , \35923 , \35924 );
xnor \U$35548 ( \35926 , \35925 , \29353 );
and \U$35549 ( \35927 , \35922 , \35926 );
and \U$35550 ( \35928 , \23136 , \29104 );
and \U$35551 ( \35929 , \23128 , \29102 );
nor \U$35552 ( \35930 , \35928 , \35929 );
xnor \U$35553 ( \35931 , \35930 , \28855 );
and \U$35554 ( \35932 , \35926 , \35931 );
and \U$35555 ( \35933 , \35922 , \35931 );
or \U$35556 ( \35934 , \35927 , \35932 , \35933 );
and \U$35557 ( \35935 , \35917 , \35934 );
and \U$35558 ( \35936 , \35901 , \35934 );
or \U$35559 ( \35937 , \35918 , \35935 , \35936 );
and \U$35560 ( \35938 , \35884 , \35937 );
and \U$35561 ( \35939 , \35839 , \35937 );
or \U$35562 ( \35940 , \35885 , \35938 , \35939 );
xor \U$35563 ( \35941 , \35608 , \35612 );
xor \U$35564 ( \35942 , \35941 , \35617 );
xor \U$35565 ( \35943 , \35637 , \35641 );
xor \U$35566 ( \35944 , \35943 , \35646 );
and \U$35567 ( \35945 , \35942 , \35944 );
xor \U$35568 ( \35946 , \35572 , \35576 );
xor \U$35569 ( \35947 , \35946 , \35581 );
and \U$35570 ( \35948 , \35944 , \35947 );
and \U$35571 ( \35949 , \35942 , \35947 );
or \U$35572 ( \35950 , \35945 , \35948 , \35949 );
nand \U$35573 ( \35951 , \32304 , \22027 );
xnor \U$35574 ( \35952 , \35951 , \21986 );
xor \U$35575 ( \35953 , \35657 , \35661 );
xor \U$35576 ( \35954 , \35953 , \35666 );
and \U$35577 ( \35955 , \35952 , \35954 );
xor \U$35578 ( \35956 , \35690 , \35694 );
xor \U$35579 ( \35957 , \35956 , \35699 );
and \U$35580 ( \35958 , \35954 , \35957 );
and \U$35581 ( \35959 , \35952 , \35957 );
or \U$35582 ( \35960 , \35955 , \35958 , \35959 );
and \U$35583 ( \35961 , \35950 , \35960 );
xor \U$35584 ( \35962 , \35673 , \35677 );
xor \U$35585 ( \35963 , \35962 , \35682 );
xor \U$35586 ( \35964 , \35556 , \35560 );
xor \U$35587 ( \35965 , \35964 , \35565 );
and \U$35588 ( \35966 , \35963 , \35965 );
xor \U$35589 ( \35967 , \35589 , \35593 );
xor \U$35590 ( \35968 , \35967 , \35598 );
and \U$35591 ( \35969 , \35965 , \35968 );
and \U$35592 ( \35970 , \35963 , \35968 );
or \U$35593 ( \35971 , \35966 , \35969 , \35970 );
and \U$35594 ( \35972 , \35960 , \35971 );
and \U$35595 ( \35973 , \35950 , \35971 );
or \U$35596 ( \35974 , \35961 , \35972 , \35973 );
and \U$35597 ( \35975 , \35940 , \35974 );
xor \U$35598 ( \35976 , \35520 , \35522 );
xor \U$35599 ( \35977 , \35976 , \35525 );
xor \U$35600 ( \35978 , \35530 , \35532 );
xor \U$35601 ( \35979 , \35978 , \35535 );
and \U$35602 ( \35980 , \35977 , \35979 );
xor \U$35603 ( \35981 , \35541 , \35543 );
xor \U$35604 ( \35982 , \35981 , \35546 );
and \U$35605 ( \35983 , \35979 , \35982 );
and \U$35606 ( \35984 , \35977 , \35982 );
or \U$35607 ( \35985 , \35980 , \35983 , \35984 );
and \U$35608 ( \35986 , \35974 , \35985 );
and \U$35609 ( \35987 , \35940 , \35985 );
or \U$35610 ( \35988 , \35975 , \35986 , \35987 );
xor \U$35611 ( \35989 , \35528 , \35538 );
xor \U$35612 ( \35990 , \35989 , \35549 );
xor \U$35613 ( \35991 , \35604 , \35652 );
xor \U$35614 ( \35992 , \35991 , \35705 );
and \U$35615 ( \35993 , \35990 , \35992 );
xor \U$35616 ( \35994 , \35711 , \35713 );
xor \U$35617 ( \35995 , \35994 , \35716 );
and \U$35618 ( \35996 , \35992 , \35995 );
and \U$35619 ( \35997 , \35990 , \35995 );
or \U$35620 ( \35998 , \35993 , \35996 , \35997 );
and \U$35621 ( \35999 , \35988 , \35998 );
xor \U$35622 ( \36000 , \35568 , \35584 );
xor \U$35623 ( \36001 , \36000 , \35601 );
xor \U$35624 ( \36002 , \35620 , \35632 );
xor \U$35625 ( \36003 , \36002 , \35649 );
and \U$35626 ( \36004 , \36001 , \36003 );
xor \U$35627 ( \36005 , \35669 , \35685 );
xor \U$35628 ( \36006 , \36005 , \35702 );
and \U$35629 ( \36007 , \36003 , \36006 );
and \U$35630 ( \36008 , \36001 , \36006 );
or \U$35631 ( \36009 , \36004 , \36007 , \36008 );
xor \U$35632 ( \36010 , \35724 , \35726 );
xor \U$35633 ( \36011 , \36010 , \35729 );
and \U$35634 ( \36012 , \36009 , \36011 );
xor \U$35635 ( \36013 , \35734 , \35736 );
and \U$35636 ( \36014 , \36011 , \36013 );
and \U$35637 ( \36015 , \36009 , \36013 );
or \U$35638 ( \36016 , \36012 , \36014 , \36015 );
and \U$35639 ( \36017 , \35998 , \36016 );
and \U$35640 ( \36018 , \35988 , \36016 );
or \U$35641 ( \36019 , \35999 , \36017 , \36018 );
xor \U$35642 ( \36020 , \35328 , \35380 );
xor \U$35643 ( \36021 , \36020 , \35433 );
xor \U$35644 ( \36022 , \35732 , \35737 );
xor \U$35645 ( \36023 , \36022 , \35740 );
and \U$35646 ( \36024 , \36021 , \36023 );
xor \U$35647 ( \36025 , \35746 , \35748 );
xor \U$35648 ( \36026 , \36025 , \35751 );
and \U$35649 ( \36027 , \36023 , \36026 );
and \U$35650 ( \36028 , \36021 , \36026 );
or \U$35651 ( \36029 , \36024 , \36027 , \36028 );
and \U$35652 ( \36030 , \36019 , \36029 );
xor \U$35653 ( \36031 , \35759 , \35761 );
xor \U$35654 ( \36032 , \36031 , \35764 );
and \U$35655 ( \36033 , \36029 , \36032 );
and \U$35656 ( \36034 , \36019 , \36032 );
or \U$35657 ( \36035 , \36030 , \36033 , \36034 );
xor \U$35658 ( \36036 , \35450 , \35468 );
xor \U$35659 ( \36037 , \36036 , \35479 );
and \U$35660 ( \36038 , \36035 , \36037 );
xor \U$35661 ( \36039 , \35757 , \35767 );
xor \U$35662 ( \36040 , \36039 , \35770 );
and \U$35663 ( \36041 , \36037 , \36040 );
and \U$35664 ( \36042 , \36035 , \36040 );
or \U$35665 ( \36043 , \36038 , \36041 , \36042 );
xor \U$35666 ( \36044 , \35773 , \35775 );
xor \U$35667 ( \36045 , \36044 , \35778 );
and \U$35668 ( \36046 , \36043 , \36045 );
and \U$35669 ( \36047 , \35787 , \36046 );
xor \U$35670 ( \36048 , \35787 , \36046 );
xor \U$35671 ( \36049 , \36043 , \36045 );
and \U$35672 ( \36050 , \25348 , \26143 );
and \U$35673 ( \36051 , \25226 , \26141 );
nor \U$35674 ( \36052 , \36050 , \36051 );
xnor \U$35675 ( \36053 , \36052 , \25911 );
and \U$35676 ( \36054 , \25609 , \25692 );
and \U$35677 ( \36055 , \25353 , \25690 );
nor \U$35678 ( \36056 , \36054 , \36055 );
xnor \U$35679 ( \36057 , \36056 , \25549 );
and \U$35680 ( \36058 , \36053 , \36057 );
and \U$35681 ( \36059 , \26108 , \25369 );
and \U$35682 ( \36060 , \25806 , \25367 );
nor \U$35683 ( \36061 , \36059 , \36060 );
xnor \U$35684 ( \36062 , \36061 , \25123 );
and \U$35685 ( \36063 , \36057 , \36062 );
and \U$35686 ( \36064 , \36053 , \36062 );
or \U$35687 ( \36065 , \36058 , \36063 , \36064 );
and \U$35688 ( \36066 , \24177 , \27572 );
and \U$35689 ( \36067 , \24003 , \27570 );
nor \U$35690 ( \36068 , \36066 , \36067 );
xnor \U$35691 ( \36069 , \36068 , \27232 );
and \U$35692 ( \36070 , \24482 , \26983 );
and \U$35693 ( \36071 , \24344 , \26981 );
nor \U$35694 ( \36072 , \36070 , \36071 );
xnor \U$35695 ( \36073 , \36072 , \26742 );
and \U$35696 ( \36074 , \36069 , \36073 );
and \U$35697 ( \36075 , \25018 , \26517 );
and \U$35698 ( \36076 , \24601 , \26515 );
nor \U$35699 ( \36077 , \36075 , \36076 );
xnor \U$35700 ( \36078 , \36077 , \26329 );
and \U$35701 ( \36079 , \36073 , \36078 );
and \U$35702 ( \36080 , \36069 , \36078 );
or \U$35703 ( \36081 , \36074 , \36079 , \36080 );
and \U$35704 ( \36082 , \36065 , \36081 );
and \U$35705 ( \36083 , \26585 , \24974 );
and \U$35706 ( \36084 , \26116 , \24972 );
nor \U$35707 ( \36085 , \36083 , \36084 );
xnor \U$35708 ( \36086 , \36085 , \24787 );
and \U$35709 ( \36087 , \26854 , \24661 );
and \U$35710 ( \36088 , \26590 , \24659 );
nor \U$35711 ( \36089 , \36087 , \36088 );
xnor \U$35712 ( \36090 , \36089 , \24456 );
and \U$35713 ( \36091 , \36086 , \36090 );
and \U$35714 ( \36092 , \27485 , \24255 );
and \U$35715 ( \36093 , \27113 , \24253 );
nor \U$35716 ( \36094 , \36092 , \36093 );
xnor \U$35717 ( \36095 , \36094 , \24106 );
and \U$35718 ( \36096 , \36090 , \36095 );
and \U$35719 ( \36097 , \36086 , \36095 );
or \U$35720 ( \36098 , \36091 , \36096 , \36097 );
and \U$35721 ( \36099 , \36081 , \36098 );
and \U$35722 ( \36100 , \36065 , \36098 );
or \U$35723 ( \36101 , \36082 , \36099 , \36100 );
and \U$35724 ( \36102 , \23379 , \29104 );
and \U$35725 ( \36103 , \23136 , \29102 );
nor \U$35726 ( \36104 , \36102 , \36103 );
xnor \U$35727 ( \36105 , \36104 , \28855 );
and \U$35728 ( \36106 , \23570 , \28575 );
and \U$35729 ( \36107 , \23384 , \28573 );
nor \U$35730 ( \36108 , \36106 , \36107 );
xnor \U$35731 ( \36109 , \36108 , \28315 );
and \U$35732 ( \36110 , \36105 , \36109 );
and \U$35733 ( \36111 , \23978 , \28081 );
and \U$35734 ( \36112 , \23714 , \28079 );
nor \U$35735 ( \36113 , \36111 , \36112 );
xnor \U$35736 ( \36114 , \36113 , \27766 );
and \U$35737 ( \36115 , \36109 , \36114 );
and \U$35738 ( \36116 , \36105 , \36114 );
or \U$35739 ( \36117 , \36110 , \36115 , \36116 );
and \U$35740 ( \36118 , \22716 , \30770 );
and \U$35741 ( \36119 , \22611 , \30768 );
nor \U$35742 ( \36120 , \36118 , \36119 );
xnor \U$35743 ( \36121 , \36120 , \30460 );
and \U$35744 ( \36122 , \22837 , \30233 );
and \U$35745 ( \36123 , \22721 , \30231 );
nor \U$35746 ( \36124 , \36122 , \36123 );
xnor \U$35747 ( \36125 , \36124 , \29862 );
and \U$35748 ( \36126 , \36121 , \36125 );
and \U$35749 ( \36127 , \23128 , \29671 );
and \U$35750 ( \36128 , \22952 , \29669 );
nor \U$35751 ( \36129 , \36127 , \36128 );
xnor \U$35752 ( \36130 , \36129 , \29353 );
and \U$35753 ( \36131 , \36125 , \36130 );
and \U$35754 ( \36132 , \36121 , \36130 );
or \U$35755 ( \36133 , \36126 , \36131 , \36132 );
and \U$35756 ( \36134 , \36117 , \36133 );
and \U$35757 ( \36135 , \22262 , \32151 );
and \U$35758 ( \36136 , \22200 , \32148 );
nor \U$35759 ( \36137 , \36135 , \36136 );
xnor \U$35760 ( \36138 , \36137 , \31096 );
and \U$35761 ( \36139 , \22523 , \31338 );
and \U$35762 ( \36140 , \22325 , \31336 );
nor \U$35763 ( \36141 , \36139 , \36140 );
xnor \U$35764 ( \36142 , \36141 , \31099 );
and \U$35765 ( \36143 , \36138 , \36142 );
and \U$35766 ( \36144 , \36142 , \22091 );
and \U$35767 ( \36145 , \36138 , \22091 );
or \U$35768 ( \36146 , \36143 , \36144 , \36145 );
and \U$35769 ( \36147 , \36133 , \36146 );
and \U$35770 ( \36148 , \36117 , \36146 );
or \U$35771 ( \36149 , \36134 , \36147 , \36148 );
and \U$35772 ( \36150 , \36101 , \36149 );
and \U$35773 ( \36151 , \27837 , \23933 );
and \U$35774 ( \36152 , \27494 , \23931 );
nor \U$35775 ( \36153 , \36151 , \36152 );
xnor \U$35776 ( \36154 , \36153 , \23791 );
and \U$35777 ( \36155 , \28342 , \23637 );
and \U$35778 ( \36156 , \28039 , \23635 );
nor \U$35779 ( \36157 , \36155 , \36156 );
xnor \U$35780 ( \36158 , \36157 , \23500 );
and \U$35781 ( \36159 , \36154 , \36158 );
and \U$35782 ( \36160 , \29040 , \23431 );
and \U$35783 ( \36161 , \28514 , \23429 );
nor \U$35784 ( \36162 , \36160 , \36161 );
xnor \U$35785 ( \36163 , \36162 , \23279 );
and \U$35786 ( \36164 , \36158 , \36163 );
and \U$35787 ( \36165 , \36154 , \36163 );
or \U$35788 ( \36166 , \36159 , \36164 , \36165 );
and \U$35789 ( \36167 , \31498 , \22497 );
and \U$35790 ( \36168 , \30895 , \22495 );
nor \U$35791 ( \36169 , \36167 , \36168 );
xnor \U$35792 ( \36170 , \36169 , \22419 );
and \U$35793 ( \36171 , \31684 , \22333 );
and \U$35794 ( \36172 , \31503 , \22331 );
nor \U$35795 ( \36173 , \36171 , \36172 );
xnor \U$35796 ( \36174 , \36173 , \22239 );
and \U$35797 ( \36175 , \36170 , \36174 );
nand \U$35798 ( \36176 , \32304 , \22161 );
xnor \U$35799 ( \36177 , \36176 , \22091 );
and \U$35800 ( \36178 , \36174 , \36177 );
and \U$35801 ( \36179 , \36170 , \36177 );
or \U$35802 ( \36180 , \36175 , \36178 , \36179 );
and \U$35803 ( \36181 , \36166 , \36180 );
and \U$35804 ( \36182 , \29710 , \23163 );
and \U$35805 ( \36183 , \29464 , \23161 );
nor \U$35806 ( \36184 , \36182 , \36183 );
xnor \U$35807 ( \36185 , \36184 , \23007 );
and \U$35808 ( \36186 , \30034 , \22891 );
and \U$35809 ( \36187 , \29715 , \22889 );
nor \U$35810 ( \36188 , \36186 , \36187 );
xnor \U$35811 ( \36189 , \36188 , \22778 );
and \U$35812 ( \36190 , \36185 , \36189 );
and \U$35813 ( \36191 , \30887 , \22697 );
and \U$35814 ( \36192 , \30318 , \22695 );
nor \U$35815 ( \36193 , \36191 , \36192 );
xnor \U$35816 ( \36194 , \36193 , \22561 );
and \U$35817 ( \36195 , \36189 , \36194 );
and \U$35818 ( \36196 , \36185 , \36194 );
or \U$35819 ( \36197 , \36190 , \36195 , \36196 );
and \U$35820 ( \36198 , \36180 , \36197 );
and \U$35821 ( \36199 , \36166 , \36197 );
or \U$35822 ( \36200 , \36181 , \36198 , \36199 );
and \U$35823 ( \36201 , \36149 , \36200 );
and \U$35824 ( \36202 , \36101 , \36200 );
or \U$35825 ( \36203 , \36150 , \36201 , \36202 );
xor \U$35826 ( \36204 , \35889 , \35893 );
xor \U$35827 ( \36205 , \36204 , \35898 );
xor \U$35828 ( \36206 , \35905 , \35909 );
xor \U$35829 ( \36207 , \36206 , \35914 );
and \U$35830 ( \36208 , \36205 , \36207 );
xor \U$35831 ( \36209 , \35922 , \35926 );
xor \U$35832 ( \36210 , \36209 , \35931 );
and \U$35833 ( \36211 , \36207 , \36210 );
and \U$35834 ( \36212 , \36205 , \36210 );
or \U$35835 ( \36213 , \36208 , \36211 , \36212 );
xor \U$35836 ( \36214 , \35791 , \35795 );
xor \U$35837 ( \36215 , \36214 , \35800 );
xor \U$35838 ( \36216 , \35807 , \35811 );
xor \U$35839 ( \36217 , \36216 , \35816 );
and \U$35840 ( \36218 , \36215 , \36217 );
xor \U$35841 ( \36219 , \35824 , \35828 );
xor \U$35842 ( \36220 , \36219 , \35833 );
and \U$35843 ( \36221 , \36217 , \36220 );
and \U$35844 ( \36222 , \36215 , \36220 );
or \U$35845 ( \36223 , \36218 , \36221 , \36222 );
and \U$35846 ( \36224 , \36213 , \36223 );
xor \U$35847 ( \36225 , \35843 , \35847 );
xor \U$35848 ( \36226 , \36225 , \35852 );
xor \U$35849 ( \36227 , \35859 , \35863 );
xor \U$35850 ( \36228 , \36227 , \35868 );
and \U$35851 ( \36229 , \36226 , \36228 );
xor \U$35852 ( \36230 , \35876 , \35880 );
and \U$35853 ( \36231 , \36228 , \36230 );
and \U$35854 ( \36232 , \36226 , \36230 );
or \U$35855 ( \36233 , \36229 , \36231 , \36232 );
and \U$35856 ( \36234 , \36223 , \36233 );
and \U$35857 ( \36235 , \36213 , \36233 );
or \U$35858 ( \36236 , \36224 , \36234 , \36235 );
and \U$35859 ( \36237 , \36203 , \36236 );
xor \U$35860 ( \36238 , \35624 , \35628 );
xor \U$35861 ( \36239 , \36238 , \21986 );
xor \U$35862 ( \36240 , \35942 , \35944 );
xor \U$35863 ( \36241 , \36240 , \35947 );
and \U$35864 ( \36242 , \36239 , \36241 );
xor \U$35865 ( \36243 , \35963 , \35965 );
xor \U$35866 ( \36244 , \36243 , \35968 );
and \U$35867 ( \36245 , \36241 , \36244 );
and \U$35868 ( \36246 , \36239 , \36244 );
or \U$35869 ( \36247 , \36242 , \36245 , \36246 );
and \U$35870 ( \36248 , \36236 , \36247 );
and \U$35871 ( \36249 , \36203 , \36247 );
or \U$35872 ( \36250 , \36237 , \36248 , \36249 );
xor \U$35873 ( \36251 , \35803 , \35819 );
xor \U$35874 ( \36252 , \36251 , \35836 );
xor \U$35875 ( \36253 , \35855 , \35871 );
xor \U$35876 ( \36254 , \36253 , \35881 );
and \U$35877 ( \36255 , \36252 , \36254 );
xor \U$35878 ( \36256 , \35952 , \35954 );
xor \U$35879 ( \36257 , \36256 , \35957 );
and \U$35880 ( \36258 , \36254 , \36257 );
and \U$35881 ( \36259 , \36252 , \36257 );
or \U$35882 ( \36260 , \36255 , \36258 , \36259 );
xor \U$35883 ( \36261 , \36001 , \36003 );
xor \U$35884 ( \36262 , \36261 , \36006 );
and \U$35885 ( \36263 , \36260 , \36262 );
xor \U$35886 ( \36264 , \35977 , \35979 );
xor \U$35887 ( \36265 , \36264 , \35982 );
and \U$35888 ( \36266 , \36262 , \36265 );
and \U$35889 ( \36267 , \36260 , \36265 );
or \U$35890 ( \36268 , \36263 , \36266 , \36267 );
and \U$35891 ( \36269 , \36250 , \36268 );
xor \U$35892 ( \36270 , \35839 , \35884 );
xor \U$35893 ( \36271 , \36270 , \35937 );
xor \U$35894 ( \36272 , \35950 , \35960 );
xor \U$35895 ( \36273 , \36272 , \35971 );
and \U$35896 ( \36274 , \36271 , \36273 );
and \U$35897 ( \36275 , \36268 , \36274 );
and \U$35898 ( \36276 , \36250 , \36274 );
or \U$35899 ( \36277 , \36269 , \36275 , \36276 );
xor \U$35900 ( \36278 , \35940 , \35974 );
xor \U$35901 ( \36279 , \36278 , \35985 );
xor \U$35902 ( \36280 , \35990 , \35992 );
xor \U$35903 ( \36281 , \36280 , \35995 );
and \U$35904 ( \36282 , \36279 , \36281 );
xor \U$35905 ( \36283 , \36009 , \36011 );
xor \U$35906 ( \36284 , \36283 , \36013 );
and \U$35907 ( \36285 , \36281 , \36284 );
and \U$35908 ( \36286 , \36279 , \36284 );
or \U$35909 ( \36287 , \36282 , \36285 , \36286 );
and \U$35910 ( \36288 , \36277 , \36287 );
xor \U$35911 ( \36289 , \35552 , \35708 );
xor \U$35912 ( \36290 , \36289 , \35719 );
and \U$35913 ( \36291 , \36287 , \36290 );
and \U$35914 ( \36292 , \36277 , \36290 );
or \U$35915 ( \36293 , \36288 , \36291 , \36292 );
xor \U$35916 ( \36294 , \35988 , \35998 );
xor \U$35917 ( \36295 , \36294 , \36016 );
xor \U$35918 ( \36296 , \36021 , \36023 );
xor \U$35919 ( \36297 , \36296 , \36026 );
and \U$35920 ( \36298 , \36295 , \36297 );
and \U$35921 ( \36299 , \36293 , \36298 );
xor \U$35922 ( \36300 , \35722 , \35743 );
xor \U$35923 ( \36301 , \36300 , \35754 );
and \U$35924 ( \36302 , \36298 , \36301 );
and \U$35925 ( \36303 , \36293 , \36301 );
or \U$35926 ( \36304 , \36299 , \36302 , \36303 );
xor \U$35927 ( \36305 , \36035 , \36037 );
xor \U$35928 ( \36306 , \36305 , \36040 );
and \U$35929 ( \36307 , \36304 , \36306 );
and \U$35930 ( \36308 , \36049 , \36307 );
xor \U$35931 ( \36309 , \36049 , \36307 );
xor \U$35932 ( \36310 , \36304 , \36306 );
xor \U$35933 ( \36311 , \36293 , \36298 );
xor \U$35934 ( \36312 , \36311 , \36301 );
xor \U$35935 ( \36313 , \36019 , \36029 );
xor \U$35936 ( \36314 , \36313 , \36032 );
and \U$35937 ( \36315 , \36312 , \36314 );
and \U$35938 ( \36316 , \36310 , \36315 );
xor \U$35939 ( \36317 , \36310 , \36315 );
xor \U$35940 ( \36318 , \36312 , \36314 );
and \U$35941 ( \36319 , \23714 , \28575 );
and \U$35942 ( \36320 , \23570 , \28573 );
nor \U$35943 ( \36321 , \36319 , \36320 );
xnor \U$35944 ( \36322 , \36321 , \28315 );
and \U$35945 ( \36323 , \24003 , \28081 );
and \U$35946 ( \36324 , \23978 , \28079 );
nor \U$35947 ( \36325 , \36323 , \36324 );
xnor \U$35948 ( \36326 , \36325 , \27766 );
and \U$35949 ( \36327 , \36322 , \36326 );
and \U$35950 ( \36328 , \24344 , \27572 );
and \U$35951 ( \36329 , \24177 , \27570 );
nor \U$35952 ( \36330 , \36328 , \36329 );
xnor \U$35953 ( \36331 , \36330 , \27232 );
and \U$35954 ( \36332 , \36326 , \36331 );
and \U$35955 ( \36333 , \36322 , \36331 );
or \U$35956 ( \36334 , \36327 , \36332 , \36333 );
and \U$35957 ( \36335 , \22325 , \32151 );
and \U$35958 ( \36336 , \22262 , \32148 );
nor \U$35959 ( \36337 , \36335 , \36336 );
xnor \U$35960 ( \36338 , \36337 , \31096 );
and \U$35961 ( \36339 , \22611 , \31338 );
and \U$35962 ( \36340 , \22523 , \31336 );
nor \U$35963 ( \36341 , \36339 , \36340 );
xnor \U$35964 ( \36342 , \36341 , \31099 );
and \U$35965 ( \36343 , \36338 , \36342 );
and \U$35966 ( \36344 , \22721 , \30770 );
and \U$35967 ( \36345 , \22716 , \30768 );
nor \U$35968 ( \36346 , \36344 , \36345 );
xnor \U$35969 ( \36347 , \36346 , \30460 );
and \U$35970 ( \36348 , \36342 , \36347 );
and \U$35971 ( \36349 , \36338 , \36347 );
or \U$35972 ( \36350 , \36343 , \36348 , \36349 );
and \U$35973 ( \36351 , \36334 , \36350 );
and \U$35974 ( \36352 , \22952 , \30233 );
and \U$35975 ( \36353 , \22837 , \30231 );
nor \U$35976 ( \36354 , \36352 , \36353 );
xnor \U$35977 ( \36355 , \36354 , \29862 );
and \U$35978 ( \36356 , \23136 , \29671 );
and \U$35979 ( \36357 , \23128 , \29669 );
nor \U$35980 ( \36358 , \36356 , \36357 );
xnor \U$35981 ( \36359 , \36358 , \29353 );
and \U$35982 ( \36360 , \36355 , \36359 );
and \U$35983 ( \36361 , \23384 , \29104 );
and \U$35984 ( \36362 , \23379 , \29102 );
nor \U$35985 ( \36363 , \36361 , \36362 );
xnor \U$35986 ( \36364 , \36363 , \28855 );
and \U$35987 ( \36365 , \36359 , \36364 );
and \U$35988 ( \36366 , \36355 , \36364 );
or \U$35989 ( \36367 , \36360 , \36365 , \36366 );
and \U$35990 ( \36368 , \36350 , \36367 );
and \U$35991 ( \36369 , \36334 , \36367 );
or \U$35992 ( \36370 , \36351 , \36368 , \36369 );
and \U$35993 ( \36371 , \25806 , \25692 );
and \U$35994 ( \36372 , \25609 , \25690 );
nor \U$35995 ( \36373 , \36371 , \36372 );
xnor \U$35996 ( \36374 , \36373 , \25549 );
and \U$35997 ( \36375 , \26116 , \25369 );
and \U$35998 ( \36376 , \26108 , \25367 );
nor \U$35999 ( \36377 , \36375 , \36376 );
xnor \U$36000 ( \36378 , \36377 , \25123 );
and \U$36001 ( \36379 , \36374 , \36378 );
and \U$36002 ( \36380 , \26590 , \24974 );
and \U$36003 ( \36381 , \26585 , \24972 );
nor \U$36004 ( \36382 , \36380 , \36381 );
xnor \U$36005 ( \36383 , \36382 , \24787 );
and \U$36006 ( \36384 , \36378 , \36383 );
and \U$36007 ( \36385 , \36374 , \36383 );
or \U$36008 ( \36386 , \36379 , \36384 , \36385 );
and \U$36009 ( \36387 , \24601 , \26983 );
and \U$36010 ( \36388 , \24482 , \26981 );
nor \U$36011 ( \36389 , \36387 , \36388 );
xnor \U$36012 ( \36390 , \36389 , \26742 );
and \U$36013 ( \36391 , \25226 , \26517 );
and \U$36014 ( \36392 , \25018 , \26515 );
nor \U$36015 ( \36393 , \36391 , \36392 );
xnor \U$36016 ( \36394 , \36393 , \26329 );
and \U$36017 ( \36395 , \36390 , \36394 );
and \U$36018 ( \36396 , \25353 , \26143 );
and \U$36019 ( \36397 , \25348 , \26141 );
nor \U$36020 ( \36398 , \36396 , \36397 );
xnor \U$36021 ( \36399 , \36398 , \25911 );
and \U$36022 ( \36400 , \36394 , \36399 );
and \U$36023 ( \36401 , \36390 , \36399 );
or \U$36024 ( \36402 , \36395 , \36400 , \36401 );
and \U$36025 ( \36403 , \36386 , \36402 );
and \U$36026 ( \36404 , \27113 , \24661 );
and \U$36027 ( \36405 , \26854 , \24659 );
nor \U$36028 ( \36406 , \36404 , \36405 );
xnor \U$36029 ( \36407 , \36406 , \24456 );
and \U$36030 ( \36408 , \27494 , \24255 );
and \U$36031 ( \36409 , \27485 , \24253 );
nor \U$36032 ( \36410 , \36408 , \36409 );
xnor \U$36033 ( \36411 , \36410 , \24106 );
and \U$36034 ( \36412 , \36407 , \36411 );
and \U$36035 ( \36413 , \28039 , \23933 );
and \U$36036 ( \36414 , \27837 , \23931 );
nor \U$36037 ( \36415 , \36413 , \36414 );
xnor \U$36038 ( \36416 , \36415 , \23791 );
and \U$36039 ( \36417 , \36411 , \36416 );
and \U$36040 ( \36418 , \36407 , \36416 );
or \U$36041 ( \36419 , \36412 , \36417 , \36418 );
and \U$36042 ( \36420 , \36402 , \36419 );
and \U$36043 ( \36421 , \36386 , \36419 );
or \U$36044 ( \36422 , \36403 , \36420 , \36421 );
and \U$36045 ( \36423 , \36370 , \36422 );
and \U$36046 ( \36424 , \30318 , \22891 );
and \U$36047 ( \36425 , \30034 , \22889 );
nor \U$36048 ( \36426 , \36424 , \36425 );
xnor \U$36049 ( \36427 , \36426 , \22778 );
and \U$36050 ( \36428 , \30895 , \22697 );
and \U$36051 ( \36429 , \30887 , \22695 );
nor \U$36052 ( \36430 , \36428 , \36429 );
xnor \U$36053 ( \36431 , \36430 , \22561 );
and \U$36054 ( \36432 , \36427 , \36431 );
and \U$36055 ( \36433 , \31503 , \22497 );
and \U$36056 ( \36434 , \31498 , \22495 );
nor \U$36057 ( \36435 , \36433 , \36434 );
xnor \U$36058 ( \36436 , \36435 , \22419 );
and \U$36059 ( \36437 , \36431 , \36436 );
and \U$36060 ( \36438 , \36427 , \36436 );
or \U$36061 ( \36439 , \36432 , \36437 , \36438 );
and \U$36062 ( \36440 , \28514 , \23637 );
and \U$36063 ( \36441 , \28342 , \23635 );
nor \U$36064 ( \36442 , \36440 , \36441 );
xnor \U$36065 ( \36443 , \36442 , \23500 );
and \U$36066 ( \36444 , \29464 , \23431 );
and \U$36067 ( \36445 , \29040 , \23429 );
nor \U$36068 ( \36446 , \36444 , \36445 );
xnor \U$36069 ( \36447 , \36446 , \23279 );
and \U$36070 ( \36448 , \36443 , \36447 );
and \U$36071 ( \36449 , \29715 , \23163 );
and \U$36072 ( \36450 , \29710 , \23161 );
nor \U$36073 ( \36451 , \36449 , \36450 );
xnor \U$36074 ( \36452 , \36451 , \23007 );
and \U$36075 ( \36453 , \36447 , \36452 );
and \U$36076 ( \36454 , \36443 , \36452 );
or \U$36077 ( \36455 , \36448 , \36453 , \36454 );
and \U$36078 ( \36456 , \36439 , \36455 );
xor \U$36079 ( \36457 , \36170 , \36174 );
xor \U$36080 ( \36458 , \36457 , \36177 );
and \U$36081 ( \36459 , \36455 , \36458 );
and \U$36082 ( \36460 , \36439 , \36458 );
or \U$36083 ( \36461 , \36456 , \36459 , \36460 );
and \U$36084 ( \36462 , \36422 , \36461 );
and \U$36085 ( \36463 , \36370 , \36461 );
or \U$36086 ( \36464 , \36423 , \36462 , \36463 );
xor \U$36087 ( \36465 , \36154 , \36158 );
xor \U$36088 ( \36466 , \36465 , \36163 );
xor \U$36089 ( \36467 , \36086 , \36090 );
xor \U$36090 ( \36468 , \36467 , \36095 );
and \U$36091 ( \36469 , \36466 , \36468 );
xor \U$36092 ( \36470 , \36185 , \36189 );
xor \U$36093 ( \36471 , \36470 , \36194 );
and \U$36094 ( \36472 , \36468 , \36471 );
and \U$36095 ( \36473 , \36466 , \36471 );
or \U$36096 ( \36474 , \36469 , \36472 , \36473 );
xor \U$36097 ( \36475 , \36053 , \36057 );
xor \U$36098 ( \36476 , \36475 , \36062 );
xor \U$36099 ( \36477 , \36069 , \36073 );
xor \U$36100 ( \36478 , \36477 , \36078 );
and \U$36101 ( \36479 , \36476 , \36478 );
xor \U$36102 ( \36480 , \36105 , \36109 );
xor \U$36103 ( \36481 , \36480 , \36114 );
and \U$36104 ( \36482 , \36478 , \36481 );
and \U$36105 ( \36483 , \36476 , \36481 );
or \U$36106 ( \36484 , \36479 , \36482 , \36483 );
and \U$36107 ( \36485 , \36474 , \36484 );
xor \U$36108 ( \36486 , \36121 , \36125 );
xor \U$36109 ( \36487 , \36486 , \36130 );
xor \U$36110 ( \36488 , \36138 , \36142 );
xor \U$36111 ( \36489 , \36488 , \22091 );
and \U$36112 ( \36490 , \36487 , \36489 );
and \U$36113 ( \36491 , \36484 , \36490 );
and \U$36114 ( \36492 , \36474 , \36490 );
or \U$36115 ( \36493 , \36485 , \36491 , \36492 );
and \U$36116 ( \36494 , \36464 , \36493 );
xor \U$36117 ( \36495 , \36205 , \36207 );
xor \U$36118 ( \36496 , \36495 , \36210 );
xor \U$36119 ( \36497 , \36215 , \36217 );
xor \U$36120 ( \36498 , \36497 , \36220 );
and \U$36121 ( \36499 , \36496 , \36498 );
xor \U$36122 ( \36500 , \36226 , \36228 );
xor \U$36123 ( \36501 , \36500 , \36230 );
and \U$36124 ( \36502 , \36498 , \36501 );
and \U$36125 ( \36503 , \36496 , \36501 );
or \U$36126 ( \36504 , \36499 , \36502 , \36503 );
and \U$36127 ( \36505 , \36493 , \36504 );
and \U$36128 ( \36506 , \36464 , \36504 );
or \U$36129 ( \36507 , \36494 , \36505 , \36506 );
xor \U$36130 ( \36508 , \36065 , \36081 );
xor \U$36131 ( \36509 , \36508 , \36098 );
xor \U$36132 ( \36510 , \36117 , \36133 );
xor \U$36133 ( \36511 , \36510 , \36146 );
and \U$36134 ( \36512 , \36509 , \36511 );
xor \U$36135 ( \36513 , \36166 , \36180 );
xor \U$36136 ( \36514 , \36513 , \36197 );
and \U$36137 ( \36515 , \36511 , \36514 );
and \U$36138 ( \36516 , \36509 , \36514 );
or \U$36139 ( \36517 , \36512 , \36515 , \36516 );
xor \U$36140 ( \36518 , \35901 , \35917 );
xor \U$36141 ( \36519 , \36518 , \35934 );
and \U$36142 ( \36520 , \36517 , \36519 );
xor \U$36143 ( \36521 , \36252 , \36254 );
xor \U$36144 ( \36522 , \36521 , \36257 );
and \U$36145 ( \36523 , \36519 , \36522 );
and \U$36146 ( \36524 , \36517 , \36522 );
or \U$36147 ( \36525 , \36520 , \36523 , \36524 );
and \U$36148 ( \36526 , \36507 , \36525 );
xor \U$36149 ( \36527 , \36101 , \36149 );
xor \U$36150 ( \36528 , \36527 , \36200 );
xor \U$36151 ( \36529 , \36213 , \36223 );
xor \U$36152 ( \36530 , \36529 , \36233 );
and \U$36153 ( \36531 , \36528 , \36530 );
xor \U$36154 ( \36532 , \36239 , \36241 );
xor \U$36155 ( \36533 , \36532 , \36244 );
and \U$36156 ( \36534 , \36530 , \36533 );
and \U$36157 ( \36535 , \36528 , \36533 );
or \U$36158 ( \36536 , \36531 , \36534 , \36535 );
and \U$36159 ( \36537 , \36525 , \36536 );
and \U$36160 ( \36538 , \36507 , \36536 );
or \U$36161 ( \36539 , \36526 , \36537 , \36538 );
xor \U$36162 ( \36540 , \36203 , \36236 );
xor \U$36163 ( \36541 , \36540 , \36247 );
xor \U$36164 ( \36542 , \36260 , \36262 );
xor \U$36165 ( \36543 , \36542 , \36265 );
and \U$36166 ( \36544 , \36541 , \36543 );
xor \U$36167 ( \36545 , \36271 , \36273 );
and \U$36168 ( \36546 , \36543 , \36545 );
and \U$36169 ( \36547 , \36541 , \36545 );
or \U$36170 ( \36548 , \36544 , \36546 , \36547 );
and \U$36171 ( \36549 , \36539 , \36548 );
xor \U$36172 ( \36550 , \36279 , \36281 );
xor \U$36173 ( \36551 , \36550 , \36284 );
and \U$36174 ( \36552 , \36548 , \36551 );
and \U$36175 ( \36553 , \36539 , \36551 );
or \U$36176 ( \36554 , \36549 , \36552 , \36553 );
xor \U$36177 ( \36555 , \36277 , \36287 );
xor \U$36178 ( \36556 , \36555 , \36290 );
and \U$36179 ( \36557 , \36554 , \36556 );
xor \U$36180 ( \36558 , \36295 , \36297 );
and \U$36181 ( \36559 , \36556 , \36558 );
and \U$36182 ( \36560 , \36554 , \36558 );
or \U$36183 ( \36561 , \36557 , \36559 , \36560 );
and \U$36184 ( \36562 , \36318 , \36561 );
xor \U$36185 ( \36563 , \36318 , \36561 );
xor \U$36186 ( \36564 , \36554 , \36556 );
xor \U$36187 ( \36565 , \36564 , \36558 );
and \U$36188 ( \36566 , \23570 , \29104 );
and \U$36189 ( \36567 , \23384 , \29102 );
nor \U$36190 ( \36568 , \36566 , \36567 );
xnor \U$36191 ( \36569 , \36568 , \28855 );
and \U$36192 ( \36570 , \23978 , \28575 );
and \U$36193 ( \36571 , \23714 , \28573 );
nor \U$36194 ( \36572 , \36570 , \36571 );
xnor \U$36195 ( \36573 , \36572 , \28315 );
and \U$36196 ( \36574 , \36569 , \36573 );
and \U$36197 ( \36575 , \24177 , \28081 );
and \U$36198 ( \36576 , \24003 , \28079 );
nor \U$36199 ( \36577 , \36575 , \36576 );
xnor \U$36200 ( \36578 , \36577 , \27766 );
and \U$36201 ( \36579 , \36573 , \36578 );
and \U$36202 ( \36580 , \36569 , \36578 );
or \U$36203 ( \36581 , \36574 , \36579 , \36580 );
and \U$36204 ( \36582 , \22837 , \30770 );
and \U$36205 ( \36583 , \22721 , \30768 );
nor \U$36206 ( \36584 , \36582 , \36583 );
xnor \U$36207 ( \36585 , \36584 , \30460 );
and \U$36208 ( \36586 , \23128 , \30233 );
and \U$36209 ( \36587 , \22952 , \30231 );
nor \U$36210 ( \36588 , \36586 , \36587 );
xnor \U$36211 ( \36589 , \36588 , \29862 );
and \U$36212 ( \36590 , \36585 , \36589 );
and \U$36213 ( \36591 , \23379 , \29671 );
and \U$36214 ( \36592 , \23136 , \29669 );
nor \U$36215 ( \36593 , \36591 , \36592 );
xnor \U$36216 ( \36594 , \36593 , \29353 );
and \U$36217 ( \36595 , \36589 , \36594 );
and \U$36218 ( \36596 , \36585 , \36594 );
or \U$36219 ( \36597 , \36590 , \36595 , \36596 );
and \U$36220 ( \36598 , \36581 , \36597 );
and \U$36221 ( \36599 , \22523 , \32151 );
and \U$36222 ( \36600 , \22325 , \32148 );
nor \U$36223 ( \36601 , \36599 , \36600 );
xnor \U$36224 ( \36602 , \36601 , \31096 );
and \U$36225 ( \36603 , \22716 , \31338 );
and \U$36226 ( \36604 , \22611 , \31336 );
nor \U$36227 ( \36605 , \36603 , \36604 );
xnor \U$36228 ( \36606 , \36605 , \31099 );
and \U$36229 ( \36607 , \36602 , \36606 );
and \U$36230 ( \36608 , \36606 , \22239 );
and \U$36231 ( \36609 , \36602 , \22239 );
or \U$36232 ( \36610 , \36607 , \36608 , \36609 );
and \U$36233 ( \36611 , \36597 , \36610 );
and \U$36234 ( \36612 , \36581 , \36610 );
or \U$36235 ( \36613 , \36598 , \36611 , \36612 );
and \U$36236 ( \36614 , \28342 , \23933 );
and \U$36237 ( \36615 , \28039 , \23931 );
nor \U$36238 ( \36616 , \36614 , \36615 );
xnor \U$36239 ( \36617 , \36616 , \23791 );
and \U$36240 ( \36618 , \29040 , \23637 );
and \U$36241 ( \36619 , \28514 , \23635 );
nor \U$36242 ( \36620 , \36618 , \36619 );
xnor \U$36243 ( \36621 , \36620 , \23500 );
and \U$36244 ( \36622 , \36617 , \36621 );
and \U$36245 ( \36623 , \29710 , \23431 );
and \U$36246 ( \36624 , \29464 , \23429 );
nor \U$36247 ( \36625 , \36623 , \36624 );
xnor \U$36248 ( \36626 , \36625 , \23279 );
and \U$36249 ( \36627 , \36621 , \36626 );
and \U$36250 ( \36628 , \36617 , \36626 );
or \U$36251 ( \36629 , \36622 , \36627 , \36628 );
and \U$36252 ( \36630 , \30034 , \23163 );
and \U$36253 ( \36631 , \29715 , \23161 );
nor \U$36254 ( \36632 , \36630 , \36631 );
xnor \U$36255 ( \36633 , \36632 , \23007 );
and \U$36256 ( \36634 , \30887 , \22891 );
and \U$36257 ( \36635 , \30318 , \22889 );
nor \U$36258 ( \36636 , \36634 , \36635 );
xnor \U$36259 ( \36637 , \36636 , \22778 );
and \U$36260 ( \36638 , \36633 , \36637 );
and \U$36261 ( \36639 , \31498 , \22697 );
and \U$36262 ( \36640 , \30895 , \22695 );
nor \U$36263 ( \36641 , \36639 , \36640 );
xnor \U$36264 ( \36642 , \36641 , \22561 );
and \U$36265 ( \36643 , \36637 , \36642 );
and \U$36266 ( \36644 , \36633 , \36642 );
or \U$36267 ( \36645 , \36638 , \36643 , \36644 );
and \U$36268 ( \36646 , \36629 , \36645 );
and \U$36269 ( \36647 , \32304 , \22333 );
and \U$36270 ( \36648 , \31684 , \22331 );
nor \U$36271 ( \36649 , \36647 , \36648 );
xnor \U$36272 ( \36650 , \36649 , \22239 );
and \U$36273 ( \36651 , \36645 , \36650 );
and \U$36274 ( \36652 , \36629 , \36650 );
or \U$36275 ( \36653 , \36646 , \36651 , \36652 );
and \U$36276 ( \36654 , \36613 , \36653 );
and \U$36277 ( \36655 , \25609 , \26143 );
and \U$36278 ( \36656 , \25353 , \26141 );
nor \U$36279 ( \36657 , \36655 , \36656 );
xnor \U$36280 ( \36658 , \36657 , \25911 );
and \U$36281 ( \36659 , \26108 , \25692 );
and \U$36282 ( \36660 , \25806 , \25690 );
nor \U$36283 ( \36661 , \36659 , \36660 );
xnor \U$36284 ( \36662 , \36661 , \25549 );
and \U$36285 ( \36663 , \36658 , \36662 );
and \U$36286 ( \36664 , \26585 , \25369 );
and \U$36287 ( \36665 , \26116 , \25367 );
nor \U$36288 ( \36666 , \36664 , \36665 );
xnor \U$36289 ( \36667 , \36666 , \25123 );
and \U$36290 ( \36668 , \36662 , \36667 );
and \U$36291 ( \36669 , \36658 , \36667 );
or \U$36292 ( \36670 , \36663 , \36668 , \36669 );
and \U$36293 ( \36671 , \24482 , \27572 );
and \U$36294 ( \36672 , \24344 , \27570 );
nor \U$36295 ( \36673 , \36671 , \36672 );
xnor \U$36296 ( \36674 , \36673 , \27232 );
and \U$36297 ( \36675 , \25018 , \26983 );
and \U$36298 ( \36676 , \24601 , \26981 );
nor \U$36299 ( \36677 , \36675 , \36676 );
xnor \U$36300 ( \36678 , \36677 , \26742 );
and \U$36301 ( \36679 , \36674 , \36678 );
and \U$36302 ( \36680 , \25348 , \26517 );
and \U$36303 ( \36681 , \25226 , \26515 );
nor \U$36304 ( \36682 , \36680 , \36681 );
xnor \U$36305 ( \36683 , \36682 , \26329 );
and \U$36306 ( \36684 , \36678 , \36683 );
and \U$36307 ( \36685 , \36674 , \36683 );
or \U$36308 ( \36686 , \36679 , \36684 , \36685 );
and \U$36309 ( \36687 , \36670 , \36686 );
and \U$36310 ( \36688 , \26854 , \24974 );
and \U$36311 ( \36689 , \26590 , \24972 );
nor \U$36312 ( \36690 , \36688 , \36689 );
xnor \U$36313 ( \36691 , \36690 , \24787 );
and \U$36314 ( \36692 , \27485 , \24661 );
and \U$36315 ( \36693 , \27113 , \24659 );
nor \U$36316 ( \36694 , \36692 , \36693 );
xnor \U$36317 ( \36695 , \36694 , \24456 );
and \U$36318 ( \36696 , \36691 , \36695 );
and \U$36319 ( \36697 , \27837 , \24255 );
and \U$36320 ( \36698 , \27494 , \24253 );
nor \U$36321 ( \36699 , \36697 , \36698 );
xnor \U$36322 ( \36700 , \36699 , \24106 );
and \U$36323 ( \36701 , \36695 , \36700 );
and \U$36324 ( \36702 , \36691 , \36700 );
or \U$36325 ( \36703 , \36696 , \36701 , \36702 );
and \U$36326 ( \36704 , \36686 , \36703 );
and \U$36327 ( \36705 , \36670 , \36703 );
or \U$36328 ( \36706 , \36687 , \36704 , \36705 );
and \U$36329 ( \36707 , \36653 , \36706 );
and \U$36330 ( \36708 , \36613 , \36706 );
or \U$36331 ( \36709 , \36654 , \36707 , \36708 );
xor \U$36332 ( \36710 , \36427 , \36431 );
xor \U$36333 ( \36711 , \36710 , \36436 );
xor \U$36334 ( \36712 , \36407 , \36411 );
xor \U$36335 ( \36713 , \36712 , \36416 );
and \U$36336 ( \36714 , \36711 , \36713 );
xor \U$36337 ( \36715 , \36443 , \36447 );
xor \U$36338 ( \36716 , \36715 , \36452 );
and \U$36339 ( \36717 , \36713 , \36716 );
and \U$36340 ( \36718 , \36711 , \36716 );
or \U$36341 ( \36719 , \36714 , \36717 , \36718 );
xor \U$36342 ( \36720 , \36374 , \36378 );
xor \U$36343 ( \36721 , \36720 , \36383 );
xor \U$36344 ( \36722 , \36390 , \36394 );
xor \U$36345 ( \36723 , \36722 , \36399 );
and \U$36346 ( \36724 , \36721 , \36723 );
xor \U$36347 ( \36725 , \36322 , \36326 );
xor \U$36348 ( \36726 , \36725 , \36331 );
and \U$36349 ( \36727 , \36723 , \36726 );
and \U$36350 ( \36728 , \36721 , \36726 );
or \U$36351 ( \36729 , \36724 , \36727 , \36728 );
and \U$36352 ( \36730 , \36719 , \36729 );
xor \U$36353 ( \36731 , \36338 , \36342 );
xor \U$36354 ( \36732 , \36731 , \36347 );
xor \U$36355 ( \36733 , \36355 , \36359 );
xor \U$36356 ( \36734 , \36733 , \36364 );
and \U$36357 ( \36735 , \36732 , \36734 );
and \U$36358 ( \36736 , \36729 , \36735 );
and \U$36359 ( \36737 , \36719 , \36735 );
or \U$36360 ( \36738 , \36730 , \36736 , \36737 );
and \U$36361 ( \36739 , \36709 , \36738 );
xor \U$36362 ( \36740 , \36466 , \36468 );
xor \U$36363 ( \36741 , \36740 , \36471 );
xor \U$36364 ( \36742 , \36476 , \36478 );
xor \U$36365 ( \36743 , \36742 , \36481 );
and \U$36366 ( \36744 , \36741 , \36743 );
xor \U$36367 ( \36745 , \36487 , \36489 );
and \U$36368 ( \36746 , \36743 , \36745 );
and \U$36369 ( \36747 , \36741 , \36745 );
or \U$36370 ( \36748 , \36744 , \36746 , \36747 );
and \U$36371 ( \36749 , \36738 , \36748 );
and \U$36372 ( \36750 , \36709 , \36748 );
or \U$36373 ( \36751 , \36739 , \36749 , \36750 );
xor \U$36374 ( \36752 , \36334 , \36350 );
xor \U$36375 ( \36753 , \36752 , \36367 );
xor \U$36376 ( \36754 , \36386 , \36402 );
xor \U$36377 ( \36755 , \36754 , \36419 );
and \U$36378 ( \36756 , \36753 , \36755 );
xor \U$36379 ( \36757 , \36439 , \36455 );
xor \U$36380 ( \36758 , \36757 , \36458 );
and \U$36381 ( \36759 , \36755 , \36758 );
and \U$36382 ( \36760 , \36753 , \36758 );
or \U$36383 ( \36761 , \36756 , \36759 , \36760 );
xor \U$36384 ( \36762 , \36509 , \36511 );
xor \U$36385 ( \36763 , \36762 , \36514 );
and \U$36386 ( \36764 , \36761 , \36763 );
xor \U$36387 ( \36765 , \36496 , \36498 );
xor \U$36388 ( \36766 , \36765 , \36501 );
and \U$36389 ( \36767 , \36763 , \36766 );
and \U$36390 ( \36768 , \36761 , \36766 );
or \U$36391 ( \36769 , \36764 , \36767 , \36768 );
and \U$36392 ( \36770 , \36751 , \36769 );
xor \U$36393 ( \36771 , \36528 , \36530 );
xor \U$36394 ( \36772 , \36771 , \36533 );
and \U$36395 ( \36773 , \36769 , \36772 );
and \U$36396 ( \36774 , \36751 , \36772 );
or \U$36397 ( \36775 , \36770 , \36773 , \36774 );
xor \U$36398 ( \36776 , \36507 , \36525 );
xor \U$36399 ( \36777 , \36776 , \36536 );
and \U$36400 ( \36778 , \36775 , \36777 );
xor \U$36401 ( \36779 , \36541 , \36543 );
xor \U$36402 ( \36780 , \36779 , \36545 );
and \U$36403 ( \36781 , \36777 , \36780 );
and \U$36404 ( \36782 , \36775 , \36780 );
or \U$36405 ( \36783 , \36778 , \36781 , \36782 );
xor \U$36406 ( \36784 , \36250 , \36268 );
xor \U$36407 ( \36785 , \36784 , \36274 );
and \U$36408 ( \36786 , \36783 , \36785 );
xor \U$36409 ( \36787 , \36539 , \36548 );
xor \U$36410 ( \36788 , \36787 , \36551 );
and \U$36411 ( \36789 , \36785 , \36788 );
and \U$36412 ( \36790 , \36783 , \36788 );
or \U$36413 ( \36791 , \36786 , \36789 , \36790 );
and \U$36414 ( \36792 , \36565 , \36791 );
xor \U$36415 ( \36793 , \36565 , \36791 );
xor \U$36416 ( \36794 , \36783 , \36785 );
xor \U$36417 ( \36795 , \36794 , \36788 );
xor \U$36418 ( \36796 , \36569 , \36573 );
xor \U$36419 ( \36797 , \36796 , \36578 );
xor \U$36420 ( \36798 , \36585 , \36589 );
xor \U$36421 ( \36799 , \36798 , \36594 );
and \U$36422 ( \36800 , \36797 , \36799 );
xor \U$36423 ( \36801 , \36602 , \36606 );
xor \U$36424 ( \36802 , \36801 , \22239 );
and \U$36425 ( \36803 , \36799 , \36802 );
and \U$36426 ( \36804 , \36797 , \36802 );
or \U$36427 ( \36805 , \36800 , \36803 , \36804 );
nand \U$36428 ( \36806 , \32304 , \22331 );
xnor \U$36429 ( \36807 , \36806 , \22239 );
xor \U$36430 ( \36808 , \36617 , \36621 );
xor \U$36431 ( \36809 , \36808 , \36626 );
and \U$36432 ( \36810 , \36807 , \36809 );
xor \U$36433 ( \36811 , \36633 , \36637 );
xor \U$36434 ( \36812 , \36811 , \36642 );
and \U$36435 ( \36813 , \36809 , \36812 );
and \U$36436 ( \36814 , \36807 , \36812 );
or \U$36437 ( \36815 , \36810 , \36813 , \36814 );
and \U$36438 ( \36816 , \36805 , \36815 );
xor \U$36439 ( \36817 , \36658 , \36662 );
xor \U$36440 ( \36818 , \36817 , \36667 );
xor \U$36441 ( \36819 , \36674 , \36678 );
xor \U$36442 ( \36820 , \36819 , \36683 );
and \U$36443 ( \36821 , \36818 , \36820 );
xor \U$36444 ( \36822 , \36691 , \36695 );
xor \U$36445 ( \36823 , \36822 , \36700 );
and \U$36446 ( \36824 , \36820 , \36823 );
and \U$36447 ( \36825 , \36818 , \36823 );
or \U$36448 ( \36826 , \36821 , \36824 , \36825 );
and \U$36449 ( \36827 , \36815 , \36826 );
and \U$36450 ( \36828 , \36805 , \36826 );
or \U$36451 ( \36829 , \36816 , \36827 , \36828 );
and \U$36452 ( \36830 , \29464 , \23637 );
and \U$36453 ( \36831 , \29040 , \23635 );
nor \U$36454 ( \36832 , \36830 , \36831 );
xnor \U$36455 ( \36833 , \36832 , \23500 );
and \U$36456 ( \36834 , \29715 , \23431 );
and \U$36457 ( \36835 , \29710 , \23429 );
nor \U$36458 ( \36836 , \36834 , \36835 );
xnor \U$36459 ( \36837 , \36836 , \23279 );
and \U$36460 ( \36838 , \36833 , \36837 );
and \U$36461 ( \36839 , \30318 , \23163 );
and \U$36462 ( \36840 , \30034 , \23161 );
nor \U$36463 ( \36841 , \36839 , \36840 );
xnor \U$36464 ( \36842 , \36841 , \23007 );
and \U$36465 ( \36843 , \36837 , \36842 );
and \U$36466 ( \36844 , \36833 , \36842 );
or \U$36467 ( \36845 , \36838 , \36843 , \36844 );
and \U$36468 ( \36846 , \30895 , \22891 );
and \U$36469 ( \36847 , \30887 , \22889 );
nor \U$36470 ( \36848 , \36846 , \36847 );
xnor \U$36471 ( \36849 , \36848 , \22778 );
and \U$36472 ( \36850 , \31503 , \22697 );
and \U$36473 ( \36851 , \31498 , \22695 );
nor \U$36474 ( \36852 , \36850 , \36851 );
xnor \U$36475 ( \36853 , \36852 , \22561 );
and \U$36476 ( \36854 , \36849 , \36853 );
and \U$36477 ( \36855 , \32304 , \22497 );
and \U$36478 ( \36856 , \31684 , \22495 );
nor \U$36479 ( \36857 , \36855 , \36856 );
xnor \U$36480 ( \36858 , \36857 , \22419 );
and \U$36481 ( \36859 , \36853 , \36858 );
and \U$36482 ( \36860 , \36849 , \36858 );
or \U$36483 ( \36861 , \36854 , \36859 , \36860 );
and \U$36484 ( \36862 , \36845 , \36861 );
and \U$36485 ( \36863 , \31684 , \22497 );
and \U$36486 ( \36864 , \31503 , \22495 );
nor \U$36487 ( \36865 , \36863 , \36864 );
xnor \U$36488 ( \36866 , \36865 , \22419 );
and \U$36489 ( \36867 , \36861 , \36866 );
and \U$36490 ( \36868 , \36845 , \36866 );
or \U$36491 ( \36869 , \36862 , \36867 , \36868 );
and \U$36492 ( \36870 , \22611 , \32151 );
and \U$36493 ( \36871 , \22523 , \32148 );
nor \U$36494 ( \36872 , \36870 , \36871 );
xnor \U$36495 ( \36873 , \36872 , \31096 );
and \U$36496 ( \36874 , \22721 , \31338 );
and \U$36497 ( \36875 , \22716 , \31336 );
nor \U$36498 ( \36876 , \36874 , \36875 );
xnor \U$36499 ( \36877 , \36876 , \31099 );
and \U$36500 ( \36878 , \36873 , \36877 );
and \U$36501 ( \36879 , \22952 , \30770 );
and \U$36502 ( \36880 , \22837 , \30768 );
nor \U$36503 ( \36881 , \36879 , \36880 );
xnor \U$36504 ( \36882 , \36881 , \30460 );
and \U$36505 ( \36883 , \36877 , \36882 );
and \U$36506 ( \36884 , \36873 , \36882 );
or \U$36507 ( \36885 , \36878 , \36883 , \36884 );
and \U$36508 ( \36886 , \23136 , \30233 );
and \U$36509 ( \36887 , \23128 , \30231 );
nor \U$36510 ( \36888 , \36886 , \36887 );
xnor \U$36511 ( \36889 , \36888 , \29862 );
and \U$36512 ( \36890 , \23384 , \29671 );
and \U$36513 ( \36891 , \23379 , \29669 );
nor \U$36514 ( \36892 , \36890 , \36891 );
xnor \U$36515 ( \36893 , \36892 , \29353 );
and \U$36516 ( \36894 , \36889 , \36893 );
and \U$36517 ( \36895 , \23714 , \29104 );
and \U$36518 ( \36896 , \23570 , \29102 );
nor \U$36519 ( \36897 , \36895 , \36896 );
xnor \U$36520 ( \36898 , \36897 , \28855 );
and \U$36521 ( \36899 , \36893 , \36898 );
and \U$36522 ( \36900 , \36889 , \36898 );
or \U$36523 ( \36901 , \36894 , \36899 , \36900 );
and \U$36524 ( \36902 , \36885 , \36901 );
and \U$36525 ( \36903 , \24003 , \28575 );
and \U$36526 ( \36904 , \23978 , \28573 );
nor \U$36527 ( \36905 , \36903 , \36904 );
xnor \U$36528 ( \36906 , \36905 , \28315 );
and \U$36529 ( \36907 , \24344 , \28081 );
and \U$36530 ( \36908 , \24177 , \28079 );
nor \U$36531 ( \36909 , \36907 , \36908 );
xnor \U$36532 ( \36910 , \36909 , \27766 );
and \U$36533 ( \36911 , \36906 , \36910 );
and \U$36534 ( \36912 , \24601 , \27572 );
and \U$36535 ( \36913 , \24482 , \27570 );
nor \U$36536 ( \36914 , \36912 , \36913 );
xnor \U$36537 ( \36915 , \36914 , \27232 );
and \U$36538 ( \36916 , \36910 , \36915 );
and \U$36539 ( \36917 , \36906 , \36915 );
or \U$36540 ( \36918 , \36911 , \36916 , \36917 );
and \U$36541 ( \36919 , \36901 , \36918 );
and \U$36542 ( \36920 , \36885 , \36918 );
or \U$36543 ( \36921 , \36902 , \36919 , \36920 );
and \U$36544 ( \36922 , \36869 , \36921 );
and \U$36545 ( \36923 , \26116 , \25692 );
and \U$36546 ( \36924 , \26108 , \25690 );
nor \U$36547 ( \36925 , \36923 , \36924 );
xnor \U$36548 ( \36926 , \36925 , \25549 );
and \U$36549 ( \36927 , \26590 , \25369 );
and \U$36550 ( \36928 , \26585 , \25367 );
nor \U$36551 ( \36929 , \36927 , \36928 );
xnor \U$36552 ( \36930 , \36929 , \25123 );
and \U$36553 ( \36931 , \36926 , \36930 );
and \U$36554 ( \36932 , \27113 , \24974 );
and \U$36555 ( \36933 , \26854 , \24972 );
nor \U$36556 ( \36934 , \36932 , \36933 );
xnor \U$36557 ( \36935 , \36934 , \24787 );
and \U$36558 ( \36936 , \36930 , \36935 );
and \U$36559 ( \36937 , \36926 , \36935 );
or \U$36560 ( \36938 , \36931 , \36936 , \36937 );
and \U$36561 ( \36939 , \27494 , \24661 );
and \U$36562 ( \36940 , \27485 , \24659 );
nor \U$36563 ( \36941 , \36939 , \36940 );
xnor \U$36564 ( \36942 , \36941 , \24456 );
and \U$36565 ( \36943 , \28039 , \24255 );
and \U$36566 ( \36944 , \27837 , \24253 );
nor \U$36567 ( \36945 , \36943 , \36944 );
xnor \U$36568 ( \36946 , \36945 , \24106 );
and \U$36569 ( \36947 , \36942 , \36946 );
and \U$36570 ( \36948 , \28514 , \23933 );
and \U$36571 ( \36949 , \28342 , \23931 );
nor \U$36572 ( \36950 , \36948 , \36949 );
xnor \U$36573 ( \36951 , \36950 , \23791 );
and \U$36574 ( \36952 , \36946 , \36951 );
and \U$36575 ( \36953 , \36942 , \36951 );
or \U$36576 ( \36954 , \36947 , \36952 , \36953 );
and \U$36577 ( \36955 , \36938 , \36954 );
and \U$36578 ( \36956 , \25226 , \26983 );
and \U$36579 ( \36957 , \25018 , \26981 );
nor \U$36580 ( \36958 , \36956 , \36957 );
xnor \U$36581 ( \36959 , \36958 , \26742 );
and \U$36582 ( \36960 , \25353 , \26517 );
and \U$36583 ( \36961 , \25348 , \26515 );
nor \U$36584 ( \36962 , \36960 , \36961 );
xnor \U$36585 ( \36963 , \36962 , \26329 );
and \U$36586 ( \36964 , \36959 , \36963 );
and \U$36587 ( \36965 , \25806 , \26143 );
and \U$36588 ( \36966 , \25609 , \26141 );
nor \U$36589 ( \36967 , \36965 , \36966 );
xnor \U$36590 ( \36968 , \36967 , \25911 );
and \U$36591 ( \36969 , \36963 , \36968 );
and \U$36592 ( \36970 , \36959 , \36968 );
or \U$36593 ( \36971 , \36964 , \36969 , \36970 );
and \U$36594 ( \36972 , \36954 , \36971 );
and \U$36595 ( \36973 , \36938 , \36971 );
or \U$36596 ( \36974 , \36955 , \36972 , \36973 );
and \U$36597 ( \36975 , \36921 , \36974 );
and \U$36598 ( \36976 , \36869 , \36974 );
or \U$36599 ( \36977 , \36922 , \36975 , \36976 );
and \U$36600 ( \36978 , \36829 , \36977 );
xor \U$36601 ( \36979 , \36711 , \36713 );
xor \U$36602 ( \36980 , \36979 , \36716 );
xor \U$36603 ( \36981 , \36721 , \36723 );
xor \U$36604 ( \36982 , \36981 , \36726 );
and \U$36605 ( \36983 , \36980 , \36982 );
xor \U$36606 ( \36984 , \36732 , \36734 );
and \U$36607 ( \36985 , \36982 , \36984 );
and \U$36608 ( \36986 , \36980 , \36984 );
or \U$36609 ( \36987 , \36983 , \36985 , \36986 );
and \U$36610 ( \36988 , \36977 , \36987 );
and \U$36611 ( \36989 , \36829 , \36987 );
or \U$36612 ( \36990 , \36978 , \36988 , \36989 );
xor \U$36613 ( \36991 , \36581 , \36597 );
xor \U$36614 ( \36992 , \36991 , \36610 );
xor \U$36615 ( \36993 , \36629 , \36645 );
xor \U$36616 ( \36994 , \36993 , \36650 );
and \U$36617 ( \36995 , \36992 , \36994 );
xor \U$36618 ( \36996 , \36670 , \36686 );
xor \U$36619 ( \36997 , \36996 , \36703 );
and \U$36620 ( \36998 , \36994 , \36997 );
and \U$36621 ( \36999 , \36992 , \36997 );
or \U$36622 ( \37000 , \36995 , \36998 , \36999 );
xor \U$36623 ( \37001 , \36753 , \36755 );
xor \U$36624 ( \37002 , \37001 , \36758 );
and \U$36625 ( \37003 , \37000 , \37002 );
xor \U$36626 ( \37004 , \36741 , \36743 );
xor \U$36627 ( \37005 , \37004 , \36745 );
and \U$36628 ( \37006 , \37002 , \37005 );
and \U$36629 ( \37007 , \37000 , \37005 );
or \U$36630 ( \37008 , \37003 , \37006 , \37007 );
and \U$36631 ( \37009 , \36990 , \37008 );
xor \U$36632 ( \37010 , \36474 , \36484 );
xor \U$36633 ( \37011 , \37010 , \36490 );
and \U$36634 ( \37012 , \37008 , \37011 );
and \U$36635 ( \37013 , \36990 , \37011 );
or \U$36636 ( \37014 , \37009 , \37012 , \37013 );
xor \U$36637 ( \37015 , \36370 , \36422 );
xor \U$36638 ( \37016 , \37015 , \36461 );
xor \U$36639 ( \37017 , \36709 , \36738 );
xor \U$36640 ( \37018 , \37017 , \36748 );
and \U$36641 ( \37019 , \37016 , \37018 );
xor \U$36642 ( \37020 , \36761 , \36763 );
xor \U$36643 ( \37021 , \37020 , \36766 );
and \U$36644 ( \37022 , \37018 , \37021 );
and \U$36645 ( \37023 , \37016 , \37021 );
or \U$36646 ( \37024 , \37019 , \37022 , \37023 );
and \U$36647 ( \37025 , \37014 , \37024 );
xor \U$36648 ( \37026 , \36517 , \36519 );
xor \U$36649 ( \37027 , \37026 , \36522 );
and \U$36650 ( \37028 , \37024 , \37027 );
and \U$36651 ( \37029 , \37014 , \37027 );
or \U$36652 ( \37030 , \37025 , \37028 , \37029 );
xor \U$36653 ( \37031 , \36464 , \36493 );
xor \U$36654 ( \37032 , \37031 , \36504 );
xor \U$36655 ( \37033 , \36751 , \36769 );
xor \U$36656 ( \37034 , \37033 , \36772 );
and \U$36657 ( \37035 , \37032 , \37034 );
and \U$36658 ( \37036 , \37030 , \37035 );
xor \U$36659 ( \37037 , \36775 , \36777 );
xor \U$36660 ( \37038 , \37037 , \36780 );
and \U$36661 ( \37039 , \37035 , \37038 );
and \U$36662 ( \37040 , \37030 , \37038 );
or \U$36663 ( \37041 , \37036 , \37039 , \37040 );
and \U$36664 ( \37042 , \36795 , \37041 );
xor \U$36665 ( \37043 , \36795 , \37041 );
xor \U$36666 ( \37044 , \37030 , \37035 );
xor \U$36667 ( \37045 , \37044 , \37038 );
and \U$36668 ( \37046 , \27485 , \24974 );
and \U$36669 ( \37047 , \27113 , \24972 );
nor \U$36670 ( \37048 , \37046 , \37047 );
xnor \U$36671 ( \37049 , \37048 , \24787 );
and \U$36672 ( \37050 , \27837 , \24661 );
and \U$36673 ( \37051 , \27494 , \24659 );
nor \U$36674 ( \37052 , \37050 , \37051 );
xnor \U$36675 ( \37053 , \37052 , \24456 );
and \U$36676 ( \37054 , \37049 , \37053 );
and \U$36677 ( \37055 , \28342 , \24255 );
and \U$36678 ( \37056 , \28039 , \24253 );
nor \U$36679 ( \37057 , \37055 , \37056 );
xnor \U$36680 ( \37058 , \37057 , \24106 );
and \U$36681 ( \37059 , \37053 , \37058 );
and \U$36682 ( \37060 , \37049 , \37058 );
or \U$36683 ( \37061 , \37054 , \37059 , \37060 );
and \U$36684 ( \37062 , \26108 , \26143 );
and \U$36685 ( \37063 , \25806 , \26141 );
nor \U$36686 ( \37064 , \37062 , \37063 );
xnor \U$36687 ( \37065 , \37064 , \25911 );
and \U$36688 ( \37066 , \26585 , \25692 );
and \U$36689 ( \37067 , \26116 , \25690 );
nor \U$36690 ( \37068 , \37066 , \37067 );
xnor \U$36691 ( \37069 , \37068 , \25549 );
and \U$36692 ( \37070 , \37065 , \37069 );
and \U$36693 ( \37071 , \26854 , \25369 );
and \U$36694 ( \37072 , \26590 , \25367 );
nor \U$36695 ( \37073 , \37071 , \37072 );
xnor \U$36696 ( \37074 , \37073 , \25123 );
and \U$36697 ( \37075 , \37069 , \37074 );
and \U$36698 ( \37076 , \37065 , \37074 );
or \U$36699 ( \37077 , \37070 , \37075 , \37076 );
and \U$36700 ( \37078 , \37061 , \37077 );
and \U$36701 ( \37079 , \25018 , \27572 );
and \U$36702 ( \37080 , \24601 , \27570 );
nor \U$36703 ( \37081 , \37079 , \37080 );
xnor \U$36704 ( \37082 , \37081 , \27232 );
and \U$36705 ( \37083 , \25348 , \26983 );
and \U$36706 ( \37084 , \25226 , \26981 );
nor \U$36707 ( \37085 , \37083 , \37084 );
xnor \U$36708 ( \37086 , \37085 , \26742 );
and \U$36709 ( \37087 , \37082 , \37086 );
and \U$36710 ( \37088 , \25609 , \26517 );
and \U$36711 ( \37089 , \25353 , \26515 );
nor \U$36712 ( \37090 , \37088 , \37089 );
xnor \U$36713 ( \37091 , \37090 , \26329 );
and \U$36714 ( \37092 , \37086 , \37091 );
and \U$36715 ( \37093 , \37082 , \37091 );
or \U$36716 ( \37094 , \37087 , \37092 , \37093 );
and \U$36717 ( \37095 , \37077 , \37094 );
and \U$36718 ( \37096 , \37061 , \37094 );
or \U$36719 ( \37097 , \37078 , \37095 , \37096 );
and \U$36720 ( \37098 , \23128 , \30770 );
and \U$36721 ( \37099 , \22952 , \30768 );
nor \U$36722 ( \37100 , \37098 , \37099 );
xnor \U$36723 ( \37101 , \37100 , \30460 );
and \U$36724 ( \37102 , \23379 , \30233 );
and \U$36725 ( \37103 , \23136 , \30231 );
nor \U$36726 ( \37104 , \37102 , \37103 );
xnor \U$36727 ( \37105 , \37104 , \29862 );
and \U$36728 ( \37106 , \37101 , \37105 );
and \U$36729 ( \37107 , \23570 , \29671 );
and \U$36730 ( \37108 , \23384 , \29669 );
nor \U$36731 ( \37109 , \37107 , \37108 );
xnor \U$36732 ( \37110 , \37109 , \29353 );
and \U$36733 ( \37111 , \37105 , \37110 );
and \U$36734 ( \37112 , \37101 , \37110 );
or \U$36735 ( \37113 , \37106 , \37111 , \37112 );
and \U$36736 ( \37114 , \22716 , \32151 );
and \U$36737 ( \37115 , \22611 , \32148 );
nor \U$36738 ( \37116 , \37114 , \37115 );
xnor \U$36739 ( \37117 , \37116 , \31096 );
and \U$36740 ( \37118 , \22837 , \31338 );
and \U$36741 ( \37119 , \22721 , \31336 );
nor \U$36742 ( \37120 , \37118 , \37119 );
xnor \U$36743 ( \37121 , \37120 , \31099 );
and \U$36744 ( \37122 , \37117 , \37121 );
and \U$36745 ( \37123 , \37121 , \22419 );
and \U$36746 ( \37124 , \37117 , \22419 );
or \U$36747 ( \37125 , \37122 , \37123 , \37124 );
and \U$36748 ( \37126 , \37113 , \37125 );
and \U$36749 ( \37127 , \23978 , \29104 );
and \U$36750 ( \37128 , \23714 , \29102 );
nor \U$36751 ( \37129 , \37127 , \37128 );
xnor \U$36752 ( \37130 , \37129 , \28855 );
and \U$36753 ( \37131 , \24177 , \28575 );
and \U$36754 ( \37132 , \24003 , \28573 );
nor \U$36755 ( \37133 , \37131 , \37132 );
xnor \U$36756 ( \37134 , \37133 , \28315 );
and \U$36757 ( \37135 , \37130 , \37134 );
and \U$36758 ( \37136 , \24482 , \28081 );
and \U$36759 ( \37137 , \24344 , \28079 );
nor \U$36760 ( \37138 , \37136 , \37137 );
xnor \U$36761 ( \37139 , \37138 , \27766 );
and \U$36762 ( \37140 , \37134 , \37139 );
and \U$36763 ( \37141 , \37130 , \37139 );
or \U$36764 ( \37142 , \37135 , \37140 , \37141 );
and \U$36765 ( \37143 , \37125 , \37142 );
and \U$36766 ( \37144 , \37113 , \37142 );
or \U$36767 ( \37145 , \37126 , \37143 , \37144 );
and \U$36768 ( \37146 , \37097 , \37145 );
and \U$36769 ( \37147 , \29040 , \23933 );
and \U$36770 ( \37148 , \28514 , \23931 );
nor \U$36771 ( \37149 , \37147 , \37148 );
xnor \U$36772 ( \37150 , \37149 , \23791 );
and \U$36773 ( \37151 , \29710 , \23637 );
and \U$36774 ( \37152 , \29464 , \23635 );
nor \U$36775 ( \37153 , \37151 , \37152 );
xnor \U$36776 ( \37154 , \37153 , \23500 );
and \U$36777 ( \37155 , \37150 , \37154 );
and \U$36778 ( \37156 , \30034 , \23431 );
and \U$36779 ( \37157 , \29715 , \23429 );
nor \U$36780 ( \37158 , \37156 , \37157 );
xnor \U$36781 ( \37159 , \37158 , \23279 );
and \U$36782 ( \37160 , \37154 , \37159 );
and \U$36783 ( \37161 , \37150 , \37159 );
or \U$36784 ( \37162 , \37155 , \37160 , \37161 );
and \U$36785 ( \37163 , \30887 , \23163 );
and \U$36786 ( \37164 , \30318 , \23161 );
nor \U$36787 ( \37165 , \37163 , \37164 );
xnor \U$36788 ( \37166 , \37165 , \23007 );
and \U$36789 ( \37167 , \31498 , \22891 );
and \U$36790 ( \37168 , \30895 , \22889 );
nor \U$36791 ( \37169 , \37167 , \37168 );
xnor \U$36792 ( \37170 , \37169 , \22778 );
and \U$36793 ( \37171 , \37166 , \37170 );
and \U$36794 ( \37172 , \31684 , \22697 );
and \U$36795 ( \37173 , \31503 , \22695 );
nor \U$36796 ( \37174 , \37172 , \37173 );
xnor \U$36797 ( \37175 , \37174 , \22561 );
and \U$36798 ( \37176 , \37170 , \37175 );
and \U$36799 ( \37177 , \37166 , \37175 );
or \U$36800 ( \37178 , \37171 , \37176 , \37177 );
and \U$36801 ( \37179 , \37162 , \37178 );
xor \U$36802 ( \37180 , \36849 , \36853 );
xor \U$36803 ( \37181 , \37180 , \36858 );
and \U$36804 ( \37182 , \37178 , \37181 );
and \U$36805 ( \37183 , \37162 , \37181 );
or \U$36806 ( \37184 , \37179 , \37182 , \37183 );
and \U$36807 ( \37185 , \37145 , \37184 );
and \U$36808 ( \37186 , \37097 , \37184 );
or \U$36809 ( \37187 , \37146 , \37185 , \37186 );
xor \U$36810 ( \37188 , \36833 , \36837 );
xor \U$36811 ( \37189 , \37188 , \36842 );
xor \U$36812 ( \37190 , \36926 , \36930 );
xor \U$36813 ( \37191 , \37190 , \36935 );
and \U$36814 ( \37192 , \37189 , \37191 );
xor \U$36815 ( \37193 , \36942 , \36946 );
xor \U$36816 ( \37194 , \37193 , \36951 );
and \U$36817 ( \37195 , \37191 , \37194 );
and \U$36818 ( \37196 , \37189 , \37194 );
or \U$36819 ( \37197 , \37192 , \37195 , \37196 );
xor \U$36820 ( \37198 , \36889 , \36893 );
xor \U$36821 ( \37199 , \37198 , \36898 );
xor \U$36822 ( \37200 , \36959 , \36963 );
xor \U$36823 ( \37201 , \37200 , \36968 );
and \U$36824 ( \37202 , \37199 , \37201 );
xor \U$36825 ( \37203 , \36906 , \36910 );
xor \U$36826 ( \37204 , \37203 , \36915 );
and \U$36827 ( \37205 , \37201 , \37204 );
and \U$36828 ( \37206 , \37199 , \37204 );
or \U$36829 ( \37207 , \37202 , \37205 , \37206 );
and \U$36830 ( \37208 , \37197 , \37207 );
xor \U$36831 ( \37209 , \36797 , \36799 );
xor \U$36832 ( \37210 , \37209 , \36802 );
and \U$36833 ( \37211 , \37207 , \37210 );
and \U$36834 ( \37212 , \37197 , \37210 );
or \U$36835 ( \37213 , \37208 , \37211 , \37212 );
and \U$36836 ( \37214 , \37187 , \37213 );
xor \U$36837 ( \37215 , \36845 , \36861 );
xor \U$36838 ( \37216 , \37215 , \36866 );
xor \U$36839 ( \37217 , \36807 , \36809 );
xor \U$36840 ( \37218 , \37217 , \36812 );
and \U$36841 ( \37219 , \37216 , \37218 );
xor \U$36842 ( \37220 , \36818 , \36820 );
xor \U$36843 ( \37221 , \37220 , \36823 );
and \U$36844 ( \37222 , \37218 , \37221 );
and \U$36845 ( \37223 , \37216 , \37221 );
or \U$36846 ( \37224 , \37219 , \37222 , \37223 );
and \U$36847 ( \37225 , \37213 , \37224 );
and \U$36848 ( \37226 , \37187 , \37224 );
or \U$36849 ( \37227 , \37214 , \37225 , \37226 );
xor \U$36850 ( \37228 , \36805 , \36815 );
xor \U$36851 ( \37229 , \37228 , \36826 );
xor \U$36852 ( \37230 , \36992 , \36994 );
xor \U$36853 ( \37231 , \37230 , \36997 );
and \U$36854 ( \37232 , \37229 , \37231 );
xor \U$36855 ( \37233 , \36980 , \36982 );
xor \U$36856 ( \37234 , \37233 , \36984 );
and \U$36857 ( \37235 , \37231 , \37234 );
and \U$36858 ( \37236 , \37229 , \37234 );
or \U$36859 ( \37237 , \37232 , \37235 , \37236 );
and \U$36860 ( \37238 , \37227 , \37237 );
xor \U$36861 ( \37239 , \36719 , \36729 );
xor \U$36862 ( \37240 , \37239 , \36735 );
and \U$36863 ( \37241 , \37237 , \37240 );
and \U$36864 ( \37242 , \37227 , \37240 );
or \U$36865 ( \37243 , \37238 , \37241 , \37242 );
xor \U$36866 ( \37244 , \36613 , \36653 );
xor \U$36867 ( \37245 , \37244 , \36706 );
xor \U$36868 ( \37246 , \36829 , \36977 );
xor \U$36869 ( \37247 , \37246 , \36987 );
and \U$36870 ( \37248 , \37245 , \37247 );
xor \U$36871 ( \37249 , \37000 , \37002 );
xor \U$36872 ( \37250 , \37249 , \37005 );
and \U$36873 ( \37251 , \37247 , \37250 );
and \U$36874 ( \37252 , \37245 , \37250 );
or \U$36875 ( \37253 , \37248 , \37251 , \37252 );
and \U$36876 ( \37254 , \37243 , \37253 );
xor \U$36877 ( \37255 , \37016 , \37018 );
xor \U$36878 ( \37256 , \37255 , \37021 );
and \U$36879 ( \37257 , \37253 , \37256 );
and \U$36880 ( \37258 , \37243 , \37256 );
or \U$36881 ( \37259 , \37254 , \37257 , \37258 );
xor \U$36882 ( \37260 , \37014 , \37024 );
xor \U$36883 ( \37261 , \37260 , \37027 );
and \U$36884 ( \37262 , \37259 , \37261 );
xor \U$36885 ( \37263 , \37032 , \37034 );
and \U$36886 ( \37264 , \37261 , \37263 );
and \U$36887 ( \37265 , \37259 , \37263 );
or \U$36888 ( \37266 , \37262 , \37264 , \37265 );
and \U$36889 ( \37267 , \37045 , \37266 );
xor \U$36890 ( \37268 , \37045 , \37266 );
xor \U$36891 ( \37269 , \37259 , \37261 );
xor \U$36892 ( \37270 , \37269 , \37263 );
and \U$36893 ( \37271 , \25353 , \26983 );
and \U$36894 ( \37272 , \25348 , \26981 );
nor \U$36895 ( \37273 , \37271 , \37272 );
xnor \U$36896 ( \37274 , \37273 , \26742 );
and \U$36897 ( \37275 , \25806 , \26517 );
and \U$36898 ( \37276 , \25609 , \26515 );
nor \U$36899 ( \37277 , \37275 , \37276 );
xnor \U$36900 ( \37278 , \37277 , \26329 );
and \U$36901 ( \37279 , \37274 , \37278 );
and \U$36902 ( \37280 , \26116 , \26143 );
and \U$36903 ( \37281 , \26108 , \26141 );
nor \U$36904 ( \37282 , \37280 , \37281 );
xnor \U$36905 ( \37283 , \37282 , \25911 );
and \U$36906 ( \37284 , \37278 , \37283 );
and \U$36907 ( \37285 , \37274 , \37283 );
or \U$36908 ( \37286 , \37279 , \37284 , \37285 );
and \U$36909 ( \37287 , \26590 , \25692 );
and \U$36910 ( \37288 , \26585 , \25690 );
nor \U$36911 ( \37289 , \37287 , \37288 );
xnor \U$36912 ( \37290 , \37289 , \25549 );
and \U$36913 ( \37291 , \27113 , \25369 );
and \U$36914 ( \37292 , \26854 , \25367 );
nor \U$36915 ( \37293 , \37291 , \37292 );
xnor \U$36916 ( \37294 , \37293 , \25123 );
and \U$36917 ( \37295 , \37290 , \37294 );
and \U$36918 ( \37296 , \27494 , \24974 );
and \U$36919 ( \37297 , \27485 , \24972 );
nor \U$36920 ( \37298 , \37296 , \37297 );
xnor \U$36921 ( \37299 , \37298 , \24787 );
and \U$36922 ( \37300 , \37294 , \37299 );
and \U$36923 ( \37301 , \37290 , \37299 );
or \U$36924 ( \37302 , \37295 , \37300 , \37301 );
and \U$36925 ( \37303 , \37286 , \37302 );
and \U$36926 ( \37304 , \28039 , \24661 );
and \U$36927 ( \37305 , \27837 , \24659 );
nor \U$36928 ( \37306 , \37304 , \37305 );
xnor \U$36929 ( \37307 , \37306 , \24456 );
and \U$36930 ( \37308 , \28514 , \24255 );
and \U$36931 ( \37309 , \28342 , \24253 );
nor \U$36932 ( \37310 , \37308 , \37309 );
xnor \U$36933 ( \37311 , \37310 , \24106 );
and \U$36934 ( \37312 , \37307 , \37311 );
and \U$36935 ( \37313 , \29464 , \23933 );
and \U$36936 ( \37314 , \29040 , \23931 );
nor \U$36937 ( \37315 , \37313 , \37314 );
xnor \U$36938 ( \37316 , \37315 , \23791 );
and \U$36939 ( \37317 , \37311 , \37316 );
and \U$36940 ( \37318 , \37307 , \37316 );
or \U$36941 ( \37319 , \37312 , \37317 , \37318 );
and \U$36942 ( \37320 , \37302 , \37319 );
and \U$36943 ( \37321 , \37286 , \37319 );
or \U$36944 ( \37322 , \37303 , \37320 , \37321 );
and \U$36945 ( \37323 , \23384 , \30233 );
and \U$36946 ( \37324 , \23379 , \30231 );
nor \U$36947 ( \37325 , \37323 , \37324 );
xnor \U$36948 ( \37326 , \37325 , \29862 );
and \U$36949 ( \37327 , \23714 , \29671 );
and \U$36950 ( \37328 , \23570 , \29669 );
nor \U$36951 ( \37329 , \37327 , \37328 );
xnor \U$36952 ( \37330 , \37329 , \29353 );
and \U$36953 ( \37331 , \37326 , \37330 );
and \U$36954 ( \37332 , \24003 , \29104 );
and \U$36955 ( \37333 , \23978 , \29102 );
nor \U$36956 ( \37334 , \37332 , \37333 );
xnor \U$36957 ( \37335 , \37334 , \28855 );
and \U$36958 ( \37336 , \37330 , \37335 );
and \U$36959 ( \37337 , \37326 , \37335 );
or \U$36960 ( \37338 , \37331 , \37336 , \37337 );
and \U$36961 ( \37339 , \24344 , \28575 );
and \U$36962 ( \37340 , \24177 , \28573 );
nor \U$36963 ( \37341 , \37339 , \37340 );
xnor \U$36964 ( \37342 , \37341 , \28315 );
and \U$36965 ( \37343 , \24601 , \28081 );
and \U$36966 ( \37344 , \24482 , \28079 );
nor \U$36967 ( \37345 , \37343 , \37344 );
xnor \U$36968 ( \37346 , \37345 , \27766 );
and \U$36969 ( \37347 , \37342 , \37346 );
and \U$36970 ( \37348 , \25226 , \27572 );
and \U$36971 ( \37349 , \25018 , \27570 );
nor \U$36972 ( \37350 , \37348 , \37349 );
xnor \U$36973 ( \37351 , \37350 , \27232 );
and \U$36974 ( \37352 , \37346 , \37351 );
and \U$36975 ( \37353 , \37342 , \37351 );
or \U$36976 ( \37354 , \37347 , \37352 , \37353 );
and \U$36977 ( \37355 , \37338 , \37354 );
and \U$36978 ( \37356 , \22721 , \32151 );
and \U$36979 ( \37357 , \22716 , \32148 );
nor \U$36980 ( \37358 , \37356 , \37357 );
xnor \U$36981 ( \37359 , \37358 , \31096 );
and \U$36982 ( \37360 , \22952 , \31338 );
and \U$36983 ( \37361 , \22837 , \31336 );
nor \U$36984 ( \37362 , \37360 , \37361 );
xnor \U$36985 ( \37363 , \37362 , \31099 );
and \U$36986 ( \37364 , \37359 , \37363 );
and \U$36987 ( \37365 , \23136 , \30770 );
and \U$36988 ( \37366 , \23128 , \30768 );
nor \U$36989 ( \37367 , \37365 , \37366 );
xnor \U$36990 ( \37368 , \37367 , \30460 );
and \U$36991 ( \37369 , \37363 , \37368 );
and \U$36992 ( \37370 , \37359 , \37368 );
or \U$36993 ( \37371 , \37364 , \37369 , \37370 );
and \U$36994 ( \37372 , \37354 , \37371 );
and \U$36995 ( \37373 , \37338 , \37371 );
or \U$36996 ( \37374 , \37355 , \37372 , \37373 );
and \U$36997 ( \37375 , \37322 , \37374 );
and \U$36998 ( \37376 , \29715 , \23637 );
and \U$36999 ( \37377 , \29710 , \23635 );
nor \U$37000 ( \37378 , \37376 , \37377 );
xnor \U$37001 ( \37379 , \37378 , \23500 );
and \U$37002 ( \37380 , \30318 , \23431 );
and \U$37003 ( \37381 , \30034 , \23429 );
nor \U$37004 ( \37382 , \37380 , \37381 );
xnor \U$37005 ( \37383 , \37382 , \23279 );
and \U$37006 ( \37384 , \37379 , \37383 );
and \U$37007 ( \37385 , \30895 , \23163 );
and \U$37008 ( \37386 , \30887 , \23161 );
nor \U$37009 ( \37387 , \37385 , \37386 );
xnor \U$37010 ( \37388 , \37387 , \23007 );
and \U$37011 ( \37389 , \37383 , \37388 );
and \U$37012 ( \37390 , \37379 , \37388 );
or \U$37013 ( \37391 , \37384 , \37389 , \37390 );
nand \U$37014 ( \37392 , \32304 , \22495 );
xnor \U$37015 ( \37393 , \37392 , \22419 );
and \U$37016 ( \37394 , \37391 , \37393 );
xor \U$37017 ( \37395 , \37166 , \37170 );
xor \U$37018 ( \37396 , \37395 , \37175 );
and \U$37019 ( \37397 , \37393 , \37396 );
and \U$37020 ( \37398 , \37391 , \37396 );
or \U$37021 ( \37399 , \37394 , \37397 , \37398 );
and \U$37022 ( \37400 , \37374 , \37399 );
and \U$37023 ( \37401 , \37322 , \37399 );
or \U$37024 ( \37402 , \37375 , \37400 , \37401 );
xor \U$37025 ( \37403 , \37049 , \37053 );
xor \U$37026 ( \37404 , \37403 , \37058 );
xor \U$37027 ( \37405 , \37150 , \37154 );
xor \U$37028 ( \37406 , \37405 , \37159 );
and \U$37029 ( \37407 , \37404 , \37406 );
xor \U$37030 ( \37408 , \37065 , \37069 );
xor \U$37031 ( \37409 , \37408 , \37074 );
and \U$37032 ( \37410 , \37406 , \37409 );
and \U$37033 ( \37411 , \37404 , \37409 );
or \U$37034 ( \37412 , \37407 , \37410 , \37411 );
xor \U$37035 ( \37413 , \37101 , \37105 );
xor \U$37036 ( \37414 , \37413 , \37110 );
xor \U$37037 ( \37415 , \37082 , \37086 );
xor \U$37038 ( \37416 , \37415 , \37091 );
and \U$37039 ( \37417 , \37414 , \37416 );
xor \U$37040 ( \37418 , \37130 , \37134 );
xor \U$37041 ( \37419 , \37418 , \37139 );
and \U$37042 ( \37420 , \37416 , \37419 );
and \U$37043 ( \37421 , \37414 , \37419 );
or \U$37044 ( \37422 , \37417 , \37420 , \37421 );
and \U$37045 ( \37423 , \37412 , \37422 );
xor \U$37046 ( \37424 , \36873 , \36877 );
xor \U$37047 ( \37425 , \37424 , \36882 );
and \U$37048 ( \37426 , \37422 , \37425 );
and \U$37049 ( \37427 , \37412 , \37425 );
or \U$37050 ( \37428 , \37423 , \37426 , \37427 );
and \U$37051 ( \37429 , \37402 , \37428 );
xor \U$37052 ( \37430 , \37189 , \37191 );
xor \U$37053 ( \37431 , \37430 , \37194 );
xor \U$37054 ( \37432 , \37199 , \37201 );
xor \U$37055 ( \37433 , \37432 , \37204 );
and \U$37056 ( \37434 , \37431 , \37433 );
xor \U$37057 ( \37435 , \37162 , \37178 );
xor \U$37058 ( \37436 , \37435 , \37181 );
and \U$37059 ( \37437 , \37433 , \37436 );
and \U$37060 ( \37438 , \37431 , \37436 );
or \U$37061 ( \37439 , \37434 , \37437 , \37438 );
and \U$37062 ( \37440 , \37428 , \37439 );
and \U$37063 ( \37441 , \37402 , \37439 );
or \U$37064 ( \37442 , \37429 , \37440 , \37441 );
xor \U$37065 ( \37443 , \36885 , \36901 );
xor \U$37066 ( \37444 , \37443 , \36918 );
xor \U$37067 ( \37445 , \36938 , \36954 );
xor \U$37068 ( \37446 , \37445 , \36971 );
and \U$37069 ( \37447 , \37444 , \37446 );
xor \U$37070 ( \37448 , \37216 , \37218 );
xor \U$37071 ( \37449 , \37448 , \37221 );
and \U$37072 ( \37450 , \37446 , \37449 );
and \U$37073 ( \37451 , \37444 , \37449 );
or \U$37074 ( \37452 , \37447 , \37450 , \37451 );
and \U$37075 ( \37453 , \37442 , \37452 );
xor \U$37076 ( \37454 , \37097 , \37145 );
xor \U$37077 ( \37455 , \37454 , \37184 );
xor \U$37078 ( \37456 , \37197 , \37207 );
xor \U$37079 ( \37457 , \37456 , \37210 );
and \U$37080 ( \37458 , \37455 , \37457 );
and \U$37081 ( \37459 , \37452 , \37458 );
and \U$37082 ( \37460 , \37442 , \37458 );
or \U$37083 ( \37461 , \37453 , \37459 , \37460 );
xor \U$37084 ( \37462 , \36869 , \36921 );
xor \U$37085 ( \37463 , \37462 , \36974 );
xor \U$37086 ( \37464 , \37187 , \37213 );
xor \U$37087 ( \37465 , \37464 , \37224 );
and \U$37088 ( \37466 , \37463 , \37465 );
xor \U$37089 ( \37467 , \37229 , \37231 );
xor \U$37090 ( \37468 , \37467 , \37234 );
and \U$37091 ( \37469 , \37465 , \37468 );
and \U$37092 ( \37470 , \37463 , \37468 );
or \U$37093 ( \37471 , \37466 , \37469 , \37470 );
and \U$37094 ( \37472 , \37461 , \37471 );
xor \U$37095 ( \37473 , \37245 , \37247 );
xor \U$37096 ( \37474 , \37473 , \37250 );
and \U$37097 ( \37475 , \37471 , \37474 );
and \U$37098 ( \37476 , \37461 , \37474 );
or \U$37099 ( \37477 , \37472 , \37475 , \37476 );
xor \U$37100 ( \37478 , \36990 , \37008 );
xor \U$37101 ( \37479 , \37478 , \37011 );
and \U$37102 ( \37480 , \37477 , \37479 );
xor \U$37103 ( \37481 , \37243 , \37253 );
xor \U$37104 ( \37482 , \37481 , \37256 );
and \U$37105 ( \37483 , \37479 , \37482 );
and \U$37106 ( \37484 , \37477 , \37482 );
or \U$37107 ( \37485 , \37480 , \37483 , \37484 );
and \U$37108 ( \37486 , \37270 , \37485 );
xor \U$37109 ( \37487 , \37270 , \37485 );
xor \U$37110 ( \37488 , \37477 , \37479 );
xor \U$37111 ( \37489 , \37488 , \37482 );
and \U$37112 ( \37490 , \22837 , \32151 );
and \U$37113 ( \37491 , \22721 , \32148 );
nor \U$37114 ( \37492 , \37490 , \37491 );
xnor \U$37115 ( \37493 , \37492 , \31096 );
and \U$37116 ( \37494 , \23128 , \31338 );
and \U$37117 ( \37495 , \22952 , \31336 );
nor \U$37118 ( \37496 , \37494 , \37495 );
xnor \U$37119 ( \37497 , \37496 , \31099 );
and \U$37120 ( \37498 , \37493 , \37497 );
and \U$37121 ( \37499 , \37497 , \22561 );
and \U$37122 ( \37500 , \37493 , \22561 );
or \U$37123 ( \37501 , \37498 , \37499 , \37500 );
and \U$37124 ( \37502 , \24177 , \29104 );
and \U$37125 ( \37503 , \24003 , \29102 );
nor \U$37126 ( \37504 , \37502 , \37503 );
xnor \U$37127 ( \37505 , \37504 , \28855 );
and \U$37128 ( \37506 , \24482 , \28575 );
and \U$37129 ( \37507 , \24344 , \28573 );
nor \U$37130 ( \37508 , \37506 , \37507 );
xnor \U$37131 ( \37509 , \37508 , \28315 );
and \U$37132 ( \37510 , \37505 , \37509 );
and \U$37133 ( \37511 , \25018 , \28081 );
and \U$37134 ( \37512 , \24601 , \28079 );
nor \U$37135 ( \37513 , \37511 , \37512 );
xnor \U$37136 ( \37514 , \37513 , \27766 );
and \U$37137 ( \37515 , \37509 , \37514 );
and \U$37138 ( \37516 , \37505 , \37514 );
or \U$37139 ( \37517 , \37510 , \37515 , \37516 );
and \U$37140 ( \37518 , \37501 , \37517 );
and \U$37141 ( \37519 , \23379 , \30770 );
and \U$37142 ( \37520 , \23136 , \30768 );
nor \U$37143 ( \37521 , \37519 , \37520 );
xnor \U$37144 ( \37522 , \37521 , \30460 );
and \U$37145 ( \37523 , \23570 , \30233 );
and \U$37146 ( \37524 , \23384 , \30231 );
nor \U$37147 ( \37525 , \37523 , \37524 );
xnor \U$37148 ( \37526 , \37525 , \29862 );
and \U$37149 ( \37527 , \37522 , \37526 );
and \U$37150 ( \37528 , \23978 , \29671 );
and \U$37151 ( \37529 , \23714 , \29669 );
nor \U$37152 ( \37530 , \37528 , \37529 );
xnor \U$37153 ( \37531 , \37530 , \29353 );
and \U$37154 ( \37532 , \37526 , \37531 );
and \U$37155 ( \37533 , \37522 , \37531 );
or \U$37156 ( \37534 , \37527 , \37532 , \37533 );
and \U$37157 ( \37535 , \37517 , \37534 );
and \U$37158 ( \37536 , \37501 , \37534 );
or \U$37159 ( \37537 , \37518 , \37535 , \37536 );
and \U$37160 ( \37538 , \25348 , \27572 );
and \U$37161 ( \37539 , \25226 , \27570 );
nor \U$37162 ( \37540 , \37538 , \37539 );
xnor \U$37163 ( \37541 , \37540 , \27232 );
and \U$37164 ( \37542 , \25609 , \26983 );
and \U$37165 ( \37543 , \25353 , \26981 );
nor \U$37166 ( \37544 , \37542 , \37543 );
xnor \U$37167 ( \37545 , \37544 , \26742 );
and \U$37168 ( \37546 , \37541 , \37545 );
and \U$37169 ( \37547 , \26108 , \26517 );
and \U$37170 ( \37548 , \25806 , \26515 );
nor \U$37171 ( \37549 , \37547 , \37548 );
xnor \U$37172 ( \37550 , \37549 , \26329 );
and \U$37173 ( \37551 , \37545 , \37550 );
and \U$37174 ( \37552 , \37541 , \37550 );
or \U$37175 ( \37553 , \37546 , \37551 , \37552 );
and \U$37176 ( \37554 , \26585 , \26143 );
and \U$37177 ( \37555 , \26116 , \26141 );
nor \U$37178 ( \37556 , \37554 , \37555 );
xnor \U$37179 ( \37557 , \37556 , \25911 );
and \U$37180 ( \37558 , \26854 , \25692 );
and \U$37181 ( \37559 , \26590 , \25690 );
nor \U$37182 ( \37560 , \37558 , \37559 );
xnor \U$37183 ( \37561 , \37560 , \25549 );
and \U$37184 ( \37562 , \37557 , \37561 );
and \U$37185 ( \37563 , \27485 , \25369 );
and \U$37186 ( \37564 , \27113 , \25367 );
nor \U$37187 ( \37565 , \37563 , \37564 );
xnor \U$37188 ( \37566 , \37565 , \25123 );
and \U$37189 ( \37567 , \37561 , \37566 );
and \U$37190 ( \37568 , \37557 , \37566 );
or \U$37191 ( \37569 , \37562 , \37567 , \37568 );
and \U$37192 ( \37570 , \37553 , \37569 );
and \U$37193 ( \37571 , \27837 , \24974 );
and \U$37194 ( \37572 , \27494 , \24972 );
nor \U$37195 ( \37573 , \37571 , \37572 );
xnor \U$37196 ( \37574 , \37573 , \24787 );
and \U$37197 ( \37575 , \28342 , \24661 );
and \U$37198 ( \37576 , \28039 , \24659 );
nor \U$37199 ( \37577 , \37575 , \37576 );
xnor \U$37200 ( \37578 , \37577 , \24456 );
and \U$37201 ( \37579 , \37574 , \37578 );
and \U$37202 ( \37580 , \29040 , \24255 );
and \U$37203 ( \37581 , \28514 , \24253 );
nor \U$37204 ( \37582 , \37580 , \37581 );
xnor \U$37205 ( \37583 , \37582 , \24106 );
and \U$37206 ( \37584 , \37578 , \37583 );
and \U$37207 ( \37585 , \37574 , \37583 );
or \U$37208 ( \37586 , \37579 , \37584 , \37585 );
and \U$37209 ( \37587 , \37569 , \37586 );
and \U$37210 ( \37588 , \37553 , \37586 );
or \U$37211 ( \37589 , \37570 , \37587 , \37588 );
and \U$37212 ( \37590 , \37537 , \37589 );
and \U$37213 ( \37591 , \31498 , \23163 );
and \U$37214 ( \37592 , \30895 , \23161 );
nor \U$37215 ( \37593 , \37591 , \37592 );
xnor \U$37216 ( \37594 , \37593 , \23007 );
and \U$37217 ( \37595 , \31684 , \22891 );
and \U$37218 ( \37596 , \31503 , \22889 );
nor \U$37219 ( \37597 , \37595 , \37596 );
xnor \U$37220 ( \37598 , \37597 , \22778 );
and \U$37221 ( \37599 , \37594 , \37598 );
nand \U$37222 ( \37600 , \32304 , \22695 );
xnor \U$37223 ( \37601 , \37600 , \22561 );
and \U$37224 ( \37602 , \37598 , \37601 );
and \U$37225 ( \37603 , \37594 , \37601 );
or \U$37226 ( \37604 , \37599 , \37602 , \37603 );
and \U$37227 ( \37605 , \29710 , \23933 );
and \U$37228 ( \37606 , \29464 , \23931 );
nor \U$37229 ( \37607 , \37605 , \37606 );
xnor \U$37230 ( \37608 , \37607 , \23791 );
and \U$37231 ( \37609 , \30034 , \23637 );
and \U$37232 ( \37610 , \29715 , \23635 );
nor \U$37233 ( \37611 , \37609 , \37610 );
xnor \U$37234 ( \37612 , \37611 , \23500 );
and \U$37235 ( \37613 , \37608 , \37612 );
and \U$37236 ( \37614 , \30887 , \23431 );
and \U$37237 ( \37615 , \30318 , \23429 );
nor \U$37238 ( \37616 , \37614 , \37615 );
xnor \U$37239 ( \37617 , \37616 , \23279 );
and \U$37240 ( \37618 , \37612 , \37617 );
and \U$37241 ( \37619 , \37608 , \37617 );
or \U$37242 ( \37620 , \37613 , \37618 , \37619 );
and \U$37243 ( \37621 , \37604 , \37620 );
and \U$37244 ( \37622 , \31503 , \22891 );
and \U$37245 ( \37623 , \31498 , \22889 );
nor \U$37246 ( \37624 , \37622 , \37623 );
xnor \U$37247 ( \37625 , \37624 , \22778 );
and \U$37248 ( \37626 , \37620 , \37625 );
and \U$37249 ( \37627 , \37604 , \37625 );
or \U$37250 ( \37628 , \37621 , \37626 , \37627 );
and \U$37251 ( \37629 , \37589 , \37628 );
and \U$37252 ( \37630 , \37537 , \37628 );
or \U$37253 ( \37631 , \37590 , \37629 , \37630 );
and \U$37254 ( \37632 , \32304 , \22697 );
and \U$37255 ( \37633 , \31684 , \22695 );
nor \U$37256 ( \37634 , \37632 , \37633 );
xnor \U$37257 ( \37635 , \37634 , \22561 );
xor \U$37258 ( \37636 , \37307 , \37311 );
xor \U$37259 ( \37637 , \37636 , \37316 );
and \U$37260 ( \37638 , \37635 , \37637 );
xor \U$37261 ( \37639 , \37379 , \37383 );
xor \U$37262 ( \37640 , \37639 , \37388 );
and \U$37263 ( \37641 , \37637 , \37640 );
and \U$37264 ( \37642 , \37635 , \37640 );
or \U$37265 ( \37643 , \37638 , \37641 , \37642 );
xor \U$37266 ( \37644 , \37274 , \37278 );
xor \U$37267 ( \37645 , \37644 , \37283 );
xor \U$37268 ( \37646 , \37290 , \37294 );
xor \U$37269 ( \37647 , \37646 , \37299 );
and \U$37270 ( \37648 , \37645 , \37647 );
xor \U$37271 ( \37649 , \37342 , \37346 );
xor \U$37272 ( \37650 , \37649 , \37351 );
and \U$37273 ( \37651 , \37647 , \37650 );
and \U$37274 ( \37652 , \37645 , \37650 );
or \U$37275 ( \37653 , \37648 , \37651 , \37652 );
and \U$37276 ( \37654 , \37643 , \37653 );
xor \U$37277 ( \37655 , \37117 , \37121 );
xor \U$37278 ( \37656 , \37655 , \22419 );
and \U$37279 ( \37657 , \37653 , \37656 );
and \U$37280 ( \37658 , \37643 , \37656 );
or \U$37281 ( \37659 , \37654 , \37657 , \37658 );
and \U$37282 ( \37660 , \37631 , \37659 );
xor \U$37283 ( \37661 , \37391 , \37393 );
xor \U$37284 ( \37662 , \37661 , \37396 );
xor \U$37285 ( \37663 , \37404 , \37406 );
xor \U$37286 ( \37664 , \37663 , \37409 );
and \U$37287 ( \37665 , \37662 , \37664 );
xor \U$37288 ( \37666 , \37414 , \37416 );
xor \U$37289 ( \37667 , \37666 , \37419 );
and \U$37290 ( \37668 , \37664 , \37667 );
and \U$37291 ( \37669 , \37662 , \37667 );
or \U$37292 ( \37670 , \37665 , \37668 , \37669 );
and \U$37293 ( \37671 , \37659 , \37670 );
and \U$37294 ( \37672 , \37631 , \37670 );
or \U$37295 ( \37673 , \37660 , \37671 , \37672 );
xor \U$37296 ( \37674 , \37061 , \37077 );
xor \U$37297 ( \37675 , \37674 , \37094 );
xor \U$37298 ( \37676 , \37113 , \37125 );
xor \U$37299 ( \37677 , \37676 , \37142 );
and \U$37300 ( \37678 , \37675 , \37677 );
xor \U$37301 ( \37679 , \37431 , \37433 );
xor \U$37302 ( \37680 , \37679 , \37436 );
and \U$37303 ( \37681 , \37677 , \37680 );
and \U$37304 ( \37682 , \37675 , \37680 );
or \U$37305 ( \37683 , \37678 , \37681 , \37682 );
and \U$37306 ( \37684 , \37673 , \37683 );
xor \U$37307 ( \37685 , \37322 , \37374 );
xor \U$37308 ( \37686 , \37685 , \37399 );
xor \U$37309 ( \37687 , \37412 , \37422 );
xor \U$37310 ( \37688 , \37687 , \37425 );
and \U$37311 ( \37689 , \37686 , \37688 );
and \U$37312 ( \37690 , \37683 , \37689 );
and \U$37313 ( \37691 , \37673 , \37689 );
or \U$37314 ( \37692 , \37684 , \37690 , \37691 );
xor \U$37315 ( \37693 , \37402 , \37428 );
xor \U$37316 ( \37694 , \37693 , \37439 );
xor \U$37317 ( \37695 , \37444 , \37446 );
xor \U$37318 ( \37696 , \37695 , \37449 );
and \U$37319 ( \37697 , \37694 , \37696 );
xor \U$37320 ( \37698 , \37455 , \37457 );
and \U$37321 ( \37699 , \37696 , \37698 );
and \U$37322 ( \37700 , \37694 , \37698 );
or \U$37323 ( \37701 , \37697 , \37699 , \37700 );
and \U$37324 ( \37702 , \37692 , \37701 );
xor \U$37325 ( \37703 , \37463 , \37465 );
xor \U$37326 ( \37704 , \37703 , \37468 );
and \U$37327 ( \37705 , \37701 , \37704 );
and \U$37328 ( \37706 , \37692 , \37704 );
or \U$37329 ( \37707 , \37702 , \37705 , \37706 );
xor \U$37330 ( \37708 , \37227 , \37237 );
xor \U$37331 ( \37709 , \37708 , \37240 );
and \U$37332 ( \37710 , \37707 , \37709 );
xor \U$37333 ( \37711 , \37461 , \37471 );
xor \U$37334 ( \37712 , \37711 , \37474 );
and \U$37335 ( \37713 , \37709 , \37712 );
and \U$37336 ( \37714 , \37707 , \37712 );
or \U$37337 ( \37715 , \37710 , \37713 , \37714 );
and \U$37338 ( \37716 , \37489 , \37715 );
xor \U$37339 ( \37717 , \37489 , \37715 );
xor \U$37340 ( \37718 , \37707 , \37709 );
xor \U$37341 ( \37719 , \37718 , \37712 );
and \U$37342 ( \37720 , \22952 , \32151 );
and \U$37343 ( \37721 , \22837 , \32148 );
nor \U$37344 ( \37722 , \37720 , \37721 );
xnor \U$37345 ( \37723 , \37722 , \31096 );
and \U$37346 ( \37724 , \23136 , \31338 );
and \U$37347 ( \37725 , \23128 , \31336 );
nor \U$37348 ( \37726 , \37724 , \37725 );
xnor \U$37349 ( \37727 , \37726 , \31099 );
and \U$37350 ( \37728 , \37723 , \37727 );
and \U$37351 ( \37729 , \23384 , \30770 );
and \U$37352 ( \37730 , \23379 , \30768 );
nor \U$37353 ( \37731 , \37729 , \37730 );
xnor \U$37354 ( \37732 , \37731 , \30460 );
and \U$37355 ( \37733 , \37727 , \37732 );
and \U$37356 ( \37734 , \37723 , \37732 );
or \U$37357 ( \37735 , \37728 , \37733 , \37734 );
and \U$37358 ( \37736 , \23714 , \30233 );
and \U$37359 ( \37737 , \23570 , \30231 );
nor \U$37360 ( \37738 , \37736 , \37737 );
xnor \U$37361 ( \37739 , \37738 , \29862 );
and \U$37362 ( \37740 , \24003 , \29671 );
and \U$37363 ( \37741 , \23978 , \29669 );
nor \U$37364 ( \37742 , \37740 , \37741 );
xnor \U$37365 ( \37743 , \37742 , \29353 );
and \U$37366 ( \37744 , \37739 , \37743 );
and \U$37367 ( \37745 , \24344 , \29104 );
and \U$37368 ( \37746 , \24177 , \29102 );
nor \U$37369 ( \37747 , \37745 , \37746 );
xnor \U$37370 ( \37748 , \37747 , \28855 );
and \U$37371 ( \37749 , \37743 , \37748 );
and \U$37372 ( \37750 , \37739 , \37748 );
or \U$37373 ( \37751 , \37744 , \37749 , \37750 );
and \U$37374 ( \37752 , \37735 , \37751 );
and \U$37375 ( \37753 , \24601 , \28575 );
and \U$37376 ( \37754 , \24482 , \28573 );
nor \U$37377 ( \37755 , \37753 , \37754 );
xnor \U$37378 ( \37756 , \37755 , \28315 );
and \U$37379 ( \37757 , \25226 , \28081 );
and \U$37380 ( \37758 , \25018 , \28079 );
nor \U$37381 ( \37759 , \37757 , \37758 );
xnor \U$37382 ( \37760 , \37759 , \27766 );
and \U$37383 ( \37761 , \37756 , \37760 );
and \U$37384 ( \37762 , \25353 , \27572 );
and \U$37385 ( \37763 , \25348 , \27570 );
nor \U$37386 ( \37764 , \37762 , \37763 );
xnor \U$37387 ( \37765 , \37764 , \27232 );
and \U$37388 ( \37766 , \37760 , \37765 );
and \U$37389 ( \37767 , \37756 , \37765 );
or \U$37390 ( \37768 , \37761 , \37766 , \37767 );
and \U$37391 ( \37769 , \37751 , \37768 );
and \U$37392 ( \37770 , \37735 , \37768 );
or \U$37393 ( \37771 , \37752 , \37769 , \37770 );
and \U$37394 ( \37772 , \27113 , \25692 );
and \U$37395 ( \37773 , \26854 , \25690 );
nor \U$37396 ( \37774 , \37772 , \37773 );
xnor \U$37397 ( \37775 , \37774 , \25549 );
and \U$37398 ( \37776 , \27494 , \25369 );
and \U$37399 ( \37777 , \27485 , \25367 );
nor \U$37400 ( \37778 , \37776 , \37777 );
xnor \U$37401 ( \37779 , \37778 , \25123 );
and \U$37402 ( \37780 , \37775 , \37779 );
and \U$37403 ( \37781 , \28039 , \24974 );
and \U$37404 ( \37782 , \27837 , \24972 );
nor \U$37405 ( \37783 , \37781 , \37782 );
xnor \U$37406 ( \37784 , \37783 , \24787 );
and \U$37407 ( \37785 , \37779 , \37784 );
and \U$37408 ( \37786 , \37775 , \37784 );
or \U$37409 ( \37787 , \37780 , \37785 , \37786 );
and \U$37410 ( \37788 , \28514 , \24661 );
and \U$37411 ( \37789 , \28342 , \24659 );
nor \U$37412 ( \37790 , \37788 , \37789 );
xnor \U$37413 ( \37791 , \37790 , \24456 );
and \U$37414 ( \37792 , \29464 , \24255 );
and \U$37415 ( \37793 , \29040 , \24253 );
nor \U$37416 ( \37794 , \37792 , \37793 );
xnor \U$37417 ( \37795 , \37794 , \24106 );
and \U$37418 ( \37796 , \37791 , \37795 );
and \U$37419 ( \37797 , \29715 , \23933 );
and \U$37420 ( \37798 , \29710 , \23931 );
nor \U$37421 ( \37799 , \37797 , \37798 );
xnor \U$37422 ( \37800 , \37799 , \23791 );
and \U$37423 ( \37801 , \37795 , \37800 );
and \U$37424 ( \37802 , \37791 , \37800 );
or \U$37425 ( \37803 , \37796 , \37801 , \37802 );
and \U$37426 ( \37804 , \37787 , \37803 );
and \U$37427 ( \37805 , \25806 , \26983 );
and \U$37428 ( \37806 , \25609 , \26981 );
nor \U$37429 ( \37807 , \37805 , \37806 );
xnor \U$37430 ( \37808 , \37807 , \26742 );
and \U$37431 ( \37809 , \26116 , \26517 );
and \U$37432 ( \37810 , \26108 , \26515 );
nor \U$37433 ( \37811 , \37809 , \37810 );
xnor \U$37434 ( \37812 , \37811 , \26329 );
and \U$37435 ( \37813 , \37808 , \37812 );
and \U$37436 ( \37814 , \26590 , \26143 );
and \U$37437 ( \37815 , \26585 , \26141 );
nor \U$37438 ( \37816 , \37814 , \37815 );
xnor \U$37439 ( \37817 , \37816 , \25911 );
and \U$37440 ( \37818 , \37812 , \37817 );
and \U$37441 ( \37819 , \37808 , \37817 );
or \U$37442 ( \37820 , \37813 , \37818 , \37819 );
and \U$37443 ( \37821 , \37803 , \37820 );
and \U$37444 ( \37822 , \37787 , \37820 );
or \U$37445 ( \37823 , \37804 , \37821 , \37822 );
and \U$37446 ( \37824 , \37771 , \37823 );
and \U$37447 ( \37825 , \30318 , \23637 );
and \U$37448 ( \37826 , \30034 , \23635 );
nor \U$37449 ( \37827 , \37825 , \37826 );
xnor \U$37450 ( \37828 , \37827 , \23500 );
and \U$37451 ( \37829 , \30895 , \23431 );
and \U$37452 ( \37830 , \30887 , \23429 );
nor \U$37453 ( \37831 , \37829 , \37830 );
xnor \U$37454 ( \37832 , \37831 , \23279 );
and \U$37455 ( \37833 , \37828 , \37832 );
and \U$37456 ( \37834 , \31503 , \23163 );
and \U$37457 ( \37835 , \31498 , \23161 );
nor \U$37458 ( \37836 , \37834 , \37835 );
xnor \U$37459 ( \37837 , \37836 , \23007 );
and \U$37460 ( \37838 , \37832 , \37837 );
and \U$37461 ( \37839 , \37828 , \37837 );
or \U$37462 ( \37840 , \37833 , \37838 , \37839 );
xor \U$37463 ( \37841 , \37594 , \37598 );
xor \U$37464 ( \37842 , \37841 , \37601 );
and \U$37465 ( \37843 , \37840 , \37842 );
xor \U$37466 ( \37844 , \37608 , \37612 );
xor \U$37467 ( \37845 , \37844 , \37617 );
and \U$37468 ( \37846 , \37842 , \37845 );
and \U$37469 ( \37847 , \37840 , \37845 );
or \U$37470 ( \37848 , \37843 , \37846 , \37847 );
and \U$37471 ( \37849 , \37823 , \37848 );
and \U$37472 ( \37850 , \37771 , \37848 );
or \U$37473 ( \37851 , \37824 , \37849 , \37850 );
xor \U$37474 ( \37852 , \37541 , \37545 );
xor \U$37475 ( \37853 , \37852 , \37550 );
xor \U$37476 ( \37854 , \37557 , \37561 );
xor \U$37477 ( \37855 , \37854 , \37566 );
and \U$37478 ( \37856 , \37853 , \37855 );
xor \U$37479 ( \37857 , \37574 , \37578 );
xor \U$37480 ( \37858 , \37857 , \37583 );
and \U$37481 ( \37859 , \37855 , \37858 );
and \U$37482 ( \37860 , \37853 , \37858 );
or \U$37483 ( \37861 , \37856 , \37859 , \37860 );
xor \U$37484 ( \37862 , \37493 , \37497 );
xor \U$37485 ( \37863 , \37862 , \22561 );
xor \U$37486 ( \37864 , \37505 , \37509 );
xor \U$37487 ( \37865 , \37864 , \37514 );
and \U$37488 ( \37866 , \37863 , \37865 );
xor \U$37489 ( \37867 , \37522 , \37526 );
xor \U$37490 ( \37868 , \37867 , \37531 );
and \U$37491 ( \37869 , \37865 , \37868 );
and \U$37492 ( \37870 , \37863 , \37868 );
or \U$37493 ( \37871 , \37866 , \37869 , \37870 );
and \U$37494 ( \37872 , \37861 , \37871 );
xor \U$37495 ( \37873 , \37326 , \37330 );
xor \U$37496 ( \37874 , \37873 , \37335 );
and \U$37497 ( \37875 , \37871 , \37874 );
and \U$37498 ( \37876 , \37861 , \37874 );
or \U$37499 ( \37877 , \37872 , \37875 , \37876 );
and \U$37500 ( \37878 , \37851 , \37877 );
xor \U$37501 ( \37879 , \37359 , \37363 );
xor \U$37502 ( \37880 , \37879 , \37368 );
xor \U$37503 ( \37881 , \37635 , \37637 );
xor \U$37504 ( \37882 , \37881 , \37640 );
and \U$37505 ( \37883 , \37880 , \37882 );
xor \U$37506 ( \37884 , \37645 , \37647 );
xor \U$37507 ( \37885 , \37884 , \37650 );
and \U$37508 ( \37886 , \37882 , \37885 );
and \U$37509 ( \37887 , \37880 , \37885 );
or \U$37510 ( \37888 , \37883 , \37886 , \37887 );
and \U$37511 ( \37889 , \37877 , \37888 );
and \U$37512 ( \37890 , \37851 , \37888 );
or \U$37513 ( \37891 , \37878 , \37889 , \37890 );
xor \U$37514 ( \37892 , \37501 , \37517 );
xor \U$37515 ( \37893 , \37892 , \37534 );
xor \U$37516 ( \37894 , \37553 , \37569 );
xor \U$37517 ( \37895 , \37894 , \37586 );
and \U$37518 ( \37896 , \37893 , \37895 );
xor \U$37519 ( \37897 , \37604 , \37620 );
xor \U$37520 ( \37898 , \37897 , \37625 );
and \U$37521 ( \37899 , \37895 , \37898 );
and \U$37522 ( \37900 , \37893 , \37898 );
or \U$37523 ( \37901 , \37896 , \37899 , \37900 );
xor \U$37524 ( \37902 , \37286 , \37302 );
xor \U$37525 ( \37903 , \37902 , \37319 );
and \U$37526 ( \37904 , \37901 , \37903 );
xor \U$37527 ( \37905 , \37338 , \37354 );
xor \U$37528 ( \37906 , \37905 , \37371 );
and \U$37529 ( \37907 , \37903 , \37906 );
and \U$37530 ( \37908 , \37901 , \37906 );
or \U$37531 ( \37909 , \37904 , \37907 , \37908 );
and \U$37532 ( \37910 , \37891 , \37909 );
xor \U$37533 ( \37911 , \37537 , \37589 );
xor \U$37534 ( \37912 , \37911 , \37628 );
xor \U$37535 ( \37913 , \37643 , \37653 );
xor \U$37536 ( \37914 , \37913 , \37656 );
and \U$37537 ( \37915 , \37912 , \37914 );
xor \U$37538 ( \37916 , \37662 , \37664 );
xor \U$37539 ( \37917 , \37916 , \37667 );
and \U$37540 ( \37918 , \37914 , \37917 );
and \U$37541 ( \37919 , \37912 , \37917 );
or \U$37542 ( \37920 , \37915 , \37918 , \37919 );
and \U$37543 ( \37921 , \37909 , \37920 );
and \U$37544 ( \37922 , \37891 , \37920 );
or \U$37545 ( \37923 , \37910 , \37921 , \37922 );
xor \U$37546 ( \37924 , \37631 , \37659 );
xor \U$37547 ( \37925 , \37924 , \37670 );
xor \U$37548 ( \37926 , \37675 , \37677 );
xor \U$37549 ( \37927 , \37926 , \37680 );
and \U$37550 ( \37928 , \37925 , \37927 );
xor \U$37551 ( \37929 , \37686 , \37688 );
and \U$37552 ( \37930 , \37927 , \37929 );
and \U$37553 ( \37931 , \37925 , \37929 );
or \U$37554 ( \37932 , \37928 , \37930 , \37931 );
and \U$37555 ( \37933 , \37923 , \37932 );
xor \U$37556 ( \37934 , \37694 , \37696 );
xor \U$37557 ( \37935 , \37934 , \37698 );
and \U$37558 ( \37936 , \37932 , \37935 );
and \U$37559 ( \37937 , \37923 , \37935 );
or \U$37560 ( \37938 , \37933 , \37936 , \37937 );
xor \U$37561 ( \37939 , \37442 , \37452 );
xor \U$37562 ( \37940 , \37939 , \37458 );
and \U$37563 ( \37941 , \37938 , \37940 );
xor \U$37564 ( \37942 , \37692 , \37701 );
xor \U$37565 ( \37943 , \37942 , \37704 );
and \U$37566 ( \37944 , \37940 , \37943 );
and \U$37567 ( \37945 , \37938 , \37943 );
or \U$37568 ( \37946 , \37941 , \37944 , \37945 );
and \U$37569 ( \37947 , \37719 , \37946 );
xor \U$37570 ( \37948 , \37719 , \37946 );
xor \U$37571 ( \37949 , \37938 , \37940 );
xor \U$37572 ( \37950 , \37949 , \37943 );
and \U$37573 ( \37951 , \28342 , \24974 );
and \U$37574 ( \37952 , \28039 , \24972 );
nor \U$37575 ( \37953 , \37951 , \37952 );
xnor \U$37576 ( \37954 , \37953 , \24787 );
and \U$37577 ( \37955 , \29040 , \24661 );
and \U$37578 ( \37956 , \28514 , \24659 );
nor \U$37579 ( \37957 , \37955 , \37956 );
xnor \U$37580 ( \37958 , \37957 , \24456 );
and \U$37581 ( \37959 , \37954 , \37958 );
and \U$37582 ( \37960 , \29710 , \24255 );
and \U$37583 ( \37961 , \29464 , \24253 );
nor \U$37584 ( \37962 , \37960 , \37961 );
xnor \U$37585 ( \37963 , \37962 , \24106 );
and \U$37586 ( \37964 , \37958 , \37963 );
and \U$37587 ( \37965 , \37954 , \37963 );
or \U$37588 ( \37966 , \37959 , \37964 , \37965 );
and \U$37589 ( \37967 , \25609 , \27572 );
and \U$37590 ( \37968 , \25353 , \27570 );
nor \U$37591 ( \37969 , \37967 , \37968 );
xnor \U$37592 ( \37970 , \37969 , \27232 );
and \U$37593 ( \37971 , \26108 , \26983 );
and \U$37594 ( \37972 , \25806 , \26981 );
nor \U$37595 ( \37973 , \37971 , \37972 );
xnor \U$37596 ( \37974 , \37973 , \26742 );
and \U$37597 ( \37975 , \37970 , \37974 );
and \U$37598 ( \37976 , \26585 , \26517 );
and \U$37599 ( \37977 , \26116 , \26515 );
nor \U$37600 ( \37978 , \37976 , \37977 );
xnor \U$37601 ( \37979 , \37978 , \26329 );
and \U$37602 ( \37980 , \37974 , \37979 );
and \U$37603 ( \37981 , \37970 , \37979 );
or \U$37604 ( \37982 , \37975 , \37980 , \37981 );
and \U$37605 ( \37983 , \37966 , \37982 );
and \U$37606 ( \37984 , \26854 , \26143 );
and \U$37607 ( \37985 , \26590 , \26141 );
nor \U$37608 ( \37986 , \37984 , \37985 );
xnor \U$37609 ( \37987 , \37986 , \25911 );
and \U$37610 ( \37988 , \27485 , \25692 );
and \U$37611 ( \37989 , \27113 , \25690 );
nor \U$37612 ( \37990 , \37988 , \37989 );
xnor \U$37613 ( \37991 , \37990 , \25549 );
and \U$37614 ( \37992 , \37987 , \37991 );
and \U$37615 ( \37993 , \27837 , \25369 );
and \U$37616 ( \37994 , \27494 , \25367 );
nor \U$37617 ( \37995 , \37993 , \37994 );
xnor \U$37618 ( \37996 , \37995 , \25123 );
and \U$37619 ( \37997 , \37991 , \37996 );
and \U$37620 ( \37998 , \37987 , \37996 );
or \U$37621 ( \37999 , \37992 , \37997 , \37998 );
and \U$37622 ( \38000 , \37982 , \37999 );
and \U$37623 ( \38001 , \37966 , \37999 );
or \U$37624 ( \38002 , \37983 , \38000 , \38001 );
and \U$37625 ( \38003 , \23128 , \32151 );
and \U$37626 ( \38004 , \22952 , \32148 );
nor \U$37627 ( \38005 , \38003 , \38004 );
xnor \U$37628 ( \38006 , \38005 , \31096 );
and \U$37629 ( \38007 , \23379 , \31338 );
and \U$37630 ( \38008 , \23136 , \31336 );
nor \U$37631 ( \38009 , \38007 , \38008 );
xnor \U$37632 ( \38010 , \38009 , \31099 );
and \U$37633 ( \38011 , \38006 , \38010 );
and \U$37634 ( \38012 , \38010 , \22778 );
and \U$37635 ( \38013 , \38006 , \22778 );
or \U$37636 ( \38014 , \38011 , \38012 , \38013 );
and \U$37637 ( \38015 , \24482 , \29104 );
and \U$37638 ( \38016 , \24344 , \29102 );
nor \U$37639 ( \38017 , \38015 , \38016 );
xnor \U$37640 ( \38018 , \38017 , \28855 );
and \U$37641 ( \38019 , \25018 , \28575 );
and \U$37642 ( \38020 , \24601 , \28573 );
nor \U$37643 ( \38021 , \38019 , \38020 );
xnor \U$37644 ( \38022 , \38021 , \28315 );
and \U$37645 ( \38023 , \38018 , \38022 );
and \U$37646 ( \38024 , \25348 , \28081 );
and \U$37647 ( \38025 , \25226 , \28079 );
nor \U$37648 ( \38026 , \38024 , \38025 );
xnor \U$37649 ( \38027 , \38026 , \27766 );
and \U$37650 ( \38028 , \38022 , \38027 );
and \U$37651 ( \38029 , \38018 , \38027 );
or \U$37652 ( \38030 , \38023 , \38028 , \38029 );
and \U$37653 ( \38031 , \38014 , \38030 );
and \U$37654 ( \38032 , \23570 , \30770 );
and \U$37655 ( \38033 , \23384 , \30768 );
nor \U$37656 ( \38034 , \38032 , \38033 );
xnor \U$37657 ( \38035 , \38034 , \30460 );
and \U$37658 ( \38036 , \23978 , \30233 );
and \U$37659 ( \38037 , \23714 , \30231 );
nor \U$37660 ( \38038 , \38036 , \38037 );
xnor \U$37661 ( \38039 , \38038 , \29862 );
and \U$37662 ( \38040 , \38035 , \38039 );
and \U$37663 ( \38041 , \24177 , \29671 );
and \U$37664 ( \38042 , \24003 , \29669 );
nor \U$37665 ( \38043 , \38041 , \38042 );
xnor \U$37666 ( \38044 , \38043 , \29353 );
and \U$37667 ( \38045 , \38039 , \38044 );
and \U$37668 ( \38046 , \38035 , \38044 );
or \U$37669 ( \38047 , \38040 , \38045 , \38046 );
and \U$37670 ( \38048 , \38030 , \38047 );
and \U$37671 ( \38049 , \38014 , \38047 );
or \U$37672 ( \38050 , \38031 , \38048 , \38049 );
and \U$37673 ( \38051 , \38002 , \38050 );
and \U$37674 ( \38052 , \30034 , \23933 );
and \U$37675 ( \38053 , \29715 , \23931 );
nor \U$37676 ( \38054 , \38052 , \38053 );
xnor \U$37677 ( \38055 , \38054 , \23791 );
and \U$37678 ( \38056 , \30887 , \23637 );
and \U$37679 ( \38057 , \30318 , \23635 );
nor \U$37680 ( \38058 , \38056 , \38057 );
xnor \U$37681 ( \38059 , \38058 , \23500 );
and \U$37682 ( \38060 , \38055 , \38059 );
and \U$37683 ( \38061 , \31498 , \23431 );
and \U$37684 ( \38062 , \30895 , \23429 );
nor \U$37685 ( \38063 , \38061 , \38062 );
xnor \U$37686 ( \38064 , \38063 , \23279 );
and \U$37687 ( \38065 , \38059 , \38064 );
and \U$37688 ( \38066 , \38055 , \38064 );
or \U$37689 ( \38067 , \38060 , \38065 , \38066 );
and \U$37690 ( \38068 , \31684 , \23163 );
and \U$37691 ( \38069 , \31503 , \23161 );
nor \U$37692 ( \38070 , \38068 , \38069 );
xnor \U$37693 ( \38071 , \38070 , \23007 );
nand \U$37694 ( \38072 , \32304 , \22889 );
xnor \U$37695 ( \38073 , \38072 , \22778 );
and \U$37696 ( \38074 , \38071 , \38073 );
and \U$37697 ( \38075 , \38067 , \38074 );
and \U$37698 ( \38076 , \32304 , \22891 );
and \U$37699 ( \38077 , \31684 , \22889 );
nor \U$37700 ( \38078 , \38076 , \38077 );
xnor \U$37701 ( \38079 , \38078 , \22778 );
and \U$37702 ( \38080 , \38074 , \38079 );
and \U$37703 ( \38081 , \38067 , \38079 );
or \U$37704 ( \38082 , \38075 , \38080 , \38081 );
and \U$37705 ( \38083 , \38050 , \38082 );
and \U$37706 ( \38084 , \38002 , \38082 );
or \U$37707 ( \38085 , \38051 , \38083 , \38084 );
xor \U$37708 ( \38086 , \37739 , \37743 );
xor \U$37709 ( \38087 , \38086 , \37748 );
xor \U$37710 ( \38088 , \37808 , \37812 );
xor \U$37711 ( \38089 , \38088 , \37817 );
and \U$37712 ( \38090 , \38087 , \38089 );
xor \U$37713 ( \38091 , \37756 , \37760 );
xor \U$37714 ( \38092 , \38091 , \37765 );
and \U$37715 ( \38093 , \38089 , \38092 );
and \U$37716 ( \38094 , \38087 , \38092 );
or \U$37717 ( \38095 , \38090 , \38093 , \38094 );
xor \U$37718 ( \38096 , \37775 , \37779 );
xor \U$37719 ( \38097 , \38096 , \37784 );
xor \U$37720 ( \38098 , \37828 , \37832 );
xor \U$37721 ( \38099 , \38098 , \37837 );
and \U$37722 ( \38100 , \38097 , \38099 );
xor \U$37723 ( \38101 , \37791 , \37795 );
xor \U$37724 ( \38102 , \38101 , \37800 );
and \U$37725 ( \38103 , \38099 , \38102 );
and \U$37726 ( \38104 , \38097 , \38102 );
or \U$37727 ( \38105 , \38100 , \38103 , \38104 );
and \U$37728 ( \38106 , \38095 , \38105 );
xor \U$37729 ( \38107 , \37863 , \37865 );
xor \U$37730 ( \38108 , \38107 , \37868 );
and \U$37731 ( \38109 , \38105 , \38108 );
and \U$37732 ( \38110 , \38095 , \38108 );
or \U$37733 ( \38111 , \38106 , \38109 , \38110 );
and \U$37734 ( \38112 , \38085 , \38111 );
xor \U$37735 ( \38113 , \37787 , \37803 );
xor \U$37736 ( \38114 , \38113 , \37820 );
xor \U$37737 ( \38115 , \37853 , \37855 );
xor \U$37738 ( \38116 , \38115 , \37858 );
and \U$37739 ( \38117 , \38114 , \38116 );
xor \U$37740 ( \38118 , \37840 , \37842 );
xor \U$37741 ( \38119 , \38118 , \37845 );
and \U$37742 ( \38120 , \38116 , \38119 );
and \U$37743 ( \38121 , \38114 , \38119 );
or \U$37744 ( \38122 , \38117 , \38120 , \38121 );
and \U$37745 ( \38123 , \38111 , \38122 );
and \U$37746 ( \38124 , \38085 , \38122 );
or \U$37747 ( \38125 , \38112 , \38123 , \38124 );
xor \U$37748 ( \38126 , \37893 , \37895 );
xor \U$37749 ( \38127 , \38126 , \37898 );
xor \U$37750 ( \38128 , \37861 , \37871 );
xor \U$37751 ( \38129 , \38128 , \37874 );
and \U$37752 ( \38130 , \38127 , \38129 );
xor \U$37753 ( \38131 , \37880 , \37882 );
xor \U$37754 ( \38132 , \38131 , \37885 );
and \U$37755 ( \38133 , \38129 , \38132 );
and \U$37756 ( \38134 , \38127 , \38132 );
or \U$37757 ( \38135 , \38130 , \38133 , \38134 );
and \U$37758 ( \38136 , \38125 , \38135 );
xor \U$37759 ( \38137 , \37912 , \37914 );
xor \U$37760 ( \38138 , \38137 , \37917 );
and \U$37761 ( \38139 , \38135 , \38138 );
and \U$37762 ( \38140 , \38125 , \38138 );
or \U$37763 ( \38141 , \38136 , \38139 , \38140 );
xor \U$37764 ( \38142 , \37891 , \37909 );
xor \U$37765 ( \38143 , \38142 , \37920 );
and \U$37766 ( \38144 , \38141 , \38143 );
xor \U$37767 ( \38145 , \37925 , \37927 );
xor \U$37768 ( \38146 , \38145 , \37929 );
and \U$37769 ( \38147 , \38143 , \38146 );
and \U$37770 ( \38148 , \38141 , \38146 );
or \U$37771 ( \38149 , \38144 , \38147 , \38148 );
xor \U$37772 ( \38150 , \37673 , \37683 );
xor \U$37773 ( \38151 , \38150 , \37689 );
and \U$37774 ( \38152 , \38149 , \38151 );
xor \U$37775 ( \38153 , \37923 , \37932 );
xor \U$37776 ( \38154 , \38153 , \37935 );
and \U$37777 ( \38155 , \38151 , \38154 );
and \U$37778 ( \38156 , \38149 , \38154 );
or \U$37779 ( \38157 , \38152 , \38155 , \38156 );
and \U$37780 ( \38158 , \37950 , \38157 );
xor \U$37781 ( \38159 , \37950 , \38157 );
xor \U$37782 ( \38160 , \38149 , \38151 );
xor \U$37783 ( \38161 , \38160 , \38154 );
and \U$37784 ( \38162 , \27494 , \25692 );
and \U$37785 ( \38163 , \27485 , \25690 );
nor \U$37786 ( \38164 , \38162 , \38163 );
xnor \U$37787 ( \38165 , \38164 , \25549 );
and \U$37788 ( \38166 , \28039 , \25369 );
and \U$37789 ( \38167 , \27837 , \25367 );
nor \U$37790 ( \38168 , \38166 , \38167 );
xnor \U$37791 ( \38169 , \38168 , \25123 );
and \U$37792 ( \38170 , \38165 , \38169 );
and \U$37793 ( \38171 , \28514 , \24974 );
and \U$37794 ( \38172 , \28342 , \24972 );
nor \U$37795 ( \38173 , \38171 , \38172 );
xnor \U$37796 ( \38174 , \38173 , \24787 );
and \U$37797 ( \38175 , \38169 , \38174 );
and \U$37798 ( \38176 , \38165 , \38174 );
or \U$37799 ( \38177 , \38170 , \38175 , \38176 );
and \U$37800 ( \38178 , \29464 , \24661 );
and \U$37801 ( \38179 , \29040 , \24659 );
nor \U$37802 ( \38180 , \38178 , \38179 );
xnor \U$37803 ( \38181 , \38180 , \24456 );
and \U$37804 ( \38182 , \29715 , \24255 );
and \U$37805 ( \38183 , \29710 , \24253 );
nor \U$37806 ( \38184 , \38182 , \38183 );
xnor \U$37807 ( \38185 , \38184 , \24106 );
and \U$37808 ( \38186 , \38181 , \38185 );
and \U$37809 ( \38187 , \30318 , \23933 );
and \U$37810 ( \38188 , \30034 , \23931 );
nor \U$37811 ( \38189 , \38187 , \38188 );
xnor \U$37812 ( \38190 , \38189 , \23791 );
and \U$37813 ( \38191 , \38185 , \38190 );
and \U$37814 ( \38192 , \38181 , \38190 );
or \U$37815 ( \38193 , \38186 , \38191 , \38192 );
and \U$37816 ( \38194 , \38177 , \38193 );
and \U$37817 ( \38195 , \26116 , \26983 );
and \U$37818 ( \38196 , \26108 , \26981 );
nor \U$37819 ( \38197 , \38195 , \38196 );
xnor \U$37820 ( \38198 , \38197 , \26742 );
and \U$37821 ( \38199 , \26590 , \26517 );
and \U$37822 ( \38200 , \26585 , \26515 );
nor \U$37823 ( \38201 , \38199 , \38200 );
xnor \U$37824 ( \38202 , \38201 , \26329 );
and \U$37825 ( \38203 , \38198 , \38202 );
and \U$37826 ( \38204 , \27113 , \26143 );
and \U$37827 ( \38205 , \26854 , \26141 );
nor \U$37828 ( \38206 , \38204 , \38205 );
xnor \U$37829 ( \38207 , \38206 , \25911 );
and \U$37830 ( \38208 , \38202 , \38207 );
and \U$37831 ( \38209 , \38198 , \38207 );
or \U$37832 ( \38210 , \38203 , \38208 , \38209 );
and \U$37833 ( \38211 , \38193 , \38210 );
and \U$37834 ( \38212 , \38177 , \38210 );
or \U$37835 ( \38213 , \38194 , \38211 , \38212 );
and \U$37836 ( \38214 , \25226 , \28575 );
and \U$37837 ( \38215 , \25018 , \28573 );
nor \U$37838 ( \38216 , \38214 , \38215 );
xnor \U$37839 ( \38217 , \38216 , \28315 );
and \U$37840 ( \38218 , \25353 , \28081 );
and \U$37841 ( \38219 , \25348 , \28079 );
nor \U$37842 ( \38220 , \38218 , \38219 );
xnor \U$37843 ( \38221 , \38220 , \27766 );
and \U$37844 ( \38222 , \38217 , \38221 );
and \U$37845 ( \38223 , \25806 , \27572 );
and \U$37846 ( \38224 , \25609 , \27570 );
nor \U$37847 ( \38225 , \38223 , \38224 );
xnor \U$37848 ( \38226 , \38225 , \27232 );
and \U$37849 ( \38227 , \38221 , \38226 );
and \U$37850 ( \38228 , \38217 , \38226 );
or \U$37851 ( \38229 , \38222 , \38227 , \38228 );
and \U$37852 ( \38230 , \24003 , \30233 );
and \U$37853 ( \38231 , \23978 , \30231 );
nor \U$37854 ( \38232 , \38230 , \38231 );
xnor \U$37855 ( \38233 , \38232 , \29862 );
and \U$37856 ( \38234 , \24344 , \29671 );
and \U$37857 ( \38235 , \24177 , \29669 );
nor \U$37858 ( \38236 , \38234 , \38235 );
xnor \U$37859 ( \38237 , \38236 , \29353 );
and \U$37860 ( \38238 , \38233 , \38237 );
and \U$37861 ( \38239 , \24601 , \29104 );
and \U$37862 ( \38240 , \24482 , \29102 );
nor \U$37863 ( \38241 , \38239 , \38240 );
xnor \U$37864 ( \38242 , \38241 , \28855 );
and \U$37865 ( \38243 , \38237 , \38242 );
and \U$37866 ( \38244 , \38233 , \38242 );
or \U$37867 ( \38245 , \38238 , \38243 , \38244 );
and \U$37868 ( \38246 , \38229 , \38245 );
and \U$37869 ( \38247 , \23136 , \32151 );
and \U$37870 ( \38248 , \23128 , \32148 );
nor \U$37871 ( \38249 , \38247 , \38248 );
xnor \U$37872 ( \38250 , \38249 , \31096 );
and \U$37873 ( \38251 , \23384 , \31338 );
and \U$37874 ( \38252 , \23379 , \31336 );
nor \U$37875 ( \38253 , \38251 , \38252 );
xnor \U$37876 ( \38254 , \38253 , \31099 );
and \U$37877 ( \38255 , \38250 , \38254 );
and \U$37878 ( \38256 , \23714 , \30770 );
and \U$37879 ( \38257 , \23570 , \30768 );
nor \U$37880 ( \38258 , \38256 , \38257 );
xnor \U$37881 ( \38259 , \38258 , \30460 );
and \U$37882 ( \38260 , \38254 , \38259 );
and \U$37883 ( \38261 , \38250 , \38259 );
or \U$37884 ( \38262 , \38255 , \38260 , \38261 );
and \U$37885 ( \38263 , \38245 , \38262 );
and \U$37886 ( \38264 , \38229 , \38262 );
or \U$37887 ( \38265 , \38246 , \38263 , \38264 );
and \U$37888 ( \38266 , \38213 , \38265 );
and \U$37889 ( \38267 , \30895 , \23637 );
and \U$37890 ( \38268 , \30887 , \23635 );
nor \U$37891 ( \38269 , \38267 , \38268 );
xnor \U$37892 ( \38270 , \38269 , \23500 );
and \U$37893 ( \38271 , \31503 , \23431 );
and \U$37894 ( \38272 , \31498 , \23429 );
nor \U$37895 ( \38273 , \38271 , \38272 );
xnor \U$37896 ( \38274 , \38273 , \23279 );
and \U$37897 ( \38275 , \38270 , \38274 );
and \U$37898 ( \38276 , \32304 , \23163 );
and \U$37899 ( \38277 , \31684 , \23161 );
nor \U$37900 ( \38278 , \38276 , \38277 );
xnor \U$37901 ( \38279 , \38278 , \23007 );
and \U$37902 ( \38280 , \38274 , \38279 );
and \U$37903 ( \38281 , \38270 , \38279 );
or \U$37904 ( \38282 , \38275 , \38280 , \38281 );
xor \U$37905 ( \38283 , \38055 , \38059 );
xor \U$37906 ( \38284 , \38283 , \38064 );
and \U$37907 ( \38285 , \38282 , \38284 );
xor \U$37908 ( \38286 , \38071 , \38073 );
and \U$37909 ( \38287 , \38284 , \38286 );
and \U$37910 ( \38288 , \38282 , \38286 );
or \U$37911 ( \38289 , \38285 , \38287 , \38288 );
and \U$37912 ( \38290 , \38265 , \38289 );
and \U$37913 ( \38291 , \38213 , \38289 );
or \U$37914 ( \38292 , \38266 , \38290 , \38291 );
xor \U$37915 ( \38293 , \38006 , \38010 );
xor \U$37916 ( \38294 , \38293 , \22778 );
xor \U$37917 ( \38295 , \38018 , \38022 );
xor \U$37918 ( \38296 , \38295 , \38027 );
and \U$37919 ( \38297 , \38294 , \38296 );
xor \U$37920 ( \38298 , \38035 , \38039 );
xor \U$37921 ( \38299 , \38298 , \38044 );
and \U$37922 ( \38300 , \38296 , \38299 );
and \U$37923 ( \38301 , \38294 , \38299 );
or \U$37924 ( \38302 , \38297 , \38300 , \38301 );
xor \U$37925 ( \38303 , \37954 , \37958 );
xor \U$37926 ( \38304 , \38303 , \37963 );
xor \U$37927 ( \38305 , \37970 , \37974 );
xor \U$37928 ( \38306 , \38305 , \37979 );
and \U$37929 ( \38307 , \38304 , \38306 );
xor \U$37930 ( \38308 , \37987 , \37991 );
xor \U$37931 ( \38309 , \38308 , \37996 );
and \U$37932 ( \38310 , \38306 , \38309 );
and \U$37933 ( \38311 , \38304 , \38309 );
or \U$37934 ( \38312 , \38307 , \38310 , \38311 );
and \U$37935 ( \38313 , \38302 , \38312 );
xor \U$37936 ( \38314 , \37723 , \37727 );
xor \U$37937 ( \38315 , \38314 , \37732 );
and \U$37938 ( \38316 , \38312 , \38315 );
and \U$37939 ( \38317 , \38302 , \38315 );
or \U$37940 ( \38318 , \38313 , \38316 , \38317 );
and \U$37941 ( \38319 , \38292 , \38318 );
xor \U$37942 ( \38320 , \38067 , \38074 );
xor \U$37943 ( \38321 , \38320 , \38079 );
xor \U$37944 ( \38322 , \38087 , \38089 );
xor \U$37945 ( \38323 , \38322 , \38092 );
and \U$37946 ( \38324 , \38321 , \38323 );
xor \U$37947 ( \38325 , \38097 , \38099 );
xor \U$37948 ( \38326 , \38325 , \38102 );
and \U$37949 ( \38327 , \38323 , \38326 );
and \U$37950 ( \38328 , \38321 , \38326 );
or \U$37951 ( \38329 , \38324 , \38327 , \38328 );
and \U$37952 ( \38330 , \38318 , \38329 );
and \U$37953 ( \38331 , \38292 , \38329 );
or \U$37954 ( \38332 , \38319 , \38330 , \38331 );
xor \U$37955 ( \38333 , \37735 , \37751 );
xor \U$37956 ( \38334 , \38333 , \37768 );
xor \U$37957 ( \38335 , \38095 , \38105 );
xor \U$37958 ( \38336 , \38335 , \38108 );
and \U$37959 ( \38337 , \38334 , \38336 );
xor \U$37960 ( \38338 , \38114 , \38116 );
xor \U$37961 ( \38339 , \38338 , \38119 );
and \U$37962 ( \38340 , \38336 , \38339 );
and \U$37963 ( \38341 , \38334 , \38339 );
or \U$37964 ( \38342 , \38337 , \38340 , \38341 );
and \U$37965 ( \38343 , \38332 , \38342 );
xor \U$37966 ( \38344 , \37771 , \37823 );
xor \U$37967 ( \38345 , \38344 , \37848 );
and \U$37968 ( \38346 , \38342 , \38345 );
and \U$37969 ( \38347 , \38332 , \38345 );
or \U$37970 ( \38348 , \38343 , \38346 , \38347 );
xor \U$37971 ( \38349 , \38085 , \38111 );
xor \U$37972 ( \38350 , \38349 , \38122 );
xor \U$37973 ( \38351 , \38127 , \38129 );
xor \U$37974 ( \38352 , \38351 , \38132 );
and \U$37975 ( \38353 , \38350 , \38352 );
and \U$37976 ( \38354 , \38348 , \38353 );
xor \U$37977 ( \38355 , \37901 , \37903 );
xor \U$37978 ( \38356 , \38355 , \37906 );
and \U$37979 ( \38357 , \38353 , \38356 );
and \U$37980 ( \38358 , \38348 , \38356 );
or \U$37981 ( \38359 , \38354 , \38357 , \38358 );
xor \U$37982 ( \38360 , \37851 , \37877 );
xor \U$37983 ( \38361 , \38360 , \37888 );
xor \U$37984 ( \38362 , \38125 , \38135 );
xor \U$37985 ( \38363 , \38362 , \38138 );
and \U$37986 ( \38364 , \38361 , \38363 );
and \U$37987 ( \38365 , \38359 , \38364 );
xor \U$37988 ( \38366 , \38141 , \38143 );
xor \U$37989 ( \38367 , \38366 , \38146 );
and \U$37990 ( \38368 , \38364 , \38367 );
and \U$37991 ( \38369 , \38359 , \38367 );
or \U$37992 ( \38370 , \38365 , \38368 , \38369 );
and \U$37993 ( \38371 , \38161 , \38370 );
xor \U$37994 ( \38372 , \38161 , \38370 );
xor \U$37995 ( \38373 , \38359 , \38364 );
xor \U$37996 ( \38374 , \38373 , \38367 );
and \U$37997 ( \38375 , \25018 , \29104 );
and \U$37998 ( \38376 , \24601 , \29102 );
nor \U$37999 ( \38377 , \38375 , \38376 );
xnor \U$38000 ( \38378 , \38377 , \28855 );
and \U$38001 ( \38379 , \25348 , \28575 );
and \U$38002 ( \38380 , \25226 , \28573 );
nor \U$38003 ( \38381 , \38379 , \38380 );
xnor \U$38004 ( \38382 , \38381 , \28315 );
and \U$38005 ( \38383 , \38378 , \38382 );
and \U$38006 ( \38384 , \25609 , \28081 );
and \U$38007 ( \38385 , \25353 , \28079 );
nor \U$38008 ( \38386 , \38384 , \38385 );
xnor \U$38009 ( \38387 , \38386 , \27766 );
and \U$38010 ( \38388 , \38382 , \38387 );
and \U$38011 ( \38389 , \38378 , \38387 );
or \U$38012 ( \38390 , \38383 , \38388 , \38389 );
and \U$38013 ( \38391 , \23978 , \30770 );
and \U$38014 ( \38392 , \23714 , \30768 );
nor \U$38015 ( \38393 , \38391 , \38392 );
xnor \U$38016 ( \38394 , \38393 , \30460 );
and \U$38017 ( \38395 , \24177 , \30233 );
and \U$38018 ( \38396 , \24003 , \30231 );
nor \U$38019 ( \38397 , \38395 , \38396 );
xnor \U$38020 ( \38398 , \38397 , \29862 );
and \U$38021 ( \38399 , \38394 , \38398 );
and \U$38022 ( \38400 , \24482 , \29671 );
and \U$38023 ( \38401 , \24344 , \29669 );
nor \U$38024 ( \38402 , \38400 , \38401 );
xnor \U$38025 ( \38403 , \38402 , \29353 );
and \U$38026 ( \38404 , \38398 , \38403 );
and \U$38027 ( \38405 , \38394 , \38403 );
or \U$38028 ( \38406 , \38399 , \38404 , \38405 );
and \U$38029 ( \38407 , \38390 , \38406 );
and \U$38030 ( \38408 , \23379 , \32151 );
and \U$38031 ( \38409 , \23136 , \32148 );
nor \U$38032 ( \38410 , \38408 , \38409 );
xnor \U$38033 ( \38411 , \38410 , \31096 );
and \U$38034 ( \38412 , \23570 , \31338 );
and \U$38035 ( \38413 , \23384 , \31336 );
nor \U$38036 ( \38414 , \38412 , \38413 );
xnor \U$38037 ( \38415 , \38414 , \31099 );
and \U$38038 ( \38416 , \38411 , \38415 );
and \U$38039 ( \38417 , \38415 , \23007 );
and \U$38040 ( \38418 , \38411 , \23007 );
or \U$38041 ( \38419 , \38416 , \38417 , \38418 );
and \U$38042 ( \38420 , \38406 , \38419 );
and \U$38043 ( \38421 , \38390 , \38419 );
or \U$38044 ( \38422 , \38407 , \38420 , \38421 );
and \U$38045 ( \38423 , \29040 , \24974 );
and \U$38046 ( \38424 , \28514 , \24972 );
nor \U$38047 ( \38425 , \38423 , \38424 );
xnor \U$38048 ( \38426 , \38425 , \24787 );
and \U$38049 ( \38427 , \29710 , \24661 );
and \U$38050 ( \38428 , \29464 , \24659 );
nor \U$38051 ( \38429 , \38427 , \38428 );
xnor \U$38052 ( \38430 , \38429 , \24456 );
and \U$38053 ( \38431 , \38426 , \38430 );
and \U$38054 ( \38432 , \30034 , \24255 );
and \U$38055 ( \38433 , \29715 , \24253 );
nor \U$38056 ( \38434 , \38432 , \38433 );
xnor \U$38057 ( \38435 , \38434 , \24106 );
and \U$38058 ( \38436 , \38430 , \38435 );
and \U$38059 ( \38437 , \38426 , \38435 );
or \U$38060 ( \38438 , \38431 , \38436 , \38437 );
and \U$38061 ( \38439 , \26108 , \27572 );
and \U$38062 ( \38440 , \25806 , \27570 );
nor \U$38063 ( \38441 , \38439 , \38440 );
xnor \U$38064 ( \38442 , \38441 , \27232 );
and \U$38065 ( \38443 , \26585 , \26983 );
and \U$38066 ( \38444 , \26116 , \26981 );
nor \U$38067 ( \38445 , \38443 , \38444 );
xnor \U$38068 ( \38446 , \38445 , \26742 );
and \U$38069 ( \38447 , \38442 , \38446 );
and \U$38070 ( \38448 , \26854 , \26517 );
and \U$38071 ( \38449 , \26590 , \26515 );
nor \U$38072 ( \38450 , \38448 , \38449 );
xnor \U$38073 ( \38451 , \38450 , \26329 );
and \U$38074 ( \38452 , \38446 , \38451 );
and \U$38075 ( \38453 , \38442 , \38451 );
or \U$38076 ( \38454 , \38447 , \38452 , \38453 );
and \U$38077 ( \38455 , \38438 , \38454 );
and \U$38078 ( \38456 , \27485 , \26143 );
and \U$38079 ( \38457 , \27113 , \26141 );
nor \U$38080 ( \38458 , \38456 , \38457 );
xnor \U$38081 ( \38459 , \38458 , \25911 );
and \U$38082 ( \38460 , \27837 , \25692 );
and \U$38083 ( \38461 , \27494 , \25690 );
nor \U$38084 ( \38462 , \38460 , \38461 );
xnor \U$38085 ( \38463 , \38462 , \25549 );
and \U$38086 ( \38464 , \38459 , \38463 );
and \U$38087 ( \38465 , \28342 , \25369 );
and \U$38088 ( \38466 , \28039 , \25367 );
nor \U$38089 ( \38467 , \38465 , \38466 );
xnor \U$38090 ( \38468 , \38467 , \25123 );
and \U$38091 ( \38469 , \38463 , \38468 );
and \U$38092 ( \38470 , \38459 , \38468 );
or \U$38093 ( \38471 , \38464 , \38469 , \38470 );
and \U$38094 ( \38472 , \38454 , \38471 );
and \U$38095 ( \38473 , \38438 , \38471 );
or \U$38096 ( \38474 , \38455 , \38472 , \38473 );
and \U$38097 ( \38475 , \38422 , \38474 );
and \U$38098 ( \38476 , \30887 , \23933 );
and \U$38099 ( \38477 , \30318 , \23931 );
nor \U$38100 ( \38478 , \38476 , \38477 );
xnor \U$38101 ( \38479 , \38478 , \23791 );
and \U$38102 ( \38480 , \31498 , \23637 );
and \U$38103 ( \38481 , \30895 , \23635 );
nor \U$38104 ( \38482 , \38480 , \38481 );
xnor \U$38105 ( \38483 , \38482 , \23500 );
and \U$38106 ( \38484 , \38479 , \38483 );
and \U$38107 ( \38485 , \31684 , \23431 );
and \U$38108 ( \38486 , \31503 , \23429 );
nor \U$38109 ( \38487 , \38485 , \38486 );
xnor \U$38110 ( \38488 , \38487 , \23279 );
and \U$38111 ( \38489 , \38483 , \38488 );
and \U$38112 ( \38490 , \38479 , \38488 );
or \U$38113 ( \38491 , \38484 , \38489 , \38490 );
xor \U$38114 ( \38492 , \38181 , \38185 );
xor \U$38115 ( \38493 , \38492 , \38190 );
and \U$38116 ( \38494 , \38491 , \38493 );
xor \U$38117 ( \38495 , \38270 , \38274 );
xor \U$38118 ( \38496 , \38495 , \38279 );
and \U$38119 ( \38497 , \38493 , \38496 );
and \U$38120 ( \38498 , \38491 , \38496 );
or \U$38121 ( \38499 , \38494 , \38497 , \38498 );
and \U$38122 ( \38500 , \38474 , \38499 );
and \U$38123 ( \38501 , \38422 , \38499 );
or \U$38124 ( \38502 , \38475 , \38500 , \38501 );
xor \U$38125 ( \38503 , \38165 , \38169 );
xor \U$38126 ( \38504 , \38503 , \38174 );
xor \U$38127 ( \38505 , \38217 , \38221 );
xor \U$38128 ( \38506 , \38505 , \38226 );
and \U$38129 ( \38507 , \38504 , \38506 );
xor \U$38130 ( \38508 , \38198 , \38202 );
xor \U$38131 ( \38509 , \38508 , \38207 );
and \U$38132 ( \38510 , \38506 , \38509 );
and \U$38133 ( \38511 , \38504 , \38509 );
or \U$38134 ( \38512 , \38507 , \38510 , \38511 );
xor \U$38135 ( \38513 , \38233 , \38237 );
xor \U$38136 ( \38514 , \38513 , \38242 );
xor \U$38137 ( \38515 , \38250 , \38254 );
xor \U$38138 ( \38516 , \38515 , \38259 );
and \U$38139 ( \38517 , \38514 , \38516 );
and \U$38140 ( \38518 , \38512 , \38517 );
xor \U$38141 ( \38519 , \38294 , \38296 );
xor \U$38142 ( \38520 , \38519 , \38299 );
and \U$38143 ( \38521 , \38517 , \38520 );
and \U$38144 ( \38522 , \38512 , \38520 );
or \U$38145 ( \38523 , \38518 , \38521 , \38522 );
and \U$38146 ( \38524 , \38502 , \38523 );
xor \U$38147 ( \38525 , \38177 , \38193 );
xor \U$38148 ( \38526 , \38525 , \38210 );
xor \U$38149 ( \38527 , \38304 , \38306 );
xor \U$38150 ( \38528 , \38527 , \38309 );
and \U$38151 ( \38529 , \38526 , \38528 );
xor \U$38152 ( \38530 , \38282 , \38284 );
xor \U$38153 ( \38531 , \38530 , \38286 );
and \U$38154 ( \38532 , \38528 , \38531 );
and \U$38155 ( \38533 , \38526 , \38531 );
or \U$38156 ( \38534 , \38529 , \38532 , \38533 );
and \U$38157 ( \38535 , \38523 , \38534 );
and \U$38158 ( \38536 , \38502 , \38534 );
or \U$38159 ( \38537 , \38524 , \38535 , \38536 );
xor \U$38160 ( \38538 , \37966 , \37982 );
xor \U$38161 ( \38539 , \38538 , \37999 );
xor \U$38162 ( \38540 , \38014 , \38030 );
xor \U$38163 ( \38541 , \38540 , \38047 );
and \U$38164 ( \38542 , \38539 , \38541 );
xor \U$38165 ( \38543 , \38321 , \38323 );
xor \U$38166 ( \38544 , \38543 , \38326 );
and \U$38167 ( \38545 , \38541 , \38544 );
and \U$38168 ( \38546 , \38539 , \38544 );
or \U$38169 ( \38547 , \38542 , \38545 , \38546 );
and \U$38170 ( \38548 , \38537 , \38547 );
xor \U$38171 ( \38549 , \38002 , \38050 );
xor \U$38172 ( \38550 , \38549 , \38082 );
and \U$38173 ( \38551 , \38547 , \38550 );
and \U$38174 ( \38552 , \38537 , \38550 );
or \U$38175 ( \38553 , \38548 , \38551 , \38552 );
xor \U$38176 ( \38554 , \38332 , \38342 );
xor \U$38177 ( \38555 , \38554 , \38345 );
and \U$38178 ( \38556 , \38553 , \38555 );
xor \U$38179 ( \38557 , \38350 , \38352 );
and \U$38180 ( \38558 , \38555 , \38557 );
and \U$38181 ( \38559 , \38553 , \38557 );
or \U$38182 ( \38560 , \38556 , \38558 , \38559 );
xor \U$38183 ( \38561 , \38348 , \38353 );
xor \U$38184 ( \38562 , \38561 , \38356 );
and \U$38185 ( \38563 , \38560 , \38562 );
xor \U$38186 ( \38564 , \38361 , \38363 );
and \U$38187 ( \38565 , \38562 , \38564 );
and \U$38188 ( \38566 , \38560 , \38564 );
or \U$38189 ( \38567 , \38563 , \38565 , \38566 );
and \U$38190 ( \38568 , \38374 , \38567 );
xor \U$38191 ( \38569 , \38374 , \38567 );
xor \U$38192 ( \38570 , \38560 , \38562 );
xor \U$38193 ( \38571 , \38570 , \38564 );
and \U$38194 ( \38572 , \23384 , \32151 );
and \U$38195 ( \38573 , \23379 , \32148 );
nor \U$38196 ( \38574 , \38572 , \38573 );
xnor \U$38197 ( \38575 , \38574 , \31096 );
and \U$38198 ( \38576 , \23714 , \31338 );
and \U$38199 ( \38577 , \23570 , \31336 );
nor \U$38200 ( \38578 , \38576 , \38577 );
xnor \U$38201 ( \38579 , \38578 , \31099 );
and \U$38202 ( \38580 , \38575 , \38579 );
and \U$38203 ( \38581 , \24003 , \30770 );
and \U$38204 ( \38582 , \23978 , \30768 );
nor \U$38205 ( \38583 , \38581 , \38582 );
xnor \U$38206 ( \38584 , \38583 , \30460 );
and \U$38207 ( \38585 , \38579 , \38584 );
and \U$38208 ( \38586 , \38575 , \38584 );
or \U$38209 ( \38587 , \38580 , \38585 , \38586 );
and \U$38210 ( \38588 , \24344 , \30233 );
and \U$38211 ( \38589 , \24177 , \30231 );
nor \U$38212 ( \38590 , \38588 , \38589 );
xnor \U$38213 ( \38591 , \38590 , \29862 );
and \U$38214 ( \38592 , \24601 , \29671 );
and \U$38215 ( \38593 , \24482 , \29669 );
nor \U$38216 ( \38594 , \38592 , \38593 );
xnor \U$38217 ( \38595 , \38594 , \29353 );
and \U$38218 ( \38596 , \38591 , \38595 );
and \U$38219 ( \38597 , \25226 , \29104 );
and \U$38220 ( \38598 , \25018 , \29102 );
nor \U$38221 ( \38599 , \38597 , \38598 );
xnor \U$38222 ( \38600 , \38599 , \28855 );
and \U$38223 ( \38601 , \38595 , \38600 );
and \U$38224 ( \38602 , \38591 , \38600 );
or \U$38225 ( \38603 , \38596 , \38601 , \38602 );
and \U$38226 ( \38604 , \38587 , \38603 );
and \U$38227 ( \38605 , \25353 , \28575 );
and \U$38228 ( \38606 , \25348 , \28573 );
nor \U$38229 ( \38607 , \38605 , \38606 );
xnor \U$38230 ( \38608 , \38607 , \28315 );
and \U$38231 ( \38609 , \25806 , \28081 );
and \U$38232 ( \38610 , \25609 , \28079 );
nor \U$38233 ( \38611 , \38609 , \38610 );
xnor \U$38234 ( \38612 , \38611 , \27766 );
and \U$38235 ( \38613 , \38608 , \38612 );
and \U$38236 ( \38614 , \26116 , \27572 );
and \U$38237 ( \38615 , \26108 , \27570 );
nor \U$38238 ( \38616 , \38614 , \38615 );
xnor \U$38239 ( \38617 , \38616 , \27232 );
and \U$38240 ( \38618 , \38612 , \38617 );
and \U$38241 ( \38619 , \38608 , \38617 );
or \U$38242 ( \38620 , \38613 , \38618 , \38619 );
and \U$38243 ( \38621 , \38603 , \38620 );
and \U$38244 ( \38622 , \38587 , \38620 );
or \U$38245 ( \38623 , \38604 , \38621 , \38622 );
and \U$38246 ( \38624 , \28039 , \25692 );
and \U$38247 ( \38625 , \27837 , \25690 );
nor \U$38248 ( \38626 , \38624 , \38625 );
xnor \U$38249 ( \38627 , \38626 , \25549 );
and \U$38250 ( \38628 , \28514 , \25369 );
and \U$38251 ( \38629 , \28342 , \25367 );
nor \U$38252 ( \38630 , \38628 , \38629 );
xnor \U$38253 ( \38631 , \38630 , \25123 );
and \U$38254 ( \38632 , \38627 , \38631 );
and \U$38255 ( \38633 , \29464 , \24974 );
and \U$38256 ( \38634 , \29040 , \24972 );
nor \U$38257 ( \38635 , \38633 , \38634 );
xnor \U$38258 ( \38636 , \38635 , \24787 );
and \U$38259 ( \38637 , \38631 , \38636 );
and \U$38260 ( \38638 , \38627 , \38636 );
or \U$38261 ( \38639 , \38632 , \38637 , \38638 );
and \U$38262 ( \38640 , \26590 , \26983 );
and \U$38263 ( \38641 , \26585 , \26981 );
nor \U$38264 ( \38642 , \38640 , \38641 );
xnor \U$38265 ( \38643 , \38642 , \26742 );
and \U$38266 ( \38644 , \27113 , \26517 );
and \U$38267 ( \38645 , \26854 , \26515 );
nor \U$38268 ( \38646 , \38644 , \38645 );
xnor \U$38269 ( \38647 , \38646 , \26329 );
and \U$38270 ( \38648 , \38643 , \38647 );
and \U$38271 ( \38649 , \27494 , \26143 );
and \U$38272 ( \38650 , \27485 , \26141 );
nor \U$38273 ( \38651 , \38649 , \38650 );
xnor \U$38274 ( \38652 , \38651 , \25911 );
and \U$38275 ( \38653 , \38647 , \38652 );
and \U$38276 ( \38654 , \38643 , \38652 );
or \U$38277 ( \38655 , \38648 , \38653 , \38654 );
and \U$38278 ( \38656 , \38639 , \38655 );
and \U$38279 ( \38657 , \29715 , \24661 );
and \U$38280 ( \38658 , \29710 , \24659 );
nor \U$38281 ( \38659 , \38657 , \38658 );
xnor \U$38282 ( \38660 , \38659 , \24456 );
and \U$38283 ( \38661 , \30318 , \24255 );
and \U$38284 ( \38662 , \30034 , \24253 );
nor \U$38285 ( \38663 , \38661 , \38662 );
xnor \U$38286 ( \38664 , \38663 , \24106 );
and \U$38287 ( \38665 , \38660 , \38664 );
and \U$38288 ( \38666 , \30895 , \23933 );
and \U$38289 ( \38667 , \30887 , \23931 );
nor \U$38290 ( \38668 , \38666 , \38667 );
xnor \U$38291 ( \38669 , \38668 , \23791 );
and \U$38292 ( \38670 , \38664 , \38669 );
and \U$38293 ( \38671 , \38660 , \38669 );
or \U$38294 ( \38672 , \38665 , \38670 , \38671 );
and \U$38295 ( \38673 , \38655 , \38672 );
and \U$38296 ( \38674 , \38639 , \38672 );
or \U$38297 ( \38675 , \38656 , \38673 , \38674 );
and \U$38298 ( \38676 , \38623 , \38675 );
nand \U$38299 ( \38677 , \32304 , \23161 );
xnor \U$38300 ( \38678 , \38677 , \23007 );
xor \U$38301 ( \38679 , \38426 , \38430 );
xor \U$38302 ( \38680 , \38679 , \38435 );
and \U$38303 ( \38681 , \38678 , \38680 );
xor \U$38304 ( \38682 , \38479 , \38483 );
xor \U$38305 ( \38683 , \38682 , \38488 );
and \U$38306 ( \38684 , \38680 , \38683 );
and \U$38307 ( \38685 , \38678 , \38683 );
or \U$38308 ( \38686 , \38681 , \38684 , \38685 );
and \U$38309 ( \38687 , \38675 , \38686 );
and \U$38310 ( \38688 , \38623 , \38686 );
or \U$38311 ( \38689 , \38676 , \38687 , \38688 );
xor \U$38312 ( \38690 , \38390 , \38406 );
xor \U$38313 ( \38691 , \38690 , \38419 );
xor \U$38314 ( \38692 , \38438 , \38454 );
xor \U$38315 ( \38693 , \38692 , \38471 );
and \U$38316 ( \38694 , \38691 , \38693 );
xor \U$38317 ( \38695 , \38491 , \38493 );
xor \U$38318 ( \38696 , \38695 , \38496 );
and \U$38319 ( \38697 , \38693 , \38696 );
and \U$38320 ( \38698 , \38691 , \38696 );
or \U$38321 ( \38699 , \38694 , \38697 , \38698 );
and \U$38322 ( \38700 , \38689 , \38699 );
xor \U$38323 ( \38701 , \38378 , \38382 );
xor \U$38324 ( \38702 , \38701 , \38387 );
xor \U$38325 ( \38703 , \38442 , \38446 );
xor \U$38326 ( \38704 , \38703 , \38451 );
and \U$38327 ( \38705 , \38702 , \38704 );
xor \U$38328 ( \38706 , \38459 , \38463 );
xor \U$38329 ( \38707 , \38706 , \38468 );
and \U$38330 ( \38708 , \38704 , \38707 );
and \U$38331 ( \38709 , \38702 , \38707 );
or \U$38332 ( \38710 , \38705 , \38708 , \38709 );
xor \U$38333 ( \38711 , \38504 , \38506 );
xor \U$38334 ( \38712 , \38711 , \38509 );
and \U$38335 ( \38713 , \38710 , \38712 );
xor \U$38336 ( \38714 , \38514 , \38516 );
and \U$38337 ( \38715 , \38712 , \38714 );
and \U$38338 ( \38716 , \38710 , \38714 );
or \U$38339 ( \38717 , \38713 , \38715 , \38716 );
and \U$38340 ( \38718 , \38699 , \38717 );
and \U$38341 ( \38719 , \38689 , \38717 );
or \U$38342 ( \38720 , \38700 , \38718 , \38719 );
xor \U$38343 ( \38721 , \38229 , \38245 );
xor \U$38344 ( \38722 , \38721 , \38262 );
xor \U$38345 ( \38723 , \38512 , \38517 );
xor \U$38346 ( \38724 , \38723 , \38520 );
and \U$38347 ( \38725 , \38722 , \38724 );
xor \U$38348 ( \38726 , \38526 , \38528 );
xor \U$38349 ( \38727 , \38726 , \38531 );
and \U$38350 ( \38728 , \38724 , \38727 );
and \U$38351 ( \38729 , \38722 , \38727 );
or \U$38352 ( \38730 , \38725 , \38728 , \38729 );
and \U$38353 ( \38731 , \38720 , \38730 );
xor \U$38354 ( \38732 , \38302 , \38312 );
xor \U$38355 ( \38733 , \38732 , \38315 );
and \U$38356 ( \38734 , \38730 , \38733 );
and \U$38357 ( \38735 , \38720 , \38733 );
or \U$38358 ( \38736 , \38731 , \38734 , \38735 );
xor \U$38359 ( \38737 , \38213 , \38265 );
xor \U$38360 ( \38738 , \38737 , \38289 );
xor \U$38361 ( \38739 , \38502 , \38523 );
xor \U$38362 ( \38740 , \38739 , \38534 );
and \U$38363 ( \38741 , \38738 , \38740 );
xor \U$38364 ( \38742 , \38539 , \38541 );
xor \U$38365 ( \38743 , \38742 , \38544 );
and \U$38366 ( \38744 , \38740 , \38743 );
and \U$38367 ( \38745 , \38738 , \38743 );
or \U$38368 ( \38746 , \38741 , \38744 , \38745 );
and \U$38369 ( \38747 , \38736 , \38746 );
xor \U$38370 ( \38748 , \38334 , \38336 );
xor \U$38371 ( \38749 , \38748 , \38339 );
and \U$38372 ( \38750 , \38746 , \38749 );
and \U$38373 ( \38751 , \38736 , \38749 );
or \U$38374 ( \38752 , \38747 , \38750 , \38751 );
xor \U$38375 ( \38753 , \38292 , \38318 );
xor \U$38376 ( \38754 , \38753 , \38329 );
xor \U$38377 ( \38755 , \38537 , \38547 );
xor \U$38378 ( \38756 , \38755 , \38550 );
and \U$38379 ( \38757 , \38754 , \38756 );
and \U$38380 ( \38758 , \38752 , \38757 );
xor \U$38381 ( \38759 , \38553 , \38555 );
xor \U$38382 ( \38760 , \38759 , \38557 );
and \U$38383 ( \38761 , \38757 , \38760 );
and \U$38384 ( \38762 , \38752 , \38760 );
or \U$38385 ( \38763 , \38758 , \38761 , \38762 );
and \U$38386 ( \38764 , \38571 , \38763 );
xor \U$38387 ( \38765 , \38571 , \38763 );
xor \U$38388 ( \38766 , \38752 , \38757 );
xor \U$38389 ( \38767 , \38766 , \38760 );
and \U$38390 ( \38768 , \23570 , \32151 );
and \U$38391 ( \38769 , \23384 , \32148 );
nor \U$38392 ( \38770 , \38768 , \38769 );
xnor \U$38393 ( \38771 , \38770 , \31096 );
and \U$38394 ( \38772 , \23978 , \31338 );
and \U$38395 ( \38773 , \23714 , \31336 );
nor \U$38396 ( \38774 , \38772 , \38773 );
xnor \U$38397 ( \38775 , \38774 , \31099 );
and \U$38398 ( \38776 , \38771 , \38775 );
and \U$38399 ( \38777 , \38775 , \23279 );
and \U$38400 ( \38778 , \38771 , \23279 );
or \U$38401 ( \38779 , \38776 , \38777 , \38778 );
and \U$38402 ( \38780 , \25348 , \29104 );
and \U$38403 ( \38781 , \25226 , \29102 );
nor \U$38404 ( \38782 , \38780 , \38781 );
xnor \U$38405 ( \38783 , \38782 , \28855 );
and \U$38406 ( \38784 , \25609 , \28575 );
and \U$38407 ( \38785 , \25353 , \28573 );
nor \U$38408 ( \38786 , \38784 , \38785 );
xnor \U$38409 ( \38787 , \38786 , \28315 );
and \U$38410 ( \38788 , \38783 , \38787 );
and \U$38411 ( \38789 , \26108 , \28081 );
and \U$38412 ( \38790 , \25806 , \28079 );
nor \U$38413 ( \38791 , \38789 , \38790 );
xnor \U$38414 ( \38792 , \38791 , \27766 );
and \U$38415 ( \38793 , \38787 , \38792 );
and \U$38416 ( \38794 , \38783 , \38792 );
or \U$38417 ( \38795 , \38788 , \38793 , \38794 );
and \U$38418 ( \38796 , \38779 , \38795 );
and \U$38419 ( \38797 , \24177 , \30770 );
and \U$38420 ( \38798 , \24003 , \30768 );
nor \U$38421 ( \38799 , \38797 , \38798 );
xnor \U$38422 ( \38800 , \38799 , \30460 );
and \U$38423 ( \38801 , \24482 , \30233 );
and \U$38424 ( \38802 , \24344 , \30231 );
nor \U$38425 ( \38803 , \38801 , \38802 );
xnor \U$38426 ( \38804 , \38803 , \29862 );
and \U$38427 ( \38805 , \38800 , \38804 );
and \U$38428 ( \38806 , \25018 , \29671 );
and \U$38429 ( \38807 , \24601 , \29669 );
nor \U$38430 ( \38808 , \38806 , \38807 );
xnor \U$38431 ( \38809 , \38808 , \29353 );
and \U$38432 ( \38810 , \38804 , \38809 );
and \U$38433 ( \38811 , \38800 , \38809 );
or \U$38434 ( \38812 , \38805 , \38810 , \38811 );
and \U$38435 ( \38813 , \38795 , \38812 );
and \U$38436 ( \38814 , \38779 , \38812 );
or \U$38437 ( \38815 , \38796 , \38813 , \38814 );
and \U$38438 ( \38816 , \31498 , \23933 );
and \U$38439 ( \38817 , \30895 , \23931 );
nor \U$38440 ( \38818 , \38816 , \38817 );
xnor \U$38441 ( \38819 , \38818 , \23791 );
and \U$38442 ( \38820 , \31684 , \23637 );
and \U$38443 ( \38821 , \31503 , \23635 );
nor \U$38444 ( \38822 , \38820 , \38821 );
xnor \U$38445 ( \38823 , \38822 , \23500 );
and \U$38446 ( \38824 , \38819 , \38823 );
nand \U$38447 ( \38825 , \32304 , \23429 );
xnor \U$38448 ( \38826 , \38825 , \23279 );
and \U$38449 ( \38827 , \38823 , \38826 );
and \U$38450 ( \38828 , \38819 , \38826 );
or \U$38451 ( \38829 , \38824 , \38827 , \38828 );
and \U$38452 ( \38830 , \31503 , \23637 );
and \U$38453 ( \38831 , \31498 , \23635 );
nor \U$38454 ( \38832 , \38830 , \38831 );
xnor \U$38455 ( \38833 , \38832 , \23500 );
and \U$38456 ( \38834 , \38829 , \38833 );
and \U$38457 ( \38835 , \32304 , \23431 );
and \U$38458 ( \38836 , \31684 , \23429 );
nor \U$38459 ( \38837 , \38835 , \38836 );
xnor \U$38460 ( \38838 , \38837 , \23279 );
and \U$38461 ( \38839 , \38833 , \38838 );
and \U$38462 ( \38840 , \38829 , \38838 );
or \U$38463 ( \38841 , \38834 , \38839 , \38840 );
and \U$38464 ( \38842 , \38815 , \38841 );
and \U$38465 ( \38843 , \26585 , \27572 );
and \U$38466 ( \38844 , \26116 , \27570 );
nor \U$38467 ( \38845 , \38843 , \38844 );
xnor \U$38468 ( \38846 , \38845 , \27232 );
and \U$38469 ( \38847 , \26854 , \26983 );
and \U$38470 ( \38848 , \26590 , \26981 );
nor \U$38471 ( \38849 , \38847 , \38848 );
xnor \U$38472 ( \38850 , \38849 , \26742 );
and \U$38473 ( \38851 , \38846 , \38850 );
and \U$38474 ( \38852 , \27485 , \26517 );
and \U$38475 ( \38853 , \27113 , \26515 );
nor \U$38476 ( \38854 , \38852 , \38853 );
xnor \U$38477 ( \38855 , \38854 , \26329 );
and \U$38478 ( \38856 , \38850 , \38855 );
and \U$38479 ( \38857 , \38846 , \38855 );
or \U$38480 ( \38858 , \38851 , \38856 , \38857 );
and \U$38481 ( \38859 , \29710 , \24974 );
and \U$38482 ( \38860 , \29464 , \24972 );
nor \U$38483 ( \38861 , \38859 , \38860 );
xnor \U$38484 ( \38862 , \38861 , \24787 );
and \U$38485 ( \38863 , \30034 , \24661 );
and \U$38486 ( \38864 , \29715 , \24659 );
nor \U$38487 ( \38865 , \38863 , \38864 );
xnor \U$38488 ( \38866 , \38865 , \24456 );
and \U$38489 ( \38867 , \38862 , \38866 );
and \U$38490 ( \38868 , \30887 , \24255 );
and \U$38491 ( \38869 , \30318 , \24253 );
nor \U$38492 ( \38870 , \38868 , \38869 );
xnor \U$38493 ( \38871 , \38870 , \24106 );
and \U$38494 ( \38872 , \38866 , \38871 );
and \U$38495 ( \38873 , \38862 , \38871 );
or \U$38496 ( \38874 , \38867 , \38872 , \38873 );
and \U$38497 ( \38875 , \38858 , \38874 );
and \U$38498 ( \38876 , \27837 , \26143 );
and \U$38499 ( \38877 , \27494 , \26141 );
nor \U$38500 ( \38878 , \38876 , \38877 );
xnor \U$38501 ( \38879 , \38878 , \25911 );
and \U$38502 ( \38880 , \28342 , \25692 );
and \U$38503 ( \38881 , \28039 , \25690 );
nor \U$38504 ( \38882 , \38880 , \38881 );
xnor \U$38505 ( \38883 , \38882 , \25549 );
and \U$38506 ( \38884 , \38879 , \38883 );
and \U$38507 ( \38885 , \29040 , \25369 );
and \U$38508 ( \38886 , \28514 , \25367 );
nor \U$38509 ( \38887 , \38885 , \38886 );
xnor \U$38510 ( \38888 , \38887 , \25123 );
and \U$38511 ( \38889 , \38883 , \38888 );
and \U$38512 ( \38890 , \38879 , \38888 );
or \U$38513 ( \38891 , \38884 , \38889 , \38890 );
and \U$38514 ( \38892 , \38874 , \38891 );
and \U$38515 ( \38893 , \38858 , \38891 );
or \U$38516 ( \38894 , \38875 , \38892 , \38893 );
and \U$38517 ( \38895 , \38841 , \38894 );
and \U$38518 ( \38896 , \38815 , \38894 );
or \U$38519 ( \38897 , \38842 , \38895 , \38896 );
xor \U$38520 ( \38898 , \38575 , \38579 );
xor \U$38521 ( \38899 , \38898 , \38584 );
xor \U$38522 ( \38900 , \38591 , \38595 );
xor \U$38523 ( \38901 , \38900 , \38600 );
and \U$38524 ( \38902 , \38899 , \38901 );
xor \U$38525 ( \38903 , \38608 , \38612 );
xor \U$38526 ( \38904 , \38903 , \38617 );
and \U$38527 ( \38905 , \38901 , \38904 );
and \U$38528 ( \38906 , \38899 , \38904 );
or \U$38529 ( \38907 , \38902 , \38905 , \38906 );
xor \U$38530 ( \38908 , \38627 , \38631 );
xor \U$38531 ( \38909 , \38908 , \38636 );
xor \U$38532 ( \38910 , \38643 , \38647 );
xor \U$38533 ( \38911 , \38910 , \38652 );
and \U$38534 ( \38912 , \38909 , \38911 );
xor \U$38535 ( \38913 , \38660 , \38664 );
xor \U$38536 ( \38914 , \38913 , \38669 );
and \U$38537 ( \38915 , \38911 , \38914 );
and \U$38538 ( \38916 , \38909 , \38914 );
or \U$38539 ( \38917 , \38912 , \38915 , \38916 );
and \U$38540 ( \38918 , \38907 , \38917 );
xor \U$38541 ( \38919 , \38394 , \38398 );
xor \U$38542 ( \38920 , \38919 , \38403 );
and \U$38543 ( \38921 , \38917 , \38920 );
and \U$38544 ( \38922 , \38907 , \38920 );
or \U$38545 ( \38923 , \38918 , \38921 , \38922 );
and \U$38546 ( \38924 , \38897 , \38923 );
xor \U$38547 ( \38925 , \38411 , \38415 );
xor \U$38548 ( \38926 , \38925 , \23007 );
xor \U$38549 ( \38927 , \38702 , \38704 );
xor \U$38550 ( \38928 , \38927 , \38707 );
and \U$38551 ( \38929 , \38926 , \38928 );
xor \U$38552 ( \38930 , \38678 , \38680 );
xor \U$38553 ( \38931 , \38930 , \38683 );
and \U$38554 ( \38932 , \38928 , \38931 );
and \U$38555 ( \38933 , \38926 , \38931 );
or \U$38556 ( \38934 , \38929 , \38932 , \38933 );
and \U$38557 ( \38935 , \38923 , \38934 );
and \U$38558 ( \38936 , \38897 , \38934 );
or \U$38559 ( \38937 , \38924 , \38935 , \38936 );
xor \U$38560 ( \38938 , \38623 , \38675 );
xor \U$38561 ( \38939 , \38938 , \38686 );
xor \U$38562 ( \38940 , \38691 , \38693 );
xor \U$38563 ( \38941 , \38940 , \38696 );
and \U$38564 ( \38942 , \38939 , \38941 );
xor \U$38565 ( \38943 , \38710 , \38712 );
xor \U$38566 ( \38944 , \38943 , \38714 );
and \U$38567 ( \38945 , \38941 , \38944 );
and \U$38568 ( \38946 , \38939 , \38944 );
or \U$38569 ( \38947 , \38942 , \38945 , \38946 );
and \U$38570 ( \38948 , \38937 , \38947 );
xor \U$38571 ( \38949 , \38422 , \38474 );
xor \U$38572 ( \38950 , \38949 , \38499 );
and \U$38573 ( \38951 , \38947 , \38950 );
and \U$38574 ( \38952 , \38937 , \38950 );
or \U$38575 ( \38953 , \38948 , \38951 , \38952 );
xor \U$38576 ( \38954 , \38689 , \38699 );
xor \U$38577 ( \38955 , \38954 , \38717 );
xor \U$38578 ( \38956 , \38722 , \38724 );
xor \U$38579 ( \38957 , \38956 , \38727 );
and \U$38580 ( \38958 , \38955 , \38957 );
and \U$38581 ( \38959 , \38953 , \38958 );
xor \U$38582 ( \38960 , \38738 , \38740 );
xor \U$38583 ( \38961 , \38960 , \38743 );
and \U$38584 ( \38962 , \38958 , \38961 );
and \U$38585 ( \38963 , \38953 , \38961 );
or \U$38586 ( \38964 , \38959 , \38962 , \38963 );
xor \U$38587 ( \38965 , \38736 , \38746 );
xor \U$38588 ( \38966 , \38965 , \38749 );
and \U$38589 ( \38967 , \38964 , \38966 );
xor \U$38590 ( \38968 , \38754 , \38756 );
and \U$38591 ( \38969 , \38966 , \38968 );
and \U$38592 ( \38970 , \38964 , \38968 );
or \U$38593 ( \38971 , \38967 , \38969 , \38970 );
and \U$38594 ( \38972 , \38767 , \38971 );
xor \U$38595 ( \38973 , \38767 , \38971 );
xor \U$38596 ( \38974 , \38964 , \38966 );
xor \U$38597 ( \38975 , \38974 , \38968 );
and \U$38598 ( \38976 , \30318 , \24661 );
and \U$38599 ( \38977 , \30034 , \24659 );
nor \U$38600 ( \38978 , \38976 , \38977 );
xnor \U$38601 ( \38979 , \38978 , \24456 );
and \U$38602 ( \38980 , \30895 , \24255 );
and \U$38603 ( \38981 , \30887 , \24253 );
nor \U$38604 ( \38982 , \38980 , \38981 );
xnor \U$38605 ( \38983 , \38982 , \24106 );
and \U$38606 ( \38984 , \38979 , \38983 );
and \U$38607 ( \38985 , \31503 , \23933 );
and \U$38608 ( \38986 , \31498 , \23931 );
nor \U$38609 ( \38987 , \38985 , \38986 );
xnor \U$38610 ( \38988 , \38987 , \23791 );
and \U$38611 ( \38989 , \38983 , \38988 );
and \U$38612 ( \38990 , \38979 , \38988 );
or \U$38613 ( \38991 , \38984 , \38989 , \38990 );
and \U$38614 ( \38992 , \27113 , \26983 );
and \U$38615 ( \38993 , \26854 , \26981 );
nor \U$38616 ( \38994 , \38992 , \38993 );
xnor \U$38617 ( \38995 , \38994 , \26742 );
and \U$38618 ( \38996 , \27494 , \26517 );
and \U$38619 ( \38997 , \27485 , \26515 );
nor \U$38620 ( \38998 , \38996 , \38997 );
xnor \U$38621 ( \38999 , \38998 , \26329 );
and \U$38622 ( \39000 , \38995 , \38999 );
and \U$38623 ( \39001 , \28039 , \26143 );
and \U$38624 ( \39002 , \27837 , \26141 );
nor \U$38625 ( \39003 , \39001 , \39002 );
xnor \U$38626 ( \39004 , \39003 , \25911 );
and \U$38627 ( \39005 , \38999 , \39004 );
and \U$38628 ( \39006 , \38995 , \39004 );
or \U$38629 ( \39007 , \39000 , \39005 , \39006 );
and \U$38630 ( \39008 , \38991 , \39007 );
and \U$38631 ( \39009 , \28514 , \25692 );
and \U$38632 ( \39010 , \28342 , \25690 );
nor \U$38633 ( \39011 , \39009 , \39010 );
xnor \U$38634 ( \39012 , \39011 , \25549 );
and \U$38635 ( \39013 , \29464 , \25369 );
and \U$38636 ( \39014 , \29040 , \25367 );
nor \U$38637 ( \39015 , \39013 , \39014 );
xnor \U$38638 ( \39016 , \39015 , \25123 );
and \U$38639 ( \39017 , \39012 , \39016 );
and \U$38640 ( \39018 , \29715 , \24974 );
and \U$38641 ( \39019 , \29710 , \24972 );
nor \U$38642 ( \39020 , \39018 , \39019 );
xnor \U$38643 ( \39021 , \39020 , \24787 );
and \U$38644 ( \39022 , \39016 , \39021 );
and \U$38645 ( \39023 , \39012 , \39021 );
or \U$38646 ( \39024 , \39017 , \39022 , \39023 );
and \U$38647 ( \39025 , \39007 , \39024 );
and \U$38648 ( \39026 , \38991 , \39024 );
or \U$38649 ( \39027 , \39008 , \39025 , \39026 );
and \U$38650 ( \39028 , \25806 , \28575 );
and \U$38651 ( \39029 , \25609 , \28573 );
nor \U$38652 ( \39030 , \39028 , \39029 );
xnor \U$38653 ( \39031 , \39030 , \28315 );
and \U$38654 ( \39032 , \26116 , \28081 );
and \U$38655 ( \39033 , \26108 , \28079 );
nor \U$38656 ( \39034 , \39032 , \39033 );
xnor \U$38657 ( \39035 , \39034 , \27766 );
and \U$38658 ( \39036 , \39031 , \39035 );
and \U$38659 ( \39037 , \26590 , \27572 );
and \U$38660 ( \39038 , \26585 , \27570 );
nor \U$38661 ( \39039 , \39037 , \39038 );
xnor \U$38662 ( \39040 , \39039 , \27232 );
and \U$38663 ( \39041 , \39035 , \39040 );
and \U$38664 ( \39042 , \39031 , \39040 );
or \U$38665 ( \39043 , \39036 , \39041 , \39042 );
and \U$38666 ( \39044 , \24601 , \30233 );
and \U$38667 ( \39045 , \24482 , \30231 );
nor \U$38668 ( \39046 , \39044 , \39045 );
xnor \U$38669 ( \39047 , \39046 , \29862 );
and \U$38670 ( \39048 , \25226 , \29671 );
and \U$38671 ( \39049 , \25018 , \29669 );
nor \U$38672 ( \39050 , \39048 , \39049 );
xnor \U$38673 ( \39051 , \39050 , \29353 );
and \U$38674 ( \39052 , \39047 , \39051 );
and \U$38675 ( \39053 , \25353 , \29104 );
and \U$38676 ( \39054 , \25348 , \29102 );
nor \U$38677 ( \39055 , \39053 , \39054 );
xnor \U$38678 ( \39056 , \39055 , \28855 );
and \U$38679 ( \39057 , \39051 , \39056 );
and \U$38680 ( \39058 , \39047 , \39056 );
or \U$38681 ( \39059 , \39052 , \39057 , \39058 );
and \U$38682 ( \39060 , \39043 , \39059 );
and \U$38683 ( \39061 , \23714 , \32151 );
and \U$38684 ( \39062 , \23570 , \32148 );
nor \U$38685 ( \39063 , \39061 , \39062 );
xnor \U$38686 ( \39064 , \39063 , \31096 );
and \U$38687 ( \39065 , \24003 , \31338 );
and \U$38688 ( \39066 , \23978 , \31336 );
nor \U$38689 ( \39067 , \39065 , \39066 );
xnor \U$38690 ( \39068 , \39067 , \31099 );
and \U$38691 ( \39069 , \39064 , \39068 );
and \U$38692 ( \39070 , \24344 , \30770 );
and \U$38693 ( \39071 , \24177 , \30768 );
nor \U$38694 ( \39072 , \39070 , \39071 );
xnor \U$38695 ( \39073 , \39072 , \30460 );
and \U$38696 ( \39074 , \39068 , \39073 );
and \U$38697 ( \39075 , \39064 , \39073 );
or \U$38698 ( \39076 , \39069 , \39074 , \39075 );
and \U$38699 ( \39077 , \39059 , \39076 );
and \U$38700 ( \39078 , \39043 , \39076 );
or \U$38701 ( \39079 , \39060 , \39077 , \39078 );
and \U$38702 ( \39080 , \39027 , \39079 );
xor \U$38703 ( \39081 , \38819 , \38823 );
xor \U$38704 ( \39082 , \39081 , \38826 );
xor \U$38705 ( \39083 , \38862 , \38866 );
xor \U$38706 ( \39084 , \39083 , \38871 );
and \U$38707 ( \39085 , \39082 , \39084 );
xor \U$38708 ( \39086 , \38879 , \38883 );
xor \U$38709 ( \39087 , \39086 , \38888 );
and \U$38710 ( \39088 , \39084 , \39087 );
and \U$38711 ( \39089 , \39082 , \39087 );
or \U$38712 ( \39090 , \39085 , \39088 , \39089 );
and \U$38713 ( \39091 , \39079 , \39090 );
and \U$38714 ( \39092 , \39027 , \39090 );
or \U$38715 ( \39093 , \39080 , \39091 , \39092 );
xor \U$38716 ( \39094 , \38779 , \38795 );
xor \U$38717 ( \39095 , \39094 , \38812 );
xor \U$38718 ( \39096 , \38829 , \38833 );
xor \U$38719 ( \39097 , \39096 , \38838 );
and \U$38720 ( \39098 , \39095 , \39097 );
xor \U$38721 ( \39099 , \38858 , \38874 );
xor \U$38722 ( \39100 , \39099 , \38891 );
and \U$38723 ( \39101 , \39097 , \39100 );
and \U$38724 ( \39102 , \39095 , \39100 );
or \U$38725 ( \39103 , \39098 , \39101 , \39102 );
and \U$38726 ( \39104 , \39093 , \39103 );
xor \U$38727 ( \39105 , \38846 , \38850 );
xor \U$38728 ( \39106 , \39105 , \38855 );
xor \U$38729 ( \39107 , \38783 , \38787 );
xor \U$38730 ( \39108 , \39107 , \38792 );
and \U$38731 ( \39109 , \39106 , \39108 );
xor \U$38732 ( \39110 , \38800 , \38804 );
xor \U$38733 ( \39111 , \39110 , \38809 );
and \U$38734 ( \39112 , \39108 , \39111 );
and \U$38735 ( \39113 , \39106 , \39111 );
or \U$38736 ( \39114 , \39109 , \39112 , \39113 );
xor \U$38737 ( \39115 , \38899 , \38901 );
xor \U$38738 ( \39116 , \39115 , \38904 );
and \U$38739 ( \39117 , \39114 , \39116 );
xor \U$38740 ( \39118 , \38909 , \38911 );
xor \U$38741 ( \39119 , \39118 , \38914 );
and \U$38742 ( \39120 , \39116 , \39119 );
and \U$38743 ( \39121 , \39114 , \39119 );
or \U$38744 ( \39122 , \39117 , \39120 , \39121 );
and \U$38745 ( \39123 , \39103 , \39122 );
and \U$38746 ( \39124 , \39093 , \39122 );
or \U$38747 ( \39125 , \39104 , \39123 , \39124 );
xor \U$38748 ( \39126 , \38587 , \38603 );
xor \U$38749 ( \39127 , \39126 , \38620 );
xor \U$38750 ( \39128 , \38639 , \38655 );
xor \U$38751 ( \39129 , \39128 , \38672 );
and \U$38752 ( \39130 , \39127 , \39129 );
xor \U$38753 ( \39131 , \38926 , \38928 );
xor \U$38754 ( \39132 , \39131 , \38931 );
and \U$38755 ( \39133 , \39129 , \39132 );
and \U$38756 ( \39134 , \39127 , \39132 );
or \U$38757 ( \39135 , \39130 , \39133 , \39134 );
and \U$38758 ( \39136 , \39125 , \39135 );
xor \U$38759 ( \39137 , \38939 , \38941 );
xor \U$38760 ( \39138 , \39137 , \38944 );
and \U$38761 ( \39139 , \39135 , \39138 );
and \U$38762 ( \39140 , \39125 , \39138 );
or \U$38763 ( \39141 , \39136 , \39139 , \39140 );
xor \U$38764 ( \39142 , \38937 , \38947 );
xor \U$38765 ( \39143 , \39142 , \38950 );
and \U$38766 ( \39144 , \39141 , \39143 );
xor \U$38767 ( \39145 , \38955 , \38957 );
and \U$38768 ( \39146 , \39143 , \39145 );
and \U$38769 ( \39147 , \39141 , \39145 );
or \U$38770 ( \39148 , \39144 , \39146 , \39147 );
xor \U$38771 ( \39149 , \38720 , \38730 );
xor \U$38772 ( \39150 , \39149 , \38733 );
and \U$38773 ( \39151 , \39148 , \39150 );
xor \U$38774 ( \39152 , \38953 , \38958 );
xor \U$38775 ( \39153 , \39152 , \38961 );
and \U$38776 ( \39154 , \39150 , \39153 );
and \U$38777 ( \39155 , \39148 , \39153 );
or \U$38778 ( \39156 , \39151 , \39154 , \39155 );
and \U$38779 ( \39157 , \38975 , \39156 );
xor \U$38780 ( \39158 , \38975 , \39156 );
xor \U$38781 ( \39159 , \39148 , \39150 );
xor \U$38782 ( \39160 , \39159 , \39153 );
and \U$38783 ( \39161 , \25609 , \29104 );
and \U$38784 ( \39162 , \25353 , \29102 );
nor \U$38785 ( \39163 , \39161 , \39162 );
xnor \U$38786 ( \39164 , \39163 , \28855 );
and \U$38787 ( \39165 , \26108 , \28575 );
and \U$38788 ( \39166 , \25806 , \28573 );
nor \U$38789 ( \39167 , \39165 , \39166 );
xnor \U$38790 ( \39168 , \39167 , \28315 );
and \U$38791 ( \39169 , \39164 , \39168 );
and \U$38792 ( \39170 , \26585 , \28081 );
and \U$38793 ( \39171 , \26116 , \28079 );
nor \U$38794 ( \39172 , \39170 , \39171 );
xnor \U$38795 ( \39173 , \39172 , \27766 );
and \U$38796 ( \39174 , \39168 , \39173 );
and \U$38797 ( \39175 , \39164 , \39173 );
or \U$38798 ( \39176 , \39169 , \39174 , \39175 );
and \U$38799 ( \39177 , \24482 , \30770 );
and \U$38800 ( \39178 , \24344 , \30768 );
nor \U$38801 ( \39179 , \39177 , \39178 );
xnor \U$38802 ( \39180 , \39179 , \30460 );
and \U$38803 ( \39181 , \25018 , \30233 );
and \U$38804 ( \39182 , \24601 , \30231 );
nor \U$38805 ( \39183 , \39181 , \39182 );
xnor \U$38806 ( \39184 , \39183 , \29862 );
and \U$38807 ( \39185 , \39180 , \39184 );
and \U$38808 ( \39186 , \25348 , \29671 );
and \U$38809 ( \39187 , \25226 , \29669 );
nor \U$38810 ( \39188 , \39186 , \39187 );
xnor \U$38811 ( \39189 , \39188 , \29353 );
and \U$38812 ( \39190 , \39184 , \39189 );
and \U$38813 ( \39191 , \39180 , \39189 );
or \U$38814 ( \39192 , \39185 , \39190 , \39191 );
and \U$38815 ( \39193 , \39176 , \39192 );
and \U$38816 ( \39194 , \23978 , \32151 );
and \U$38817 ( \39195 , \23714 , \32148 );
nor \U$38818 ( \39196 , \39194 , \39195 );
xnor \U$38819 ( \39197 , \39196 , \31096 );
and \U$38820 ( \39198 , \24177 , \31338 );
and \U$38821 ( \39199 , \24003 , \31336 );
nor \U$38822 ( \39200 , \39198 , \39199 );
xnor \U$38823 ( \39201 , \39200 , \31099 );
and \U$38824 ( \39202 , \39197 , \39201 );
and \U$38825 ( \39203 , \39201 , \23500 );
and \U$38826 ( \39204 , \39197 , \23500 );
or \U$38827 ( \39205 , \39202 , \39203 , \39204 );
and \U$38828 ( \39206 , \39192 , \39205 );
and \U$38829 ( \39207 , \39176 , \39205 );
or \U$38830 ( \39208 , \39193 , \39206 , \39207 );
and \U$38831 ( \39209 , \30034 , \24974 );
and \U$38832 ( \39210 , \29715 , \24972 );
nor \U$38833 ( \39211 , \39209 , \39210 );
xnor \U$38834 ( \39212 , \39211 , \24787 );
and \U$38835 ( \39213 , \30887 , \24661 );
and \U$38836 ( \39214 , \30318 , \24659 );
nor \U$38837 ( \39215 , \39213 , \39214 );
xnor \U$38838 ( \39216 , \39215 , \24456 );
and \U$38839 ( \39217 , \39212 , \39216 );
and \U$38840 ( \39218 , \31498 , \24255 );
and \U$38841 ( \39219 , \30895 , \24253 );
nor \U$38842 ( \39220 , \39218 , \39219 );
xnor \U$38843 ( \39221 , \39220 , \24106 );
and \U$38844 ( \39222 , \39216 , \39221 );
and \U$38845 ( \39223 , \39212 , \39221 );
or \U$38846 ( \39224 , \39217 , \39222 , \39223 );
and \U$38847 ( \39225 , \26854 , \27572 );
and \U$38848 ( \39226 , \26590 , \27570 );
nor \U$38849 ( \39227 , \39225 , \39226 );
xnor \U$38850 ( \39228 , \39227 , \27232 );
and \U$38851 ( \39229 , \27485 , \26983 );
and \U$38852 ( \39230 , \27113 , \26981 );
nor \U$38853 ( \39231 , \39229 , \39230 );
xnor \U$38854 ( \39232 , \39231 , \26742 );
and \U$38855 ( \39233 , \39228 , \39232 );
and \U$38856 ( \39234 , \27837 , \26517 );
and \U$38857 ( \39235 , \27494 , \26515 );
nor \U$38858 ( \39236 , \39234 , \39235 );
xnor \U$38859 ( \39237 , \39236 , \26329 );
and \U$38860 ( \39238 , \39232 , \39237 );
and \U$38861 ( \39239 , \39228 , \39237 );
or \U$38862 ( \39240 , \39233 , \39238 , \39239 );
and \U$38863 ( \39241 , \39224 , \39240 );
and \U$38864 ( \39242 , \28342 , \26143 );
and \U$38865 ( \39243 , \28039 , \26141 );
nor \U$38866 ( \39244 , \39242 , \39243 );
xnor \U$38867 ( \39245 , \39244 , \25911 );
and \U$38868 ( \39246 , \29040 , \25692 );
and \U$38869 ( \39247 , \28514 , \25690 );
nor \U$38870 ( \39248 , \39246 , \39247 );
xnor \U$38871 ( \39249 , \39248 , \25549 );
and \U$38872 ( \39250 , \39245 , \39249 );
and \U$38873 ( \39251 , \29710 , \25369 );
and \U$38874 ( \39252 , \29464 , \25367 );
nor \U$38875 ( \39253 , \39251 , \39252 );
xnor \U$38876 ( \39254 , \39253 , \25123 );
and \U$38877 ( \39255 , \39249 , \39254 );
and \U$38878 ( \39256 , \39245 , \39254 );
or \U$38879 ( \39257 , \39250 , \39255 , \39256 );
and \U$38880 ( \39258 , \39240 , \39257 );
and \U$38881 ( \39259 , \39224 , \39257 );
or \U$38882 ( \39260 , \39241 , \39258 , \39259 );
and \U$38883 ( \39261 , \39208 , \39260 );
and \U$38884 ( \39262 , \32304 , \23637 );
and \U$38885 ( \39263 , \31684 , \23635 );
nor \U$38886 ( \39264 , \39262 , \39263 );
xnor \U$38887 ( \39265 , \39264 , \23500 );
xor \U$38888 ( \39266 , \38979 , \38983 );
xor \U$38889 ( \39267 , \39266 , \38988 );
and \U$38890 ( \39268 , \39265 , \39267 );
xor \U$38891 ( \39269 , \39012 , \39016 );
xor \U$38892 ( \39270 , \39269 , \39021 );
and \U$38893 ( \39271 , \39267 , \39270 );
and \U$38894 ( \39272 , \39265 , \39270 );
or \U$38895 ( \39273 , \39268 , \39271 , \39272 );
and \U$38896 ( \39274 , \39260 , \39273 );
and \U$38897 ( \39275 , \39208 , \39273 );
or \U$38898 ( \39276 , \39261 , \39274 , \39275 );
xor \U$38899 ( \39277 , \39031 , \39035 );
xor \U$38900 ( \39278 , \39277 , \39040 );
xor \U$38901 ( \39279 , \38995 , \38999 );
xor \U$38902 ( \39280 , \39279 , \39004 );
and \U$38903 ( \39281 , \39278 , \39280 );
xor \U$38904 ( \39282 , \39047 , \39051 );
xor \U$38905 ( \39283 , \39282 , \39056 );
and \U$38906 ( \39284 , \39280 , \39283 );
and \U$38907 ( \39285 , \39278 , \39283 );
or \U$38908 ( \39286 , \39281 , \39284 , \39285 );
xor \U$38909 ( \39287 , \38771 , \38775 );
xor \U$38910 ( \39288 , \39287 , \23279 );
and \U$38911 ( \39289 , \39286 , \39288 );
xor \U$38912 ( \39290 , \39106 , \39108 );
xor \U$38913 ( \39291 , \39290 , \39111 );
and \U$38914 ( \39292 , \39288 , \39291 );
and \U$38915 ( \39293 , \39286 , \39291 );
or \U$38916 ( \39294 , \39289 , \39292 , \39293 );
and \U$38917 ( \39295 , \39276 , \39294 );
xor \U$38918 ( \39296 , \38991 , \39007 );
xor \U$38919 ( \39297 , \39296 , \39024 );
xor \U$38920 ( \39298 , \39043 , \39059 );
xor \U$38921 ( \39299 , \39298 , \39076 );
and \U$38922 ( \39300 , \39297 , \39299 );
xor \U$38923 ( \39301 , \39082 , \39084 );
xor \U$38924 ( \39302 , \39301 , \39087 );
and \U$38925 ( \39303 , \39299 , \39302 );
and \U$38926 ( \39304 , \39297 , \39302 );
or \U$38927 ( \39305 , \39300 , \39303 , \39304 );
and \U$38928 ( \39306 , \39294 , \39305 );
and \U$38929 ( \39307 , \39276 , \39305 );
or \U$38930 ( \39308 , \39295 , \39306 , \39307 );
xor \U$38931 ( \39309 , \39027 , \39079 );
xor \U$38932 ( \39310 , \39309 , \39090 );
xor \U$38933 ( \39311 , \39095 , \39097 );
xor \U$38934 ( \39312 , \39311 , \39100 );
and \U$38935 ( \39313 , \39310 , \39312 );
xor \U$38936 ( \39314 , \39114 , \39116 );
xor \U$38937 ( \39315 , \39314 , \39119 );
and \U$38938 ( \39316 , \39312 , \39315 );
and \U$38939 ( \39317 , \39310 , \39315 );
or \U$38940 ( \39318 , \39313 , \39316 , \39317 );
and \U$38941 ( \39319 , \39308 , \39318 );
xor \U$38942 ( \39320 , \38907 , \38917 );
xor \U$38943 ( \39321 , \39320 , \38920 );
and \U$38944 ( \39322 , \39318 , \39321 );
and \U$38945 ( \39323 , \39308 , \39321 );
or \U$38946 ( \39324 , \39319 , \39322 , \39323 );
xor \U$38947 ( \39325 , \38815 , \38841 );
xor \U$38948 ( \39326 , \39325 , \38894 );
xor \U$38949 ( \39327 , \39093 , \39103 );
xor \U$38950 ( \39328 , \39327 , \39122 );
and \U$38951 ( \39329 , \39326 , \39328 );
xor \U$38952 ( \39330 , \39127 , \39129 );
xor \U$38953 ( \39331 , \39330 , \39132 );
and \U$38954 ( \39332 , \39328 , \39331 );
and \U$38955 ( \39333 , \39326 , \39331 );
or \U$38956 ( \39334 , \39329 , \39332 , \39333 );
and \U$38957 ( \39335 , \39324 , \39334 );
xor \U$38958 ( \39336 , \38897 , \38923 );
xor \U$38959 ( \39337 , \39336 , \38934 );
and \U$38960 ( \39338 , \39334 , \39337 );
and \U$38961 ( \39339 , \39324 , \39337 );
or \U$38962 ( \39340 , \39335 , \39338 , \39339 );
xor \U$38963 ( \39341 , \39141 , \39143 );
xor \U$38964 ( \39342 , \39341 , \39145 );
and \U$38965 ( \39343 , \39340 , \39342 );
and \U$38966 ( \39344 , \39160 , \39343 );
xor \U$38967 ( \39345 , \39160 , \39343 );
xor \U$38968 ( \39346 , \39340 , \39342 );
and \U$38969 ( \39347 , \24003 , \32151 );
and \U$38970 ( \39348 , \23978 , \32148 );
nor \U$38971 ( \39349 , \39347 , \39348 );
xnor \U$38972 ( \39350 , \39349 , \31096 );
and \U$38973 ( \39351 , \24344 , \31338 );
and \U$38974 ( \39352 , \24177 , \31336 );
nor \U$38975 ( \39353 , \39351 , \39352 );
xnor \U$38976 ( \39354 , \39353 , \31099 );
and \U$38977 ( \39355 , \39350 , \39354 );
and \U$38978 ( \39356 , \24601 , \30770 );
and \U$38979 ( \39357 , \24482 , \30768 );
nor \U$38980 ( \39358 , \39356 , \39357 );
xnor \U$38981 ( \39359 , \39358 , \30460 );
and \U$38982 ( \39360 , \39354 , \39359 );
and \U$38983 ( \39361 , \39350 , \39359 );
or \U$38984 ( \39362 , \39355 , \39360 , \39361 );
and \U$38985 ( \39363 , \25226 , \30233 );
and \U$38986 ( \39364 , \25018 , \30231 );
nor \U$38987 ( \39365 , \39363 , \39364 );
xnor \U$38988 ( \39366 , \39365 , \29862 );
and \U$38989 ( \39367 , \25353 , \29671 );
and \U$38990 ( \39368 , \25348 , \29669 );
nor \U$38991 ( \39369 , \39367 , \39368 );
xnor \U$38992 ( \39370 , \39369 , \29353 );
and \U$38993 ( \39371 , \39366 , \39370 );
and \U$38994 ( \39372 , \25806 , \29104 );
and \U$38995 ( \39373 , \25609 , \29102 );
nor \U$38996 ( \39374 , \39372 , \39373 );
xnor \U$38997 ( \39375 , \39374 , \28855 );
and \U$38998 ( \39376 , \39370 , \39375 );
and \U$38999 ( \39377 , \39366 , \39375 );
or \U$39000 ( \39378 , \39371 , \39376 , \39377 );
and \U$39001 ( \39379 , \39362 , \39378 );
and \U$39002 ( \39380 , \26116 , \28575 );
and \U$39003 ( \39381 , \26108 , \28573 );
nor \U$39004 ( \39382 , \39380 , \39381 );
xnor \U$39005 ( \39383 , \39382 , \28315 );
and \U$39006 ( \39384 , \26590 , \28081 );
and \U$39007 ( \39385 , \26585 , \28079 );
nor \U$39008 ( \39386 , \39384 , \39385 );
xnor \U$39009 ( \39387 , \39386 , \27766 );
and \U$39010 ( \39388 , \39383 , \39387 );
and \U$39011 ( \39389 , \27113 , \27572 );
and \U$39012 ( \39390 , \26854 , \27570 );
nor \U$39013 ( \39391 , \39389 , \39390 );
xnor \U$39014 ( \39392 , \39391 , \27232 );
and \U$39015 ( \39393 , \39387 , \39392 );
and \U$39016 ( \39394 , \39383 , \39392 );
or \U$39017 ( \39395 , \39388 , \39393 , \39394 );
and \U$39018 ( \39396 , \39378 , \39395 );
and \U$39019 ( \39397 , \39362 , \39395 );
or \U$39020 ( \39398 , \39379 , \39396 , \39397 );
and \U$39021 ( \39399 , \30895 , \24661 );
and \U$39022 ( \39400 , \30887 , \24659 );
nor \U$39023 ( \39401 , \39399 , \39400 );
xnor \U$39024 ( \39402 , \39401 , \24456 );
and \U$39025 ( \39403 , \31503 , \24255 );
and \U$39026 ( \39404 , \31498 , \24253 );
nor \U$39027 ( \39405 , \39403 , \39404 );
xnor \U$39028 ( \39406 , \39405 , \24106 );
and \U$39029 ( \39407 , \39402 , \39406 );
and \U$39030 ( \39408 , \32304 , \23933 );
and \U$39031 ( \39409 , \31684 , \23931 );
nor \U$39032 ( \39410 , \39408 , \39409 );
xnor \U$39033 ( \39411 , \39410 , \23791 );
and \U$39034 ( \39412 , \39406 , \39411 );
and \U$39035 ( \39413 , \39402 , \39411 );
or \U$39036 ( \39414 , \39407 , \39412 , \39413 );
and \U$39037 ( \39415 , \29464 , \25692 );
and \U$39038 ( \39416 , \29040 , \25690 );
nor \U$39039 ( \39417 , \39415 , \39416 );
xnor \U$39040 ( \39418 , \39417 , \25549 );
and \U$39041 ( \39419 , \29715 , \25369 );
and \U$39042 ( \39420 , \29710 , \25367 );
nor \U$39043 ( \39421 , \39419 , \39420 );
xnor \U$39044 ( \39422 , \39421 , \25123 );
and \U$39045 ( \39423 , \39418 , \39422 );
and \U$39046 ( \39424 , \30318 , \24974 );
and \U$39047 ( \39425 , \30034 , \24972 );
nor \U$39048 ( \39426 , \39424 , \39425 );
xnor \U$39049 ( \39427 , \39426 , \24787 );
and \U$39050 ( \39428 , \39422 , \39427 );
and \U$39051 ( \39429 , \39418 , \39427 );
or \U$39052 ( \39430 , \39423 , \39428 , \39429 );
and \U$39053 ( \39431 , \39414 , \39430 );
and \U$39054 ( \39432 , \27494 , \26983 );
and \U$39055 ( \39433 , \27485 , \26981 );
nor \U$39056 ( \39434 , \39432 , \39433 );
xnor \U$39057 ( \39435 , \39434 , \26742 );
and \U$39058 ( \39436 , \28039 , \26517 );
and \U$39059 ( \39437 , \27837 , \26515 );
nor \U$39060 ( \39438 , \39436 , \39437 );
xnor \U$39061 ( \39439 , \39438 , \26329 );
and \U$39062 ( \39440 , \39435 , \39439 );
and \U$39063 ( \39441 , \28514 , \26143 );
and \U$39064 ( \39442 , \28342 , \26141 );
nor \U$39065 ( \39443 , \39441 , \39442 );
xnor \U$39066 ( \39444 , \39443 , \25911 );
and \U$39067 ( \39445 , \39439 , \39444 );
and \U$39068 ( \39446 , \39435 , \39444 );
or \U$39069 ( \39447 , \39440 , \39445 , \39446 );
and \U$39070 ( \39448 , \39430 , \39447 );
and \U$39071 ( \39449 , \39414 , \39447 );
or \U$39072 ( \39450 , \39431 , \39448 , \39449 );
and \U$39073 ( \39451 , \39398 , \39450 );
and \U$39074 ( \39452 , \31684 , \23933 );
and \U$39075 ( \39453 , \31503 , \23931 );
nor \U$39076 ( \39454 , \39452 , \39453 );
xnor \U$39077 ( \39455 , \39454 , \23791 );
nand \U$39078 ( \39456 , \32304 , \23635 );
xnor \U$39079 ( \39457 , \39456 , \23500 );
and \U$39080 ( \39458 , \39455 , \39457 );
xor \U$39081 ( \39459 , \39212 , \39216 );
xor \U$39082 ( \39460 , \39459 , \39221 );
and \U$39083 ( \39461 , \39457 , \39460 );
and \U$39084 ( \39462 , \39455 , \39460 );
or \U$39085 ( \39463 , \39458 , \39461 , \39462 );
and \U$39086 ( \39464 , \39450 , \39463 );
and \U$39087 ( \39465 , \39398 , \39463 );
or \U$39088 ( \39466 , \39451 , \39464 , \39465 );
xor \U$39089 ( \39467 , \39164 , \39168 );
xor \U$39090 ( \39468 , \39467 , \39173 );
xor \U$39091 ( \39469 , \39228 , \39232 );
xor \U$39092 ( \39470 , \39469 , \39237 );
and \U$39093 ( \39471 , \39468 , \39470 );
xor \U$39094 ( \39472 , \39245 , \39249 );
xor \U$39095 ( \39473 , \39472 , \39254 );
and \U$39096 ( \39474 , \39470 , \39473 );
and \U$39097 ( \39475 , \39468 , \39473 );
or \U$39098 ( \39476 , \39471 , \39474 , \39475 );
xor \U$39099 ( \39477 , \39180 , \39184 );
xor \U$39100 ( \39478 , \39477 , \39189 );
xor \U$39101 ( \39479 , \39197 , \39201 );
xor \U$39102 ( \39480 , \39479 , \23500 );
and \U$39103 ( \39481 , \39478 , \39480 );
and \U$39104 ( \39482 , \39476 , \39481 );
xor \U$39105 ( \39483 , \39064 , \39068 );
xor \U$39106 ( \39484 , \39483 , \39073 );
and \U$39107 ( \39485 , \39481 , \39484 );
and \U$39108 ( \39486 , \39476 , \39484 );
or \U$39109 ( \39487 , \39482 , \39485 , \39486 );
and \U$39110 ( \39488 , \39466 , \39487 );
xor \U$39111 ( \39489 , \39224 , \39240 );
xor \U$39112 ( \39490 , \39489 , \39257 );
xor \U$39113 ( \39491 , \39278 , \39280 );
xor \U$39114 ( \39492 , \39491 , \39283 );
and \U$39115 ( \39493 , \39490 , \39492 );
xor \U$39116 ( \39494 , \39265 , \39267 );
xor \U$39117 ( \39495 , \39494 , \39270 );
and \U$39118 ( \39496 , \39492 , \39495 );
and \U$39119 ( \39497 , \39490 , \39495 );
or \U$39120 ( \39498 , \39493 , \39496 , \39497 );
and \U$39121 ( \39499 , \39487 , \39498 );
and \U$39122 ( \39500 , \39466 , \39498 );
or \U$39123 ( \39501 , \39488 , \39499 , \39500 );
xor \U$39124 ( \39502 , \39208 , \39260 );
xor \U$39125 ( \39503 , \39502 , \39273 );
xor \U$39126 ( \39504 , \39286 , \39288 );
xor \U$39127 ( \39505 , \39504 , \39291 );
and \U$39128 ( \39506 , \39503 , \39505 );
xor \U$39129 ( \39507 , \39297 , \39299 );
xor \U$39130 ( \39508 , \39507 , \39302 );
and \U$39131 ( \39509 , \39505 , \39508 );
and \U$39132 ( \39510 , \39503 , \39508 );
or \U$39133 ( \39511 , \39506 , \39509 , \39510 );
and \U$39134 ( \39512 , \39501 , \39511 );
xor \U$39135 ( \39513 , \39310 , \39312 );
xor \U$39136 ( \39514 , \39513 , \39315 );
and \U$39137 ( \39515 , \39511 , \39514 );
and \U$39138 ( \39516 , \39501 , \39514 );
or \U$39139 ( \39517 , \39512 , \39515 , \39516 );
xor \U$39140 ( \39518 , \39308 , \39318 );
xor \U$39141 ( \39519 , \39518 , \39321 );
and \U$39142 ( \39520 , \39517 , \39519 );
xor \U$39143 ( \39521 , \39326 , \39328 );
xor \U$39144 ( \39522 , \39521 , \39331 );
and \U$39145 ( \39523 , \39519 , \39522 );
and \U$39146 ( \39524 , \39517 , \39522 );
or \U$39147 ( \39525 , \39520 , \39523 , \39524 );
xor \U$39148 ( \39526 , \39324 , \39334 );
xor \U$39149 ( \39527 , \39526 , \39337 );
and \U$39150 ( \39528 , \39525 , \39527 );
xor \U$39151 ( \39529 , \39125 , \39135 );
xor \U$39152 ( \39530 , \39529 , \39138 );
and \U$39153 ( \39531 , \39527 , \39530 );
and \U$39154 ( \39532 , \39525 , \39530 );
or \U$39155 ( \39533 , \39528 , \39531 , \39532 );
and \U$39156 ( \39534 , \39346 , \39533 );
xor \U$39157 ( \39535 , \39346 , \39533 );
xor \U$39158 ( \39536 , \39525 , \39527 );
xor \U$39159 ( \39537 , \39536 , \39530 );
and \U$39160 ( \39538 , \24177 , \32151 );
and \U$39161 ( \39539 , \24003 , \32148 );
nor \U$39162 ( \39540 , \39538 , \39539 );
xnor \U$39163 ( \39541 , \39540 , \31096 );
and \U$39164 ( \39542 , \24482 , \31338 );
and \U$39165 ( \39543 , \24344 , \31336 );
nor \U$39166 ( \39544 , \39542 , \39543 );
xnor \U$39167 ( \39545 , \39544 , \31099 );
and \U$39168 ( \39546 , \39541 , \39545 );
and \U$39169 ( \39547 , \39545 , \23791 );
and \U$39170 ( \39548 , \39541 , \23791 );
or \U$39171 ( \39549 , \39546 , \39547 , \39548 );
and \U$39172 ( \39550 , \25018 , \30770 );
and \U$39173 ( \39551 , \24601 , \30768 );
nor \U$39174 ( \39552 , \39550 , \39551 );
xnor \U$39175 ( \39553 , \39552 , \30460 );
and \U$39176 ( \39554 , \25348 , \30233 );
and \U$39177 ( \39555 , \25226 , \30231 );
nor \U$39178 ( \39556 , \39554 , \39555 );
xnor \U$39179 ( \39557 , \39556 , \29862 );
and \U$39180 ( \39558 , \39553 , \39557 );
and \U$39181 ( \39559 , \25609 , \29671 );
and \U$39182 ( \39560 , \25353 , \29669 );
nor \U$39183 ( \39561 , \39559 , \39560 );
xnor \U$39184 ( \39562 , \39561 , \29353 );
and \U$39185 ( \39563 , \39557 , \39562 );
and \U$39186 ( \39564 , \39553 , \39562 );
or \U$39187 ( \39565 , \39558 , \39563 , \39564 );
and \U$39188 ( \39566 , \39549 , \39565 );
and \U$39189 ( \39567 , \26108 , \29104 );
and \U$39190 ( \39568 , \25806 , \29102 );
nor \U$39191 ( \39569 , \39567 , \39568 );
xnor \U$39192 ( \39570 , \39569 , \28855 );
and \U$39193 ( \39571 , \26585 , \28575 );
and \U$39194 ( \39572 , \26116 , \28573 );
nor \U$39195 ( \39573 , \39571 , \39572 );
xnor \U$39196 ( \39574 , \39573 , \28315 );
and \U$39197 ( \39575 , \39570 , \39574 );
and \U$39198 ( \39576 , \26854 , \28081 );
and \U$39199 ( \39577 , \26590 , \28079 );
nor \U$39200 ( \39578 , \39576 , \39577 );
xnor \U$39201 ( \39579 , \39578 , \27766 );
and \U$39202 ( \39580 , \39574 , \39579 );
and \U$39203 ( \39581 , \39570 , \39579 );
or \U$39204 ( \39582 , \39575 , \39580 , \39581 );
and \U$39205 ( \39583 , \39565 , \39582 );
and \U$39206 ( \39584 , \39549 , \39582 );
or \U$39207 ( \39585 , \39566 , \39583 , \39584 );
and \U$39208 ( \39586 , \27485 , \27572 );
and \U$39209 ( \39587 , \27113 , \27570 );
nor \U$39210 ( \39588 , \39586 , \39587 );
xnor \U$39211 ( \39589 , \39588 , \27232 );
and \U$39212 ( \39590 , \27837 , \26983 );
and \U$39213 ( \39591 , \27494 , \26981 );
nor \U$39214 ( \39592 , \39590 , \39591 );
xnor \U$39215 ( \39593 , \39592 , \26742 );
and \U$39216 ( \39594 , \39589 , \39593 );
and \U$39217 ( \39595 , \28342 , \26517 );
and \U$39218 ( \39596 , \28039 , \26515 );
nor \U$39219 ( \39597 , \39595 , \39596 );
xnor \U$39220 ( \39598 , \39597 , \26329 );
and \U$39221 ( \39599 , \39593 , \39598 );
and \U$39222 ( \39600 , \39589 , \39598 );
or \U$39223 ( \39601 , \39594 , \39599 , \39600 );
and \U$39224 ( \39602 , \29040 , \26143 );
and \U$39225 ( \39603 , \28514 , \26141 );
nor \U$39226 ( \39604 , \39602 , \39603 );
xnor \U$39227 ( \39605 , \39604 , \25911 );
and \U$39228 ( \39606 , \29710 , \25692 );
and \U$39229 ( \39607 , \29464 , \25690 );
nor \U$39230 ( \39608 , \39606 , \39607 );
xnor \U$39231 ( \39609 , \39608 , \25549 );
and \U$39232 ( \39610 , \39605 , \39609 );
and \U$39233 ( \39611 , \30034 , \25369 );
and \U$39234 ( \39612 , \29715 , \25367 );
nor \U$39235 ( \39613 , \39611 , \39612 );
xnor \U$39236 ( \39614 , \39613 , \25123 );
and \U$39237 ( \39615 , \39609 , \39614 );
and \U$39238 ( \39616 , \39605 , \39614 );
or \U$39239 ( \39617 , \39610 , \39615 , \39616 );
and \U$39240 ( \39618 , \39601 , \39617 );
and \U$39241 ( \39619 , \30887 , \24974 );
and \U$39242 ( \39620 , \30318 , \24972 );
nor \U$39243 ( \39621 , \39619 , \39620 );
xnor \U$39244 ( \39622 , \39621 , \24787 );
and \U$39245 ( \39623 , \31498 , \24661 );
and \U$39246 ( \39624 , \30895 , \24659 );
nor \U$39247 ( \39625 , \39623 , \39624 );
xnor \U$39248 ( \39626 , \39625 , \24456 );
and \U$39249 ( \39627 , \39622 , \39626 );
and \U$39250 ( \39628 , \31684 , \24255 );
and \U$39251 ( \39629 , \31503 , \24253 );
nor \U$39252 ( \39630 , \39628 , \39629 );
xnor \U$39253 ( \39631 , \39630 , \24106 );
and \U$39254 ( \39632 , \39626 , \39631 );
and \U$39255 ( \39633 , \39622 , \39631 );
or \U$39256 ( \39634 , \39627 , \39632 , \39633 );
and \U$39257 ( \39635 , \39617 , \39634 );
and \U$39258 ( \39636 , \39601 , \39634 );
or \U$39259 ( \39637 , \39618 , \39635 , \39636 );
and \U$39260 ( \39638 , \39585 , \39637 );
xor \U$39261 ( \39639 , \39402 , \39406 );
xor \U$39262 ( \39640 , \39639 , \39411 );
xor \U$39263 ( \39641 , \39418 , \39422 );
xor \U$39264 ( \39642 , \39641 , \39427 );
and \U$39265 ( \39643 , \39640 , \39642 );
xor \U$39266 ( \39644 , \39435 , \39439 );
xor \U$39267 ( \39645 , \39644 , \39444 );
and \U$39268 ( \39646 , \39642 , \39645 );
and \U$39269 ( \39647 , \39640 , \39645 );
or \U$39270 ( \39648 , \39643 , \39646 , \39647 );
and \U$39271 ( \39649 , \39637 , \39648 );
and \U$39272 ( \39650 , \39585 , \39648 );
or \U$39273 ( \39651 , \39638 , \39649 , \39650 );
xor \U$39274 ( \39652 , \39362 , \39378 );
xor \U$39275 ( \39653 , \39652 , \39395 );
xor \U$39276 ( \39654 , \39414 , \39430 );
xor \U$39277 ( \39655 , \39654 , \39447 );
and \U$39278 ( \39656 , \39653 , \39655 );
xor \U$39279 ( \39657 , \39455 , \39457 );
xor \U$39280 ( \39658 , \39657 , \39460 );
and \U$39281 ( \39659 , \39655 , \39658 );
and \U$39282 ( \39660 , \39653 , \39658 );
or \U$39283 ( \39661 , \39656 , \39659 , \39660 );
and \U$39284 ( \39662 , \39651 , \39661 );
xor \U$39285 ( \39663 , \39350 , \39354 );
xor \U$39286 ( \39664 , \39663 , \39359 );
xor \U$39287 ( \39665 , \39366 , \39370 );
xor \U$39288 ( \39666 , \39665 , \39375 );
and \U$39289 ( \39667 , \39664 , \39666 );
xor \U$39290 ( \39668 , \39383 , \39387 );
xor \U$39291 ( \39669 , \39668 , \39392 );
and \U$39292 ( \39670 , \39666 , \39669 );
and \U$39293 ( \39671 , \39664 , \39669 );
or \U$39294 ( \39672 , \39667 , \39670 , \39671 );
xor \U$39295 ( \39673 , \39468 , \39470 );
xor \U$39296 ( \39674 , \39673 , \39473 );
and \U$39297 ( \39675 , \39672 , \39674 );
xor \U$39298 ( \39676 , \39478 , \39480 );
and \U$39299 ( \39677 , \39674 , \39676 );
and \U$39300 ( \39678 , \39672 , \39676 );
or \U$39301 ( \39679 , \39675 , \39677 , \39678 );
and \U$39302 ( \39680 , \39661 , \39679 );
and \U$39303 ( \39681 , \39651 , \39679 );
or \U$39304 ( \39682 , \39662 , \39680 , \39681 );
xor \U$39305 ( \39683 , \39176 , \39192 );
xor \U$39306 ( \39684 , \39683 , \39205 );
xor \U$39307 ( \39685 , \39476 , \39481 );
xor \U$39308 ( \39686 , \39685 , \39484 );
and \U$39309 ( \39687 , \39684 , \39686 );
xor \U$39310 ( \39688 , \39490 , \39492 );
xor \U$39311 ( \39689 , \39688 , \39495 );
and \U$39312 ( \39690 , \39686 , \39689 );
and \U$39313 ( \39691 , \39684 , \39689 );
or \U$39314 ( \39692 , \39687 , \39690 , \39691 );
and \U$39315 ( \39693 , \39682 , \39692 );
xor \U$39316 ( \39694 , \39503 , \39505 );
xor \U$39317 ( \39695 , \39694 , \39508 );
and \U$39318 ( \39696 , \39692 , \39695 );
and \U$39319 ( \39697 , \39682 , \39695 );
or \U$39320 ( \39698 , \39693 , \39696 , \39697 );
xor \U$39321 ( \39699 , \39276 , \39294 );
xor \U$39322 ( \39700 , \39699 , \39305 );
and \U$39323 ( \39701 , \39698 , \39700 );
xor \U$39324 ( \39702 , \39501 , \39511 );
xor \U$39325 ( \39703 , \39702 , \39514 );
and \U$39326 ( \39704 , \39700 , \39703 );
and \U$39327 ( \39705 , \39698 , \39703 );
or \U$39328 ( \39706 , \39701 , \39704 , \39705 );
xor \U$39329 ( \39707 , \39517 , \39519 );
xor \U$39330 ( \39708 , \39707 , \39522 );
and \U$39331 ( \39709 , \39706 , \39708 );
and \U$39332 ( \39710 , \39537 , \39709 );
xor \U$39333 ( \39711 , \39537 , \39709 );
xor \U$39334 ( \39712 , \39706 , \39708 );
and \U$39335 ( \39713 , \26590 , \28575 );
and \U$39336 ( \39714 , \26585 , \28573 );
nor \U$39337 ( \39715 , \39713 , \39714 );
xnor \U$39338 ( \39716 , \39715 , \28315 );
and \U$39339 ( \39717 , \27113 , \28081 );
and \U$39340 ( \39718 , \26854 , \28079 );
nor \U$39341 ( \39719 , \39717 , \39718 );
xnor \U$39342 ( \39720 , \39719 , \27766 );
and \U$39343 ( \39721 , \39716 , \39720 );
and \U$39344 ( \39722 , \27494 , \27572 );
and \U$39345 ( \39723 , \27485 , \27570 );
nor \U$39346 ( \39724 , \39722 , \39723 );
xnor \U$39347 ( \39725 , \39724 , \27232 );
and \U$39348 ( \39726 , \39720 , \39725 );
and \U$39349 ( \39727 , \39716 , \39725 );
or \U$39350 ( \39728 , \39721 , \39726 , \39727 );
and \U$39351 ( \39729 , \24344 , \32151 );
and \U$39352 ( \39730 , \24177 , \32148 );
nor \U$39353 ( \39731 , \39729 , \39730 );
xnor \U$39354 ( \39732 , \39731 , \31096 );
and \U$39355 ( \39733 , \24601 , \31338 );
and \U$39356 ( \39734 , \24482 , \31336 );
nor \U$39357 ( \39735 , \39733 , \39734 );
xnor \U$39358 ( \39736 , \39735 , \31099 );
and \U$39359 ( \39737 , \39732 , \39736 );
and \U$39360 ( \39738 , \25226 , \30770 );
and \U$39361 ( \39739 , \25018 , \30768 );
nor \U$39362 ( \39740 , \39738 , \39739 );
xnor \U$39363 ( \39741 , \39740 , \30460 );
and \U$39364 ( \39742 , \39736 , \39741 );
and \U$39365 ( \39743 , \39732 , \39741 );
or \U$39366 ( \39744 , \39737 , \39742 , \39743 );
and \U$39367 ( \39745 , \39728 , \39744 );
and \U$39368 ( \39746 , \25353 , \30233 );
and \U$39369 ( \39747 , \25348 , \30231 );
nor \U$39370 ( \39748 , \39746 , \39747 );
xnor \U$39371 ( \39749 , \39748 , \29862 );
and \U$39372 ( \39750 , \25806 , \29671 );
and \U$39373 ( \39751 , \25609 , \29669 );
nor \U$39374 ( \39752 , \39750 , \39751 );
xnor \U$39375 ( \39753 , \39752 , \29353 );
and \U$39376 ( \39754 , \39749 , \39753 );
and \U$39377 ( \39755 , \26116 , \29104 );
and \U$39378 ( \39756 , \26108 , \29102 );
nor \U$39379 ( \39757 , \39755 , \39756 );
xnor \U$39380 ( \39758 , \39757 , \28855 );
and \U$39381 ( \39759 , \39753 , \39758 );
and \U$39382 ( \39760 , \39749 , \39758 );
or \U$39383 ( \39761 , \39754 , \39759 , \39760 );
and \U$39384 ( \39762 , \39744 , \39761 );
and \U$39385 ( \39763 , \39728 , \39761 );
or \U$39386 ( \39764 , \39745 , \39762 , \39763 );
and \U$39387 ( \39765 , \29715 , \25692 );
and \U$39388 ( \39766 , \29710 , \25690 );
nor \U$39389 ( \39767 , \39765 , \39766 );
xnor \U$39390 ( \39768 , \39767 , \25549 );
and \U$39391 ( \39769 , \30318 , \25369 );
and \U$39392 ( \39770 , \30034 , \25367 );
nor \U$39393 ( \39771 , \39769 , \39770 );
xnor \U$39394 ( \39772 , \39771 , \25123 );
and \U$39395 ( \39773 , \39768 , \39772 );
and \U$39396 ( \39774 , \30895 , \24974 );
and \U$39397 ( \39775 , \30887 , \24972 );
nor \U$39398 ( \39776 , \39774 , \39775 );
xnor \U$39399 ( \39777 , \39776 , \24787 );
and \U$39400 ( \39778 , \39772 , \39777 );
and \U$39401 ( \39779 , \39768 , \39777 );
or \U$39402 ( \39780 , \39773 , \39778 , \39779 );
and \U$39403 ( \39781 , \28039 , \26983 );
and \U$39404 ( \39782 , \27837 , \26981 );
nor \U$39405 ( \39783 , \39781 , \39782 );
xnor \U$39406 ( \39784 , \39783 , \26742 );
and \U$39407 ( \39785 , \28514 , \26517 );
and \U$39408 ( \39786 , \28342 , \26515 );
nor \U$39409 ( \39787 , \39785 , \39786 );
xnor \U$39410 ( \39788 , \39787 , \26329 );
and \U$39411 ( \39789 , \39784 , \39788 );
and \U$39412 ( \39790 , \29464 , \26143 );
and \U$39413 ( \39791 , \29040 , \26141 );
nor \U$39414 ( \39792 , \39790 , \39791 );
xnor \U$39415 ( \39793 , \39792 , \25911 );
and \U$39416 ( \39794 , \39788 , \39793 );
and \U$39417 ( \39795 , \39784 , \39793 );
or \U$39418 ( \39796 , \39789 , \39794 , \39795 );
and \U$39419 ( \39797 , \39780 , \39796 );
and \U$39420 ( \39798 , \31503 , \24661 );
and \U$39421 ( \39799 , \31498 , \24659 );
nor \U$39422 ( \39800 , \39798 , \39799 );
xnor \U$39423 ( \39801 , \39800 , \24456 );
and \U$39424 ( \39802 , \32304 , \24255 );
and \U$39425 ( \39803 , \31684 , \24253 );
nor \U$39426 ( \39804 , \39802 , \39803 );
xnor \U$39427 ( \39805 , \39804 , \24106 );
and \U$39428 ( \39806 , \39801 , \39805 );
and \U$39429 ( \39807 , \39796 , \39806 );
and \U$39430 ( \39808 , \39780 , \39806 );
or \U$39431 ( \39809 , \39797 , \39807 , \39808 );
and \U$39432 ( \39810 , \39764 , \39809 );
nand \U$39433 ( \39811 , \32304 , \23931 );
xnor \U$39434 ( \39812 , \39811 , \23791 );
xor \U$39435 ( \39813 , \39605 , \39609 );
xor \U$39436 ( \39814 , \39813 , \39614 );
and \U$39437 ( \39815 , \39812 , \39814 );
xor \U$39438 ( \39816 , \39622 , \39626 );
xor \U$39439 ( \39817 , \39816 , \39631 );
and \U$39440 ( \39818 , \39814 , \39817 );
and \U$39441 ( \39819 , \39812 , \39817 );
or \U$39442 ( \39820 , \39815 , \39818 , \39819 );
and \U$39443 ( \39821 , \39809 , \39820 );
and \U$39444 ( \39822 , \39764 , \39820 );
or \U$39445 ( \39823 , \39810 , \39821 , \39822 );
xor \U$39446 ( \39824 , \39553 , \39557 );
xor \U$39447 ( \39825 , \39824 , \39562 );
xor \U$39448 ( \39826 , \39589 , \39593 );
xor \U$39449 ( \39827 , \39826 , \39598 );
and \U$39450 ( \39828 , \39825 , \39827 );
xor \U$39451 ( \39829 , \39570 , \39574 );
xor \U$39452 ( \39830 , \39829 , \39579 );
and \U$39453 ( \39831 , \39827 , \39830 );
and \U$39454 ( \39832 , \39825 , \39830 );
or \U$39455 ( \39833 , \39828 , \39831 , \39832 );
xor \U$39456 ( \39834 , \39640 , \39642 );
xor \U$39457 ( \39835 , \39834 , \39645 );
and \U$39458 ( \39836 , \39833 , \39835 );
xor \U$39459 ( \39837 , \39664 , \39666 );
xor \U$39460 ( \39838 , \39837 , \39669 );
and \U$39461 ( \39839 , \39835 , \39838 );
and \U$39462 ( \39840 , \39833 , \39838 );
or \U$39463 ( \39841 , \39836 , \39839 , \39840 );
and \U$39464 ( \39842 , \39823 , \39841 );
xor \U$39465 ( \39843 , \39549 , \39565 );
xor \U$39466 ( \39844 , \39843 , \39582 );
xor \U$39467 ( \39845 , \39601 , \39617 );
xor \U$39468 ( \39846 , \39845 , \39634 );
and \U$39469 ( \39847 , \39844 , \39846 );
and \U$39470 ( \39848 , \39841 , \39847 );
and \U$39471 ( \39849 , \39823 , \39847 );
or \U$39472 ( \39850 , \39842 , \39848 , \39849 );
xor \U$39473 ( \39851 , \39585 , \39637 );
xor \U$39474 ( \39852 , \39851 , \39648 );
xor \U$39475 ( \39853 , \39653 , \39655 );
xor \U$39476 ( \39854 , \39853 , \39658 );
and \U$39477 ( \39855 , \39852 , \39854 );
xor \U$39478 ( \39856 , \39672 , \39674 );
xor \U$39479 ( \39857 , \39856 , \39676 );
and \U$39480 ( \39858 , \39854 , \39857 );
and \U$39481 ( \39859 , \39852 , \39857 );
or \U$39482 ( \39860 , \39855 , \39858 , \39859 );
and \U$39483 ( \39861 , \39850 , \39860 );
xor \U$39484 ( \39862 , \39398 , \39450 );
xor \U$39485 ( \39863 , \39862 , \39463 );
and \U$39486 ( \39864 , \39860 , \39863 );
and \U$39487 ( \39865 , \39850 , \39863 );
or \U$39488 ( \39866 , \39861 , \39864 , \39865 );
xor \U$39489 ( \39867 , \39651 , \39661 );
xor \U$39490 ( \39868 , \39867 , \39679 );
xor \U$39491 ( \39869 , \39684 , \39686 );
xor \U$39492 ( \39870 , \39869 , \39689 );
and \U$39493 ( \39871 , \39868 , \39870 );
and \U$39494 ( \39872 , \39866 , \39871 );
xor \U$39495 ( \39873 , \39466 , \39487 );
xor \U$39496 ( \39874 , \39873 , \39498 );
and \U$39497 ( \39875 , \39871 , \39874 );
and \U$39498 ( \39876 , \39866 , \39874 );
or \U$39499 ( \39877 , \39872 , \39875 , \39876 );
xor \U$39500 ( \39878 , \39698 , \39700 );
xor \U$39501 ( \39879 , \39878 , \39703 );
and \U$39502 ( \39880 , \39877 , \39879 );
and \U$39503 ( \39881 , \39712 , \39880 );
xor \U$39504 ( \39882 , \39712 , \39880 );
xor \U$39505 ( \39883 , \39877 , \39879 );
xor \U$39506 ( \39884 , \39866 , \39871 );
xor \U$39507 ( \39885 , \39884 , \39874 );
xor \U$39508 ( \39886 , \39682 , \39692 );
xor \U$39509 ( \39887 , \39886 , \39695 );
and \U$39510 ( \39888 , \39885 , \39887 );
and \U$39511 ( \39889 , \39883 , \39888 );
xor \U$39512 ( \39890 , \39883 , \39888 );
xor \U$39513 ( \39891 , \39885 , \39887 );
and \U$39514 ( \39892 , \29710 , \26143 );
and \U$39515 ( \39893 , \29464 , \26141 );
nor \U$39516 ( \39894 , \39892 , \39893 );
xnor \U$39517 ( \39895 , \39894 , \25911 );
and \U$39518 ( \39896 , \30034 , \25692 );
and \U$39519 ( \39897 , \29715 , \25690 );
nor \U$39520 ( \39898 , \39896 , \39897 );
xnor \U$39521 ( \39899 , \39898 , \25549 );
and \U$39522 ( \39900 , \39895 , \39899 );
and \U$39523 ( \39901 , \30887 , \25369 );
and \U$39524 ( \39902 , \30318 , \25367 );
nor \U$39525 ( \39903 , \39901 , \39902 );
xnor \U$39526 ( \39904 , \39903 , \25123 );
and \U$39527 ( \39905 , \39899 , \39904 );
and \U$39528 ( \39906 , \39895 , \39904 );
or \U$39529 ( \39907 , \39900 , \39905 , \39906 );
and \U$39530 ( \39908 , \31498 , \24974 );
and \U$39531 ( \39909 , \30895 , \24972 );
nor \U$39532 ( \39910 , \39908 , \39909 );
xnor \U$39533 ( \39911 , \39910 , \24787 );
and \U$39534 ( \39912 , \31684 , \24661 );
and \U$39535 ( \39913 , \31503 , \24659 );
nor \U$39536 ( \39914 , \39912 , \39913 );
xnor \U$39537 ( \39915 , \39914 , \24456 );
and \U$39538 ( \39916 , \39911 , \39915 );
nand \U$39539 ( \39917 , \32304 , \24253 );
xnor \U$39540 ( \39918 , \39917 , \24106 );
and \U$39541 ( \39919 , \39915 , \39918 );
and \U$39542 ( \39920 , \39911 , \39918 );
or \U$39543 ( \39921 , \39916 , \39919 , \39920 );
and \U$39544 ( \39922 , \39907 , \39921 );
and \U$39545 ( \39923 , \27837 , \27572 );
and \U$39546 ( \39924 , \27494 , \27570 );
nor \U$39547 ( \39925 , \39923 , \39924 );
xnor \U$39548 ( \39926 , \39925 , \27232 );
and \U$39549 ( \39927 , \28342 , \26983 );
and \U$39550 ( \39928 , \28039 , \26981 );
nor \U$39551 ( \39929 , \39927 , \39928 );
xnor \U$39552 ( \39930 , \39929 , \26742 );
and \U$39553 ( \39931 , \39926 , \39930 );
and \U$39554 ( \39932 , \29040 , \26517 );
and \U$39555 ( \39933 , \28514 , \26515 );
nor \U$39556 ( \39934 , \39932 , \39933 );
xnor \U$39557 ( \39935 , \39934 , \26329 );
and \U$39558 ( \39936 , \39930 , \39935 );
and \U$39559 ( \39937 , \39926 , \39935 );
or \U$39560 ( \39938 , \39931 , \39936 , \39937 );
and \U$39561 ( \39939 , \39921 , \39938 );
and \U$39562 ( \39940 , \39907 , \39938 );
or \U$39563 ( \39941 , \39922 , \39939 , \39940 );
and \U$39564 ( \39942 , \26585 , \29104 );
and \U$39565 ( \39943 , \26116 , \29102 );
nor \U$39566 ( \39944 , \39942 , \39943 );
xnor \U$39567 ( \39945 , \39944 , \28855 );
and \U$39568 ( \39946 , \26854 , \28575 );
and \U$39569 ( \39947 , \26590 , \28573 );
nor \U$39570 ( \39948 , \39946 , \39947 );
xnor \U$39571 ( \39949 , \39948 , \28315 );
and \U$39572 ( \39950 , \39945 , \39949 );
and \U$39573 ( \39951 , \27485 , \28081 );
and \U$39574 ( \39952 , \27113 , \28079 );
nor \U$39575 ( \39953 , \39951 , \39952 );
xnor \U$39576 ( \39954 , \39953 , \27766 );
and \U$39577 ( \39955 , \39949 , \39954 );
and \U$39578 ( \39956 , \39945 , \39954 );
or \U$39579 ( \39957 , \39950 , \39955 , \39956 );
and \U$39580 ( \39958 , \24482 , \32151 );
and \U$39581 ( \39959 , \24344 , \32148 );
nor \U$39582 ( \39960 , \39958 , \39959 );
xnor \U$39583 ( \39961 , \39960 , \31096 );
and \U$39584 ( \39962 , \25018 , \31338 );
and \U$39585 ( \39963 , \24601 , \31336 );
nor \U$39586 ( \39964 , \39962 , \39963 );
xnor \U$39587 ( \39965 , \39964 , \31099 );
and \U$39588 ( \39966 , \39961 , \39965 );
and \U$39589 ( \39967 , \39965 , \24106 );
and \U$39590 ( \39968 , \39961 , \24106 );
or \U$39591 ( \39969 , \39966 , \39967 , \39968 );
and \U$39592 ( \39970 , \39957 , \39969 );
and \U$39593 ( \39971 , \25348 , \30770 );
and \U$39594 ( \39972 , \25226 , \30768 );
nor \U$39595 ( \39973 , \39971 , \39972 );
xnor \U$39596 ( \39974 , \39973 , \30460 );
and \U$39597 ( \39975 , \25609 , \30233 );
and \U$39598 ( \39976 , \25353 , \30231 );
nor \U$39599 ( \39977 , \39975 , \39976 );
xnor \U$39600 ( \39978 , \39977 , \29862 );
and \U$39601 ( \39979 , \39974 , \39978 );
and \U$39602 ( \39980 , \26108 , \29671 );
and \U$39603 ( \39981 , \25806 , \29669 );
nor \U$39604 ( \39982 , \39980 , \39981 );
xnor \U$39605 ( \39983 , \39982 , \29353 );
and \U$39606 ( \39984 , \39978 , \39983 );
and \U$39607 ( \39985 , \39974 , \39983 );
or \U$39608 ( \39986 , \39979 , \39984 , \39985 );
and \U$39609 ( \39987 , \39969 , \39986 );
and \U$39610 ( \39988 , \39957 , \39986 );
or \U$39611 ( \39989 , \39970 , \39987 , \39988 );
and \U$39612 ( \39990 , \39941 , \39989 );
xor \U$39613 ( \39991 , \39768 , \39772 );
xor \U$39614 ( \39992 , \39991 , \39777 );
xor \U$39615 ( \39993 , \39784 , \39788 );
xor \U$39616 ( \39994 , \39993 , \39793 );
and \U$39617 ( \39995 , \39992 , \39994 );
xor \U$39618 ( \39996 , \39801 , \39805 );
and \U$39619 ( \39997 , \39994 , \39996 );
and \U$39620 ( \39998 , \39992 , \39996 );
or \U$39621 ( \39999 , \39995 , \39997 , \39998 );
and \U$39622 ( \40000 , \39989 , \39999 );
and \U$39623 ( \40001 , \39941 , \39999 );
or \U$39624 ( \40002 , \39990 , \40000 , \40001 );
xor \U$39625 ( \40003 , \39716 , \39720 );
xor \U$39626 ( \40004 , \40003 , \39725 );
xor \U$39627 ( \40005 , \39732 , \39736 );
xor \U$39628 ( \40006 , \40005 , \39741 );
and \U$39629 ( \40007 , \40004 , \40006 );
xor \U$39630 ( \40008 , \39749 , \39753 );
xor \U$39631 ( \40009 , \40008 , \39758 );
and \U$39632 ( \40010 , \40006 , \40009 );
and \U$39633 ( \40011 , \40004 , \40009 );
or \U$39634 ( \40012 , \40007 , \40010 , \40011 );
xor \U$39635 ( \40013 , \39541 , \39545 );
xor \U$39636 ( \40014 , \40013 , \23791 );
and \U$39637 ( \40015 , \40012 , \40014 );
xor \U$39638 ( \40016 , \39825 , \39827 );
xor \U$39639 ( \40017 , \40016 , \39830 );
and \U$39640 ( \40018 , \40014 , \40017 );
and \U$39641 ( \40019 , \40012 , \40017 );
or \U$39642 ( \40020 , \40015 , \40018 , \40019 );
and \U$39643 ( \40021 , \40002 , \40020 );
xor \U$39644 ( \40022 , \39728 , \39744 );
xor \U$39645 ( \40023 , \40022 , \39761 );
xor \U$39646 ( \40024 , \39780 , \39796 );
xor \U$39647 ( \40025 , \40024 , \39806 );
and \U$39648 ( \40026 , \40023 , \40025 );
xor \U$39649 ( \40027 , \39812 , \39814 );
xor \U$39650 ( \40028 , \40027 , \39817 );
and \U$39651 ( \40029 , \40025 , \40028 );
and \U$39652 ( \40030 , \40023 , \40028 );
or \U$39653 ( \40031 , \40026 , \40029 , \40030 );
and \U$39654 ( \40032 , \40020 , \40031 );
and \U$39655 ( \40033 , \40002 , \40031 );
or \U$39656 ( \40034 , \40021 , \40032 , \40033 );
xor \U$39657 ( \40035 , \39764 , \39809 );
xor \U$39658 ( \40036 , \40035 , \39820 );
xor \U$39659 ( \40037 , \39833 , \39835 );
xor \U$39660 ( \40038 , \40037 , \39838 );
and \U$39661 ( \40039 , \40036 , \40038 );
xor \U$39662 ( \40040 , \39844 , \39846 );
and \U$39663 ( \40041 , \40038 , \40040 );
and \U$39664 ( \40042 , \40036 , \40040 );
or \U$39665 ( \40043 , \40039 , \40041 , \40042 );
and \U$39666 ( \40044 , \40034 , \40043 );
xor \U$39667 ( \40045 , \39852 , \39854 );
xor \U$39668 ( \40046 , \40045 , \39857 );
and \U$39669 ( \40047 , \40043 , \40046 );
and \U$39670 ( \40048 , \40034 , \40046 );
or \U$39671 ( \40049 , \40044 , \40047 , \40048 );
xor \U$39672 ( \40050 , \39850 , \39860 );
xor \U$39673 ( \40051 , \40050 , \39863 );
and \U$39674 ( \40052 , \40049 , \40051 );
xor \U$39675 ( \40053 , \39868 , \39870 );
and \U$39676 ( \40054 , \40051 , \40053 );
and \U$39677 ( \40055 , \40049 , \40053 );
or \U$39678 ( \40056 , \40052 , \40054 , \40055 );
and \U$39679 ( \40057 , \39891 , \40056 );
xor \U$39680 ( \40058 , \39891 , \40056 );
xor \U$39681 ( \40059 , \40049 , \40051 );
xor \U$39682 ( \40060 , \40059 , \40053 );
and \U$39683 ( \40061 , \25806 , \30233 );
and \U$39684 ( \40062 , \25609 , \30231 );
nor \U$39685 ( \40063 , \40061 , \40062 );
xnor \U$39686 ( \40064 , \40063 , \29862 );
and \U$39687 ( \40065 , \26116 , \29671 );
and \U$39688 ( \40066 , \26108 , \29669 );
nor \U$39689 ( \40067 , \40065 , \40066 );
xnor \U$39690 ( \40068 , \40067 , \29353 );
and \U$39691 ( \40069 , \40064 , \40068 );
and \U$39692 ( \40070 , \26590 , \29104 );
and \U$39693 ( \40071 , \26585 , \29102 );
nor \U$39694 ( \40072 , \40070 , \40071 );
xnor \U$39695 ( \40073 , \40072 , \28855 );
and \U$39696 ( \40074 , \40068 , \40073 );
and \U$39697 ( \40075 , \40064 , \40073 );
or \U$39698 ( \40076 , \40069 , \40074 , \40075 );
and \U$39699 ( \40077 , \24601 , \32151 );
and \U$39700 ( \40078 , \24482 , \32148 );
nor \U$39701 ( \40079 , \40077 , \40078 );
xnor \U$39702 ( \40080 , \40079 , \31096 );
and \U$39703 ( \40081 , \25226 , \31338 );
and \U$39704 ( \40082 , \25018 , \31336 );
nor \U$39705 ( \40083 , \40081 , \40082 );
xnor \U$39706 ( \40084 , \40083 , \31099 );
and \U$39707 ( \40085 , \40080 , \40084 );
and \U$39708 ( \40086 , \25353 , \30770 );
and \U$39709 ( \40087 , \25348 , \30768 );
nor \U$39710 ( \40088 , \40086 , \40087 );
xnor \U$39711 ( \40089 , \40088 , \30460 );
and \U$39712 ( \40090 , \40084 , \40089 );
and \U$39713 ( \40091 , \40080 , \40089 );
or \U$39714 ( \40092 , \40085 , \40090 , \40091 );
and \U$39715 ( \40093 , \40076 , \40092 );
and \U$39716 ( \40094 , \27113 , \28575 );
and \U$39717 ( \40095 , \26854 , \28573 );
nor \U$39718 ( \40096 , \40094 , \40095 );
xnor \U$39719 ( \40097 , \40096 , \28315 );
and \U$39720 ( \40098 , \27494 , \28081 );
and \U$39721 ( \40099 , \27485 , \28079 );
nor \U$39722 ( \40100 , \40098 , \40099 );
xnor \U$39723 ( \40101 , \40100 , \27766 );
and \U$39724 ( \40102 , \40097 , \40101 );
and \U$39725 ( \40103 , \28039 , \27572 );
and \U$39726 ( \40104 , \27837 , \27570 );
nor \U$39727 ( \40105 , \40103 , \40104 );
xnor \U$39728 ( \40106 , \40105 , \27232 );
and \U$39729 ( \40107 , \40101 , \40106 );
and \U$39730 ( \40108 , \40097 , \40106 );
or \U$39731 ( \40109 , \40102 , \40107 , \40108 );
and \U$39732 ( \40110 , \40092 , \40109 );
and \U$39733 ( \40111 , \40076 , \40109 );
or \U$39734 ( \40112 , \40093 , \40110 , \40111 );
xor \U$39735 ( \40113 , \39895 , \39899 );
xor \U$39736 ( \40114 , \40113 , \39904 );
xor \U$39737 ( \40115 , \39945 , \39949 );
xor \U$39738 ( \40116 , \40115 , \39954 );
and \U$39739 ( \40117 , \40114 , \40116 );
xor \U$39740 ( \40118 , \39926 , \39930 );
xor \U$39741 ( \40119 , \40118 , \39935 );
and \U$39742 ( \40120 , \40116 , \40119 );
and \U$39743 ( \40121 , \40114 , \40119 );
or \U$39744 ( \40122 , \40117 , \40120 , \40121 );
and \U$39745 ( \40123 , \40112 , \40122 );
and \U$39746 ( \40124 , \28514 , \26983 );
and \U$39747 ( \40125 , \28342 , \26981 );
nor \U$39748 ( \40126 , \40124 , \40125 );
xnor \U$39749 ( \40127 , \40126 , \26742 );
and \U$39750 ( \40128 , \29464 , \26517 );
and \U$39751 ( \40129 , \29040 , \26515 );
nor \U$39752 ( \40130 , \40128 , \40129 );
xnor \U$39753 ( \40131 , \40130 , \26329 );
and \U$39754 ( \40132 , \40127 , \40131 );
and \U$39755 ( \40133 , \29715 , \26143 );
and \U$39756 ( \40134 , \29710 , \26141 );
nor \U$39757 ( \40135 , \40133 , \40134 );
xnor \U$39758 ( \40136 , \40135 , \25911 );
and \U$39759 ( \40137 , \40131 , \40136 );
and \U$39760 ( \40138 , \40127 , \40136 );
or \U$39761 ( \40139 , \40132 , \40137 , \40138 );
and \U$39762 ( \40140 , \30318 , \25692 );
and \U$39763 ( \40141 , \30034 , \25690 );
nor \U$39764 ( \40142 , \40140 , \40141 );
xnor \U$39765 ( \40143 , \40142 , \25549 );
and \U$39766 ( \40144 , \30895 , \25369 );
and \U$39767 ( \40145 , \30887 , \25367 );
nor \U$39768 ( \40146 , \40144 , \40145 );
xnor \U$39769 ( \40147 , \40146 , \25123 );
and \U$39770 ( \40148 , \40143 , \40147 );
and \U$39771 ( \40149 , \31503 , \24974 );
and \U$39772 ( \40150 , \31498 , \24972 );
nor \U$39773 ( \40151 , \40149 , \40150 );
xnor \U$39774 ( \40152 , \40151 , \24787 );
and \U$39775 ( \40153 , \40147 , \40152 );
and \U$39776 ( \40154 , \40143 , \40152 );
or \U$39777 ( \40155 , \40148 , \40153 , \40154 );
and \U$39778 ( \40156 , \40139 , \40155 );
xor \U$39779 ( \40157 , \39911 , \39915 );
xor \U$39780 ( \40158 , \40157 , \39918 );
and \U$39781 ( \40159 , \40155 , \40158 );
and \U$39782 ( \40160 , \40139 , \40158 );
or \U$39783 ( \40161 , \40156 , \40159 , \40160 );
and \U$39784 ( \40162 , \40122 , \40161 );
and \U$39785 ( \40163 , \40112 , \40161 );
or \U$39786 ( \40164 , \40123 , \40162 , \40163 );
xor \U$39787 ( \40165 , \39907 , \39921 );
xor \U$39788 ( \40166 , \40165 , \39938 );
xor \U$39789 ( \40167 , \40004 , \40006 );
xor \U$39790 ( \40168 , \40167 , \40009 );
and \U$39791 ( \40169 , \40166 , \40168 );
xor \U$39792 ( \40170 , \39992 , \39994 );
xor \U$39793 ( \40171 , \40170 , \39996 );
and \U$39794 ( \40172 , \40168 , \40171 );
and \U$39795 ( \40173 , \40166 , \40171 );
or \U$39796 ( \40174 , \40169 , \40172 , \40173 );
and \U$39797 ( \40175 , \40164 , \40174 );
xor \U$39798 ( \40176 , \40023 , \40025 );
xor \U$39799 ( \40177 , \40176 , \40028 );
and \U$39800 ( \40178 , \40174 , \40177 );
and \U$39801 ( \40179 , \40164 , \40177 );
or \U$39802 ( \40180 , \40175 , \40178 , \40179 );
xor \U$39803 ( \40181 , \40002 , \40020 );
xor \U$39804 ( \40182 , \40181 , \40031 );
and \U$39805 ( \40183 , \40180 , \40182 );
xor \U$39806 ( \40184 , \40036 , \40038 );
xor \U$39807 ( \40185 , \40184 , \40040 );
and \U$39808 ( \40186 , \40182 , \40185 );
and \U$39809 ( \40187 , \40180 , \40185 );
or \U$39810 ( \40188 , \40183 , \40186 , \40187 );
xor \U$39811 ( \40189 , \39823 , \39841 );
xor \U$39812 ( \40190 , \40189 , \39847 );
and \U$39813 ( \40191 , \40188 , \40190 );
xor \U$39814 ( \40192 , \40034 , \40043 );
xor \U$39815 ( \40193 , \40192 , \40046 );
and \U$39816 ( \40194 , \40190 , \40193 );
and \U$39817 ( \40195 , \40188 , \40193 );
or \U$39818 ( \40196 , \40191 , \40194 , \40195 );
and \U$39819 ( \40197 , \40060 , \40196 );
xor \U$39820 ( \40198 , \40060 , \40196 );
xor \U$39821 ( \40199 , \40188 , \40190 );
xor \U$39822 ( \40200 , \40199 , \40193 );
and \U$39823 ( \40201 , \25609 , \30770 );
and \U$39824 ( \40202 , \25353 , \30768 );
nor \U$39825 ( \40203 , \40201 , \40202 );
xnor \U$39826 ( \40204 , \40203 , \30460 );
and \U$39827 ( \40205 , \26108 , \30233 );
and \U$39828 ( \40206 , \25806 , \30231 );
nor \U$39829 ( \40207 , \40205 , \40206 );
xnor \U$39830 ( \40208 , \40207 , \29862 );
and \U$39831 ( \40209 , \40204 , \40208 );
and \U$39832 ( \40210 , \26585 , \29671 );
and \U$39833 ( \40211 , \26116 , \29669 );
nor \U$39834 ( \40212 , \40210 , \40211 );
xnor \U$39835 ( \40213 , \40212 , \29353 );
and \U$39836 ( \40214 , \40208 , \40213 );
and \U$39837 ( \40215 , \40204 , \40213 );
or \U$39838 ( \40216 , \40209 , \40214 , \40215 );
and \U$39839 ( \40217 , \26854 , \29104 );
and \U$39840 ( \40218 , \26590 , \29102 );
nor \U$39841 ( \40219 , \40217 , \40218 );
xnor \U$39842 ( \40220 , \40219 , \28855 );
and \U$39843 ( \40221 , \27485 , \28575 );
and \U$39844 ( \40222 , \27113 , \28573 );
nor \U$39845 ( \40223 , \40221 , \40222 );
xnor \U$39846 ( \40224 , \40223 , \28315 );
and \U$39847 ( \40225 , \40220 , \40224 );
and \U$39848 ( \40226 , \27837 , \28081 );
and \U$39849 ( \40227 , \27494 , \28079 );
nor \U$39850 ( \40228 , \40226 , \40227 );
xnor \U$39851 ( \40229 , \40228 , \27766 );
and \U$39852 ( \40230 , \40224 , \40229 );
and \U$39853 ( \40231 , \40220 , \40229 );
or \U$39854 ( \40232 , \40225 , \40230 , \40231 );
and \U$39855 ( \40233 , \40216 , \40232 );
and \U$39856 ( \40234 , \25018 , \32151 );
and \U$39857 ( \40235 , \24601 , \32148 );
nor \U$39858 ( \40236 , \40234 , \40235 );
xnor \U$39859 ( \40237 , \40236 , \31096 );
and \U$39860 ( \40238 , \25348 , \31338 );
and \U$39861 ( \40239 , \25226 , \31336 );
nor \U$39862 ( \40240 , \40238 , \40239 );
xnor \U$39863 ( \40241 , \40240 , \31099 );
and \U$39864 ( \40242 , \40237 , \40241 );
and \U$39865 ( \40243 , \40241 , \24456 );
and \U$39866 ( \40244 , \40237 , \24456 );
or \U$39867 ( \40245 , \40242 , \40243 , \40244 );
and \U$39868 ( \40246 , \40232 , \40245 );
and \U$39869 ( \40247 , \40216 , \40245 );
or \U$39870 ( \40248 , \40233 , \40246 , \40247 );
and \U$39871 ( \40249 , \30034 , \26143 );
and \U$39872 ( \40250 , \29715 , \26141 );
nor \U$39873 ( \40251 , \40249 , \40250 );
xnor \U$39874 ( \40252 , \40251 , \25911 );
and \U$39875 ( \40253 , \30887 , \25692 );
and \U$39876 ( \40254 , \30318 , \25690 );
nor \U$39877 ( \40255 , \40253 , \40254 );
xnor \U$39878 ( \40256 , \40255 , \25549 );
and \U$39879 ( \40257 , \40252 , \40256 );
and \U$39880 ( \40258 , \31498 , \25369 );
and \U$39881 ( \40259 , \30895 , \25367 );
nor \U$39882 ( \40260 , \40258 , \40259 );
xnor \U$39883 ( \40261 , \40260 , \25123 );
and \U$39884 ( \40262 , \40256 , \40261 );
and \U$39885 ( \40263 , \40252 , \40261 );
or \U$39886 ( \40264 , \40257 , \40262 , \40263 );
and \U$39887 ( \40265 , \28342 , \27572 );
and \U$39888 ( \40266 , \28039 , \27570 );
nor \U$39889 ( \40267 , \40265 , \40266 );
xnor \U$39890 ( \40268 , \40267 , \27232 );
and \U$39891 ( \40269 , \29040 , \26983 );
and \U$39892 ( \40270 , \28514 , \26981 );
nor \U$39893 ( \40271 , \40269 , \40270 );
xnor \U$39894 ( \40272 , \40271 , \26742 );
and \U$39895 ( \40273 , \40268 , \40272 );
and \U$39896 ( \40274 , \29710 , \26517 );
and \U$39897 ( \40275 , \29464 , \26515 );
nor \U$39898 ( \40276 , \40274 , \40275 );
xnor \U$39899 ( \40277 , \40276 , \26329 );
and \U$39900 ( \40278 , \40272 , \40277 );
and \U$39901 ( \40279 , \40268 , \40277 );
or \U$39902 ( \40280 , \40273 , \40278 , \40279 );
and \U$39903 ( \40281 , \40264 , \40280 );
and \U$39904 ( \40282 , \32304 , \24661 );
and \U$39905 ( \40283 , \31684 , \24659 );
nor \U$39906 ( \40284 , \40282 , \40283 );
xnor \U$39907 ( \40285 , \40284 , \24456 );
and \U$39908 ( \40286 , \40280 , \40285 );
and \U$39909 ( \40287 , \40264 , \40285 );
or \U$39910 ( \40288 , \40281 , \40286 , \40287 );
and \U$39911 ( \40289 , \40248 , \40288 );
xor \U$39912 ( \40290 , \40127 , \40131 );
xor \U$39913 ( \40291 , \40290 , \40136 );
xor \U$39914 ( \40292 , \40143 , \40147 );
xor \U$39915 ( \40293 , \40292 , \40152 );
and \U$39916 ( \40294 , \40291 , \40293 );
xor \U$39917 ( \40295 , \40097 , \40101 );
xor \U$39918 ( \40296 , \40295 , \40106 );
and \U$39919 ( \40297 , \40293 , \40296 );
and \U$39920 ( \40298 , \40291 , \40296 );
or \U$39921 ( \40299 , \40294 , \40297 , \40298 );
and \U$39922 ( \40300 , \40288 , \40299 );
and \U$39923 ( \40301 , \40248 , \40299 );
or \U$39924 ( \40302 , \40289 , \40300 , \40301 );
xor \U$39925 ( \40303 , \39961 , \39965 );
xor \U$39926 ( \40304 , \40303 , \24106 );
xor \U$39927 ( \40305 , \39974 , \39978 );
xor \U$39928 ( \40306 , \40305 , \39983 );
and \U$39929 ( \40307 , \40304 , \40306 );
xor \U$39930 ( \40308 , \40114 , \40116 );
xor \U$39931 ( \40309 , \40308 , \40119 );
and \U$39932 ( \40310 , \40306 , \40309 );
and \U$39933 ( \40311 , \40304 , \40309 );
or \U$39934 ( \40312 , \40307 , \40310 , \40311 );
and \U$39935 ( \40313 , \40302 , \40312 );
xor \U$39936 ( \40314 , \40076 , \40092 );
xor \U$39937 ( \40315 , \40314 , \40109 );
xor \U$39938 ( \40316 , \40139 , \40155 );
xor \U$39939 ( \40317 , \40316 , \40158 );
and \U$39940 ( \40318 , \40315 , \40317 );
and \U$39941 ( \40319 , \40312 , \40318 );
and \U$39942 ( \40320 , \40302 , \40318 );
or \U$39943 ( \40321 , \40313 , \40319 , \40320 );
xor \U$39944 ( \40322 , \39957 , \39969 );
xor \U$39945 ( \40323 , \40322 , \39986 );
xor \U$39946 ( \40324 , \40112 , \40122 );
xor \U$39947 ( \40325 , \40324 , \40161 );
and \U$39948 ( \40326 , \40323 , \40325 );
xor \U$39949 ( \40327 , \40166 , \40168 );
xor \U$39950 ( \40328 , \40327 , \40171 );
and \U$39951 ( \40329 , \40325 , \40328 );
and \U$39952 ( \40330 , \40323 , \40328 );
or \U$39953 ( \40331 , \40326 , \40329 , \40330 );
and \U$39954 ( \40332 , \40321 , \40331 );
xor \U$39955 ( \40333 , \40012 , \40014 );
xor \U$39956 ( \40334 , \40333 , \40017 );
and \U$39957 ( \40335 , \40331 , \40334 );
and \U$39958 ( \40336 , \40321 , \40334 );
or \U$39959 ( \40337 , \40332 , \40335 , \40336 );
xor \U$39960 ( \40338 , \39941 , \39989 );
xor \U$39961 ( \40339 , \40338 , \39999 );
xor \U$39962 ( \40340 , \40164 , \40174 );
xor \U$39963 ( \40341 , \40340 , \40177 );
and \U$39964 ( \40342 , \40339 , \40341 );
and \U$39965 ( \40343 , \40337 , \40342 );
xor \U$39966 ( \40344 , \40180 , \40182 );
xor \U$39967 ( \40345 , \40344 , \40185 );
and \U$39968 ( \40346 , \40342 , \40345 );
and \U$39969 ( \40347 , \40337 , \40345 );
or \U$39970 ( \40348 , \40343 , \40346 , \40347 );
and \U$39971 ( \40349 , \40200 , \40348 );
xor \U$39972 ( \40350 , \40200 , \40348 );
xor \U$39973 ( \40351 , \40337 , \40342 );
xor \U$39974 ( \40352 , \40351 , \40345 );
and \U$39975 ( \40353 , \27494 , \28575 );
and \U$39976 ( \40354 , \27485 , \28573 );
nor \U$39977 ( \40355 , \40353 , \40354 );
xnor \U$39978 ( \40356 , \40355 , \28315 );
and \U$39979 ( \40357 , \28039 , \28081 );
and \U$39980 ( \40358 , \27837 , \28079 );
nor \U$39981 ( \40359 , \40357 , \40358 );
xnor \U$39982 ( \40360 , \40359 , \27766 );
and \U$39983 ( \40361 , \40356 , \40360 );
and \U$39984 ( \40362 , \28514 , \27572 );
and \U$39985 ( \40363 , \28342 , \27570 );
nor \U$39986 ( \40364 , \40362 , \40363 );
xnor \U$39987 ( \40365 , \40364 , \27232 );
and \U$39988 ( \40366 , \40360 , \40365 );
and \U$39989 ( \40367 , \40356 , \40365 );
or \U$39990 ( \40368 , \40361 , \40366 , \40367 );
and \U$39991 ( \40369 , \26116 , \30233 );
and \U$39992 ( \40370 , \26108 , \30231 );
nor \U$39993 ( \40371 , \40369 , \40370 );
xnor \U$39994 ( \40372 , \40371 , \29862 );
and \U$39995 ( \40373 , \26590 , \29671 );
and \U$39996 ( \40374 , \26585 , \29669 );
nor \U$39997 ( \40375 , \40373 , \40374 );
xnor \U$39998 ( \40376 , \40375 , \29353 );
and \U$39999 ( \40377 , \40372 , \40376 );
and \U$40000 ( \40378 , \27113 , \29104 );
and \U$40001 ( \40379 , \26854 , \29102 );
nor \U$40002 ( \40380 , \40378 , \40379 );
xnor \U$40003 ( \40381 , \40380 , \28855 );
and \U$40004 ( \40382 , \40376 , \40381 );
and \U$40005 ( \40383 , \40372 , \40381 );
or \U$40006 ( \40384 , \40377 , \40382 , \40383 );
and \U$40007 ( \40385 , \40368 , \40384 );
and \U$40008 ( \40386 , \25226 , \32151 );
and \U$40009 ( \40387 , \25018 , \32148 );
nor \U$40010 ( \40388 , \40386 , \40387 );
xnor \U$40011 ( \40389 , \40388 , \31096 );
and \U$40012 ( \40390 , \25353 , \31338 );
and \U$40013 ( \40391 , \25348 , \31336 );
nor \U$40014 ( \40392 , \40390 , \40391 );
xnor \U$40015 ( \40393 , \40392 , \31099 );
and \U$40016 ( \40394 , \40389 , \40393 );
and \U$40017 ( \40395 , \25806 , \30770 );
and \U$40018 ( \40396 , \25609 , \30768 );
nor \U$40019 ( \40397 , \40395 , \40396 );
xnor \U$40020 ( \40398 , \40397 , \30460 );
and \U$40021 ( \40399 , \40393 , \40398 );
and \U$40022 ( \40400 , \40389 , \40398 );
or \U$40023 ( \40401 , \40394 , \40399 , \40400 );
and \U$40024 ( \40402 , \40384 , \40401 );
and \U$40025 ( \40403 , \40368 , \40401 );
or \U$40026 ( \40404 , \40385 , \40402 , \40403 );
and \U$40027 ( \40405 , \30895 , \25692 );
and \U$40028 ( \40406 , \30887 , \25690 );
nor \U$40029 ( \40407 , \40405 , \40406 );
xnor \U$40030 ( \40408 , \40407 , \25549 );
and \U$40031 ( \40409 , \31503 , \25369 );
and \U$40032 ( \40410 , \31498 , \25367 );
nor \U$40033 ( \40411 , \40409 , \40410 );
xnor \U$40034 ( \40412 , \40411 , \25123 );
and \U$40035 ( \40413 , \40408 , \40412 );
and \U$40036 ( \40414 , \32304 , \24974 );
and \U$40037 ( \40415 , \31684 , \24972 );
nor \U$40038 ( \40416 , \40414 , \40415 );
xnor \U$40039 ( \40417 , \40416 , \24787 );
and \U$40040 ( \40418 , \40412 , \40417 );
and \U$40041 ( \40419 , \40408 , \40417 );
or \U$40042 ( \40420 , \40413 , \40418 , \40419 );
and \U$40043 ( \40421 , \29464 , \26983 );
and \U$40044 ( \40422 , \29040 , \26981 );
nor \U$40045 ( \40423 , \40421 , \40422 );
xnor \U$40046 ( \40424 , \40423 , \26742 );
and \U$40047 ( \40425 , \29715 , \26517 );
and \U$40048 ( \40426 , \29710 , \26515 );
nor \U$40049 ( \40427 , \40425 , \40426 );
xnor \U$40050 ( \40428 , \40427 , \26329 );
and \U$40051 ( \40429 , \40424 , \40428 );
and \U$40052 ( \40430 , \30318 , \26143 );
and \U$40053 ( \40431 , \30034 , \26141 );
nor \U$40054 ( \40432 , \40430 , \40431 );
xnor \U$40055 ( \40433 , \40432 , \25911 );
and \U$40056 ( \40434 , \40428 , \40433 );
and \U$40057 ( \40435 , \40424 , \40433 );
or \U$40058 ( \40436 , \40429 , \40434 , \40435 );
and \U$40059 ( \40437 , \40420 , \40436 );
and \U$40060 ( \40438 , \31684 , \24974 );
and \U$40061 ( \40439 , \31503 , \24972 );
nor \U$40062 ( \40440 , \40438 , \40439 );
xnor \U$40063 ( \40441 , \40440 , \24787 );
and \U$40064 ( \40442 , \40436 , \40441 );
and \U$40065 ( \40443 , \40420 , \40441 );
or \U$40066 ( \40444 , \40437 , \40442 , \40443 );
and \U$40067 ( \40445 , \40404 , \40444 );
nand \U$40068 ( \40446 , \32304 , \24659 );
xnor \U$40069 ( \40447 , \40446 , \24456 );
xor \U$40070 ( \40448 , \40252 , \40256 );
xor \U$40071 ( \40449 , \40448 , \40261 );
and \U$40072 ( \40450 , \40447 , \40449 );
xor \U$40073 ( \40451 , \40268 , \40272 );
xor \U$40074 ( \40452 , \40451 , \40277 );
and \U$40075 ( \40453 , \40449 , \40452 );
and \U$40076 ( \40454 , \40447 , \40452 );
or \U$40077 ( \40455 , \40450 , \40453 , \40454 );
and \U$40078 ( \40456 , \40444 , \40455 );
and \U$40079 ( \40457 , \40404 , \40455 );
or \U$40080 ( \40458 , \40445 , \40456 , \40457 );
xor \U$40081 ( \40459 , \40204 , \40208 );
xor \U$40082 ( \40460 , \40459 , \40213 );
xor \U$40083 ( \40461 , \40220 , \40224 );
xor \U$40084 ( \40462 , \40461 , \40229 );
and \U$40085 ( \40463 , \40460 , \40462 );
xor \U$40086 ( \40464 , \40237 , \40241 );
xor \U$40087 ( \40465 , \40464 , \24456 );
and \U$40088 ( \40466 , \40462 , \40465 );
and \U$40089 ( \40467 , \40460 , \40465 );
or \U$40090 ( \40468 , \40463 , \40466 , \40467 );
xor \U$40091 ( \40469 , \40064 , \40068 );
xor \U$40092 ( \40470 , \40469 , \40073 );
and \U$40093 ( \40471 , \40468 , \40470 );
xor \U$40094 ( \40472 , \40080 , \40084 );
xor \U$40095 ( \40473 , \40472 , \40089 );
and \U$40096 ( \40474 , \40470 , \40473 );
and \U$40097 ( \40475 , \40468 , \40473 );
or \U$40098 ( \40476 , \40471 , \40474 , \40475 );
and \U$40099 ( \40477 , \40458 , \40476 );
xor \U$40100 ( \40478 , \40216 , \40232 );
xor \U$40101 ( \40479 , \40478 , \40245 );
xor \U$40102 ( \40480 , \40264 , \40280 );
xor \U$40103 ( \40481 , \40480 , \40285 );
and \U$40104 ( \40482 , \40479 , \40481 );
xor \U$40105 ( \40483 , \40291 , \40293 );
xor \U$40106 ( \40484 , \40483 , \40296 );
and \U$40107 ( \40485 , \40481 , \40484 );
and \U$40108 ( \40486 , \40479 , \40484 );
or \U$40109 ( \40487 , \40482 , \40485 , \40486 );
and \U$40110 ( \40488 , \40476 , \40487 );
and \U$40111 ( \40489 , \40458 , \40487 );
or \U$40112 ( \40490 , \40477 , \40488 , \40489 );
xor \U$40113 ( \40491 , \40248 , \40288 );
xor \U$40114 ( \40492 , \40491 , \40299 );
xor \U$40115 ( \40493 , \40304 , \40306 );
xor \U$40116 ( \40494 , \40493 , \40309 );
and \U$40117 ( \40495 , \40492 , \40494 );
xor \U$40118 ( \40496 , \40315 , \40317 );
and \U$40119 ( \40497 , \40494 , \40496 );
and \U$40120 ( \40498 , \40492 , \40496 );
or \U$40121 ( \40499 , \40495 , \40497 , \40498 );
and \U$40122 ( \40500 , \40490 , \40499 );
xor \U$40123 ( \40501 , \40323 , \40325 );
xor \U$40124 ( \40502 , \40501 , \40328 );
and \U$40125 ( \40503 , \40499 , \40502 );
and \U$40126 ( \40504 , \40490 , \40502 );
or \U$40127 ( \40505 , \40500 , \40503 , \40504 );
xor \U$40128 ( \40506 , \40321 , \40331 );
xor \U$40129 ( \40507 , \40506 , \40334 );
and \U$40130 ( \40508 , \40505 , \40507 );
xor \U$40131 ( \40509 , \40339 , \40341 );
and \U$40132 ( \40510 , \40507 , \40509 );
and \U$40133 ( \40511 , \40505 , \40509 );
or \U$40134 ( \40512 , \40508 , \40510 , \40511 );
and \U$40135 ( \40513 , \40352 , \40512 );
xor \U$40136 ( \40514 , \40352 , \40512 );
xor \U$40137 ( \40515 , \40505 , \40507 );
xor \U$40138 ( \40516 , \40515 , \40509 );
and \U$40139 ( \40517 , \27485 , \29104 );
and \U$40140 ( \40518 , \27113 , \29102 );
nor \U$40141 ( \40519 , \40517 , \40518 );
xnor \U$40142 ( \40520 , \40519 , \28855 );
and \U$40143 ( \40521 , \27837 , \28575 );
and \U$40144 ( \40522 , \27494 , \28573 );
nor \U$40145 ( \40523 , \40521 , \40522 );
xnor \U$40146 ( \40524 , \40523 , \28315 );
and \U$40147 ( \40525 , \40520 , \40524 );
and \U$40148 ( \40526 , \28342 , \28081 );
and \U$40149 ( \40527 , \28039 , \28079 );
nor \U$40150 ( \40528 , \40526 , \40527 );
xnor \U$40151 ( \40529 , \40528 , \27766 );
and \U$40152 ( \40530 , \40524 , \40529 );
and \U$40153 ( \40531 , \40520 , \40529 );
or \U$40154 ( \40532 , \40525 , \40530 , \40531 );
and \U$40155 ( \40533 , \26108 , \30770 );
and \U$40156 ( \40534 , \25806 , \30768 );
nor \U$40157 ( \40535 , \40533 , \40534 );
xnor \U$40158 ( \40536 , \40535 , \30460 );
and \U$40159 ( \40537 , \26585 , \30233 );
and \U$40160 ( \40538 , \26116 , \30231 );
nor \U$40161 ( \40539 , \40537 , \40538 );
xnor \U$40162 ( \40540 , \40539 , \29862 );
and \U$40163 ( \40541 , \40536 , \40540 );
and \U$40164 ( \40542 , \26854 , \29671 );
and \U$40165 ( \40543 , \26590 , \29669 );
nor \U$40166 ( \40544 , \40542 , \40543 );
xnor \U$40167 ( \40545 , \40544 , \29353 );
and \U$40168 ( \40546 , \40540 , \40545 );
and \U$40169 ( \40547 , \40536 , \40545 );
or \U$40170 ( \40548 , \40541 , \40546 , \40547 );
and \U$40171 ( \40549 , \40532 , \40548 );
and \U$40172 ( \40550 , \25348 , \32151 );
and \U$40173 ( \40551 , \25226 , \32148 );
nor \U$40174 ( \40552 , \40550 , \40551 );
xnor \U$40175 ( \40553 , \40552 , \31096 );
and \U$40176 ( \40554 , \25609 , \31338 );
and \U$40177 ( \40555 , \25353 , \31336 );
nor \U$40178 ( \40556 , \40554 , \40555 );
xnor \U$40179 ( \40557 , \40556 , \31099 );
and \U$40180 ( \40558 , \40553 , \40557 );
and \U$40181 ( \40559 , \40557 , \24787 );
and \U$40182 ( \40560 , \40553 , \24787 );
or \U$40183 ( \40561 , \40558 , \40559 , \40560 );
and \U$40184 ( \40562 , \40548 , \40561 );
and \U$40185 ( \40563 , \40532 , \40561 );
or \U$40186 ( \40564 , \40549 , \40562 , \40563 );
and \U$40187 ( \40565 , \29040 , \27572 );
and \U$40188 ( \40566 , \28514 , \27570 );
nor \U$40189 ( \40567 , \40565 , \40566 );
xnor \U$40190 ( \40568 , \40567 , \27232 );
and \U$40191 ( \40569 , \29710 , \26983 );
and \U$40192 ( \40570 , \29464 , \26981 );
nor \U$40193 ( \40571 , \40569 , \40570 );
xnor \U$40194 ( \40572 , \40571 , \26742 );
and \U$40195 ( \40573 , \40568 , \40572 );
and \U$40196 ( \40574 , \30034 , \26517 );
and \U$40197 ( \40575 , \29715 , \26515 );
nor \U$40198 ( \40576 , \40574 , \40575 );
xnor \U$40199 ( \40577 , \40576 , \26329 );
and \U$40200 ( \40578 , \40572 , \40577 );
and \U$40201 ( \40579 , \40568 , \40577 );
or \U$40202 ( \40580 , \40573 , \40578 , \40579 );
and \U$40203 ( \40581 , \30887 , \26143 );
and \U$40204 ( \40582 , \30318 , \26141 );
nor \U$40205 ( \40583 , \40581 , \40582 );
xnor \U$40206 ( \40584 , \40583 , \25911 );
and \U$40207 ( \40585 , \31498 , \25692 );
and \U$40208 ( \40586 , \30895 , \25690 );
nor \U$40209 ( \40587 , \40585 , \40586 );
xnor \U$40210 ( \40588 , \40587 , \25549 );
and \U$40211 ( \40589 , \40584 , \40588 );
and \U$40212 ( \40590 , \31684 , \25369 );
and \U$40213 ( \40591 , \31503 , \25367 );
nor \U$40214 ( \40592 , \40590 , \40591 );
xnor \U$40215 ( \40593 , \40592 , \25123 );
and \U$40216 ( \40594 , \40588 , \40593 );
and \U$40217 ( \40595 , \40584 , \40593 );
or \U$40218 ( \40596 , \40589 , \40594 , \40595 );
and \U$40219 ( \40597 , \40580 , \40596 );
xor \U$40220 ( \40598 , \40408 , \40412 );
xor \U$40221 ( \40599 , \40598 , \40417 );
and \U$40222 ( \40600 , \40596 , \40599 );
and \U$40223 ( \40601 , \40580 , \40599 );
or \U$40224 ( \40602 , \40597 , \40600 , \40601 );
and \U$40225 ( \40603 , \40564 , \40602 );
xor \U$40226 ( \40604 , \40356 , \40360 );
xor \U$40227 ( \40605 , \40604 , \40365 );
xor \U$40228 ( \40606 , \40372 , \40376 );
xor \U$40229 ( \40607 , \40606 , \40381 );
and \U$40230 ( \40608 , \40605 , \40607 );
xor \U$40231 ( \40609 , \40424 , \40428 );
xor \U$40232 ( \40610 , \40609 , \40433 );
and \U$40233 ( \40611 , \40607 , \40610 );
and \U$40234 ( \40612 , \40605 , \40610 );
or \U$40235 ( \40613 , \40608 , \40611 , \40612 );
and \U$40236 ( \40614 , \40602 , \40613 );
and \U$40237 ( \40615 , \40564 , \40613 );
or \U$40238 ( \40616 , \40603 , \40614 , \40615 );
xor \U$40239 ( \40617 , \40420 , \40436 );
xor \U$40240 ( \40618 , \40617 , \40441 );
xor \U$40241 ( \40619 , \40460 , \40462 );
xor \U$40242 ( \40620 , \40619 , \40465 );
and \U$40243 ( \40621 , \40618 , \40620 );
xor \U$40244 ( \40622 , \40447 , \40449 );
xor \U$40245 ( \40623 , \40622 , \40452 );
and \U$40246 ( \40624 , \40620 , \40623 );
and \U$40247 ( \40625 , \40618 , \40623 );
or \U$40248 ( \40626 , \40621 , \40624 , \40625 );
and \U$40249 ( \40627 , \40616 , \40626 );
xor \U$40250 ( \40628 , \40479 , \40481 );
xor \U$40251 ( \40629 , \40628 , \40484 );
and \U$40252 ( \40630 , \40626 , \40629 );
and \U$40253 ( \40631 , \40616 , \40629 );
or \U$40254 ( \40632 , \40627 , \40630 , \40631 );
xor \U$40255 ( \40633 , \40404 , \40444 );
xor \U$40256 ( \40634 , \40633 , \40455 );
xor \U$40257 ( \40635 , \40468 , \40470 );
xor \U$40258 ( \40636 , \40635 , \40473 );
and \U$40259 ( \40637 , \40634 , \40636 );
and \U$40260 ( \40638 , \40632 , \40637 );
xor \U$40261 ( \40639 , \40492 , \40494 );
xor \U$40262 ( \40640 , \40639 , \40496 );
and \U$40263 ( \40641 , \40637 , \40640 );
and \U$40264 ( \40642 , \40632 , \40640 );
or \U$40265 ( \40643 , \40638 , \40641 , \40642 );
xor \U$40266 ( \40644 , \40302 , \40312 );
xor \U$40267 ( \40645 , \40644 , \40318 );
and \U$40268 ( \40646 , \40643 , \40645 );
xor \U$40269 ( \40647 , \40490 , \40499 );
xor \U$40270 ( \40648 , \40647 , \40502 );
and \U$40271 ( \40649 , \40645 , \40648 );
and \U$40272 ( \40650 , \40643 , \40648 );
or \U$40273 ( \40651 , \40646 , \40649 , \40650 );
and \U$40274 ( \40652 , \40516 , \40651 );
xor \U$40275 ( \40653 , \40516 , \40651 );
xor \U$40276 ( \40654 , \40643 , \40645 );
xor \U$40277 ( \40655 , \40654 , \40648 );
and \U$40278 ( \40656 , \25353 , \32151 );
and \U$40279 ( \40657 , \25348 , \32148 );
nor \U$40280 ( \40658 , \40656 , \40657 );
xnor \U$40281 ( \40659 , \40658 , \31096 );
and \U$40282 ( \40660 , \25806 , \31338 );
and \U$40283 ( \40661 , \25609 , \31336 );
nor \U$40284 ( \40662 , \40660 , \40661 );
xnor \U$40285 ( \40663 , \40662 , \31099 );
and \U$40286 ( \40664 , \40659 , \40663 );
and \U$40287 ( \40665 , \26116 , \30770 );
and \U$40288 ( \40666 , \26108 , \30768 );
nor \U$40289 ( \40667 , \40665 , \40666 );
xnor \U$40290 ( \40668 , \40667 , \30460 );
and \U$40291 ( \40669 , \40663 , \40668 );
and \U$40292 ( \40670 , \40659 , \40668 );
or \U$40293 ( \40671 , \40664 , \40669 , \40670 );
and \U$40294 ( \40672 , \28039 , \28575 );
and \U$40295 ( \40673 , \27837 , \28573 );
nor \U$40296 ( \40674 , \40672 , \40673 );
xnor \U$40297 ( \40675 , \40674 , \28315 );
and \U$40298 ( \40676 , \28514 , \28081 );
and \U$40299 ( \40677 , \28342 , \28079 );
nor \U$40300 ( \40678 , \40676 , \40677 );
xnor \U$40301 ( \40679 , \40678 , \27766 );
and \U$40302 ( \40680 , \40675 , \40679 );
and \U$40303 ( \40681 , \29464 , \27572 );
and \U$40304 ( \40682 , \29040 , \27570 );
nor \U$40305 ( \40683 , \40681 , \40682 );
xnor \U$40306 ( \40684 , \40683 , \27232 );
and \U$40307 ( \40685 , \40679 , \40684 );
and \U$40308 ( \40686 , \40675 , \40684 );
or \U$40309 ( \40687 , \40680 , \40685 , \40686 );
and \U$40310 ( \40688 , \40671 , \40687 );
and \U$40311 ( \40689 , \26590 , \30233 );
and \U$40312 ( \40690 , \26585 , \30231 );
nor \U$40313 ( \40691 , \40689 , \40690 );
xnor \U$40314 ( \40692 , \40691 , \29862 );
and \U$40315 ( \40693 , \27113 , \29671 );
and \U$40316 ( \40694 , \26854 , \29669 );
nor \U$40317 ( \40695 , \40693 , \40694 );
xnor \U$40318 ( \40696 , \40695 , \29353 );
and \U$40319 ( \40697 , \40692 , \40696 );
and \U$40320 ( \40698 , \27494 , \29104 );
and \U$40321 ( \40699 , \27485 , \29102 );
nor \U$40322 ( \40700 , \40698 , \40699 );
xnor \U$40323 ( \40701 , \40700 , \28855 );
and \U$40324 ( \40702 , \40696 , \40701 );
and \U$40325 ( \40703 , \40692 , \40701 );
or \U$40326 ( \40704 , \40697 , \40702 , \40703 );
and \U$40327 ( \40705 , \40687 , \40704 );
and \U$40328 ( \40706 , \40671 , \40704 );
or \U$40329 ( \40707 , \40688 , \40705 , \40706 );
xor \U$40330 ( \40708 , \40520 , \40524 );
xor \U$40331 ( \40709 , \40708 , \40529 );
xor \U$40332 ( \40710 , \40536 , \40540 );
xor \U$40333 ( \40711 , \40710 , \40545 );
and \U$40334 ( \40712 , \40709 , \40711 );
xor \U$40335 ( \40713 , \40568 , \40572 );
xor \U$40336 ( \40714 , \40713 , \40577 );
and \U$40337 ( \40715 , \40711 , \40714 );
and \U$40338 ( \40716 , \40709 , \40714 );
or \U$40339 ( \40717 , \40712 , \40715 , \40716 );
and \U$40340 ( \40718 , \40707 , \40717 );
and \U$40341 ( \40719 , \29715 , \26983 );
and \U$40342 ( \40720 , \29710 , \26981 );
nor \U$40343 ( \40721 , \40719 , \40720 );
xnor \U$40344 ( \40722 , \40721 , \26742 );
and \U$40345 ( \40723 , \30318 , \26517 );
and \U$40346 ( \40724 , \30034 , \26515 );
nor \U$40347 ( \40725 , \40723 , \40724 );
xnor \U$40348 ( \40726 , \40725 , \26329 );
and \U$40349 ( \40727 , \40722 , \40726 );
and \U$40350 ( \40728 , \30895 , \26143 );
and \U$40351 ( \40729 , \30887 , \26141 );
nor \U$40352 ( \40730 , \40728 , \40729 );
xnor \U$40353 ( \40731 , \40730 , \25911 );
and \U$40354 ( \40732 , \40726 , \40731 );
and \U$40355 ( \40733 , \40722 , \40731 );
or \U$40356 ( \40734 , \40727 , \40732 , \40733 );
nand \U$40357 ( \40735 , \32304 , \24972 );
xnor \U$40358 ( \40736 , \40735 , \24787 );
and \U$40359 ( \40737 , \40734 , \40736 );
xor \U$40360 ( \40738 , \40584 , \40588 );
xor \U$40361 ( \40739 , \40738 , \40593 );
and \U$40362 ( \40740 , \40736 , \40739 );
and \U$40363 ( \40741 , \40734 , \40739 );
or \U$40364 ( \40742 , \40737 , \40740 , \40741 );
and \U$40365 ( \40743 , \40717 , \40742 );
and \U$40366 ( \40744 , \40707 , \40742 );
or \U$40367 ( \40745 , \40718 , \40743 , \40744 );
xor \U$40368 ( \40746 , \40389 , \40393 );
xor \U$40369 ( \40747 , \40746 , \40398 );
xor \U$40370 ( \40748 , \40580 , \40596 );
xor \U$40371 ( \40749 , \40748 , \40599 );
and \U$40372 ( \40750 , \40747 , \40749 );
xor \U$40373 ( \40751 , \40605 , \40607 );
xor \U$40374 ( \40752 , \40751 , \40610 );
and \U$40375 ( \40753 , \40749 , \40752 );
and \U$40376 ( \40754 , \40747 , \40752 );
or \U$40377 ( \40755 , \40750 , \40753 , \40754 );
and \U$40378 ( \40756 , \40745 , \40755 );
xor \U$40379 ( \40757 , \40368 , \40384 );
xor \U$40380 ( \40758 , \40757 , \40401 );
and \U$40381 ( \40759 , \40755 , \40758 );
and \U$40382 ( \40760 , \40745 , \40758 );
or \U$40383 ( \40761 , \40756 , \40759 , \40760 );
xor \U$40384 ( \40762 , \40616 , \40626 );
xor \U$40385 ( \40763 , \40762 , \40629 );
and \U$40386 ( \40764 , \40761 , \40763 );
xor \U$40387 ( \40765 , \40634 , \40636 );
and \U$40388 ( \40766 , \40763 , \40765 );
and \U$40389 ( \40767 , \40761 , \40765 );
or \U$40390 ( \40768 , \40764 , \40766 , \40767 );
xor \U$40391 ( \40769 , \40458 , \40476 );
xor \U$40392 ( \40770 , \40769 , \40487 );
and \U$40393 ( \40771 , \40768 , \40770 );
xor \U$40394 ( \40772 , \40632 , \40637 );
xor \U$40395 ( \40773 , \40772 , \40640 );
and \U$40396 ( \40774 , \40770 , \40773 );
and \U$40397 ( \40775 , \40768 , \40773 );
or \U$40398 ( \40776 , \40771 , \40774 , \40775 );
and \U$40399 ( \40777 , \40655 , \40776 );
xor \U$40400 ( \40778 , \40655 , \40776 );
xor \U$40401 ( \40779 , \40768 , \40770 );
xor \U$40402 ( \40780 , \40779 , \40773 );
and \U$40403 ( \40781 , \29710 , \27572 );
and \U$40404 ( \40782 , \29464 , \27570 );
nor \U$40405 ( \40783 , \40781 , \40782 );
xnor \U$40406 ( \40784 , \40783 , \27232 );
and \U$40407 ( \40785 , \30034 , \26983 );
and \U$40408 ( \40786 , \29715 , \26981 );
nor \U$40409 ( \40787 , \40785 , \40786 );
xnor \U$40410 ( \40788 , \40787 , \26742 );
and \U$40411 ( \40789 , \40784 , \40788 );
and \U$40412 ( \40790 , \30887 , \26517 );
and \U$40413 ( \40791 , \30318 , \26515 );
nor \U$40414 ( \40792 , \40790 , \40791 );
xnor \U$40415 ( \40793 , \40792 , \26329 );
and \U$40416 ( \40794 , \40788 , \40793 );
and \U$40417 ( \40795 , \40784 , \40793 );
or \U$40418 ( \40796 , \40789 , \40794 , \40795 );
and \U$40419 ( \40797 , \31498 , \26143 );
and \U$40420 ( \40798 , \30895 , \26141 );
nor \U$40421 ( \40799 , \40797 , \40798 );
xnor \U$40422 ( \40800 , \40799 , \25911 );
and \U$40423 ( \40801 , \31684 , \25692 );
and \U$40424 ( \40802 , \31503 , \25690 );
nor \U$40425 ( \40803 , \40801 , \40802 );
xnor \U$40426 ( \40804 , \40803 , \25549 );
and \U$40427 ( \40805 , \40800 , \40804 );
nand \U$40428 ( \40806 , \32304 , \25367 );
xnor \U$40429 ( \40807 , \40806 , \25123 );
and \U$40430 ( \40808 , \40804 , \40807 );
and \U$40431 ( \40809 , \40800 , \40807 );
or \U$40432 ( \40810 , \40805 , \40808 , \40809 );
and \U$40433 ( \40811 , \40796 , \40810 );
and \U$40434 ( \40812 , \31503 , \25692 );
and \U$40435 ( \40813 , \31498 , \25690 );
nor \U$40436 ( \40814 , \40812 , \40813 );
xnor \U$40437 ( \40815 , \40814 , \25549 );
and \U$40438 ( \40816 , \40810 , \40815 );
and \U$40439 ( \40817 , \40796 , \40815 );
or \U$40440 ( \40818 , \40811 , \40816 , \40817 );
and \U$40441 ( \40819 , \27837 , \29104 );
and \U$40442 ( \40820 , \27494 , \29102 );
nor \U$40443 ( \40821 , \40819 , \40820 );
xnor \U$40444 ( \40822 , \40821 , \28855 );
and \U$40445 ( \40823 , \28342 , \28575 );
and \U$40446 ( \40824 , \28039 , \28573 );
nor \U$40447 ( \40825 , \40823 , \40824 );
xnor \U$40448 ( \40826 , \40825 , \28315 );
and \U$40449 ( \40827 , \40822 , \40826 );
and \U$40450 ( \40828 , \29040 , \28081 );
and \U$40451 ( \40829 , \28514 , \28079 );
nor \U$40452 ( \40830 , \40828 , \40829 );
xnor \U$40453 ( \40831 , \40830 , \27766 );
and \U$40454 ( \40832 , \40826 , \40831 );
and \U$40455 ( \40833 , \40822 , \40831 );
or \U$40456 ( \40834 , \40827 , \40832 , \40833 );
and \U$40457 ( \40835 , \25609 , \32151 );
and \U$40458 ( \40836 , \25353 , \32148 );
nor \U$40459 ( \40837 , \40835 , \40836 );
xnor \U$40460 ( \40838 , \40837 , \31096 );
and \U$40461 ( \40839 , \26108 , \31338 );
and \U$40462 ( \40840 , \25806 , \31336 );
nor \U$40463 ( \40841 , \40839 , \40840 );
xnor \U$40464 ( \40842 , \40841 , \31099 );
and \U$40465 ( \40843 , \40838 , \40842 );
and \U$40466 ( \40844 , \40842 , \25123 );
and \U$40467 ( \40845 , \40838 , \25123 );
or \U$40468 ( \40846 , \40843 , \40844 , \40845 );
and \U$40469 ( \40847 , \40834 , \40846 );
and \U$40470 ( \40848 , \26585 , \30770 );
and \U$40471 ( \40849 , \26116 , \30768 );
nor \U$40472 ( \40850 , \40848 , \40849 );
xnor \U$40473 ( \40851 , \40850 , \30460 );
and \U$40474 ( \40852 , \26854 , \30233 );
and \U$40475 ( \40853 , \26590 , \30231 );
nor \U$40476 ( \40854 , \40852 , \40853 );
xnor \U$40477 ( \40855 , \40854 , \29862 );
and \U$40478 ( \40856 , \40851 , \40855 );
and \U$40479 ( \40857 , \27485 , \29671 );
and \U$40480 ( \40858 , \27113 , \29669 );
nor \U$40481 ( \40859 , \40857 , \40858 );
xnor \U$40482 ( \40860 , \40859 , \29353 );
and \U$40483 ( \40861 , \40855 , \40860 );
and \U$40484 ( \40862 , \40851 , \40860 );
or \U$40485 ( \40863 , \40856 , \40861 , \40862 );
and \U$40486 ( \40864 , \40846 , \40863 );
and \U$40487 ( \40865 , \40834 , \40863 );
or \U$40488 ( \40866 , \40847 , \40864 , \40865 );
and \U$40489 ( \40867 , \40818 , \40866 );
and \U$40490 ( \40868 , \32304 , \25369 );
and \U$40491 ( \40869 , \31684 , \25367 );
nor \U$40492 ( \40870 , \40868 , \40869 );
xnor \U$40493 ( \40871 , \40870 , \25123 );
xor \U$40494 ( \40872 , \40722 , \40726 );
xor \U$40495 ( \40873 , \40872 , \40731 );
and \U$40496 ( \40874 , \40871 , \40873 );
xor \U$40497 ( \40875 , \40675 , \40679 );
xor \U$40498 ( \40876 , \40875 , \40684 );
and \U$40499 ( \40877 , \40873 , \40876 );
and \U$40500 ( \40878 , \40871 , \40876 );
or \U$40501 ( \40879 , \40874 , \40877 , \40878 );
and \U$40502 ( \40880 , \40866 , \40879 );
and \U$40503 ( \40881 , \40818 , \40879 );
or \U$40504 ( \40882 , \40867 , \40880 , \40881 );
xor \U$40505 ( \40883 , \40553 , \40557 );
xor \U$40506 ( \40884 , \40883 , \24787 );
xor \U$40507 ( \40885 , \40709 , \40711 );
xor \U$40508 ( \40886 , \40885 , \40714 );
and \U$40509 ( \40887 , \40884 , \40886 );
xor \U$40510 ( \40888 , \40734 , \40736 );
xor \U$40511 ( \40889 , \40888 , \40739 );
and \U$40512 ( \40890 , \40886 , \40889 );
and \U$40513 ( \40891 , \40884 , \40889 );
or \U$40514 ( \40892 , \40887 , \40890 , \40891 );
and \U$40515 ( \40893 , \40882 , \40892 );
xor \U$40516 ( \40894 , \40532 , \40548 );
xor \U$40517 ( \40895 , \40894 , \40561 );
and \U$40518 ( \40896 , \40892 , \40895 );
and \U$40519 ( \40897 , \40882 , \40895 );
or \U$40520 ( \40898 , \40893 , \40896 , \40897 );
xor \U$40521 ( \40899 , \40707 , \40717 );
xor \U$40522 ( \40900 , \40899 , \40742 );
xor \U$40523 ( \40901 , \40747 , \40749 );
xor \U$40524 ( \40902 , \40901 , \40752 );
and \U$40525 ( \40903 , \40900 , \40902 );
and \U$40526 ( \40904 , \40898 , \40903 );
xor \U$40527 ( \40905 , \40618 , \40620 );
xor \U$40528 ( \40906 , \40905 , \40623 );
and \U$40529 ( \40907 , \40903 , \40906 );
and \U$40530 ( \40908 , \40898 , \40906 );
or \U$40531 ( \40909 , \40904 , \40907 , \40908 );
xor \U$40532 ( \40910 , \40564 , \40602 );
xor \U$40533 ( \40911 , \40910 , \40613 );
xor \U$40534 ( \40912 , \40745 , \40755 );
xor \U$40535 ( \40913 , \40912 , \40758 );
and \U$40536 ( \40914 , \40911 , \40913 );
and \U$40537 ( \40915 , \40909 , \40914 );
xor \U$40538 ( \40916 , \40761 , \40763 );
xor \U$40539 ( \40917 , \40916 , \40765 );
and \U$40540 ( \40918 , \40914 , \40917 );
and \U$40541 ( \40919 , \40909 , \40917 );
or \U$40542 ( \40920 , \40915 , \40918 , \40919 );
and \U$40543 ( \40921 , \40780 , \40920 );
xor \U$40544 ( \40922 , \40780 , \40920 );
xor \U$40545 ( \40923 , \40909 , \40914 );
xor \U$40546 ( \40924 , \40923 , \40917 );
and \U$40547 ( \40925 , \27113 , \30233 );
and \U$40548 ( \40926 , \26854 , \30231 );
nor \U$40549 ( \40927 , \40925 , \40926 );
xnor \U$40550 ( \40928 , \40927 , \29862 );
and \U$40551 ( \40929 , \27494 , \29671 );
and \U$40552 ( \40930 , \27485 , \29669 );
nor \U$40553 ( \40931 , \40929 , \40930 );
xnor \U$40554 ( \40932 , \40931 , \29353 );
and \U$40555 ( \40933 , \40928 , \40932 );
and \U$40556 ( \40934 , \28039 , \29104 );
and \U$40557 ( \40935 , \27837 , \29102 );
nor \U$40558 ( \40936 , \40934 , \40935 );
xnor \U$40559 ( \40937 , \40936 , \28855 );
and \U$40560 ( \40938 , \40932 , \40937 );
and \U$40561 ( \40939 , \40928 , \40937 );
or \U$40562 ( \40940 , \40933 , \40938 , \40939 );
and \U$40563 ( \40941 , \25806 , \32151 );
and \U$40564 ( \40942 , \25609 , \32148 );
nor \U$40565 ( \40943 , \40941 , \40942 );
xnor \U$40566 ( \40944 , \40943 , \31096 );
and \U$40567 ( \40945 , \26116 , \31338 );
and \U$40568 ( \40946 , \26108 , \31336 );
nor \U$40569 ( \40947 , \40945 , \40946 );
xnor \U$40570 ( \40948 , \40947 , \31099 );
and \U$40571 ( \40949 , \40944 , \40948 );
and \U$40572 ( \40950 , \26590 , \30770 );
and \U$40573 ( \40951 , \26585 , \30768 );
nor \U$40574 ( \40952 , \40950 , \40951 );
xnor \U$40575 ( \40953 , \40952 , \30460 );
and \U$40576 ( \40954 , \40948 , \40953 );
and \U$40577 ( \40955 , \40944 , \40953 );
or \U$40578 ( \40956 , \40949 , \40954 , \40955 );
and \U$40579 ( \40957 , \40940 , \40956 );
and \U$40580 ( \40958 , \28514 , \28575 );
and \U$40581 ( \40959 , \28342 , \28573 );
nor \U$40582 ( \40960 , \40958 , \40959 );
xnor \U$40583 ( \40961 , \40960 , \28315 );
and \U$40584 ( \40962 , \29464 , \28081 );
and \U$40585 ( \40963 , \29040 , \28079 );
nor \U$40586 ( \40964 , \40962 , \40963 );
xnor \U$40587 ( \40965 , \40964 , \27766 );
and \U$40588 ( \40966 , \40961 , \40965 );
and \U$40589 ( \40967 , \29715 , \27572 );
and \U$40590 ( \40968 , \29710 , \27570 );
nor \U$40591 ( \40969 , \40967 , \40968 );
xnor \U$40592 ( \40970 , \40969 , \27232 );
and \U$40593 ( \40971 , \40965 , \40970 );
and \U$40594 ( \40972 , \40961 , \40970 );
or \U$40595 ( \40973 , \40966 , \40971 , \40972 );
and \U$40596 ( \40974 , \40956 , \40973 );
and \U$40597 ( \40975 , \40940 , \40973 );
or \U$40598 ( \40976 , \40957 , \40974 , \40975 );
xor \U$40599 ( \40977 , \40822 , \40826 );
xor \U$40600 ( \40978 , \40977 , \40831 );
xor \U$40601 ( \40979 , \40838 , \40842 );
xor \U$40602 ( \40980 , \40979 , \25123 );
and \U$40603 ( \40981 , \40978 , \40980 );
xor \U$40604 ( \40982 , \40851 , \40855 );
xor \U$40605 ( \40983 , \40982 , \40860 );
and \U$40606 ( \40984 , \40980 , \40983 );
and \U$40607 ( \40985 , \40978 , \40983 );
or \U$40608 ( \40986 , \40981 , \40984 , \40985 );
and \U$40609 ( \40987 , \40976 , \40986 );
and \U$40610 ( \40988 , \30318 , \26983 );
and \U$40611 ( \40989 , \30034 , \26981 );
nor \U$40612 ( \40990 , \40988 , \40989 );
xnor \U$40613 ( \40991 , \40990 , \26742 );
and \U$40614 ( \40992 , \30895 , \26517 );
and \U$40615 ( \40993 , \30887 , \26515 );
nor \U$40616 ( \40994 , \40992 , \40993 );
xnor \U$40617 ( \40995 , \40994 , \26329 );
and \U$40618 ( \40996 , \40991 , \40995 );
and \U$40619 ( \40997 , \31503 , \26143 );
and \U$40620 ( \40998 , \31498 , \26141 );
nor \U$40621 ( \40999 , \40997 , \40998 );
xnor \U$40622 ( \41000 , \40999 , \25911 );
and \U$40623 ( \41001 , \40995 , \41000 );
and \U$40624 ( \41002 , \40991 , \41000 );
or \U$40625 ( \41003 , \40996 , \41001 , \41002 );
xor \U$40626 ( \41004 , \40784 , \40788 );
xor \U$40627 ( \41005 , \41004 , \40793 );
and \U$40628 ( \41006 , \41003 , \41005 );
xor \U$40629 ( \41007 , \40800 , \40804 );
xor \U$40630 ( \41008 , \41007 , \40807 );
and \U$40631 ( \41009 , \41005 , \41008 );
and \U$40632 ( \41010 , \41003 , \41008 );
or \U$40633 ( \41011 , \41006 , \41009 , \41010 );
and \U$40634 ( \41012 , \40986 , \41011 );
and \U$40635 ( \41013 , \40976 , \41011 );
or \U$40636 ( \41014 , \40987 , \41012 , \41013 );
xor \U$40637 ( \41015 , \40659 , \40663 );
xor \U$40638 ( \41016 , \41015 , \40668 );
xor \U$40639 ( \41017 , \40692 , \40696 );
xor \U$40640 ( \41018 , \41017 , \40701 );
and \U$40641 ( \41019 , \41016 , \41018 );
xor \U$40642 ( \41020 , \40871 , \40873 );
xor \U$40643 ( \41021 , \41020 , \40876 );
and \U$40644 ( \41022 , \41018 , \41021 );
and \U$40645 ( \41023 , \41016 , \41021 );
or \U$40646 ( \41024 , \41019 , \41022 , \41023 );
and \U$40647 ( \41025 , \41014 , \41024 );
xor \U$40648 ( \41026 , \40671 , \40687 );
xor \U$40649 ( \41027 , \41026 , \40704 );
and \U$40650 ( \41028 , \41024 , \41027 );
and \U$40651 ( \41029 , \41014 , \41027 );
or \U$40652 ( \41030 , \41025 , \41028 , \41029 );
xor \U$40653 ( \41031 , \40882 , \40892 );
xor \U$40654 ( \41032 , \41031 , \40895 );
and \U$40655 ( \41033 , \41030 , \41032 );
xor \U$40656 ( \41034 , \40900 , \40902 );
and \U$40657 ( \41035 , \41032 , \41034 );
and \U$40658 ( \41036 , \41030 , \41034 );
or \U$40659 ( \41037 , \41033 , \41035 , \41036 );
xor \U$40660 ( \41038 , \40898 , \40903 );
xor \U$40661 ( \41039 , \41038 , \40906 );
and \U$40662 ( \41040 , \41037 , \41039 );
xor \U$40663 ( \41041 , \40911 , \40913 );
and \U$40664 ( \41042 , \41039 , \41041 );
and \U$40665 ( \41043 , \41037 , \41041 );
or \U$40666 ( \41044 , \41040 , \41042 , \41043 );
and \U$40667 ( \41045 , \40924 , \41044 );
xor \U$40668 ( \41046 , \40924 , \41044 );
xor \U$40669 ( \41047 , \41037 , \41039 );
xor \U$40670 ( \41048 , \41047 , \41041 );
and \U$40671 ( \41049 , \26854 , \30770 );
and \U$40672 ( \41050 , \26590 , \30768 );
nor \U$40673 ( \41051 , \41049 , \41050 );
xnor \U$40674 ( \41052 , \41051 , \30460 );
and \U$40675 ( \41053 , \27485 , \30233 );
and \U$40676 ( \41054 , \27113 , \30231 );
nor \U$40677 ( \41055 , \41053 , \41054 );
xnor \U$40678 ( \41056 , \41055 , \29862 );
and \U$40679 ( \41057 , \41052 , \41056 );
and \U$40680 ( \41058 , \27837 , \29671 );
and \U$40681 ( \41059 , \27494 , \29669 );
nor \U$40682 ( \41060 , \41058 , \41059 );
xnor \U$40683 ( \41061 , \41060 , \29353 );
and \U$40684 ( \41062 , \41056 , \41061 );
and \U$40685 ( \41063 , \41052 , \41061 );
or \U$40686 ( \41064 , \41057 , \41062 , \41063 );
and \U$40687 ( \41065 , \26108 , \32151 );
and \U$40688 ( \41066 , \25806 , \32148 );
nor \U$40689 ( \41067 , \41065 , \41066 );
xnor \U$40690 ( \41068 , \41067 , \31096 );
and \U$40691 ( \41069 , \26585 , \31338 );
and \U$40692 ( \41070 , \26116 , \31336 );
nor \U$40693 ( \41071 , \41069 , \41070 );
xnor \U$40694 ( \41072 , \41071 , \31099 );
and \U$40695 ( \41073 , \41068 , \41072 );
and \U$40696 ( \41074 , \41072 , \25549 );
and \U$40697 ( \41075 , \41068 , \25549 );
or \U$40698 ( \41076 , \41073 , \41074 , \41075 );
and \U$40699 ( \41077 , \41064 , \41076 );
and \U$40700 ( \41078 , \28342 , \29104 );
and \U$40701 ( \41079 , \28039 , \29102 );
nor \U$40702 ( \41080 , \41078 , \41079 );
xnor \U$40703 ( \41081 , \41080 , \28855 );
and \U$40704 ( \41082 , \29040 , \28575 );
and \U$40705 ( \41083 , \28514 , \28573 );
nor \U$40706 ( \41084 , \41082 , \41083 );
xnor \U$40707 ( \41085 , \41084 , \28315 );
and \U$40708 ( \41086 , \41081 , \41085 );
and \U$40709 ( \41087 , \29710 , \28081 );
and \U$40710 ( \41088 , \29464 , \28079 );
nor \U$40711 ( \41089 , \41087 , \41088 );
xnor \U$40712 ( \41090 , \41089 , \27766 );
and \U$40713 ( \41091 , \41085 , \41090 );
and \U$40714 ( \41092 , \41081 , \41090 );
or \U$40715 ( \41093 , \41086 , \41091 , \41092 );
and \U$40716 ( \41094 , \41076 , \41093 );
and \U$40717 ( \41095 , \41064 , \41093 );
or \U$40718 ( \41096 , \41077 , \41094 , \41095 );
and \U$40719 ( \41097 , \30034 , \27572 );
and \U$40720 ( \41098 , \29715 , \27570 );
nor \U$40721 ( \41099 , \41097 , \41098 );
xnor \U$40722 ( \41100 , \41099 , \27232 );
and \U$40723 ( \41101 , \30887 , \26983 );
and \U$40724 ( \41102 , \30318 , \26981 );
nor \U$40725 ( \41103 , \41101 , \41102 );
xnor \U$40726 ( \41104 , \41103 , \26742 );
and \U$40727 ( \41105 , \41100 , \41104 );
and \U$40728 ( \41106 , \31498 , \26517 );
and \U$40729 ( \41107 , \30895 , \26515 );
nor \U$40730 ( \41108 , \41106 , \41107 );
xnor \U$40731 ( \41109 , \41108 , \26329 );
and \U$40732 ( \41110 , \41104 , \41109 );
and \U$40733 ( \41111 , \41100 , \41109 );
or \U$40734 ( \41112 , \41105 , \41110 , \41111 );
and \U$40735 ( \41113 , \31684 , \26143 );
and \U$40736 ( \41114 , \31503 , \26141 );
nor \U$40737 ( \41115 , \41113 , \41114 );
xnor \U$40738 ( \41116 , \41115 , \25911 );
nand \U$40739 ( \41117 , \32304 , \25690 );
xnor \U$40740 ( \41118 , \41117 , \25549 );
and \U$40741 ( \41119 , \41116 , \41118 );
and \U$40742 ( \41120 , \41112 , \41119 );
and \U$40743 ( \41121 , \32304 , \25692 );
and \U$40744 ( \41122 , \31684 , \25690 );
nor \U$40745 ( \41123 , \41121 , \41122 );
xnor \U$40746 ( \41124 , \41123 , \25549 );
and \U$40747 ( \41125 , \41119 , \41124 );
and \U$40748 ( \41126 , \41112 , \41124 );
or \U$40749 ( \41127 , \41120 , \41125 , \41126 );
and \U$40750 ( \41128 , \41096 , \41127 );
xor \U$40751 ( \41129 , \40928 , \40932 );
xor \U$40752 ( \41130 , \41129 , \40937 );
xor \U$40753 ( \41131 , \40991 , \40995 );
xor \U$40754 ( \41132 , \41131 , \41000 );
and \U$40755 ( \41133 , \41130 , \41132 );
xor \U$40756 ( \41134 , \40961 , \40965 );
xor \U$40757 ( \41135 , \41134 , \40970 );
and \U$40758 ( \41136 , \41132 , \41135 );
and \U$40759 ( \41137 , \41130 , \41135 );
or \U$40760 ( \41138 , \41133 , \41136 , \41137 );
and \U$40761 ( \41139 , \41127 , \41138 );
and \U$40762 ( \41140 , \41096 , \41138 );
or \U$40763 ( \41141 , \41128 , \41139 , \41140 );
xor \U$40764 ( \41142 , \40940 , \40956 );
xor \U$40765 ( \41143 , \41142 , \40973 );
xor \U$40766 ( \41144 , \40978 , \40980 );
xor \U$40767 ( \41145 , \41144 , \40983 );
and \U$40768 ( \41146 , \41143 , \41145 );
xor \U$40769 ( \41147 , \41003 , \41005 );
xor \U$40770 ( \41148 , \41147 , \41008 );
and \U$40771 ( \41149 , \41145 , \41148 );
and \U$40772 ( \41150 , \41143 , \41148 );
or \U$40773 ( \41151 , \41146 , \41149 , \41150 );
and \U$40774 ( \41152 , \41141 , \41151 );
xor \U$40775 ( \41153 , \40796 , \40810 );
xor \U$40776 ( \41154 , \41153 , \40815 );
and \U$40777 ( \41155 , \41151 , \41154 );
and \U$40778 ( \41156 , \41141 , \41154 );
or \U$40779 ( \41157 , \41152 , \41155 , \41156 );
xor \U$40780 ( \41158 , \40834 , \40846 );
xor \U$40781 ( \41159 , \41158 , \40863 );
xor \U$40782 ( \41160 , \40976 , \40986 );
xor \U$40783 ( \41161 , \41160 , \41011 );
and \U$40784 ( \41162 , \41159 , \41161 );
xor \U$40785 ( \41163 , \41016 , \41018 );
xor \U$40786 ( \41164 , \41163 , \41021 );
and \U$40787 ( \41165 , \41161 , \41164 );
and \U$40788 ( \41166 , \41159 , \41164 );
or \U$40789 ( \41167 , \41162 , \41165 , \41166 );
and \U$40790 ( \41168 , \41157 , \41167 );
xor \U$40791 ( \41169 , \40884 , \40886 );
xor \U$40792 ( \41170 , \41169 , \40889 );
and \U$40793 ( \41171 , \41167 , \41170 );
and \U$40794 ( \41172 , \41157 , \41170 );
or \U$40795 ( \41173 , \41168 , \41171 , \41172 );
xor \U$40796 ( \41174 , \40818 , \40866 );
xor \U$40797 ( \41175 , \41174 , \40879 );
xor \U$40798 ( \41176 , \41014 , \41024 );
xor \U$40799 ( \41177 , \41176 , \41027 );
and \U$40800 ( \41178 , \41175 , \41177 );
and \U$40801 ( \41179 , \41173 , \41178 );
xor \U$40802 ( \41180 , \41030 , \41032 );
xor \U$40803 ( \41181 , \41180 , \41034 );
and \U$40804 ( \41182 , \41178 , \41181 );
and \U$40805 ( \41183 , \41173 , \41181 );
or \U$40806 ( \41184 , \41179 , \41182 , \41183 );
and \U$40807 ( \41185 , \41048 , \41184 );
xor \U$40808 ( \41186 , \41048 , \41184 );
xor \U$40809 ( \41187 , \41173 , \41178 );
xor \U$40810 ( \41188 , \41187 , \41181 );
and \U$40811 ( \41189 , \27494 , \30233 );
and \U$40812 ( \41190 , \27485 , \30231 );
nor \U$40813 ( \41191 , \41189 , \41190 );
xnor \U$40814 ( \41192 , \41191 , \29862 );
and \U$40815 ( \41193 , \28039 , \29671 );
and \U$40816 ( \41194 , \27837 , \29669 );
nor \U$40817 ( \41195 , \41193 , \41194 );
xnor \U$40818 ( \41196 , \41195 , \29353 );
and \U$40819 ( \41197 , \41192 , \41196 );
and \U$40820 ( \41198 , \28514 , \29104 );
and \U$40821 ( \41199 , \28342 , \29102 );
nor \U$40822 ( \41200 , \41198 , \41199 );
xnor \U$40823 ( \41201 , \41200 , \28855 );
and \U$40824 ( \41202 , \41196 , \41201 );
and \U$40825 ( \41203 , \41192 , \41201 );
or \U$40826 ( \41204 , \41197 , \41202 , \41203 );
and \U$40827 ( \41205 , \29464 , \28575 );
and \U$40828 ( \41206 , \29040 , \28573 );
nor \U$40829 ( \41207 , \41205 , \41206 );
xnor \U$40830 ( \41208 , \41207 , \28315 );
and \U$40831 ( \41209 , \29715 , \28081 );
and \U$40832 ( \41210 , \29710 , \28079 );
nor \U$40833 ( \41211 , \41209 , \41210 );
xnor \U$40834 ( \41212 , \41211 , \27766 );
and \U$40835 ( \41213 , \41208 , \41212 );
and \U$40836 ( \41214 , \30318 , \27572 );
and \U$40837 ( \41215 , \30034 , \27570 );
nor \U$40838 ( \41216 , \41214 , \41215 );
xnor \U$40839 ( \41217 , \41216 , \27232 );
and \U$40840 ( \41218 , \41212 , \41217 );
and \U$40841 ( \41219 , \41208 , \41217 );
or \U$40842 ( \41220 , \41213 , \41218 , \41219 );
and \U$40843 ( \41221 , \41204 , \41220 );
and \U$40844 ( \41222 , \26116 , \32151 );
and \U$40845 ( \41223 , \26108 , \32148 );
nor \U$40846 ( \41224 , \41222 , \41223 );
xnor \U$40847 ( \41225 , \41224 , \31096 );
and \U$40848 ( \41226 , \26590 , \31338 );
and \U$40849 ( \41227 , \26585 , \31336 );
nor \U$40850 ( \41228 , \41226 , \41227 );
xnor \U$40851 ( \41229 , \41228 , \31099 );
and \U$40852 ( \41230 , \41225 , \41229 );
and \U$40853 ( \41231 , \27113 , \30770 );
and \U$40854 ( \41232 , \26854 , \30768 );
nor \U$40855 ( \41233 , \41231 , \41232 );
xnor \U$40856 ( \41234 , \41233 , \30460 );
and \U$40857 ( \41235 , \41229 , \41234 );
and \U$40858 ( \41236 , \41225 , \41234 );
or \U$40859 ( \41237 , \41230 , \41235 , \41236 );
and \U$40860 ( \41238 , \41220 , \41237 );
and \U$40861 ( \41239 , \41204 , \41237 );
or \U$40862 ( \41240 , \41221 , \41238 , \41239 );
xor \U$40863 ( \41241 , \41052 , \41056 );
xor \U$40864 ( \41242 , \41241 , \41061 );
xor \U$40865 ( \41243 , \41068 , \41072 );
xor \U$40866 ( \41244 , \41243 , \25549 );
and \U$40867 ( \41245 , \41242 , \41244 );
xor \U$40868 ( \41246 , \41081 , \41085 );
xor \U$40869 ( \41247 , \41246 , \41090 );
and \U$40870 ( \41248 , \41244 , \41247 );
and \U$40871 ( \41249 , \41242 , \41247 );
or \U$40872 ( \41250 , \41245 , \41248 , \41249 );
and \U$40873 ( \41251 , \41240 , \41250 );
and \U$40874 ( \41252 , \30895 , \26983 );
and \U$40875 ( \41253 , \30887 , \26981 );
nor \U$40876 ( \41254 , \41252 , \41253 );
xnor \U$40877 ( \41255 , \41254 , \26742 );
and \U$40878 ( \41256 , \31503 , \26517 );
and \U$40879 ( \41257 , \31498 , \26515 );
nor \U$40880 ( \41258 , \41256 , \41257 );
xnor \U$40881 ( \41259 , \41258 , \26329 );
and \U$40882 ( \41260 , \41255 , \41259 );
and \U$40883 ( \41261 , \32304 , \26143 );
and \U$40884 ( \41262 , \31684 , \26141 );
nor \U$40885 ( \41263 , \41261 , \41262 );
xnor \U$40886 ( \41264 , \41263 , \25911 );
and \U$40887 ( \41265 , \41259 , \41264 );
and \U$40888 ( \41266 , \41255 , \41264 );
or \U$40889 ( \41267 , \41260 , \41265 , \41266 );
xor \U$40890 ( \41268 , \41100 , \41104 );
xor \U$40891 ( \41269 , \41268 , \41109 );
and \U$40892 ( \41270 , \41267 , \41269 );
xor \U$40893 ( \41271 , \41116 , \41118 );
and \U$40894 ( \41272 , \41269 , \41271 );
and \U$40895 ( \41273 , \41267 , \41271 );
or \U$40896 ( \41274 , \41270 , \41272 , \41273 );
and \U$40897 ( \41275 , \41250 , \41274 );
and \U$40898 ( \41276 , \41240 , \41274 );
or \U$40899 ( \41277 , \41251 , \41275 , \41276 );
xor \U$40900 ( \41278 , \40944 , \40948 );
xor \U$40901 ( \41279 , \41278 , \40953 );
xor \U$40902 ( \41280 , \41112 , \41119 );
xor \U$40903 ( \41281 , \41280 , \41124 );
and \U$40904 ( \41282 , \41279 , \41281 );
xor \U$40905 ( \41283 , \41130 , \41132 );
xor \U$40906 ( \41284 , \41283 , \41135 );
and \U$40907 ( \41285 , \41281 , \41284 );
and \U$40908 ( \41286 , \41279 , \41284 );
or \U$40909 ( \41287 , \41282 , \41285 , \41286 );
and \U$40910 ( \41288 , \41277 , \41287 );
xor \U$40911 ( \41289 , \41143 , \41145 );
xor \U$40912 ( \41290 , \41289 , \41148 );
and \U$40913 ( \41291 , \41287 , \41290 );
and \U$40914 ( \41292 , \41277 , \41290 );
or \U$40915 ( \41293 , \41288 , \41291 , \41292 );
xor \U$40916 ( \41294 , \41141 , \41151 );
xor \U$40917 ( \41295 , \41294 , \41154 );
and \U$40918 ( \41296 , \41293 , \41295 );
xor \U$40919 ( \41297 , \41159 , \41161 );
xor \U$40920 ( \41298 , \41297 , \41164 );
and \U$40921 ( \41299 , \41295 , \41298 );
and \U$40922 ( \41300 , \41293 , \41298 );
or \U$40923 ( \41301 , \41296 , \41299 , \41300 );
xor \U$40924 ( \41302 , \41157 , \41167 );
xor \U$40925 ( \41303 , \41302 , \41170 );
and \U$40926 ( \41304 , \41301 , \41303 );
xor \U$40927 ( \41305 , \41175 , \41177 );
and \U$40928 ( \41306 , \41303 , \41305 );
and \U$40929 ( \41307 , \41301 , \41305 );
or \U$40930 ( \41308 , \41304 , \41306 , \41307 );
and \U$40931 ( \41309 , \41188 , \41308 );
xor \U$40932 ( \41310 , \41188 , \41308 );
xor \U$40933 ( \41311 , \41301 , \41303 );
xor \U$40934 ( \41312 , \41311 , \41305 );
and \U$40935 ( \41313 , \27485 , \30770 );
and \U$40936 ( \41314 , \27113 , \30768 );
nor \U$40937 ( \41315 , \41313 , \41314 );
xnor \U$40938 ( \41316 , \41315 , \30460 );
and \U$40939 ( \41317 , \27837 , \30233 );
and \U$40940 ( \41318 , \27494 , \30231 );
nor \U$40941 ( \41319 , \41317 , \41318 );
xnor \U$40942 ( \41320 , \41319 , \29862 );
and \U$40943 ( \41321 , \41316 , \41320 );
and \U$40944 ( \41322 , \28342 , \29671 );
and \U$40945 ( \41323 , \28039 , \29669 );
nor \U$40946 ( \41324 , \41322 , \41323 );
xnor \U$40947 ( \41325 , \41324 , \29353 );
and \U$40948 ( \41326 , \41320 , \41325 );
and \U$40949 ( \41327 , \41316 , \41325 );
or \U$40950 ( \41328 , \41321 , \41326 , \41327 );
and \U$40951 ( \41329 , \29040 , \29104 );
and \U$40952 ( \41330 , \28514 , \29102 );
nor \U$40953 ( \41331 , \41329 , \41330 );
xnor \U$40954 ( \41332 , \41331 , \28855 );
and \U$40955 ( \41333 , \29710 , \28575 );
and \U$40956 ( \41334 , \29464 , \28573 );
nor \U$40957 ( \41335 , \41333 , \41334 );
xnor \U$40958 ( \41336 , \41335 , \28315 );
and \U$40959 ( \41337 , \41332 , \41336 );
and \U$40960 ( \41338 , \30034 , \28081 );
and \U$40961 ( \41339 , \29715 , \28079 );
nor \U$40962 ( \41340 , \41338 , \41339 );
xnor \U$40963 ( \41341 , \41340 , \27766 );
and \U$40964 ( \41342 , \41336 , \41341 );
and \U$40965 ( \41343 , \41332 , \41341 );
or \U$40966 ( \41344 , \41337 , \41342 , \41343 );
and \U$40967 ( \41345 , \41328 , \41344 );
and \U$40968 ( \41346 , \26585 , \32151 );
and \U$40969 ( \41347 , \26116 , \32148 );
nor \U$40970 ( \41348 , \41346 , \41347 );
xnor \U$40971 ( \41349 , \41348 , \31096 );
and \U$40972 ( \41350 , \26854 , \31338 );
and \U$40973 ( \41351 , \26590 , \31336 );
nor \U$40974 ( \41352 , \41350 , \41351 );
xnor \U$40975 ( \41353 , \41352 , \31099 );
and \U$40976 ( \41354 , \41349 , \41353 );
and \U$40977 ( \41355 , \41353 , \25911 );
and \U$40978 ( \41356 , \41349 , \25911 );
or \U$40979 ( \41357 , \41354 , \41355 , \41356 );
and \U$40980 ( \41358 , \41344 , \41357 );
and \U$40981 ( \41359 , \41328 , \41357 );
or \U$40982 ( \41360 , \41345 , \41358 , \41359 );
and \U$40983 ( \41361 , \30887 , \27572 );
and \U$40984 ( \41362 , \30318 , \27570 );
nor \U$40985 ( \41363 , \41361 , \41362 );
xnor \U$40986 ( \41364 , \41363 , \27232 );
and \U$40987 ( \41365 , \31498 , \26983 );
and \U$40988 ( \41366 , \30895 , \26981 );
nor \U$40989 ( \41367 , \41365 , \41366 );
xnor \U$40990 ( \41368 , \41367 , \26742 );
and \U$40991 ( \41369 , \41364 , \41368 );
and \U$40992 ( \41370 , \31684 , \26517 );
and \U$40993 ( \41371 , \31503 , \26515 );
nor \U$40994 ( \41372 , \41370 , \41371 );
xnor \U$40995 ( \41373 , \41372 , \26329 );
and \U$40996 ( \41374 , \41368 , \41373 );
and \U$40997 ( \41375 , \41364 , \41373 );
or \U$40998 ( \41376 , \41369 , \41374 , \41375 );
xor \U$40999 ( \41377 , \41208 , \41212 );
xor \U$41000 ( \41378 , \41377 , \41217 );
and \U$41001 ( \41379 , \41376 , \41378 );
xor \U$41002 ( \41380 , \41255 , \41259 );
xor \U$41003 ( \41381 , \41380 , \41264 );
and \U$41004 ( \41382 , \41378 , \41381 );
and \U$41005 ( \41383 , \41376 , \41381 );
or \U$41006 ( \41384 , \41379 , \41382 , \41383 );
and \U$41007 ( \41385 , \41360 , \41384 );
xor \U$41008 ( \41386 , \41192 , \41196 );
xor \U$41009 ( \41387 , \41386 , \41201 );
xor \U$41010 ( \41388 , \41225 , \41229 );
xor \U$41011 ( \41389 , \41388 , \41234 );
and \U$41012 ( \41390 , \41387 , \41389 );
and \U$41013 ( \41391 , \41384 , \41390 );
and \U$41014 ( \41392 , \41360 , \41390 );
or \U$41015 ( \41393 , \41385 , \41391 , \41392 );
xor \U$41016 ( \41394 , \41204 , \41220 );
xor \U$41017 ( \41395 , \41394 , \41237 );
xor \U$41018 ( \41396 , \41242 , \41244 );
xor \U$41019 ( \41397 , \41396 , \41247 );
and \U$41020 ( \41398 , \41395 , \41397 );
xor \U$41021 ( \41399 , \41267 , \41269 );
xor \U$41022 ( \41400 , \41399 , \41271 );
and \U$41023 ( \41401 , \41397 , \41400 );
and \U$41024 ( \41402 , \41395 , \41400 );
or \U$41025 ( \41403 , \41398 , \41401 , \41402 );
and \U$41026 ( \41404 , \41393 , \41403 );
xor \U$41027 ( \41405 , \41064 , \41076 );
xor \U$41028 ( \41406 , \41405 , \41093 );
and \U$41029 ( \41407 , \41403 , \41406 );
and \U$41030 ( \41408 , \41393 , \41406 );
or \U$41031 ( \41409 , \41404 , \41407 , \41408 );
xor \U$41032 ( \41410 , \41240 , \41250 );
xor \U$41033 ( \41411 , \41410 , \41274 );
xor \U$41034 ( \41412 , \41279 , \41281 );
xor \U$41035 ( \41413 , \41412 , \41284 );
and \U$41036 ( \41414 , \41411 , \41413 );
and \U$41037 ( \41415 , \41409 , \41414 );
xor \U$41038 ( \41416 , \41096 , \41127 );
xor \U$41039 ( \41417 , \41416 , \41138 );
and \U$41040 ( \41418 , \41414 , \41417 );
and \U$41041 ( \41419 , \41409 , \41417 );
or \U$41042 ( \41420 , \41415 , \41418 , \41419 );
xor \U$41043 ( \41421 , \41293 , \41295 );
xor \U$41044 ( \41422 , \41421 , \41298 );
and \U$41045 ( \41423 , \41420 , \41422 );
and \U$41046 ( \41424 , \41312 , \41423 );
xor \U$41047 ( \41425 , \41312 , \41423 );
xor \U$41048 ( \41426 , \41420 , \41422 );
xor \U$41049 ( \41427 , \41409 , \41414 );
xor \U$41050 ( \41428 , \41427 , \41417 );
xor \U$41051 ( \41429 , \41277 , \41287 );
xor \U$41052 ( \41430 , \41429 , \41290 );
and \U$41053 ( \41431 , \41428 , \41430 );
and \U$41054 ( \41432 , \41426 , \41431 );
xor \U$41055 ( \41433 , \41426 , \41431 );
xor \U$41056 ( \41434 , \41428 , \41430 );
and \U$41057 ( \41435 , \26590 , \32151 );
and \U$41058 ( \41436 , \26585 , \32148 );
nor \U$41059 ( \41437 , \41435 , \41436 );
xnor \U$41060 ( \41438 , \41437 , \31096 );
and \U$41061 ( \41439 , \27113 , \31338 );
and \U$41062 ( \41440 , \26854 , \31336 );
nor \U$41063 ( \41441 , \41439 , \41440 );
xnor \U$41064 ( \41442 , \41441 , \31099 );
and \U$41065 ( \41443 , \41438 , \41442 );
and \U$41066 ( \41444 , \27494 , \30770 );
and \U$41067 ( \41445 , \27485 , \30768 );
nor \U$41068 ( \41446 , \41444 , \41445 );
xnor \U$41069 ( \41447 , \41446 , \30460 );
and \U$41070 ( \41448 , \41442 , \41447 );
and \U$41071 ( \41449 , \41438 , \41447 );
or \U$41072 ( \41450 , \41443 , \41448 , \41449 );
and \U$41073 ( \41451 , \29715 , \28575 );
and \U$41074 ( \41452 , \29710 , \28573 );
nor \U$41075 ( \41453 , \41451 , \41452 );
xnor \U$41076 ( \41454 , \41453 , \28315 );
and \U$41077 ( \41455 , \30318 , \28081 );
and \U$41078 ( \41456 , \30034 , \28079 );
nor \U$41079 ( \41457 , \41455 , \41456 );
xnor \U$41080 ( \41458 , \41457 , \27766 );
and \U$41081 ( \41459 , \41454 , \41458 );
and \U$41082 ( \41460 , \30895 , \27572 );
and \U$41083 ( \41461 , \30887 , \27570 );
nor \U$41084 ( \41462 , \41460 , \41461 );
xnor \U$41085 ( \41463 , \41462 , \27232 );
and \U$41086 ( \41464 , \41458 , \41463 );
and \U$41087 ( \41465 , \41454 , \41463 );
or \U$41088 ( \41466 , \41459 , \41464 , \41465 );
and \U$41089 ( \41467 , \41450 , \41466 );
and \U$41090 ( \41468 , \28039 , \30233 );
and \U$41091 ( \41469 , \27837 , \30231 );
nor \U$41092 ( \41470 , \41468 , \41469 );
xnor \U$41093 ( \41471 , \41470 , \29862 );
and \U$41094 ( \41472 , \28514 , \29671 );
and \U$41095 ( \41473 , \28342 , \29669 );
nor \U$41096 ( \41474 , \41472 , \41473 );
xnor \U$41097 ( \41475 , \41474 , \29353 );
and \U$41098 ( \41476 , \41471 , \41475 );
and \U$41099 ( \41477 , \29464 , \29104 );
and \U$41100 ( \41478 , \29040 , \29102 );
nor \U$41101 ( \41479 , \41477 , \41478 );
xnor \U$41102 ( \41480 , \41479 , \28855 );
and \U$41103 ( \41481 , \41475 , \41480 );
and \U$41104 ( \41482 , \41471 , \41480 );
or \U$41105 ( \41483 , \41476 , \41481 , \41482 );
and \U$41106 ( \41484 , \41466 , \41483 );
and \U$41107 ( \41485 , \41450 , \41483 );
or \U$41108 ( \41486 , \41467 , \41484 , \41485 );
nand \U$41109 ( \41487 , \32304 , \26141 );
xnor \U$41110 ( \41488 , \41487 , \25911 );
xor \U$41111 ( \41489 , \41332 , \41336 );
xor \U$41112 ( \41490 , \41489 , \41341 );
and \U$41113 ( \41491 , \41488 , \41490 );
xor \U$41114 ( \41492 , \41364 , \41368 );
xor \U$41115 ( \41493 , \41492 , \41373 );
and \U$41116 ( \41494 , \41490 , \41493 );
and \U$41117 ( \41495 , \41488 , \41493 );
or \U$41118 ( \41496 , \41491 , \41494 , \41495 );
and \U$41119 ( \41497 , \41486 , \41496 );
xor \U$41120 ( \41498 , \41316 , \41320 );
xor \U$41121 ( \41499 , \41498 , \41325 );
xor \U$41122 ( \41500 , \41349 , \41353 );
xor \U$41123 ( \41501 , \41500 , \25911 );
and \U$41124 ( \41502 , \41499 , \41501 );
and \U$41125 ( \41503 , \41496 , \41502 );
and \U$41126 ( \41504 , \41486 , \41502 );
or \U$41127 ( \41505 , \41497 , \41503 , \41504 );
xor \U$41128 ( \41506 , \41328 , \41344 );
xor \U$41129 ( \41507 , \41506 , \41357 );
xor \U$41130 ( \41508 , \41376 , \41378 );
xor \U$41131 ( \41509 , \41508 , \41381 );
and \U$41132 ( \41510 , \41507 , \41509 );
xor \U$41133 ( \41511 , \41387 , \41389 );
and \U$41134 ( \41512 , \41509 , \41511 );
and \U$41135 ( \41513 , \41507 , \41511 );
or \U$41136 ( \41514 , \41510 , \41512 , \41513 );
and \U$41137 ( \41515 , \41505 , \41514 );
xor \U$41138 ( \41516 , \41395 , \41397 );
xor \U$41139 ( \41517 , \41516 , \41400 );
and \U$41140 ( \41518 , \41514 , \41517 );
and \U$41141 ( \41519 , \41505 , \41517 );
or \U$41142 ( \41520 , \41515 , \41518 , \41519 );
xor \U$41143 ( \41521 , \41393 , \41403 );
xor \U$41144 ( \41522 , \41521 , \41406 );
and \U$41145 ( \41523 , \41520 , \41522 );
xor \U$41146 ( \41524 , \41411 , \41413 );
and \U$41147 ( \41525 , \41522 , \41524 );
and \U$41148 ( \41526 , \41520 , \41524 );
or \U$41149 ( \41527 , \41523 , \41525 , \41526 );
and \U$41150 ( \41528 , \41434 , \41527 );
xor \U$41151 ( \41529 , \41434 , \41527 );
xor \U$41152 ( \41530 , \41520 , \41522 );
xor \U$41153 ( \41531 , \41530 , \41524 );
and \U$41154 ( \41532 , \31498 , \27572 );
and \U$41155 ( \41533 , \30895 , \27570 );
nor \U$41156 ( \41534 , \41532 , \41533 );
xnor \U$41157 ( \41535 , \41534 , \27232 );
and \U$41158 ( \41536 , \31684 , \26983 );
and \U$41159 ( \41537 , \31503 , \26981 );
nor \U$41160 ( \41538 , \41536 , \41537 );
xnor \U$41161 ( \41539 , \41538 , \26742 );
and \U$41162 ( \41540 , \41535 , \41539 );
nand \U$41163 ( \41541 , \32304 , \26515 );
xnor \U$41164 ( \41542 , \41541 , \26329 );
and \U$41165 ( \41543 , \41539 , \41542 );
and \U$41166 ( \41544 , \41535 , \41542 );
or \U$41167 ( \41545 , \41540 , \41543 , \41544 );
and \U$41168 ( \41546 , \31503 , \26983 );
and \U$41169 ( \41547 , \31498 , \26981 );
nor \U$41170 ( \41548 , \41546 , \41547 );
xnor \U$41171 ( \41549 , \41548 , \26742 );
and \U$41172 ( \41550 , \41545 , \41549 );
and \U$41173 ( \41551 , \32304 , \26517 );
and \U$41174 ( \41552 , \31684 , \26515 );
nor \U$41175 ( \41553 , \41551 , \41552 );
xnor \U$41176 ( \41554 , \41553 , \26329 );
and \U$41177 ( \41555 , \41549 , \41554 );
and \U$41178 ( \41556 , \41545 , \41554 );
or \U$41179 ( \41557 , \41550 , \41555 , \41556 );
and \U$41180 ( \41558 , \26854 , \32151 );
and \U$41181 ( \41559 , \26590 , \32148 );
nor \U$41182 ( \41560 , \41558 , \41559 );
xnor \U$41183 ( \41561 , \41560 , \31096 );
and \U$41184 ( \41562 , \27485 , \31338 );
and \U$41185 ( \41563 , \27113 , \31336 );
nor \U$41186 ( \41564 , \41562 , \41563 );
xnor \U$41187 ( \41565 , \41564 , \31099 );
and \U$41188 ( \41566 , \41561 , \41565 );
and \U$41189 ( \41567 , \41565 , \26329 );
and \U$41190 ( \41568 , \41561 , \26329 );
or \U$41191 ( \41569 , \41566 , \41567 , \41568 );
and \U$41192 ( \41570 , \27837 , \30770 );
and \U$41193 ( \41571 , \27494 , \30768 );
nor \U$41194 ( \41572 , \41570 , \41571 );
xnor \U$41195 ( \41573 , \41572 , \30460 );
and \U$41196 ( \41574 , \28342 , \30233 );
and \U$41197 ( \41575 , \28039 , \30231 );
nor \U$41198 ( \41576 , \41574 , \41575 );
xnor \U$41199 ( \41577 , \41576 , \29862 );
and \U$41200 ( \41578 , \41573 , \41577 );
and \U$41201 ( \41579 , \29040 , \29671 );
and \U$41202 ( \41580 , \28514 , \29669 );
nor \U$41203 ( \41581 , \41579 , \41580 );
xnor \U$41204 ( \41582 , \41581 , \29353 );
and \U$41205 ( \41583 , \41577 , \41582 );
and \U$41206 ( \41584 , \41573 , \41582 );
or \U$41207 ( \41585 , \41578 , \41583 , \41584 );
and \U$41208 ( \41586 , \41569 , \41585 );
and \U$41209 ( \41587 , \29710 , \29104 );
and \U$41210 ( \41588 , \29464 , \29102 );
nor \U$41211 ( \41589 , \41587 , \41588 );
xnor \U$41212 ( \41590 , \41589 , \28855 );
and \U$41213 ( \41591 , \30034 , \28575 );
and \U$41214 ( \41592 , \29715 , \28573 );
nor \U$41215 ( \41593 , \41591 , \41592 );
xnor \U$41216 ( \41594 , \41593 , \28315 );
and \U$41217 ( \41595 , \41590 , \41594 );
and \U$41218 ( \41596 , \30887 , \28081 );
and \U$41219 ( \41597 , \30318 , \28079 );
nor \U$41220 ( \41598 , \41596 , \41597 );
xnor \U$41221 ( \41599 , \41598 , \27766 );
and \U$41222 ( \41600 , \41594 , \41599 );
and \U$41223 ( \41601 , \41590 , \41599 );
or \U$41224 ( \41602 , \41595 , \41600 , \41601 );
and \U$41225 ( \41603 , \41585 , \41602 );
and \U$41226 ( \41604 , \41569 , \41602 );
or \U$41227 ( \41605 , \41586 , \41603 , \41604 );
and \U$41228 ( \41606 , \41557 , \41605 );
xor \U$41229 ( \41607 , \41438 , \41442 );
xor \U$41230 ( \41608 , \41607 , \41447 );
xor \U$41231 ( \41609 , \41454 , \41458 );
xor \U$41232 ( \41610 , \41609 , \41463 );
and \U$41233 ( \41611 , \41608 , \41610 );
xor \U$41234 ( \41612 , \41471 , \41475 );
xor \U$41235 ( \41613 , \41612 , \41480 );
and \U$41236 ( \41614 , \41610 , \41613 );
and \U$41237 ( \41615 , \41608 , \41613 );
or \U$41238 ( \41616 , \41611 , \41614 , \41615 );
and \U$41239 ( \41617 , \41605 , \41616 );
and \U$41240 ( \41618 , \41557 , \41616 );
or \U$41241 ( \41619 , \41606 , \41617 , \41618 );
xor \U$41242 ( \41620 , \41450 , \41466 );
xor \U$41243 ( \41621 , \41620 , \41483 );
xor \U$41244 ( \41622 , \41488 , \41490 );
xor \U$41245 ( \41623 , \41622 , \41493 );
and \U$41246 ( \41624 , \41621 , \41623 );
xor \U$41247 ( \41625 , \41499 , \41501 );
and \U$41248 ( \41626 , \41623 , \41625 );
and \U$41249 ( \41627 , \41621 , \41625 );
or \U$41250 ( \41628 , \41624 , \41626 , \41627 );
and \U$41251 ( \41629 , \41619 , \41628 );
xor \U$41252 ( \41630 , \41507 , \41509 );
xor \U$41253 ( \41631 , \41630 , \41511 );
and \U$41254 ( \41632 , \41628 , \41631 );
and \U$41255 ( \41633 , \41619 , \41631 );
or \U$41256 ( \41634 , \41629 , \41632 , \41633 );
xor \U$41257 ( \41635 , \41360 , \41384 );
xor \U$41258 ( \41636 , \41635 , \41390 );
and \U$41259 ( \41637 , \41634 , \41636 );
xor \U$41260 ( \41638 , \41505 , \41514 );
xor \U$41261 ( \41639 , \41638 , \41517 );
and \U$41262 ( \41640 , \41636 , \41639 );
and \U$41263 ( \41641 , \41634 , \41639 );
or \U$41264 ( \41642 , \41637 , \41640 , \41641 );
and \U$41265 ( \41643 , \41531 , \41642 );
xor \U$41266 ( \41644 , \41531 , \41642 );
xor \U$41267 ( \41645 , \41634 , \41636 );
xor \U$41268 ( \41646 , \41645 , \41639 );
and \U$41269 ( \41647 , \30318 , \28575 );
and \U$41270 ( \41648 , \30034 , \28573 );
nor \U$41271 ( \41649 , \41647 , \41648 );
xnor \U$41272 ( \41650 , \41649 , \28315 );
and \U$41273 ( \41651 , \30895 , \28081 );
and \U$41274 ( \41652 , \30887 , \28079 );
nor \U$41275 ( \41653 , \41651 , \41652 );
xnor \U$41276 ( \41654 , \41653 , \27766 );
and \U$41277 ( \41655 , \41650 , \41654 );
and \U$41278 ( \41656 , \31503 , \27572 );
and \U$41279 ( \41657 , \31498 , \27570 );
nor \U$41280 ( \41658 , \41656 , \41657 );
xnor \U$41281 ( \41659 , \41658 , \27232 );
and \U$41282 ( \41660 , \41654 , \41659 );
and \U$41283 ( \41661 , \41650 , \41659 );
or \U$41284 ( \41662 , \41655 , \41660 , \41661 );
and \U$41285 ( \41663 , \27113 , \32151 );
and \U$41286 ( \41664 , \26854 , \32148 );
nor \U$41287 ( \41665 , \41663 , \41664 );
xnor \U$41288 ( \41666 , \41665 , \31096 );
and \U$41289 ( \41667 , \27494 , \31338 );
and \U$41290 ( \41668 , \27485 , \31336 );
nor \U$41291 ( \41669 , \41667 , \41668 );
xnor \U$41292 ( \41670 , \41669 , \31099 );
and \U$41293 ( \41671 , \41666 , \41670 );
and \U$41294 ( \41672 , \28039 , \30770 );
and \U$41295 ( \41673 , \27837 , \30768 );
nor \U$41296 ( \41674 , \41672 , \41673 );
xnor \U$41297 ( \41675 , \41674 , \30460 );
and \U$41298 ( \41676 , \41670 , \41675 );
and \U$41299 ( \41677 , \41666 , \41675 );
or \U$41300 ( \41678 , \41671 , \41676 , \41677 );
and \U$41301 ( \41679 , \41662 , \41678 );
and \U$41302 ( \41680 , \28514 , \30233 );
and \U$41303 ( \41681 , \28342 , \30231 );
nor \U$41304 ( \41682 , \41680 , \41681 );
xnor \U$41305 ( \41683 , \41682 , \29862 );
and \U$41306 ( \41684 , \29464 , \29671 );
and \U$41307 ( \41685 , \29040 , \29669 );
nor \U$41308 ( \41686 , \41684 , \41685 );
xnor \U$41309 ( \41687 , \41686 , \29353 );
and \U$41310 ( \41688 , \41683 , \41687 );
and \U$41311 ( \41689 , \29715 , \29104 );
and \U$41312 ( \41690 , \29710 , \29102 );
nor \U$41313 ( \41691 , \41689 , \41690 );
xnor \U$41314 ( \41692 , \41691 , \28855 );
and \U$41315 ( \41693 , \41687 , \41692 );
and \U$41316 ( \41694 , \41683 , \41692 );
or \U$41317 ( \41695 , \41688 , \41693 , \41694 );
and \U$41318 ( \41696 , \41678 , \41695 );
and \U$41319 ( \41697 , \41662 , \41695 );
or \U$41320 ( \41698 , \41679 , \41696 , \41697 );
xor \U$41321 ( \41699 , \41573 , \41577 );
xor \U$41322 ( \41700 , \41699 , \41582 );
xor \U$41323 ( \41701 , \41535 , \41539 );
xor \U$41324 ( \41702 , \41701 , \41542 );
and \U$41325 ( \41703 , \41700 , \41702 );
xor \U$41326 ( \41704 , \41590 , \41594 );
xor \U$41327 ( \41705 , \41704 , \41599 );
and \U$41328 ( \41706 , \41702 , \41705 );
and \U$41329 ( \41707 , \41700 , \41705 );
or \U$41330 ( \41708 , \41703 , \41706 , \41707 );
and \U$41331 ( \41709 , \41698 , \41708 );
xor \U$41332 ( \41710 , \41608 , \41610 );
xor \U$41333 ( \41711 , \41710 , \41613 );
and \U$41334 ( \41712 , \41708 , \41711 );
and \U$41335 ( \41713 , \41698 , \41711 );
or \U$41336 ( \41714 , \41709 , \41712 , \41713 );
xor \U$41337 ( \41715 , \41557 , \41605 );
xor \U$41338 ( \41716 , \41715 , \41616 );
and \U$41339 ( \41717 , \41714 , \41716 );
xor \U$41340 ( \41718 , \41621 , \41623 );
xor \U$41341 ( \41719 , \41718 , \41625 );
and \U$41342 ( \41720 , \41716 , \41719 );
and \U$41343 ( \41721 , \41714 , \41719 );
or \U$41344 ( \41722 , \41717 , \41720 , \41721 );
xor \U$41345 ( \41723 , \41486 , \41496 );
xor \U$41346 ( \41724 , \41723 , \41502 );
and \U$41347 ( \41725 , \41722 , \41724 );
xor \U$41348 ( \41726 , \41619 , \41628 );
xor \U$41349 ( \41727 , \41726 , \41631 );
and \U$41350 ( \41728 , \41724 , \41727 );
and \U$41351 ( \41729 , \41722 , \41727 );
or \U$41352 ( \41730 , \41725 , \41728 , \41729 );
and \U$41353 ( \41731 , \41646 , \41730 );
xor \U$41354 ( \41732 , \41646 , \41730 );
xor \U$41355 ( \41733 , \41722 , \41724 );
xor \U$41356 ( \41734 , \41733 , \41727 );
and \U$41357 ( \41735 , \27485 , \32151 );
and \U$41358 ( \41736 , \27113 , \32148 );
nor \U$41359 ( \41737 , \41735 , \41736 );
xnor \U$41360 ( \41738 , \41737 , \31096 );
and \U$41361 ( \41739 , \27837 , \31338 );
and \U$41362 ( \41740 , \27494 , \31336 );
nor \U$41363 ( \41741 , \41739 , \41740 );
xnor \U$41364 ( \41742 , \41741 , \31099 );
and \U$41365 ( \41743 , \41738 , \41742 );
and \U$41366 ( \41744 , \41742 , \26742 );
and \U$41367 ( \41745 , \41738 , \26742 );
or \U$41368 ( \41746 , \41743 , \41744 , \41745 );
and \U$41369 ( \41747 , \30034 , \29104 );
and \U$41370 ( \41748 , \29715 , \29102 );
nor \U$41371 ( \41749 , \41747 , \41748 );
xnor \U$41372 ( \41750 , \41749 , \28855 );
and \U$41373 ( \41751 , \30887 , \28575 );
and \U$41374 ( \41752 , \30318 , \28573 );
nor \U$41375 ( \41753 , \41751 , \41752 );
xnor \U$41376 ( \41754 , \41753 , \28315 );
and \U$41377 ( \41755 , \41750 , \41754 );
and \U$41378 ( \41756 , \31498 , \28081 );
and \U$41379 ( \41757 , \30895 , \28079 );
nor \U$41380 ( \41758 , \41756 , \41757 );
xnor \U$41381 ( \41759 , \41758 , \27766 );
and \U$41382 ( \41760 , \41754 , \41759 );
and \U$41383 ( \41761 , \41750 , \41759 );
or \U$41384 ( \41762 , \41755 , \41760 , \41761 );
and \U$41385 ( \41763 , \41746 , \41762 );
and \U$41386 ( \41764 , \28342 , \30770 );
and \U$41387 ( \41765 , \28039 , \30768 );
nor \U$41388 ( \41766 , \41764 , \41765 );
xnor \U$41389 ( \41767 , \41766 , \30460 );
and \U$41390 ( \41768 , \29040 , \30233 );
and \U$41391 ( \41769 , \28514 , \30231 );
nor \U$41392 ( \41770 , \41768 , \41769 );
xnor \U$41393 ( \41771 , \41770 , \29862 );
and \U$41394 ( \41772 , \41767 , \41771 );
and \U$41395 ( \41773 , \29710 , \29671 );
and \U$41396 ( \41774 , \29464 , \29669 );
nor \U$41397 ( \41775 , \41773 , \41774 );
xnor \U$41398 ( \41776 , \41775 , \29353 );
and \U$41399 ( \41777 , \41771 , \41776 );
and \U$41400 ( \41778 , \41767 , \41776 );
or \U$41401 ( \41779 , \41772 , \41777 , \41778 );
and \U$41402 ( \41780 , \41762 , \41779 );
and \U$41403 ( \41781 , \41746 , \41779 );
or \U$41404 ( \41782 , \41763 , \41780 , \41781 );
and \U$41405 ( \41783 , \32304 , \26983 );
and \U$41406 ( \41784 , \31684 , \26981 );
nor \U$41407 ( \41785 , \41783 , \41784 );
xnor \U$41408 ( \41786 , \41785 , \26742 );
xor \U$41409 ( \41787 , \41650 , \41654 );
xor \U$41410 ( \41788 , \41787 , \41659 );
and \U$41411 ( \41789 , \41786 , \41788 );
xor \U$41412 ( \41790 , \41683 , \41687 );
xor \U$41413 ( \41791 , \41790 , \41692 );
and \U$41414 ( \41792 , \41788 , \41791 );
and \U$41415 ( \41793 , \41786 , \41791 );
or \U$41416 ( \41794 , \41789 , \41792 , \41793 );
and \U$41417 ( \41795 , \41782 , \41794 );
xor \U$41418 ( \41796 , \41561 , \41565 );
xor \U$41419 ( \41797 , \41796 , \26329 );
and \U$41420 ( \41798 , \41794 , \41797 );
and \U$41421 ( \41799 , \41782 , \41797 );
or \U$41422 ( \41800 , \41795 , \41798 , \41799 );
xor \U$41423 ( \41801 , \41662 , \41678 );
xor \U$41424 ( \41802 , \41801 , \41695 );
xor \U$41425 ( \41803 , \41700 , \41702 );
xor \U$41426 ( \41804 , \41803 , \41705 );
and \U$41427 ( \41805 , \41802 , \41804 );
and \U$41428 ( \41806 , \41800 , \41805 );
xor \U$41429 ( \41807 , \41545 , \41549 );
xor \U$41430 ( \41808 , \41807 , \41554 );
and \U$41431 ( \41809 , \41805 , \41808 );
and \U$41432 ( \41810 , \41800 , \41808 );
or \U$41433 ( \41811 , \41806 , \41809 , \41810 );
xor \U$41434 ( \41812 , \41569 , \41585 );
xor \U$41435 ( \41813 , \41812 , \41602 );
xor \U$41436 ( \41814 , \41698 , \41708 );
xor \U$41437 ( \41815 , \41814 , \41711 );
and \U$41438 ( \41816 , \41813 , \41815 );
and \U$41439 ( \41817 , \41811 , \41816 );
xor \U$41440 ( \41818 , \41714 , \41716 );
xor \U$41441 ( \41819 , \41818 , \41719 );
and \U$41442 ( \41820 , \41816 , \41819 );
and \U$41443 ( \41821 , \41811 , \41819 );
or \U$41444 ( \41822 , \41817 , \41820 , \41821 );
and \U$41445 ( \41823 , \41734 , \41822 );
xor \U$41446 ( \41824 , \41734 , \41822 );
xor \U$41447 ( \41825 , \41811 , \41816 );
xor \U$41448 ( \41826 , \41825 , \41819 );
and \U$41449 ( \41827 , \29464 , \30233 );
and \U$41450 ( \41828 , \29040 , \30231 );
nor \U$41451 ( \41829 , \41827 , \41828 );
xnor \U$41452 ( \41830 , \41829 , \29862 );
and \U$41453 ( \41831 , \29715 , \29671 );
and \U$41454 ( \41832 , \29710 , \29669 );
nor \U$41455 ( \41833 , \41831 , \41832 );
xnor \U$41456 ( \41834 , \41833 , \29353 );
and \U$41457 ( \41835 , \41830 , \41834 );
and \U$41458 ( \41836 , \30318 , \29104 );
and \U$41459 ( \41837 , \30034 , \29102 );
nor \U$41460 ( \41838 , \41836 , \41837 );
xnor \U$41461 ( \41839 , \41838 , \28855 );
and \U$41462 ( \41840 , \41834 , \41839 );
and \U$41463 ( \41841 , \41830 , \41839 );
or \U$41464 ( \41842 , \41835 , \41840 , \41841 );
and \U$41465 ( \41843 , \27494 , \32151 );
and \U$41466 ( \41844 , \27485 , \32148 );
nor \U$41467 ( \41845 , \41843 , \41844 );
xnor \U$41468 ( \41846 , \41845 , \31096 );
and \U$41469 ( \41847 , \28039 , \31338 );
and \U$41470 ( \41848 , \27837 , \31336 );
nor \U$41471 ( \41849 , \41847 , \41848 );
xnor \U$41472 ( \41850 , \41849 , \31099 );
and \U$41473 ( \41851 , \41846 , \41850 );
and \U$41474 ( \41852 , \28514 , \30770 );
and \U$41475 ( \41853 , \28342 , \30768 );
nor \U$41476 ( \41854 , \41852 , \41853 );
xnor \U$41477 ( \41855 , \41854 , \30460 );
and \U$41478 ( \41856 , \41850 , \41855 );
and \U$41479 ( \41857 , \41846 , \41855 );
or \U$41480 ( \41858 , \41851 , \41856 , \41857 );
and \U$41481 ( \41859 , \41842 , \41858 );
and \U$41482 ( \41860 , \30895 , \28575 );
and \U$41483 ( \41861 , \30887 , \28573 );
nor \U$41484 ( \41862 , \41860 , \41861 );
xnor \U$41485 ( \41863 , \41862 , \28315 );
and \U$41486 ( \41864 , \31503 , \28081 );
and \U$41487 ( \41865 , \31498 , \28079 );
nor \U$41488 ( \41866 , \41864 , \41865 );
xnor \U$41489 ( \41867 , \41866 , \27766 );
and \U$41490 ( \41868 , \41863 , \41867 );
and \U$41491 ( \41869 , \32304 , \27572 );
and \U$41492 ( \41870 , \31684 , \27570 );
nor \U$41493 ( \41871 , \41869 , \41870 );
xnor \U$41494 ( \41872 , \41871 , \27232 );
and \U$41495 ( \41873 , \41867 , \41872 );
and \U$41496 ( \41874 , \41863 , \41872 );
or \U$41497 ( \41875 , \41868 , \41873 , \41874 );
and \U$41498 ( \41876 , \41858 , \41875 );
and \U$41499 ( \41877 , \41842 , \41875 );
or \U$41500 ( \41878 , \41859 , \41876 , \41877 );
and \U$41501 ( \41879 , \31684 , \27572 );
and \U$41502 ( \41880 , \31503 , \27570 );
nor \U$41503 ( \41881 , \41879 , \41880 );
xnor \U$41504 ( \41882 , \41881 , \27232 );
nand \U$41505 ( \41883 , \32304 , \26981 );
xnor \U$41506 ( \41884 , \41883 , \26742 );
and \U$41507 ( \41885 , \41882 , \41884 );
xor \U$41508 ( \41886 , \41750 , \41754 );
xor \U$41509 ( \41887 , \41886 , \41759 );
and \U$41510 ( \41888 , \41884 , \41887 );
and \U$41511 ( \41889 , \41882 , \41887 );
or \U$41512 ( \41890 , \41885 , \41888 , \41889 );
and \U$41513 ( \41891 , \41878 , \41890 );
xor \U$41514 ( \41892 , \41666 , \41670 );
xor \U$41515 ( \41893 , \41892 , \41675 );
and \U$41516 ( \41894 , \41890 , \41893 );
and \U$41517 ( \41895 , \41878 , \41893 );
or \U$41518 ( \41896 , \41891 , \41894 , \41895 );
xor \U$41519 ( \41897 , \41782 , \41794 );
xor \U$41520 ( \41898 , \41897 , \41797 );
and \U$41521 ( \41899 , \41896 , \41898 );
xor \U$41522 ( \41900 , \41802 , \41804 );
and \U$41523 ( \41901 , \41898 , \41900 );
and \U$41524 ( \41902 , \41896 , \41900 );
or \U$41525 ( \41903 , \41899 , \41901 , \41902 );
xor \U$41526 ( \41904 , \41800 , \41805 );
xor \U$41527 ( \41905 , \41904 , \41808 );
and \U$41528 ( \41906 , \41903 , \41905 );
xor \U$41529 ( \41907 , \41813 , \41815 );
and \U$41530 ( \41908 , \41905 , \41907 );
and \U$41531 ( \41909 , \41903 , \41907 );
or \U$41532 ( \41910 , \41906 , \41908 , \41909 );
and \U$41533 ( \41911 , \41826 , \41910 );
xor \U$41534 ( \41912 , \41826 , \41910 );
xor \U$41535 ( \41913 , \41903 , \41905 );
xor \U$41536 ( \41914 , \41913 , \41907 );
and \U$41537 ( \41915 , \29040 , \30770 );
and \U$41538 ( \41916 , \28514 , \30768 );
nor \U$41539 ( \41917 , \41915 , \41916 );
xnor \U$41540 ( \41918 , \41917 , \30460 );
and \U$41541 ( \41919 , \29710 , \30233 );
and \U$41542 ( \41920 , \29464 , \30231 );
nor \U$41543 ( \41921 , \41919 , \41920 );
xnor \U$41544 ( \41922 , \41921 , \29862 );
and \U$41545 ( \41923 , \41918 , \41922 );
and \U$41546 ( \41924 , \30034 , \29671 );
and \U$41547 ( \41925 , \29715 , \29669 );
nor \U$41548 ( \41926 , \41924 , \41925 );
xnor \U$41549 ( \41927 , \41926 , \29353 );
and \U$41550 ( \41928 , \41922 , \41927 );
and \U$41551 ( \41929 , \41918 , \41927 );
or \U$41552 ( \41930 , \41923 , \41928 , \41929 );
and \U$41553 ( \41931 , \27837 , \32151 );
and \U$41554 ( \41932 , \27494 , \32148 );
nor \U$41555 ( \41933 , \41931 , \41932 );
xnor \U$41556 ( \41934 , \41933 , \31096 );
and \U$41557 ( \41935 , \28342 , \31338 );
and \U$41558 ( \41936 , \28039 , \31336 );
nor \U$41559 ( \41937 , \41935 , \41936 );
xnor \U$41560 ( \41938 , \41937 , \31099 );
and \U$41561 ( \41939 , \41934 , \41938 );
and \U$41562 ( \41940 , \41938 , \27232 );
and \U$41563 ( \41941 , \41934 , \27232 );
or \U$41564 ( \41942 , \41939 , \41940 , \41941 );
and \U$41565 ( \41943 , \41930 , \41942 );
and \U$41566 ( \41944 , \30887 , \29104 );
and \U$41567 ( \41945 , \30318 , \29102 );
nor \U$41568 ( \41946 , \41944 , \41945 );
xnor \U$41569 ( \41947 , \41946 , \28855 );
and \U$41570 ( \41948 , \31498 , \28575 );
and \U$41571 ( \41949 , \30895 , \28573 );
nor \U$41572 ( \41950 , \41948 , \41949 );
xnor \U$41573 ( \41951 , \41950 , \28315 );
and \U$41574 ( \41952 , \41947 , \41951 );
and \U$41575 ( \41953 , \31684 , \28081 );
and \U$41576 ( \41954 , \31503 , \28079 );
nor \U$41577 ( \41955 , \41953 , \41954 );
xnor \U$41578 ( \41956 , \41955 , \27766 );
and \U$41579 ( \41957 , \41951 , \41956 );
and \U$41580 ( \41958 , \41947 , \41956 );
or \U$41581 ( \41959 , \41952 , \41957 , \41958 );
and \U$41582 ( \41960 , \41942 , \41959 );
and \U$41583 ( \41961 , \41930 , \41959 );
or \U$41584 ( \41962 , \41943 , \41960 , \41961 );
xor \U$41585 ( \41963 , \41830 , \41834 );
xor \U$41586 ( \41964 , \41963 , \41839 );
xor \U$41587 ( \41965 , \41846 , \41850 );
xor \U$41588 ( \41966 , \41965 , \41855 );
and \U$41589 ( \41967 , \41964 , \41966 );
xor \U$41590 ( \41968 , \41863 , \41867 );
xor \U$41591 ( \41969 , \41968 , \41872 );
and \U$41592 ( \41970 , \41966 , \41969 );
and \U$41593 ( \41971 , \41964 , \41969 );
or \U$41594 ( \41972 , \41967 , \41970 , \41971 );
and \U$41595 ( \41973 , \41962 , \41972 );
xor \U$41596 ( \41974 , \41767 , \41771 );
xor \U$41597 ( \41975 , \41974 , \41776 );
and \U$41598 ( \41976 , \41972 , \41975 );
and \U$41599 ( \41977 , \41962 , \41975 );
or \U$41600 ( \41978 , \41973 , \41976 , \41977 );
xor \U$41601 ( \41979 , \41738 , \41742 );
xor \U$41602 ( \41980 , \41979 , \26742 );
xor \U$41603 ( \41981 , \41842 , \41858 );
xor \U$41604 ( \41982 , \41981 , \41875 );
and \U$41605 ( \41983 , \41980 , \41982 );
xor \U$41606 ( \41984 , \41882 , \41884 );
xor \U$41607 ( \41985 , \41984 , \41887 );
and \U$41608 ( \41986 , \41982 , \41985 );
and \U$41609 ( \41987 , \41980 , \41985 );
or \U$41610 ( \41988 , \41983 , \41986 , \41987 );
and \U$41611 ( \41989 , \41978 , \41988 );
xor \U$41612 ( \41990 , \41786 , \41788 );
xor \U$41613 ( \41991 , \41990 , \41791 );
and \U$41614 ( \41992 , \41988 , \41991 );
and \U$41615 ( \41993 , \41978 , \41991 );
or \U$41616 ( \41994 , \41989 , \41992 , \41993 );
xor \U$41617 ( \41995 , \41746 , \41762 );
xor \U$41618 ( \41996 , \41995 , \41779 );
xor \U$41619 ( \41997 , \41878 , \41890 );
xor \U$41620 ( \41998 , \41997 , \41893 );
and \U$41621 ( \41999 , \41996 , \41998 );
and \U$41622 ( \42000 , \41994 , \41999 );
xor \U$41623 ( \42001 , \41896 , \41898 );
xor \U$41624 ( \42002 , \42001 , \41900 );
and \U$41625 ( \42003 , \41999 , \42002 );
and \U$41626 ( \42004 , \41994 , \42002 );
or \U$41627 ( \42005 , \42000 , \42003 , \42004 );
and \U$41628 ( \42006 , \41914 , \42005 );
xor \U$41629 ( \42007 , \41914 , \42005 );
xor \U$41630 ( \42008 , \41994 , \41999 );
xor \U$41631 ( \42009 , \42008 , \42002 );
and \U$41632 ( \42010 , \28039 , \32151 );
and \U$41633 ( \42011 , \27837 , \32148 );
nor \U$41634 ( \42012 , \42010 , \42011 );
xnor \U$41635 ( \42013 , \42012 , \31096 );
and \U$41636 ( \42014 , \28514 , \31338 );
and \U$41637 ( \42015 , \28342 , \31336 );
nor \U$41638 ( \42016 , \42014 , \42015 );
xnor \U$41639 ( \42017 , \42016 , \31099 );
and \U$41640 ( \42018 , \42013 , \42017 );
and \U$41641 ( \42019 , \29464 , \30770 );
and \U$41642 ( \42020 , \29040 , \30768 );
nor \U$41643 ( \42021 , \42019 , \42020 );
xnor \U$41644 ( \42022 , \42021 , \30460 );
and \U$41645 ( \42023 , \42017 , \42022 );
and \U$41646 ( \42024 , \42013 , \42022 );
or \U$41647 ( \42025 , \42018 , \42023 , \42024 );
and \U$41648 ( \42026 , \29715 , \30233 );
and \U$41649 ( \42027 , \29710 , \30231 );
nor \U$41650 ( \42028 , \42026 , \42027 );
xnor \U$41651 ( \42029 , \42028 , \29862 );
and \U$41652 ( \42030 , \30318 , \29671 );
and \U$41653 ( \42031 , \30034 , \29669 );
nor \U$41654 ( \42032 , \42030 , \42031 );
xnor \U$41655 ( \42033 , \42032 , \29353 );
and \U$41656 ( \42034 , \42029 , \42033 );
and \U$41657 ( \42035 , \30895 , \29104 );
and \U$41658 ( \42036 , \30887 , \29102 );
nor \U$41659 ( \42037 , \42035 , \42036 );
xnor \U$41660 ( \42038 , \42037 , \28855 );
and \U$41661 ( \42039 , \42033 , \42038 );
and \U$41662 ( \42040 , \42029 , \42038 );
or \U$41663 ( \42041 , \42034 , \42039 , \42040 );
and \U$41664 ( \42042 , \42025 , \42041 );
and \U$41665 ( \42043 , \31503 , \28575 );
and \U$41666 ( \42044 , \31498 , \28573 );
nor \U$41667 ( \42045 , \42043 , \42044 );
xnor \U$41668 ( \42046 , \42045 , \28315 );
and \U$41669 ( \42047 , \32304 , \28081 );
and \U$41670 ( \42048 , \31684 , \28079 );
nor \U$41671 ( \42049 , \42047 , \42048 );
xnor \U$41672 ( \42050 , \42049 , \27766 );
and \U$41673 ( \42051 , \42046 , \42050 );
and \U$41674 ( \42052 , \42041 , \42051 );
and \U$41675 ( \42053 , \42025 , \42051 );
or \U$41676 ( \42054 , \42042 , \42052 , \42053 );
nand \U$41677 ( \42055 , \32304 , \27570 );
xnor \U$41678 ( \42056 , \42055 , \27232 );
xor \U$41679 ( \42057 , \41918 , \41922 );
xor \U$41680 ( \42058 , \42057 , \41927 );
and \U$41681 ( \42059 , \42056 , \42058 );
xor \U$41682 ( \42060 , \41947 , \41951 );
xor \U$41683 ( \42061 , \42060 , \41956 );
and \U$41684 ( \42062 , \42058 , \42061 );
and \U$41685 ( \42063 , \42056 , \42061 );
or \U$41686 ( \42064 , \42059 , \42062 , \42063 );
and \U$41687 ( \42065 , \42054 , \42064 );
xor \U$41688 ( \42066 , \41964 , \41966 );
xor \U$41689 ( \42067 , \42066 , \41969 );
and \U$41690 ( \42068 , \42064 , \42067 );
and \U$41691 ( \42069 , \42054 , \42067 );
or \U$41692 ( \42070 , \42065 , \42068 , \42069 );
xor \U$41693 ( \42071 , \41962 , \41972 );
xor \U$41694 ( \42072 , \42071 , \41975 );
and \U$41695 ( \42073 , \42070 , \42072 );
xor \U$41696 ( \42074 , \41980 , \41982 );
xor \U$41697 ( \42075 , \42074 , \41985 );
and \U$41698 ( \42076 , \42072 , \42075 );
and \U$41699 ( \42077 , \42070 , \42075 );
or \U$41700 ( \42078 , \42073 , \42076 , \42077 );
xor \U$41701 ( \42079 , \41978 , \41988 );
xor \U$41702 ( \42080 , \42079 , \41991 );
and \U$41703 ( \42081 , \42078 , \42080 );
xor \U$41704 ( \42082 , \41996 , \41998 );
and \U$41705 ( \42083 , \42080 , \42082 );
and \U$41706 ( \42084 , \42078 , \42082 );
or \U$41707 ( \42085 , \42081 , \42083 , \42084 );
and \U$41708 ( \42086 , \42009 , \42085 );
xor \U$41709 ( \42087 , \42009 , \42085 );
xor \U$41710 ( \42088 , \42078 , \42080 );
xor \U$41711 ( \42089 , \42088 , \42082 );
and \U$41712 ( \42090 , \31498 , \29104 );
and \U$41713 ( \42091 , \30895 , \29102 );
nor \U$41714 ( \42092 , \42090 , \42091 );
xnor \U$41715 ( \42093 , \42092 , \28855 );
and \U$41716 ( \42094 , \31684 , \28575 );
and \U$41717 ( \42095 , \31503 , \28573 );
nor \U$41718 ( \42096 , \42094 , \42095 );
xnor \U$41719 ( \42097 , \42096 , \28315 );
and \U$41720 ( \42098 , \42093 , \42097 );
nand \U$41721 ( \42099 , \32304 , \28079 );
xnor \U$41722 ( \42100 , \42099 , \27766 );
and \U$41723 ( \42101 , \42097 , \42100 );
and \U$41724 ( \42102 , \42093 , \42100 );
or \U$41725 ( \42103 , \42098 , \42101 , \42102 );
and \U$41726 ( \42104 , \28342 , \32151 );
and \U$41727 ( \42105 , \28039 , \32148 );
nor \U$41728 ( \42106 , \42104 , \42105 );
xnor \U$41729 ( \42107 , \42106 , \31096 );
and \U$41730 ( \42108 , \29040 , \31338 );
and \U$41731 ( \42109 , \28514 , \31336 );
nor \U$41732 ( \42110 , \42108 , \42109 );
xnor \U$41733 ( \42111 , \42110 , \31099 );
and \U$41734 ( \42112 , \42107 , \42111 );
and \U$41735 ( \42113 , \42111 , \27766 );
and \U$41736 ( \42114 , \42107 , \27766 );
or \U$41737 ( \42115 , \42112 , \42113 , \42114 );
and \U$41738 ( \42116 , \42103 , \42115 );
and \U$41739 ( \42117 , \29710 , \30770 );
and \U$41740 ( \42118 , \29464 , \30768 );
nor \U$41741 ( \42119 , \42117 , \42118 );
xnor \U$41742 ( \42120 , \42119 , \30460 );
and \U$41743 ( \42121 , \30034 , \30233 );
and \U$41744 ( \42122 , \29715 , \30231 );
nor \U$41745 ( \42123 , \42121 , \42122 );
xnor \U$41746 ( \42124 , \42123 , \29862 );
and \U$41747 ( \42125 , \42120 , \42124 );
and \U$41748 ( \42126 , \30887 , \29671 );
and \U$41749 ( \42127 , \30318 , \29669 );
nor \U$41750 ( \42128 , \42126 , \42127 );
xnor \U$41751 ( \42129 , \42128 , \29353 );
and \U$41752 ( \42130 , \42124 , \42129 );
and \U$41753 ( \42131 , \42120 , \42129 );
or \U$41754 ( \42132 , \42125 , \42130 , \42131 );
and \U$41755 ( \42133 , \42115 , \42132 );
and \U$41756 ( \42134 , \42103 , \42132 );
or \U$41757 ( \42135 , \42116 , \42133 , \42134 );
xor \U$41758 ( \42136 , \42013 , \42017 );
xor \U$41759 ( \42137 , \42136 , \42022 );
xor \U$41760 ( \42138 , \42029 , \42033 );
xor \U$41761 ( \42139 , \42138 , \42038 );
and \U$41762 ( \42140 , \42137 , \42139 );
xor \U$41763 ( \42141 , \42046 , \42050 );
and \U$41764 ( \42142 , \42139 , \42141 );
and \U$41765 ( \42143 , \42137 , \42141 );
or \U$41766 ( \42144 , \42140 , \42142 , \42143 );
and \U$41767 ( \42145 , \42135 , \42144 );
xor \U$41768 ( \42146 , \41934 , \41938 );
xor \U$41769 ( \42147 , \42146 , \27232 );
and \U$41770 ( \42148 , \42144 , \42147 );
and \U$41771 ( \42149 , \42135 , \42147 );
or \U$41772 ( \42150 , \42145 , \42148 , \42149 );
xor \U$41773 ( \42151 , \42025 , \42041 );
xor \U$41774 ( \42152 , \42151 , \42051 );
xor \U$41775 ( \42153 , \42056 , \42058 );
xor \U$41776 ( \42154 , \42153 , \42061 );
and \U$41777 ( \42155 , \42152 , \42154 );
and \U$41778 ( \42156 , \42150 , \42155 );
xor \U$41779 ( \42157 , \41930 , \41942 );
xor \U$41780 ( \42158 , \42157 , \41959 );
and \U$41781 ( \42159 , \42155 , \42158 );
and \U$41782 ( \42160 , \42150 , \42158 );
or \U$41783 ( \42161 , \42156 , \42159 , \42160 );
xor \U$41784 ( \42162 , \42070 , \42072 );
xor \U$41785 ( \42163 , \42162 , \42075 );
and \U$41786 ( \42164 , \42161 , \42163 );
and \U$41787 ( \42165 , \42089 , \42164 );
xor \U$41788 ( \42166 , \42089 , \42164 );
xor \U$41789 ( \42167 , \42161 , \42163 );
xor \U$41790 ( \42168 , \42150 , \42155 );
xor \U$41791 ( \42169 , \42168 , \42158 );
xor \U$41792 ( \42170 , \42054 , \42064 );
xor \U$41793 ( \42171 , \42170 , \42067 );
and \U$41794 ( \42172 , \42169 , \42171 );
and \U$41795 ( \42173 , \42167 , \42172 );
xor \U$41796 ( \42174 , \42167 , \42172 );
xor \U$41797 ( \42175 , \42169 , \42171 );
and \U$41798 ( \42176 , \28514 , \32151 );
and \U$41799 ( \42177 , \28342 , \32148 );
nor \U$41800 ( \42178 , \42176 , \42177 );
xnor \U$41801 ( \42179 , \42178 , \31096 );
and \U$41802 ( \42180 , \29464 , \31338 );
and \U$41803 ( \42181 , \29040 , \31336 );
nor \U$41804 ( \42182 , \42180 , \42181 );
xnor \U$41805 ( \42183 , \42182 , \31099 );
and \U$41806 ( \42184 , \42179 , \42183 );
and \U$41807 ( \42185 , \29715 , \30770 );
and \U$41808 ( \42186 , \29710 , \30768 );
nor \U$41809 ( \42187 , \42185 , \42186 );
xnor \U$41810 ( \42188 , \42187 , \30460 );
and \U$41811 ( \42189 , \42183 , \42188 );
and \U$41812 ( \42190 , \42179 , \42188 );
or \U$41813 ( \42191 , \42184 , \42189 , \42190 );
and \U$41814 ( \42192 , \30318 , \30233 );
and \U$41815 ( \42193 , \30034 , \30231 );
nor \U$41816 ( \42194 , \42192 , \42193 );
xnor \U$41817 ( \42195 , \42194 , \29862 );
and \U$41818 ( \42196 , \30895 , \29671 );
and \U$41819 ( \42197 , \30887 , \29669 );
nor \U$41820 ( \42198 , \42196 , \42197 );
xnor \U$41821 ( \42199 , \42198 , \29353 );
and \U$41822 ( \42200 , \42195 , \42199 );
and \U$41823 ( \42201 , \31503 , \29104 );
and \U$41824 ( \42202 , \31498 , \29102 );
nor \U$41825 ( \42203 , \42201 , \42202 );
xnor \U$41826 ( \42204 , \42203 , \28855 );
and \U$41827 ( \42205 , \42199 , \42204 );
and \U$41828 ( \42206 , \42195 , \42204 );
or \U$41829 ( \42207 , \42200 , \42205 , \42206 );
and \U$41830 ( \42208 , \42191 , \42207 );
xor \U$41831 ( \42209 , \42093 , \42097 );
xor \U$41832 ( \42210 , \42209 , \42100 );
and \U$41833 ( \42211 , \42207 , \42210 );
and \U$41834 ( \42212 , \42191 , \42210 );
or \U$41835 ( \42213 , \42208 , \42211 , \42212 );
xor \U$41836 ( \42214 , \42107 , \42111 );
xor \U$41837 ( \42215 , \42214 , \27766 );
xor \U$41838 ( \42216 , \42120 , \42124 );
xor \U$41839 ( \42217 , \42216 , \42129 );
and \U$41840 ( \42218 , \42215 , \42217 );
and \U$41841 ( \42219 , \42213 , \42218 );
xor \U$41842 ( \42220 , \42137 , \42139 );
xor \U$41843 ( \42221 , \42220 , \42141 );
and \U$41844 ( \42222 , \42218 , \42221 );
and \U$41845 ( \42223 , \42213 , \42221 );
or \U$41846 ( \42224 , \42219 , \42222 , \42223 );
xor \U$41847 ( \42225 , \42135 , \42144 );
xor \U$41848 ( \42226 , \42225 , \42147 );
and \U$41849 ( \42227 , \42224 , \42226 );
xor \U$41850 ( \42228 , \42152 , \42154 );
and \U$41851 ( \42229 , \42226 , \42228 );
and \U$41852 ( \42230 , \42224 , \42228 );
or \U$41853 ( \42231 , \42227 , \42229 , \42230 );
and \U$41854 ( \42232 , \42175 , \42231 );
xor \U$41855 ( \42233 , \42175 , \42231 );
xor \U$41856 ( \42234 , \42224 , \42226 );
xor \U$41857 ( \42235 , \42234 , \42228 );
and \U$41858 ( \42236 , \29040 , \32151 );
and \U$41859 ( \42237 , \28514 , \32148 );
nor \U$41860 ( \42238 , \42236 , \42237 );
xnor \U$41861 ( \42239 , \42238 , \31096 );
and \U$41862 ( \42240 , \29710 , \31338 );
and \U$41863 ( \42241 , \29464 , \31336 );
nor \U$41864 ( \42242 , \42240 , \42241 );
xnor \U$41865 ( \42243 , \42242 , \31099 );
and \U$41866 ( \42244 , \42239 , \42243 );
and \U$41867 ( \42245 , \42243 , \28315 );
and \U$41868 ( \42246 , \42239 , \28315 );
or \U$41869 ( \42247 , \42244 , \42245 , \42246 );
and \U$41870 ( \42248 , \30034 , \30770 );
and \U$41871 ( \42249 , \29715 , \30768 );
nor \U$41872 ( \42250 , \42248 , \42249 );
xnor \U$41873 ( \42251 , \42250 , \30460 );
and \U$41874 ( \42252 , \30887 , \30233 );
and \U$41875 ( \42253 , \30318 , \30231 );
nor \U$41876 ( \42254 , \42252 , \42253 );
xnor \U$41877 ( \42255 , \42254 , \29862 );
and \U$41878 ( \42256 , \42251 , \42255 );
and \U$41879 ( \42257 , \31498 , \29671 );
and \U$41880 ( \42258 , \30895 , \29669 );
nor \U$41881 ( \42259 , \42257 , \42258 );
xnor \U$41882 ( \42260 , \42259 , \29353 );
and \U$41883 ( \42261 , \42255 , \42260 );
and \U$41884 ( \42262 , \42251 , \42260 );
or \U$41885 ( \42263 , \42256 , \42261 , \42262 );
and \U$41886 ( \42264 , \42247 , \42263 );
and \U$41887 ( \42265 , \32304 , \28575 );
and \U$41888 ( \42266 , \31684 , \28573 );
nor \U$41889 ( \42267 , \42265 , \42266 );
xnor \U$41890 ( \42268 , \42267 , \28315 );
and \U$41891 ( \42269 , \42263 , \42268 );
and \U$41892 ( \42270 , \42247 , \42268 );
or \U$41893 ( \42271 , \42264 , \42269 , \42270 );
xor \U$41894 ( \42272 , \42191 , \42207 );
xor \U$41895 ( \42273 , \42272 , \42210 );
and \U$41896 ( \42274 , \42271 , \42273 );
xor \U$41897 ( \42275 , \42215 , \42217 );
and \U$41898 ( \42276 , \42273 , \42275 );
and \U$41899 ( \42277 , \42271 , \42275 );
or \U$41900 ( \42278 , \42274 , \42276 , \42277 );
xor \U$41901 ( \42279 , \42103 , \42115 );
xor \U$41902 ( \42280 , \42279 , \42132 );
and \U$41903 ( \42281 , \42278 , \42280 );
xor \U$41904 ( \42282 , \42213 , \42218 );
xor \U$41905 ( \42283 , \42282 , \42221 );
and \U$41906 ( \42284 , \42280 , \42283 );
and \U$41907 ( \42285 , \42278 , \42283 );
or \U$41908 ( \42286 , \42281 , \42284 , \42285 );
and \U$41909 ( \42287 , \42235 , \42286 );
xor \U$41910 ( \42288 , \42235 , \42286 );
xor \U$41911 ( \42289 , \42278 , \42280 );
xor \U$41912 ( \42290 , \42289 , \42283 );
and \U$41913 ( \42291 , \30895 , \30233 );
and \U$41914 ( \42292 , \30887 , \30231 );
nor \U$41915 ( \42293 , \42291 , \42292 );
xnor \U$41916 ( \42294 , \42293 , \29862 );
and \U$41917 ( \42295 , \31503 , \29671 );
and \U$41918 ( \42296 , \31498 , \29669 );
nor \U$41919 ( \42297 , \42295 , \42296 );
xnor \U$41920 ( \42298 , \42297 , \29353 );
and \U$41921 ( \42299 , \42294 , \42298 );
and \U$41922 ( \42300 , \32304 , \29104 );
and \U$41923 ( \42301 , \31684 , \29102 );
nor \U$41924 ( \42302 , \42300 , \42301 );
xnor \U$41925 ( \42303 , \42302 , \28855 );
and \U$41926 ( \42304 , \42298 , \42303 );
and \U$41927 ( \42305 , \42294 , \42303 );
or \U$41928 ( \42306 , \42299 , \42304 , \42305 );
and \U$41929 ( \42307 , \29464 , \32151 );
and \U$41930 ( \42308 , \29040 , \32148 );
nor \U$41931 ( \42309 , \42307 , \42308 );
xnor \U$41932 ( \42310 , \42309 , \31096 );
and \U$41933 ( \42311 , \29715 , \31338 );
and \U$41934 ( \42312 , \29710 , \31336 );
nor \U$41935 ( \42313 , \42311 , \42312 );
xnor \U$41936 ( \42314 , \42313 , \31099 );
and \U$41937 ( \42315 , \42310 , \42314 );
and \U$41938 ( \42316 , \30318 , \30770 );
and \U$41939 ( \42317 , \30034 , \30768 );
nor \U$41940 ( \42318 , \42316 , \42317 );
xnor \U$41941 ( \42319 , \42318 , \30460 );
and \U$41942 ( \42320 , \42314 , \42319 );
and \U$41943 ( \42321 , \42310 , \42319 );
or \U$41944 ( \42322 , \42315 , \42320 , \42321 );
and \U$41945 ( \42323 , \42306 , \42322 );
and \U$41946 ( \42324 , \31684 , \29104 );
and \U$41947 ( \42325 , \31503 , \29102 );
nor \U$41948 ( \42326 , \42324 , \42325 );
xnor \U$41949 ( \42327 , \42326 , \28855 );
and \U$41950 ( \42328 , \42322 , \42327 );
and \U$41951 ( \42329 , \42306 , \42327 );
or \U$41952 ( \42330 , \42323 , \42328 , \42329 );
nand \U$41953 ( \42331 , \32304 , \28573 );
xnor \U$41954 ( \42332 , \42331 , \28315 );
xor \U$41955 ( \42333 , \42239 , \42243 );
xor \U$41956 ( \42334 , \42333 , \28315 );
and \U$41957 ( \42335 , \42332 , \42334 );
xor \U$41958 ( \42336 , \42251 , \42255 );
xor \U$41959 ( \42337 , \42336 , \42260 );
and \U$41960 ( \42338 , \42334 , \42337 );
and \U$41961 ( \42339 , \42332 , \42337 );
or \U$41962 ( \42340 , \42335 , \42338 , \42339 );
and \U$41963 ( \42341 , \42330 , \42340 );
xor \U$41964 ( \42342 , \42195 , \42199 );
xor \U$41965 ( \42343 , \42342 , \42204 );
and \U$41966 ( \42344 , \42340 , \42343 );
and \U$41967 ( \42345 , \42330 , \42343 );
or \U$41968 ( \42346 , \42341 , \42344 , \42345 );
xor \U$41969 ( \42347 , \42179 , \42183 );
xor \U$41970 ( \42348 , \42347 , \42188 );
xor \U$41971 ( \42349 , \42247 , \42263 );
xor \U$41972 ( \42350 , \42349 , \42268 );
and \U$41973 ( \42351 , \42348 , \42350 );
and \U$41974 ( \42352 , \42346 , \42351 );
xor \U$41975 ( \42353 , \42271 , \42273 );
xor \U$41976 ( \42354 , \42353 , \42275 );
and \U$41977 ( \42355 , \42351 , \42354 );
and \U$41978 ( \42356 , \42346 , \42354 );
or \U$41979 ( \42357 , \42352 , \42355 , \42356 );
and \U$41980 ( \42358 , \42290 , \42357 );
xor \U$41981 ( \42359 , \42290 , \42357 );
xor \U$41982 ( \42360 , \42346 , \42351 );
xor \U$41983 ( \42361 , \42360 , \42354 );
and \U$41984 ( \42362 , \30887 , \30770 );
and \U$41985 ( \42363 , \30318 , \30768 );
nor \U$41986 ( \42364 , \42362 , \42363 );
xnor \U$41987 ( \42365 , \42364 , \30460 );
and \U$41988 ( \42366 , \31498 , \30233 );
and \U$41989 ( \42367 , \30895 , \30231 );
nor \U$41990 ( \42368 , \42366 , \42367 );
xnor \U$41991 ( \42369 , \42368 , \29862 );
and \U$41992 ( \42370 , \42365 , \42369 );
and \U$41993 ( \42371 , \31684 , \29671 );
and \U$41994 ( \42372 , \31503 , \29669 );
nor \U$41995 ( \42373 , \42371 , \42372 );
xnor \U$41996 ( \42374 , \42373 , \29353 );
and \U$41997 ( \42375 , \42369 , \42374 );
and \U$41998 ( \42376 , \42365 , \42374 );
or \U$41999 ( \42377 , \42370 , \42375 , \42376 );
and \U$42000 ( \42378 , \29710 , \32151 );
and \U$42001 ( \42379 , \29464 , \32148 );
nor \U$42002 ( \42380 , \42378 , \42379 );
xnor \U$42003 ( \42381 , \42380 , \31096 );
and \U$42004 ( \42382 , \30034 , \31338 );
and \U$42005 ( \42383 , \29715 , \31336 );
nor \U$42006 ( \42384 , \42382 , \42383 );
xnor \U$42007 ( \42385 , \42384 , \31099 );
and \U$42008 ( \42386 , \42381 , \42385 );
and \U$42009 ( \42387 , \42385 , \28855 );
and \U$42010 ( \42388 , \42381 , \28855 );
or \U$42011 ( \42389 , \42386 , \42387 , \42388 );
and \U$42012 ( \42390 , \42377 , \42389 );
xor \U$42013 ( \42391 , \42294 , \42298 );
xor \U$42014 ( \42392 , \42391 , \42303 );
and \U$42015 ( \42393 , \42389 , \42392 );
and \U$42016 ( \42394 , \42377 , \42392 );
or \U$42017 ( \42395 , \42390 , \42393 , \42394 );
xor \U$42018 ( \42396 , \42306 , \42322 );
xor \U$42019 ( \42397 , \42396 , \42327 );
and \U$42020 ( \42398 , \42395 , \42397 );
xor \U$42021 ( \42399 , \42332 , \42334 );
xor \U$42022 ( \42400 , \42399 , \42337 );
and \U$42023 ( \42401 , \42397 , \42400 );
and \U$42024 ( \42402 , \42395 , \42400 );
or \U$42025 ( \42403 , \42398 , \42401 , \42402 );
xor \U$42026 ( \42404 , \42330 , \42340 );
xor \U$42027 ( \42405 , \42404 , \42343 );
and \U$42028 ( \42406 , \42403 , \42405 );
xor \U$42029 ( \42407 , \42348 , \42350 );
and \U$42030 ( \42408 , \42405 , \42407 );
and \U$42031 ( \42409 , \42403 , \42407 );
or \U$42032 ( \42410 , \42406 , \42408 , \42409 );
and \U$42033 ( \42411 , \42361 , \42410 );
xor \U$42034 ( \42412 , \42361 , \42410 );
xor \U$42035 ( \42413 , \42403 , \42405 );
xor \U$42036 ( \42414 , \42413 , \42407 );
and \U$42037 ( \42415 , \29715 , \32151 );
and \U$42038 ( \42416 , \29710 , \32148 );
nor \U$42039 ( \42417 , \42415 , \42416 );
xnor \U$42040 ( \42418 , \42417 , \31096 );
and \U$42041 ( \42419 , \30318 , \31338 );
and \U$42042 ( \42420 , \30034 , \31336 );
nor \U$42043 ( \42421 , \42419 , \42420 );
xnor \U$42044 ( \42422 , \42421 , \31099 );
and \U$42045 ( \42423 , \42418 , \42422 );
and \U$42046 ( \42424 , \30895 , \30770 );
and \U$42047 ( \42425 , \30887 , \30768 );
nor \U$42048 ( \42426 , \42424 , \42425 );
xnor \U$42049 ( \42427 , \42426 , \30460 );
and \U$42050 ( \42428 , \42422 , \42427 );
and \U$42051 ( \42429 , \42418 , \42427 );
or \U$42052 ( \42430 , \42423 , \42428 , \42429 );
nand \U$42053 ( \42431 , \32304 , \29102 );
xnor \U$42054 ( \42432 , \42431 , \28855 );
and \U$42055 ( \42433 , \42430 , \42432 );
xor \U$42056 ( \42434 , \42365 , \42369 );
xor \U$42057 ( \42435 , \42434 , \42374 );
and \U$42058 ( \42436 , \42432 , \42435 );
and \U$42059 ( \42437 , \42430 , \42435 );
or \U$42060 ( \42438 , \42433 , \42436 , \42437 );
xor \U$42061 ( \42439 , \42310 , \42314 );
xor \U$42062 ( \42440 , \42439 , \42319 );
and \U$42063 ( \42441 , \42438 , \42440 );
xor \U$42064 ( \42442 , \42377 , \42389 );
xor \U$42065 ( \42443 , \42442 , \42392 );
and \U$42066 ( \42444 , \42440 , \42443 );
and \U$42067 ( \42445 , \42438 , \42443 );
or \U$42068 ( \42446 , \42441 , \42444 , \42445 );
xor \U$42069 ( \42447 , \42395 , \42397 );
xor \U$42070 ( \42448 , \42447 , \42400 );
and \U$42071 ( \42449 , \42446 , \42448 );
and \U$42072 ( \42450 , \42414 , \42449 );
xor \U$42073 ( \42451 , \42414 , \42449 );
xor \U$42074 ( \42452 , \42446 , \42448 );
and \U$42075 ( \42453 , \31498 , \30770 );
and \U$42076 ( \42454 , \30895 , \30768 );
nor \U$42077 ( \42455 , \42453 , \42454 );
xnor \U$42078 ( \42456 , \42455 , \30460 );
and \U$42079 ( \42457 , \31684 , \30233 );
and \U$42080 ( \42458 , \31503 , \30231 );
nor \U$42081 ( \42459 , \42457 , \42458 );
xnor \U$42082 ( \42460 , \42459 , \29862 );
and \U$42083 ( \42461 , \42456 , \42460 );
nand \U$42084 ( \42462 , \32304 , \29669 );
xnor \U$42085 ( \42463 , \42462 , \29353 );
and \U$42086 ( \42464 , \42460 , \42463 );
and \U$42087 ( \42465 , \42456 , \42463 );
or \U$42088 ( \42466 , \42461 , \42464 , \42465 );
and \U$42089 ( \42467 , \30034 , \32151 );
and \U$42090 ( \42468 , \29715 , \32148 );
nor \U$42091 ( \42469 , \42467 , \42468 );
xnor \U$42092 ( \42470 , \42469 , \31096 );
and \U$42093 ( \42471 , \30887 , \31338 );
and \U$42094 ( \42472 , \30318 , \31336 );
nor \U$42095 ( \42473 , \42471 , \42472 );
xnor \U$42096 ( \42474 , \42473 , \31099 );
and \U$42097 ( \42475 , \42470 , \42474 );
and \U$42098 ( \42476 , \42474 , \29353 );
and \U$42099 ( \42477 , \42470 , \29353 );
or \U$42100 ( \42478 , \42475 , \42476 , \42477 );
and \U$42101 ( \42479 , \42466 , \42478 );
and \U$42102 ( \42480 , \31503 , \30233 );
and \U$42103 ( \42481 , \31498 , \30231 );
nor \U$42104 ( \42482 , \42480 , \42481 );
xnor \U$42105 ( \42483 , \42482 , \29862 );
and \U$42106 ( \42484 , \42478 , \42483 );
and \U$42107 ( \42485 , \42466 , \42483 );
or \U$42108 ( \42486 , \42479 , \42484 , \42485 );
and \U$42109 ( \42487 , \32304 , \29671 );
and \U$42110 ( \42488 , \31684 , \29669 );
nor \U$42111 ( \42489 , \42487 , \42488 );
xnor \U$42112 ( \42490 , \42489 , \29353 );
xor \U$42113 ( \42491 , \42418 , \42422 );
xor \U$42114 ( \42492 , \42491 , \42427 );
and \U$42115 ( \42493 , \42490 , \42492 );
and \U$42116 ( \42494 , \42486 , \42493 );
xor \U$42117 ( \42495 , \42381 , \42385 );
xor \U$42118 ( \42496 , \42495 , \28855 );
and \U$42119 ( \42497 , \42493 , \42496 );
and \U$42120 ( \42498 , \42486 , \42496 );
or \U$42121 ( \42499 , \42494 , \42497 , \42498 );
xor \U$42122 ( \42500 , \42438 , \42440 );
xor \U$42123 ( \42501 , \42500 , \42443 );
and \U$42124 ( \42502 , \42499 , \42501 );
and \U$42125 ( \42503 , \42452 , \42502 );
xor \U$42126 ( \42504 , \42452 , \42502 );
xor \U$42127 ( \42505 , \42499 , \42501 );
xor \U$42128 ( \42506 , \42430 , \42432 );
xor \U$42129 ( \42507 , \42506 , \42435 );
xor \U$42130 ( \42508 , \42486 , \42493 );
xor \U$42131 ( \42509 , \42508 , \42496 );
and \U$42132 ( \42510 , \42507 , \42509 );
and \U$42133 ( \42511 , \42505 , \42510 );
xor \U$42134 ( \42512 , \42505 , \42510 );
xor \U$42135 ( \42513 , \42507 , \42509 );
and \U$42136 ( \42514 , \30318 , \32151 );
and \U$42137 ( \42515 , \30034 , \32148 );
nor \U$42138 ( \42516 , \42514 , \42515 );
xnor \U$42139 ( \42517 , \42516 , \31096 );
and \U$42140 ( \42518 , \30895 , \31338 );
and \U$42141 ( \42519 , \30887 , \31336 );
nor \U$42142 ( \42520 , \42518 , \42519 );
xnor \U$42143 ( \42521 , \42520 , \31099 );
and \U$42144 ( \42522 , \42517 , \42521 );
and \U$42145 ( \42523 , \31503 , \30770 );
and \U$42146 ( \42524 , \31498 , \30768 );
nor \U$42147 ( \42525 , \42523 , \42524 );
xnor \U$42148 ( \42526 , \42525 , \30460 );
and \U$42149 ( \42527 , \42521 , \42526 );
and \U$42150 ( \42528 , \42517 , \42526 );
or \U$42151 ( \42529 , \42522 , \42527 , \42528 );
xor \U$42152 ( \42530 , \42456 , \42460 );
xor \U$42153 ( \42531 , \42530 , \42463 );
and \U$42154 ( \42532 , \42529 , \42531 );
xor \U$42155 ( \42533 , \42470 , \42474 );
xor \U$42156 ( \42534 , \42533 , \29353 );
and \U$42157 ( \42535 , \42531 , \42534 );
and \U$42158 ( \42536 , \42529 , \42534 );
or \U$42159 ( \42537 , \42532 , \42535 , \42536 );
xor \U$42160 ( \42538 , \42466 , \42478 );
xor \U$42161 ( \42539 , \42538 , \42483 );
and \U$42162 ( \42540 , \42537 , \42539 );
xor \U$42163 ( \42541 , \42490 , \42492 );
and \U$42164 ( \42542 , \42539 , \42541 );
and \U$42165 ( \42543 , \42537 , \42541 );
or \U$42166 ( \42544 , \42540 , \42542 , \42543 );
and \U$42167 ( \42545 , \42513 , \42544 );
xor \U$42168 ( \42546 , \42513 , \42544 );
xor \U$42169 ( \42547 , \42537 , \42539 );
xor \U$42170 ( \42548 , \42547 , \42541 );
and \U$42171 ( \42549 , \30887 , \32151 );
and \U$42172 ( \42550 , \30318 , \32148 );
nor \U$42173 ( \42551 , \42549 , \42550 );
xnor \U$42174 ( \42552 , \42551 , \31096 );
and \U$42175 ( \42553 , \31498 , \31338 );
and \U$42176 ( \42554 , \30895 , \31336 );
nor \U$42177 ( \42555 , \42553 , \42554 );
xnor \U$42178 ( \42556 , \42555 , \31099 );
and \U$42179 ( \42557 , \42552 , \42556 );
and \U$42180 ( \42558 , \42556 , \29862 );
and \U$42181 ( \42559 , \42552 , \29862 );
or \U$42182 ( \42560 , \42557 , \42558 , \42559 );
and \U$42183 ( \42561 , \31684 , \30770 );
and \U$42184 ( \42562 , \31503 , \30768 );
nor \U$42185 ( \42563 , \42561 , \42562 );
xnor \U$42186 ( \42564 , \42563 , \30460 );
nand \U$42187 ( \42565 , \32304 , \30231 );
xnor \U$42188 ( \42566 , \42565 , \29862 );
and \U$42189 ( \42567 , \42564 , \42566 );
and \U$42190 ( \42568 , \42560 , \42567 );
and \U$42191 ( \42569 , \32304 , \30233 );
and \U$42192 ( \42570 , \31684 , \30231 );
nor \U$42193 ( \42571 , \42569 , \42570 );
xnor \U$42194 ( \42572 , \42571 , \29862 );
and \U$42195 ( \42573 , \42567 , \42572 );
and \U$42196 ( \42574 , \42560 , \42572 );
or \U$42197 ( \42575 , \42568 , \42573 , \42574 );
xor \U$42198 ( \42576 , \42529 , \42531 );
xor \U$42199 ( \42577 , \42576 , \42534 );
and \U$42200 ( \42578 , \42575 , \42577 );
and \U$42201 ( \42579 , \42548 , \42578 );
xor \U$42202 ( \42580 , \42548 , \42578 );
xor \U$42203 ( \42581 , \42575 , \42577 );
xor \U$42204 ( \42582 , \42517 , \42521 );
xor \U$42205 ( \42583 , \42582 , \42526 );
xor \U$42206 ( \42584 , \42560 , \42567 );
xor \U$42207 ( \42585 , \42584 , \42572 );
and \U$42208 ( \42586 , \42583 , \42585 );
and \U$42209 ( \42587 , \42581 , \42586 );
xor \U$42210 ( \42588 , \42581 , \42586 );
xor \U$42211 ( \42589 , \42583 , \42585 );
and \U$42212 ( \42590 , \30895 , \32151 );
and \U$42213 ( \42591 , \30887 , \32148 );
nor \U$42214 ( \42592 , \42590 , \42591 );
xnor \U$42215 ( \42593 , \42592 , \31096 );
and \U$42216 ( \42594 , \31503 , \31338 );
and \U$42217 ( \42595 , \31498 , \31336 );
nor \U$42218 ( \42596 , \42594 , \42595 );
xnor \U$42219 ( \42597 , \42596 , \31099 );
and \U$42220 ( \42598 , \42593 , \42597 );
and \U$42221 ( \42599 , \32304 , \30770 );
and \U$42222 ( \42600 , \31684 , \30768 );
nor \U$42223 ( \42601 , \42599 , \42600 );
xnor \U$42224 ( \42602 , \42601 , \30460 );
and \U$42225 ( \42603 , \42597 , \42602 );
and \U$42226 ( \42604 , \42593 , \42602 );
or \U$42227 ( \42605 , \42598 , \42603 , \42604 );
xor \U$42228 ( \42606 , \42552 , \42556 );
xor \U$42229 ( \42607 , \42606 , \29862 );
and \U$42230 ( \42608 , \42605 , \42607 );
xor \U$42231 ( \42609 , \42564 , \42566 );
and \U$42232 ( \42610 , \42607 , \42609 );
and \U$42233 ( \42611 , \42605 , \42609 );
or \U$42234 ( \42612 , \42608 , \42610 , \42611 );
and \U$42235 ( \42613 , \42589 , \42612 );
xor \U$42236 ( \42614 , \42589 , \42612 );
xor \U$42237 ( \42615 , \42605 , \42607 );
xor \U$42238 ( \42616 , \42615 , \42609 );
and \U$42239 ( \42617 , \31498 , \32151 );
and \U$42240 ( \42618 , \30895 , \32148 );
nor \U$42241 ( \42619 , \42617 , \42618 );
xnor \U$42242 ( \42620 , \42619 , \31096 );
and \U$42243 ( \42621 , \31684 , \31338 );
and \U$42244 ( \42622 , \31503 , \31336 );
nor \U$42245 ( \42623 , \42621 , \42622 );
xnor \U$42246 ( \42624 , \42623 , \31099 );
and \U$42247 ( \42625 , \42620 , \42624 );
and \U$42248 ( \42626 , \42624 , \30460 );
and \U$42249 ( \42627 , \42620 , \30460 );
or \U$42250 ( \42628 , \42625 , \42626 , \42627 );
xor \U$42251 ( \42629 , \42593 , \42597 );
xor \U$42252 ( \42630 , \42629 , \42602 );
and \U$42253 ( \42631 , \42628 , \42630 );
and \U$42254 ( \42632 , \42616 , \42631 );
xor \U$42255 ( \42633 , \42616 , \42631 );
xor \U$42256 ( \42634 , \42628 , \42630 );
nand \U$42257 ( \42635 , \32304 , \30768 );
xnor \U$42258 ( \42636 , \42635 , \30460 );
xor \U$42259 ( \42637 , \42620 , \42624 );
xor \U$42260 ( \42638 , \42637 , \30460 );
and \U$42261 ( \42639 , \42636 , \42638 );
and \U$42262 ( \42640 , \42634 , \42639 );
xor \U$42263 ( \42641 , \42634 , \42639 );
xor \U$42264 ( \42642 , \42636 , \42638 );
and \U$42265 ( \42643 , \31503 , \32151 );
and \U$42266 ( \42644 , \31498 , \32148 );
nor \U$42267 ( \42645 , \42643 , \42644 );
xnor \U$42268 ( \42646 , \42645 , \31096 );
and \U$42269 ( \42647 , \32304 , \31338 );
and \U$42270 ( \42648 , \31684 , \31336 );
nor \U$42271 ( \42649 , \42647 , \42648 );
xnor \U$42272 ( \42650 , \42649 , \31099 );
and \U$42273 ( \42651 , \42646 , \42650 );
and \U$42274 ( \42652 , \42642 , \42651 );
xor \U$42275 ( \42653 , \42642 , \42651 );
xor \U$42276 ( \42654 , \42646 , \42650 );
and \U$42277 ( \42655 , \31684 , \32151 );
and \U$42278 ( \42656 , \31503 , \32148 );
nor \U$42279 ( \42657 , \42655 , \42656 );
xnor \U$42280 ( \42658 , \42657 , \31096 );
and \U$42281 ( \42659 , \42658 , \31099 );
and \U$42282 ( \42660 , \42654 , \42659 );
xor \U$42283 ( \42661 , \42654 , \42659 );
nand \U$42284 ( \42662 , \32304 , \31336 );
xnor \U$42285 ( \42663 , \42662 , \31099 );
xor \U$42286 ( \42664 , \42658 , \31099 );
and \U$42287 ( \42665 , \42663 , \42664 );
xor \U$42288 ( \42666 , \42663 , \42664 );
and \U$42289 ( \42667 , \32304 , \32151 );
and \U$42290 ( \42668 , \31684 , \32148 );
nor \U$42291 ( \42669 , \42667 , \42668 );
xnor \U$42292 ( \42670 , \42669 , \31096 );
nand \U$42293 ( \42671 , \32304 , \32148 );
xnor \U$42294 ( \42672 , \42671 , \31096 );
and \U$42295 ( \42673 , \42672 , \31096 );
and \U$42296 ( \42674 , \42670 , \42673 );
and \U$42297 ( \42675 , \42666 , \42674 );
or \U$42298 ( \42676 , \42665 , \42675 );
and \U$42299 ( \42677 , \42661 , \42676 );
or \U$42300 ( \42678 , \42660 , \42677 );
and \U$42301 ( \42679 , \42653 , \42678 );
or \U$42302 ( \42680 , \42652 , \42679 );
and \U$42303 ( \42681 , \42641 , \42680 );
or \U$42304 ( \42682 , \42640 , \42681 );
and \U$42305 ( \42683 , \42633 , \42682 );
or \U$42306 ( \42684 , \42632 , \42683 );
and \U$42307 ( \42685 , \42614 , \42684 );
or \U$42308 ( \42686 , \42613 , \42685 );
and \U$42309 ( \42687 , \42588 , \42686 );
or \U$42310 ( \42688 , \42587 , \42687 );
and \U$42311 ( \42689 , \42580 , \42688 );
or \U$42312 ( \42690 , \42579 , \42689 );
and \U$42313 ( \42691 , \42546 , \42690 );
or \U$42314 ( \42692 , \42545 , \42691 );
and \U$42315 ( \42693 , \42512 , \42692 );
or \U$42316 ( \42694 , \42511 , \42693 );
and \U$42317 ( \42695 , \42504 , \42694 );
or \U$42318 ( \42696 , \42503 , \42695 );
and \U$42319 ( \42697 , \42451 , \42696 );
or \U$42320 ( \42698 , \42450 , \42697 );
and \U$42321 ( \42699 , \42412 , \42698 );
or \U$42322 ( \42700 , \42411 , \42699 );
and \U$42323 ( \42701 , \42359 , \42700 );
or \U$42324 ( \42702 , \42358 , \42701 );
and \U$42325 ( \42703 , \42288 , \42702 );
or \U$42326 ( \42704 , \42287 , \42703 );
and \U$42327 ( \42705 , \42233 , \42704 );
or \U$42328 ( \42706 , \42232 , \42705 );
and \U$42329 ( \42707 , \42174 , \42706 );
or \U$42330 ( \42708 , \42173 , \42707 );
and \U$42331 ( \42709 , \42166 , \42708 );
or \U$42332 ( \42710 , \42165 , \42709 );
and \U$42333 ( \42711 , \42087 , \42710 );
or \U$42334 ( \42712 , \42086 , \42711 );
and \U$42335 ( \42713 , \42007 , \42712 );
or \U$42336 ( \42714 , \42006 , \42713 );
and \U$42337 ( \42715 , \41912 , \42714 );
or \U$42338 ( \42716 , \41911 , \42715 );
and \U$42339 ( \42717 , \41824 , \42716 );
or \U$42340 ( \42718 , \41823 , \42717 );
and \U$42341 ( \42719 , \41732 , \42718 );
or \U$42342 ( \42720 , \41731 , \42719 );
and \U$42343 ( \42721 , \41644 , \42720 );
or \U$42344 ( \42722 , \41643 , \42721 );
and \U$42345 ( \42723 , \41529 , \42722 );
or \U$42346 ( \42724 , \41528 , \42723 );
and \U$42347 ( \42725 , \41433 , \42724 );
or \U$42348 ( \42726 , \41432 , \42725 );
and \U$42349 ( \42727 , \41425 , \42726 );
or \U$42350 ( \42728 , \41424 , \42727 );
and \U$42351 ( \42729 , \41310 , \42728 );
or \U$42352 ( \42730 , \41309 , \42729 );
and \U$42353 ( \42731 , \41186 , \42730 );
or \U$42354 ( \42732 , \41185 , \42731 );
and \U$42355 ( \42733 , \41046 , \42732 );
or \U$42356 ( \42734 , \41045 , \42733 );
and \U$42357 ( \42735 , \40922 , \42734 );
or \U$42358 ( \42736 , \40921 , \42735 );
and \U$42359 ( \42737 , \40778 , \42736 );
or \U$42360 ( \42738 , \40777 , \42737 );
and \U$42361 ( \42739 , \40653 , \42738 );
or \U$42362 ( \42740 , \40652 , \42739 );
and \U$42363 ( \42741 , \40514 , \42740 );
or \U$42364 ( \42742 , \40513 , \42741 );
and \U$42365 ( \42743 , \40350 , \42742 );
or \U$42366 ( \42744 , \40349 , \42743 );
and \U$42367 ( \42745 , \40198 , \42744 );
or \U$42368 ( \42746 , \40197 , \42745 );
and \U$42369 ( \42747 , \40058 , \42746 );
or \U$42370 ( \42748 , \40057 , \42747 );
and \U$42371 ( \42749 , \39890 , \42748 );
or \U$42372 ( \42750 , \39889 , \42749 );
and \U$42373 ( \42751 , \39882 , \42750 );
or \U$42374 ( \42752 , \39881 , \42751 );
and \U$42375 ( \42753 , \39711 , \42752 );
or \U$42376 ( \42754 , \39710 , \42753 );
and \U$42377 ( \42755 , \39535 , \42754 );
or \U$42378 ( \42756 , \39534 , \42755 );
and \U$42379 ( \42757 , \39345 , \42756 );
or \U$42380 ( \42758 , \39344 , \42757 );
and \U$42381 ( \42759 , \39158 , \42758 );
or \U$42382 ( \42760 , \39157 , \42759 );
and \U$42383 ( \42761 , \38973 , \42760 );
or \U$42384 ( \42762 , \38972 , \42761 );
and \U$42385 ( \42763 , \38765 , \42762 );
or \U$42386 ( \42764 , \38764 , \42763 );
and \U$42387 ( \42765 , \38569 , \42764 );
or \U$42388 ( \42766 , \38568 , \42765 );
and \U$42389 ( \42767 , \38372 , \42766 );
or \U$42390 ( \42768 , \38371 , \42767 );
and \U$42391 ( \42769 , \38159 , \42768 );
or \U$42392 ( \42770 , \38158 , \42769 );
and \U$42393 ( \42771 , \37948 , \42770 );
or \U$42394 ( \42772 , \37947 , \42771 );
and \U$42395 ( \42773 , \37717 , \42772 );
or \U$42396 ( \42774 , \37716 , \42773 );
and \U$42397 ( \42775 , \37487 , \42774 );
or \U$42398 ( \42776 , \37486 , \42775 );
and \U$42399 ( \42777 , \37268 , \42776 );
or \U$42400 ( \42778 , \37267 , \42777 );
and \U$42401 ( \42779 , \37043 , \42778 );
or \U$42402 ( \42780 , \37042 , \42779 );
and \U$42403 ( \42781 , \36793 , \42780 );
or \U$42404 ( \42782 , \36792 , \42781 );
and \U$42405 ( \42783 , \36563 , \42782 );
or \U$42406 ( \42784 , \36562 , \42783 );
and \U$42407 ( \42785 , \36317 , \42784 );
or \U$42408 ( \42786 , \36316 , \42785 );
and \U$42409 ( \42787 , \36309 , \42786 );
or \U$42410 ( \42788 , \36308 , \42787 );
and \U$42411 ( \42789 , \36048 , \42788 );
or \U$42412 ( \42790 , \36047 , \42789 );
and \U$42413 ( \42791 , \35786 , \42790 );
or \U$42414 ( \42792 , \35785 , \42791 );
and \U$42415 ( \42793 , \35516 , \42792 );
or \U$42416 ( \42794 , \35515 , \42793 );
and \U$42417 ( \42795 , \35239 , \42794 );
or \U$42418 ( \42796 , \35238 , \42795 );
and \U$42419 ( \42797 , \34963 , \42796 );
or \U$42420 ( \42798 , \34962 , \42797 );
and \U$42421 ( \42799 , \34692 , \42798 );
or \U$42422 ( \42800 , \34691 , \42799 );
and \U$42423 ( \42801 , \34389 , \42800 );
or \U$42424 ( \42802 , \34388 , \42801 );
and \U$42425 ( \42803 , \34110 , \42802 );
or \U$42426 ( \42804 , \34109 , \42803 );
and \U$42427 ( \42805 , \33825 , \42804 );
or \U$42428 ( \42806 , \33824 , \42805 );
and \U$42429 ( \42807 , \33509 , \42806 );
or \U$42430 ( \42808 , \33508 , \42807 );
and \U$42431 ( \42809 , \33209 , \42808 );
or \U$42432 ( \42810 , \33208 , \42809 );
and \U$42433 ( \42811 , \32893 , \42810 );
or \U$42434 ( \42812 , \32892 , \42811 );
and \U$42435 ( \42813 , \32575 , \42812 );
or \U$42436 ( \42814 , \32574 , \42813 );
and \U$42437 ( \42815 , \32264 , \42814 );
or \U$42438 ( \42816 , \32263 , \42815 );
and \U$42439 ( \42817 , \31951 , \42816 );
or \U$42440 ( \42818 , \31950 , \42817 );
and \U$42441 ( \42819 , \31635 , \42818 );
or \U$42442 ( \42820 , \31634 , \42819 );
and \U$42443 ( \42821 , \31317 , \42820 );
or \U$42444 ( \42822 , \31316 , \42821 );
and \U$42445 ( \42823 , \31008 , \42822 );
or \U$42446 ( \42824 , \31007 , \42823 );
and \U$42447 ( \42825 , \30712 , \42824 );
or \U$42448 ( \42826 , \30711 , \42825 );
and \U$42449 ( \42827 , \30411 , \42826 );
or \U$42450 ( \42828 , \30410 , \42827 );
and \U$42451 ( \42829 , \30123 , \42828 );
or \U$42452 ( \42830 , \30122 , \42829 );
and \U$42453 ( \42831 , \29840 , \42830 );
or \U$42454 ( \42832 , \29839 , \42831 );
and \U$42455 ( \42833 , \29545 , \42832 );
or \U$42456 ( \42834 , \29544 , \42833 );
and \U$42457 ( \42835 , \29279 , \42834 );
or \U$42458 ( \42836 , \29278 , \42835 );
and \U$42459 ( \42837 , \29013 , \42836 );
or \U$42460 ( \42838 , \29012 , \42837 );
and \U$42461 ( \42839 , \28752 , \42838 );
or \U$42462 ( \42840 , \28751 , \42839 );
and \U$42463 ( \42841 , \28487 , \42840 );
or \U$42464 ( \42842 , \28486 , \42841 );
and \U$42465 ( \42843 , \28224 , \42842 );
or \U$42466 ( \42844 , \28223 , \42843 );
and \U$42467 ( \42845 , \27967 , \42844 );
or \U$42468 ( \42846 , \27966 , \42845 );
and \U$42469 ( \42847 , \27711 , \42846 );
or \U$42470 ( \42848 , \27710 , \42847 );
and \U$42471 ( \42849 , \27458 , \42848 );
or \U$42472 ( \42850 , \27457 , \42849 );
and \U$42473 ( \42851 , \27210 , \42850 );
or \U$42474 ( \42852 , \27209 , \42851 );
and \U$42475 ( \42853 , \26978 , \42852 );
or \U$42476 ( \42854 , \26977 , \42853 );
and \U$42477 ( \42855 , \26735 , \42854 );
or \U$42478 ( \42856 , \26734 , \42855 );
and \U$42479 ( \42857 , \26306 , \42856 );
or \U$42480 ( \42858 , \26305 , \42857 );
and \U$42481 ( \42859 , \26096 , \42858 );
or \U$42482 ( \42860 , \26095 , \42859 );
and \U$42483 ( \42861 , \25889 , \42860 );
or \U$42484 ( \42862 , \25888 , \42861 );
and \U$42485 ( \42863 , \25687 , \42862 );
or \U$42486 ( \42864 , \25686 , \42863 );
and \U$42487 ( \42865 , \25491 , \42864 );
or \U$42488 ( \42866 , \25490 , \42865 );
and \U$42489 ( \42867 , \25294 , \42866 );
or \U$42490 ( \42868 , \25293 , \42867 );
and \U$42491 ( \42869 , \25117 , \42868 );
or \U$42492 ( \42870 , \25116 , \42869 );
and \U$42493 ( \42871 , \24936 , \42870 );
or \U$42494 ( \42872 , \24935 , \42871 );
and \U$42495 ( \42873 , \24765 , \42872 );
or \U$42496 ( \42874 , \24764 , \42873 );
and \U$42497 ( \42875 , \24590 , \42874 );
or \U$42498 ( \42876 , \24589 , \42875 );
and \U$42499 ( \42877 , \24417 , \42876 );
or \U$42500 ( \42878 , \24416 , \42877 );
and \U$42501 ( \42879 , \24250 , \42878 );
or \U$42502 ( \42880 , \24249 , \42879 );
and \U$42503 ( \42881 , \24084 , \42880 );
or \U$42504 ( \42882 , \24083 , \42881 );
and \U$42505 ( \42883 , \23911 , \42882 );
or \U$42506 ( \42884 , \23910 , \42883 );
and \U$42507 ( \42885 , \23631 , \42884 );
or \U$42508 ( \42886 , \23630 , \42885 );
and \U$42509 ( \42887 , \23494 , \42886 );
or \U$42510 ( \42888 , \23493 , \42887 );
and \U$42511 ( \42889 , \23361 , \42888 );
or \U$42512 ( \42890 , \23360 , \42889 );
and \U$42513 ( \42891 , \23240 , \42890 );
or \U$42514 ( \42892 , \23239 , \42891 );
and \U$42515 ( \42893 , \23117 , \42892 );
or \U$42516 ( \42894 , \23116 , \42893 );
and \U$42517 ( \42895 , \23001 , \42894 );
or \U$42518 ( \42896 , \23000 , \42895 );
and \U$42519 ( \42897 , \22886 , \42896 );
or \U$42520 ( \42898 , \22885 , \42897 );
and \U$42521 ( \42899 , \22772 , \42898 );
or \U$42522 ( \42900 , \22771 , \42899 );
and \U$42523 ( \42901 , \22658 , \42900 );
or \U$42524 ( \42902 , \22657 , \42901 );
and \U$42525 ( \42903 , \22476 , \42902 );
or \U$42526 ( \42904 , \22475 , \42903 );
and \U$42527 ( \42905 , \22397 , \42904 );
or \U$42528 ( \42906 , \22396 , \42905 );
and \U$42529 ( \42907 , \22314 , \42906 );
or \U$42530 ( \42908 , \22313 , \42907 );
and \U$42531 ( \42909 , \22233 , \42908 );
or \U$42532 ( \42910 , \22232 , \42909 );
and \U$42533 ( \42911 , \22158 , \42910 );
or \U$42534 ( \42912 , \22157 , \42911 );
and \U$42535 ( \42913 , \22084 , \42912 );
or \U$42536 ( \42914 , \22083 , \42913 );
and \U$42537 ( \42915 , \21964 , \42914 );
or \U$42538 ( \42916 , \21963 , \42915 );
and \U$42539 ( \42917 , \21911 , \42916 );
or \U$42540 ( \42918 , \21910 , \42917 );
and \U$42541 ( \42919 , \21861 , \42918 );
or \U$42542 ( \42920 , \21860 , \42919 );
and \U$42543 ( \42921 , \21809 , \42920 );
or \U$42544 ( \42922 , \21808 , \42921 );
and \U$42545 ( \42923 , \21739 , \42922 );
or \U$42546 ( \42924 , \21738 , \42923 );
xor \U$42547 ( \42925 , \21692 , \42924 );
buf gaee1_GF_PartitionCandidate( \42926_nGaee1 , \42925 );
buf \U$42548 ( \42927 , \42926_nGaee1 );
xor \U$42549 ( \42928 , \21652 , \42927 );
xor \U$42550 ( \42929 , \464 , \21647 );
buf gaeaa_GF_PartitionCandidate( \42930_nGaeaa , \42929 );
buf \U$42551 ( \42931 , \42930_nGaeaa );
xor \U$42552 ( \42932 , \21739 , \42922 );
buf gaebf_GF_PartitionCandidate( \42933_nGaebf , \42932 );
buf \U$42553 ( \42934 , \42933_nGaebf );
and \U$42554 ( \42935 , \42931 , \42934 );
xor \U$42555 ( \42936 , \534 , \21645 );
buf gae73_GF_PartitionCandidate( \42937_nGae73 , \42936 );
buf \U$42556 ( \42938 , \42937_nGae73 );
xor \U$42557 ( \42939 , \21809 , \42920 );
buf gae8d_GF_PartitionCandidate( \42940_nGae8d , \42939 );
buf \U$42558 ( \42941 , \42940_nGae8d );
and \U$42559 ( \42942 , \42938 , \42941 );
xor \U$42560 ( \42943 , \586 , \21643 );
buf gae30_GF_PartitionCandidate( \42944_nGae30 , \42943 );
buf \U$42561 ( \42945 , \42944_nGae30 );
xor \U$42562 ( \42946 , \21861 , \42918 );
buf gae51_GF_PartitionCandidate( \42947_nGae51 , \42946 );
buf \U$42563 ( \42948 , \42947_nGae51 );
and \U$42564 ( \42949 , \42945 , \42948 );
xor \U$42565 ( \42950 , \636 , \21641 );
buf gade1_GF_PartitionCandidate( \42951_nGade1 , \42950 );
buf \U$42566 ( \42952 , \42951_nGade1 );
xor \U$42567 ( \42953 , \21911 , \42916 );
buf gae07_GF_PartitionCandidate( \42954_nGae07 , \42953 );
buf \U$42568 ( \42955 , \42954_nGae07 );
and \U$42569 ( \42956 , \42952 , \42955 );
xor \U$42570 ( \42957 , \689 , \21639 );
buf gad8a_GF_PartitionCandidate( \42958_nGad8a , \42957 );
buf \U$42571 ( \42959 , \42958_nGad8a );
xor \U$42572 ( \42960 , \21964 , \42914 );
buf gadb3_GF_PartitionCandidate( \42961_nGadb3 , \42960 );
buf \U$42573 ( \42962 , \42961_nGadb3 );
and \U$42574 ( \42963 , \42959 , \42962 );
xor \U$42575 ( \42964 , \809 , \21637 );
buf gad2b_GF_PartitionCandidate( \42965_nGad2b , \42964 );
buf \U$42576 ( \42966 , \42965_nGad2b );
xor \U$42577 ( \42967 , \22084 , \42912 );
buf gad59_GF_PartitionCandidate( \42968_nGad59 , \42967 );
buf \U$42578 ( \42969 , \42968_nGad59 );
and \U$42579 ( \42970 , \42966 , \42969 );
xor \U$42580 ( \42971 , \883 , \21635 );
buf gacc0_GF_PartitionCandidate( \42972_nGacc0 , \42971 );
buf \U$42581 ( \42973 , \42972_nGacc0 );
xor \U$42582 ( \42974 , \22158 , \42910 );
buf gacf5_GF_PartitionCandidate( \42975_nGacf5 , \42974 );
buf \U$42583 ( \42976 , \42975_nGacf5 );
and \U$42584 ( \42977 , \42973 , \42976 );
xor \U$42585 ( \42978 , \958 , \21633 );
buf gac4c_GF_PartitionCandidate( \42979_nGac4c , \42978 );
buf \U$42586 ( \42980 , \42979_nGac4c );
xor \U$42587 ( \42981 , \22233 , \42908 );
buf gac83_GF_PartitionCandidate( \42982_nGac83 , \42981 );
buf \U$42588 ( \42983 , \42982_nGac83 );
and \U$42589 ( \42984 , \42980 , \42983 );
xor \U$42590 ( \42985 , \1039 , \21631 );
buf gabce_GF_PartitionCandidate( \42986_nGabce , \42985 );
buf \U$42591 ( \42987 , \42986_nGabce );
xor \U$42592 ( \42988 , \22314 , \42906 );
buf gac0d_GF_PartitionCandidate( \42989_nGac0d , \42988 );
buf \U$42593 ( \42990 , \42989_nGac0d );
and \U$42594 ( \42991 , \42987 , \42990 );
xor \U$42595 ( \42992 , \1122 , \21629 );
buf gab43_GF_PartitionCandidate( \42993_nGab43 , \42992 );
buf \U$42596 ( \42994 , \42993_nGab43 );
xor \U$42597 ( \42995 , \22397 , \42904 );
buf gab87_GF_PartitionCandidate( \42996_nGab87 , \42995 );
buf \U$42598 ( \42997 , \42996_nGab87 );
and \U$42599 ( \42998 , \42994 , \42997 );
xor \U$42600 ( \42999 , \1201 , \21627 );
buf gaab0_GF_PartitionCandidate( \43000_nGaab0 , \42999 );
buf \U$42601 ( \43001 , \43000_nGaab0 );
xor \U$42602 ( \43002 , \22476 , \42902 );
buf gaaf7_GF_PartitionCandidate( \43003_nGaaf7 , \43002 );
buf \U$42603 ( \43004 , \43003_nGaaf7 );
and \U$42604 ( \43005 , \43001 , \43004 );
xor \U$42605 ( \43006 , \1383 , \21625 );
buf gaa15_GF_PartitionCandidate( \43007_nGaa15 , \43006 );
buf \U$42606 ( \43008 , \43007_nGaa15 );
xor \U$42607 ( \43009 , \22658 , \42900 );
buf gaa61_GF_PartitionCandidate( \43010_nGaa61 , \43009 );
buf \U$42608 ( \43011 , \43010_nGaa61 );
and \U$42609 ( \43012 , \43008 , \43011 );
xor \U$42610 ( \43013 , \1497 , \21623 );
buf ga96e_GF_PartitionCandidate( \43014_nGa96e , \43013 );
buf \U$42611 ( \43015 , \43014_nGa96e );
xor \U$42612 ( \43016 , \22772 , \42898 );
buf ga9c1_GF_PartitionCandidate( \43017_nGa9c1 , \43016 );
buf \U$42613 ( \43018 , \43017_nGa9c1 );
and \U$42614 ( \43019 , \43015 , \43018 );
xor \U$42615 ( \43020 , \1611 , \21621 );
buf ga8be_GF_PartitionCandidate( \43021_nGa8be , \43020 );
buf \U$42616 ( \43022 , \43021_nGa8be );
xor \U$42617 ( \43023 , \22886 , \42896 );
buf ga913_GF_PartitionCandidate( \43024_nGa913 , \43023 );
buf \U$42618 ( \43025 , \43024_nGa913 );
and \U$42619 ( \43026 , \43022 , \43025 );
xor \U$42620 ( \43027 , \1726 , \21619 );
buf ga804_GF_PartitionCandidate( \43028_nGa804 , \43027 );
buf \U$42621 ( \43029 , \43028_nGa804 );
xor \U$42622 ( \43030 , \23001 , \42894 );
buf ga861_GF_PartitionCandidate( \43031_nGa861 , \43030 );
buf \U$42623 ( \43032 , \43031_nGa861 );
and \U$42624 ( \43033 , \43029 , \43032 );
xor \U$42625 ( \43034 , \1842 , \21617 );
buf ga740_GF_PartitionCandidate( \43035_nGa740 , \43034 );
buf \U$42626 ( \43036 , \43035_nGa740 );
xor \U$42627 ( \43037 , \23117 , \42892 );
buf ga79f_GF_PartitionCandidate( \43038_nGa79f , \43037 );
buf \U$42628 ( \43039 , \43038_nGa79f );
and \U$42629 ( \43040 , \43036 , \43039 );
xor \U$42630 ( \43041 , \1965 , \21615 );
buf ga672_GF_PartitionCandidate( \43042_nGa672 , \43041 );
buf \U$42631 ( \43043 , \43042_nGa672 );
xor \U$42632 ( \43044 , \23240 , \42890 );
buf ga6d9_GF_PartitionCandidate( \43045_nGa6d9 , \43044 );
buf \U$42633 ( \43046 , \43045_nGa6d9 );
and \U$42634 ( \43047 , \43043 , \43046 );
xor \U$42635 ( \43048 , \2086 , \21613 );
buf ga59a_GF_PartitionCandidate( \43049_nGa59a , \43048 );
buf \U$42636 ( \43050 , \43049_nGa59a );
xor \U$42637 ( \43051 , \23361 , \42888 );
buf ga603_GF_PartitionCandidate( \43052_nGa603 , \43051 );
buf \U$42638 ( \43053 , \43052_nGa603 );
and \U$42639 ( \43054 , \43050 , \43053 );
xor \U$42640 ( \43055 , \2219 , \21611 );
buf ga4bb_GF_PartitionCandidate( \43056_nGa4bb , \43055 );
buf \U$42641 ( \43057 , \43056_nGa4bb );
xor \U$42642 ( \43058 , \23494 , \42886 );
buf ga529_GF_PartitionCandidate( \43059_nGa529 , \43058 );
buf \U$42643 ( \43060 , \43059_nGa529 );
and \U$42644 ( \43061 , \43057 , \43060 );
xor \U$42645 ( \43062 , \2356 , \21609 );
buf ga3d1_GF_PartitionCandidate( \43063_nGa3d1 , \43062 );
buf \U$42646 ( \43064 , \43063_nGa3d1 );
xor \U$42647 ( \43065 , \23631 , \42884 );
buf ga445_GF_PartitionCandidate( \43066_nGa445 , \43065 );
buf \U$42648 ( \43067 , \43066_nGa445 );
and \U$42649 ( \43068 , \43064 , \43067 );
xor \U$42650 ( \43069 , \2636 , \21607 );
buf ga2da_GF_PartitionCandidate( \43070_nGa2da , \43069 );
buf \U$42651 ( \43071 , \43070_nGa2da );
xor \U$42652 ( \43072 , \23911 , \42882 );
buf ga355_GF_PartitionCandidate( \43073_nGa355 , \43072 );
buf \U$42653 ( \43074 , \43073_nGa355 );
and \U$42654 ( \43075 , \43071 , \43074 );
xor \U$42655 ( \43076 , \2809 , \21605 );
buf ga1d7_GF_PartitionCandidate( \43077_nGa1d7 , \43076 );
buf \U$42656 ( \43078 , \43077_nGa1d7 );
xor \U$42657 ( \43079 , \24084 , \42880 );
buf ga257_GF_PartitionCandidate( \43080_nGa257 , \43079 );
buf \U$42658 ( \43081 , \43080_nGa257 );
and \U$42659 ( \43082 , \43078 , \43081 );
xor \U$42660 ( \43083 , \2975 , \21603 );
buf ga0c9_GF_PartitionCandidate( \43084_nGa0c9 , \43083 );
buf \U$42661 ( \43085 , \43084_nGa0c9 );
xor \U$42662 ( \43086 , \24250 , \42878 );
buf ga14f_GF_PartitionCandidate( \43087_nGa14f , \43086 );
buf \U$42663 ( \43088 , \43087_nGa14f );
and \U$42664 ( \43089 , \43085 , \43088 );
xor \U$42665 ( \43090 , \3142 , \21601 );
buf g9fb4_GF_PartitionCandidate( \43091_nG9fb4 , \43090 );
buf \U$42666 ( \43092 , \43091_nG9fb4 );
xor \U$42667 ( \43093 , \24417 , \42876 );
buf ga03b_GF_PartitionCandidate( \43094_nGa03b , \43093 );
buf \U$42668 ( \43095 , \43094_nGa03b );
and \U$42669 ( \43096 , \43092 , \43095 );
xor \U$42670 ( \43097 , \3315 , \21599 );
buf g9e96_GF_PartitionCandidate( \43098_nG9e96 , \43097 );
buf \U$42671 ( \43099 , \43098_nG9e96 );
xor \U$42672 ( \43100 , \24590 , \42874 );
buf g9f25_GF_PartitionCandidate( \43101_nG9f25 , \43100 );
buf \U$42673 ( \43102 , \43101_nG9f25 );
and \U$42674 ( \43103 , \43099 , \43102 );
xor \U$42675 ( \43104 , \3490 , \21597 );
buf g9d6b_GF_PartitionCandidate( \43105_nG9d6b , \43104 );
buf \U$42676 ( \43106 , \43105_nG9d6b );
xor \U$42677 ( \43107 , \24765 , \42872 );
buf g9dff_GF_PartitionCandidate( \43108_nG9dff , \43107 );
buf \U$42678 ( \43109 , \43108_nG9dff );
and \U$42679 ( \43110 , \43106 , \43109 );
xor \U$42680 ( \43111 , \3661 , \21595 );
buf g9c34_GF_PartitionCandidate( \43112_nG9c34 , \43111 );
buf \U$42681 ( \43113 , \43112_nG9c34 );
xor \U$42682 ( \43114 , \24936 , \42870 );
buf g9ccf_GF_PartitionCandidate( \43115_nG9ccf , \43114 );
buf \U$42683 ( \43116 , \43115_nG9ccf );
and \U$42684 ( \43117 , \43113 , \43116 );
xor \U$42685 ( \43118 , \3842 , \21593 );
buf g9af1_GF_PartitionCandidate( \43119_nG9af1 , \43118 );
buf \U$42686 ( \43120 , \43119_nG9af1 );
xor \U$42687 ( \43121 , \25117 , \42868 );
buf g9b91_GF_PartitionCandidate( \43122_nG9b91 , \43121 );
buf \U$42688 ( \43123 , \43122_nG9b91 );
and \U$42689 ( \43124 , \43120 , \43123 );
xor \U$42690 ( \43125 , \4019 , \21591 );
buf g99a6_GF_PartitionCandidate( \43126_nG99a6 , \43125 );
buf \U$42691 ( \43127 , \43126_nG99a6 );
xor \U$42692 ( \43128 , \25294 , \42866 );
buf g9a49_GF_PartitionCandidate( \43129_nG9a49 , \43128 );
buf \U$42693 ( \43130 , \43129_nG9a49 );
and \U$42694 ( \43131 , \43127 , \43130 );
xor \U$42695 ( \43132 , \4216 , \21589 );
buf g9856_GF_PartitionCandidate( \43133_nG9856 , \43132 );
buf \U$42696 ( \43134 , \43133_nG9856 );
xor \U$42697 ( \43135 , \25491 , \42864 );
buf g98fb_GF_PartitionCandidate( \43136_nG98fb , \43135 );
buf \U$42698 ( \43137 , \43136_nG98fb );
and \U$42699 ( \43138 , \43134 , \43137 );
xor \U$42700 ( \43139 , \4412 , \21587 );
buf g96ff_GF_PartitionCandidate( \43140_nG96ff , \43139 );
buf \U$42701 ( \43141 , \43140_nG96ff );
xor \U$42702 ( \43142 , \25687 , \42862 );
buf g97a9_GF_PartitionCandidate( \43143_nG97a9 , \43142 );
buf \U$42703 ( \43144 , \43143_nG97a9 );
and \U$42704 ( \43145 , \43141 , \43144 );
xor \U$42705 ( \43146 , \4614 , \21585 );
buf g95a0_GF_PartitionCandidate( \43147_nG95a0 , \43146 );
buf \U$42706 ( \43148 , \43147_nG95a0 );
xor \U$42707 ( \43149 , \25889 , \42860 );
buf g964d_GF_PartitionCandidate( \43150_nG964d , \43149 );
buf \U$42708 ( \43151 , \43150_nG964d );
and \U$42709 ( \43152 , \43148 , \43151 );
xor \U$42710 ( \43153 , \4821 , \21583 );
buf g9436_GF_PartitionCandidate( \43154_nG9436 , \43153 );
buf \U$42711 ( \43155 , \43154_nG9436 );
xor \U$42712 ( \43156 , \26096 , \42858 );
buf g94eb_GF_PartitionCandidate( \43157_nG94eb , \43156 );
buf \U$42713 ( \43158 , \43157_nG94eb );
and \U$42714 ( \43159 , \43155 , \43158 );
xor \U$42715 ( \43160 , \5031 , \21581 );
buf g92bf_GF_PartitionCandidate( \43161_nG92bf , \43160 );
buf \U$42716 ( \43162 , \43161_nG92bf );
xor \U$42717 ( \43163 , \26306 , \42856 );
buf g9379_GF_PartitionCandidate( \43164_nG9379 , \43163 );
buf \U$42718 ( \43165 , \43164_nG9379 );
and \U$42719 ( \43166 , \43162 , \43165 );
xor \U$42720 ( \43167 , \5460 , \21579 );
buf g913c_GF_PartitionCandidate( \43168_nG913c , \43167 );
buf \U$42721 ( \43169 , \43168_nG913c );
xor \U$42722 ( \43170 , \26735 , \42854 );
buf g91fd_GF_PartitionCandidate( \43171_nG91fd , \43170 );
buf \U$42723 ( \43172 , \43171_nG91fd );
and \U$42724 ( \43173 , \43169 , \43172 );
xor \U$42725 ( \43174 , \5703 , \21577 );
buf g8fb0_GF_PartitionCandidate( \43175_nG8fb0 , \43174 );
buf \U$42726 ( \43176 , \43175_nG8fb0 );
xor \U$42727 ( \43177 , \26978 , \42852 );
buf g9073_GF_PartitionCandidate( \43178_nG9073 , \43177 );
buf \U$42728 ( \43179 , \43178_nG9073 );
and \U$42729 ( \43180 , \43176 , \43179 );
xor \U$42730 ( \43181 , \5935 , \21575 );
buf g8e1a_GF_PartitionCandidate( \43182_nG8e1a , \43181 );
buf \U$42731 ( \43183 , \43182_nG8e1a );
xor \U$42732 ( \43184 , \27210 , \42850 );
buf g8ee5_GF_PartitionCandidate( \43185_nG8ee5 , \43184 );
buf \U$42733 ( \43186 , \43185_nG8ee5 );
and \U$42734 ( \43187 , \43183 , \43186 );
xor \U$42735 ( \43188 , \6183 , \21573 );
buf g8c7a_GF_PartitionCandidate( \43189_nG8c7a , \43188 );
buf \U$42736 ( \43190 , \43189_nG8c7a );
xor \U$42737 ( \43191 , \27458 , \42848 );
buf g8d47_GF_PartitionCandidate( \43192_nG8d47 , \43191 );
buf \U$42738 ( \43193 , \43192_nG8d47 );
and \U$42739 ( \43194 , \43190 , \43193 );
xor \U$42740 ( \43195 , \6436 , \21571 );
buf g8ad0_GF_PartitionCandidate( \43196_nG8ad0 , \43195 );
buf \U$42741 ( \43197 , \43196_nG8ad0 );
xor \U$42742 ( \43198 , \27711 , \42846 );
buf g8ba5_GF_PartitionCandidate( \43199_nG8ba5 , \43198 );
buf \U$42743 ( \43200 , \43199_nG8ba5 );
and \U$42744 ( \43201 , \43197 , \43200 );
xor \U$42745 ( \43202 , \6692 , \21569 );
buf g8919_GF_PartitionCandidate( \43203_nG8919 , \43202 );
buf \U$42746 ( \43204 , \43203_nG8919 );
xor \U$42747 ( \43205 , \27967 , \42844 );
buf g89f3_GF_PartitionCandidate( \43206_nG89f3 , \43205 );
buf \U$42748 ( \43207 , \43206_nG89f3 );
and \U$42749 ( \43208 , \43204 , \43207 );
xor \U$42750 ( \43209 , \6949 , \21567 );
buf g8757_GF_PartitionCandidate( \43210_nG8757 , \43209 );
buf \U$42751 ( \43211 , \43210_nG8757 );
xor \U$42752 ( \43212 , \28224 , \42842 );
buf g8837_GF_PartitionCandidate( \43213_nG8837 , \43212 );
buf \U$42753 ( \43214 , \43213_nG8837 );
and \U$42754 ( \43215 , \43211 , \43214 );
xor \U$42755 ( \43216 , \7212 , \21565 );
buf g858b_GF_PartitionCandidate( \43217_nG858b , \43216 );
buf \U$42756 ( \43218 , \43217_nG858b );
xor \U$42757 ( \43219 , \28487 , \42840 );
buf g866f_GF_PartitionCandidate( \43220_nG866f , \43219 );
buf \U$42758 ( \43221 , \43220_nG866f );
and \U$42759 ( \43222 , \43218 , \43221 );
xor \U$42760 ( \43223 , \7477 , \21563 );
buf g83b4_GF_PartitionCandidate( \43224_nG83b4 , \43223 );
buf \U$42761 ( \43225 , \43224_nG83b4 );
xor \U$42762 ( \43226 , \28752 , \42838 );
buf g849f_GF_PartitionCandidate( \43227_nG849f , \43226 );
buf \U$42763 ( \43228 , \43227_nG849f );
and \U$42764 ( \43229 , \43225 , \43228 );
xor \U$42765 ( \43230 , \7738 , \21561 );
buf g81d4_GF_PartitionCandidate( \43231_nG81d4 , \43230 );
buf \U$42766 ( \43232 , \43231_nG81d4 );
xor \U$42767 ( \43233 , \29013 , \42836 );
buf g82c1_GF_PartitionCandidate( \43234_nG82c1 , \43233 );
buf \U$42768 ( \43235 , \43234_nG82c1 );
and \U$42769 ( \43236 , \43232 , \43235 );
xor \U$42770 ( \43237 , \8004 , \21559 );
buf g7fea_GF_PartitionCandidate( \43238_nG7fea , \43237 );
buf \U$42771 ( \43239 , \43238_nG7fea );
xor \U$42772 ( \43240 , \29279 , \42834 );
buf g80df_GF_PartitionCandidate( \43241_nG80df , \43240 );
buf \U$42773 ( \43242 , \43241_nG80df );
and \U$42774 ( \43243 , \43239 , \43242 );
xor \U$42775 ( \43244 , \8270 , \21557 );
buf g7df3_GF_PartitionCandidate( \43245_nG7df3 , \43244 );
buf \U$42776 ( \43246 , \43245_nG7df3 );
xor \U$42777 ( \43247 , \29545 , \42832 );
buf g7eed_GF_PartitionCandidate( \43248_nG7eed , \43247 );
buf \U$42778 ( \43249 , \43248_nG7eed );
and \U$42779 ( \43250 , \43246 , \43249 );
xor \U$42780 ( \43251 , \8565 , \21555 );
buf g7bf4_GF_PartitionCandidate( \43252_nG7bf4 , \43251 );
buf \U$42781 ( \43253 , \43252_nG7bf4 );
xor \U$42782 ( \43254 , \29840 , \42830 );
buf g7cf1_GF_PartitionCandidate( \43255_nG7cf1 , \43254 );
buf \U$42783 ( \43256 , \43255_nG7cf1 );
and \U$42784 ( \43257 , \43253 , \43256 );
xor \U$42785 ( \43258 , \8848 , \21553 );
buf g79f0_GF_PartitionCandidate( \43259_nG79f0 , \43258 );
buf \U$42786 ( \43260 , \43259_nG79f0 );
xor \U$42787 ( \43261 , \30123 , \42828 );
buf g7aef_GF_PartitionCandidate( \43262_nG7aef , \43261 );
buf \U$42788 ( \43263 , \43262_nG7aef );
and \U$42789 ( \43264 , \43260 , \43263 );
xor \U$42790 ( \43265 , \9136 , \21551 );
buf g77e5_GF_PartitionCandidate( \43266_nG77e5 , \43265 );
buf \U$42791 ( \43267 , \43266_nG77e5 );
xor \U$42792 ( \43268 , \30411 , \42826 );
buf g78e9_GF_PartitionCandidate( \43269_nG78e9 , \43268 );
buf \U$42793 ( \43270 , \43269_nG78e9 );
and \U$42794 ( \43271 , \43267 , \43270 );
xor \U$42795 ( \43272 , \9437 , \21549 );
buf g75cf_GF_PartitionCandidate( \43273_nG75cf , \43272 );
buf \U$42796 ( \43274 , \43273_nG75cf );
xor \U$42797 ( \43275 , \30712 , \42824 );
buf g76d9_GF_PartitionCandidate( \43276_nG76d9 , \43275 );
buf \U$42798 ( \43277 , \43276_nG76d9 );
and \U$42799 ( \43278 , \43274 , \43277 );
xor \U$42800 ( \43279 , \9733 , \21547 );
buf g73af_GF_PartitionCandidate( \43280_nG73af , \43279 );
buf \U$42801 ( \43281 , \43280_nG73af );
xor \U$42802 ( \43282 , \31008 , \42822 );
buf g74bd_GF_PartitionCandidate( \43283_nG74bd , \43282 );
buf \U$42803 ( \43284 , \43283_nG74bd );
and \U$42804 ( \43285 , \43281 , \43284 );
xor \U$42805 ( \43286 , \10042 , \21545 );
buf g7188_GF_PartitionCandidate( \43287_nG7188 , \43286 );
buf \U$42806 ( \43288 , \43287_nG7188 );
xor \U$42807 ( \43289 , \31317 , \42820 );
buf g7299_GF_PartitionCandidate( \43290_nG7299 , \43289 );
buf \U$42808 ( \43291 , \43290_nG7299 );
and \U$42809 ( \43292 , \43288 , \43291 );
xor \U$42810 ( \43293 , \10360 , \21543 );
buf g6f56_GF_PartitionCandidate( \43294_nG6f56 , \43293 );
buf \U$42811 ( \43295 , \43294_nG6f56 );
xor \U$42812 ( \43296 , \31635 , \42818 );
buf g706f_GF_PartitionCandidate( \43297_nG706f , \43296 );
buf \U$42813 ( \43298 , \43297_nG706f );
and \U$42814 ( \43299 , \43295 , \43298 );
xor \U$42815 ( \43300 , \10676 , \21541 );
buf g6d1a_GF_PartitionCandidate( \43301_nG6d1a , \43300 );
buf \U$42816 ( \43302 , \43301_nG6d1a );
xor \U$42817 ( \43303 , \31951 , \42816 );
buf g6e35_GF_PartitionCandidate( \43304_nG6e35 , \43303 );
buf \U$42818 ( \43305 , \43304_nG6e35 );
and \U$42819 ( \43306 , \43302 , \43305 );
xor \U$42820 ( \43307 , \10989 , \21539 );
buf g6ad4_GF_PartitionCandidate( \43308_nG6ad4 , \43307 );
buf \U$42821 ( \43309 , \43308_nG6ad4 );
xor \U$42822 ( \43310 , \32264 , \42814 );
buf g6bf7_GF_PartitionCandidate( \43311_nG6bf7 , \43310 );
buf \U$42823 ( \43312 , \43311_nG6bf7 );
and \U$42824 ( \43313 , \43309 , \43312 );
xor \U$42825 ( \43314 , \11300 , \21537 );
buf g6881_GF_PartitionCandidate( \43315_nG6881 , \43314 );
buf \U$42826 ( \43316 , \43315_nG6881 );
xor \U$42827 ( \43317 , \32575 , \42812 );
buf g69a9_GF_PartitionCandidate( \43318_nG69a9 , \43317 );
buf \U$42828 ( \43319 , \43318_nG69a9 );
and \U$42829 ( \43320 , \43316 , \43319 );
xor \U$42830 ( \43321 , \11618 , \21535 );
buf g6622_GF_PartitionCandidate( \43322_nG6622 , \43321 );
buf \U$42831 ( \43323 , \43322_nG6622 );
xor \U$42832 ( \43324 , \32893 , \42810 );
buf g6751_GF_PartitionCandidate( \43325_nG6751 , \43324 );
buf \U$42833 ( \43326 , \43325_nG6751 );
and \U$42834 ( \43327 , \43323 , \43326 );
xor \U$42835 ( \43328 , \11934 , \21533 );
buf g63b7_GF_PartitionCandidate( \43329_nG63b7 , \43328 );
buf \U$42836 ( \43330 , \43329_nG63b7 );
xor \U$42837 ( \43331 , \33209 , \42808 );
buf g64eb_GF_PartitionCandidate( \43332_nG64eb , \43331 );
buf \U$42838 ( \43333 , \43332_nG64eb );
and \U$42839 ( \43334 , \43330 , \43333 );
xor \U$42840 ( \43335 , \12234 , \21531 );
buf g6144_GF_PartitionCandidate( \43336_nG6144 , \43335 );
buf \U$42841 ( \43337 , \43336_nG6144 );
xor \U$42842 ( \43338 , \33509 , \42806 );
buf g627b_GF_PartitionCandidate( \43339_nG627b , \43338 );
buf \U$42843 ( \43340 , \43339_nG627b );
and \U$42844 ( \43341 , \43337 , \43340 );
xor \U$42845 ( \43342 , \12550 , \21529 );
buf g5ec9_GF_PartitionCandidate( \43343_nG5ec9 , \43342 );
buf \U$42846 ( \43344 , \43343_nG5ec9 );
xor \U$42847 ( \43345 , \33825 , \42804 );
buf g6005_GF_PartitionCandidate( \43346_nG6005 , \43345 );
buf \U$42848 ( \43347 , \43346_nG6005 );
and \U$42849 ( \43348 , \43344 , \43347 );
xor \U$42850 ( \43349 , \12835 , \21527 );
buf g5c48_GF_PartitionCandidate( \43350_nG5c48 , \43349 );
buf \U$42851 ( \43351 , \43350_nG5c48 );
xor \U$42852 ( \43352 , \34110 , \42802 );
buf g5d85_GF_PartitionCandidate( \43353_nG5d85 , \43352 );
buf \U$42853 ( \43354 , \43353_nG5d85 );
and \U$42854 ( \43355 , \43351 , \43354 );
xor \U$42855 ( \43356 , \13114 , \21525 );
buf g59c5_GF_PartitionCandidate( \43357_nG59c5 , \43356 );
buf \U$42856 ( \43358 , \43357_nG59c5 );
xor \U$42857 ( \43359 , \34389 , \42800 );
buf g5b03_GF_PartitionCandidate( \43360_nG5b03 , \43359 );
buf \U$42858 ( \43361 , \43360_nG5b03 );
and \U$42859 ( \43362 , \43358 , \43361 );
xor \U$42860 ( \43363 , \13417 , \21523 );
buf g5740_GF_PartitionCandidate( \43364_nG5740 , \43363 );
buf \U$42861 ( \43365 , \43364_nG5740 );
xor \U$42862 ( \43366 , \34692 , \42798 );
buf g587f_GF_PartitionCandidate( \43367_nG587f , \43366 );
buf \U$42863 ( \43368 , \43367_nG587f );
and \U$42864 ( \43369 , \43365 , \43368 );
xor \U$42865 ( \43370 , \13688 , \21521 );
buf g54b8_GF_PartitionCandidate( \43371_nG54b8 , \43370 );
buf \U$42866 ( \43372 , \43371_nG54b8 );
xor \U$42867 ( \43373 , \34963 , \42796 );
buf g55f9_GF_PartitionCandidate( \43374_nG55f9 , \43373 );
buf \U$42868 ( \43375 , \43374_nG55f9 );
and \U$42869 ( \43376 , \43372 , \43375 );
xor \U$42870 ( \43377 , \13964 , \21519 );
buf g5231_GF_PartitionCandidate( \43378_nG5231 , \43377 );
buf \U$42871 ( \43379 , \43378_nG5231 );
xor \U$42872 ( \43380 , \35239 , \42794 );
buf g536f_GF_PartitionCandidate( \43381_nG536f , \43380 );
buf \U$42873 ( \43382 , \43381_nG536f );
and \U$42874 ( \43383 , \43379 , \43382 );
xor \U$42875 ( \43384 , \14241 , \21517 );
buf g4fb4_GF_PartitionCandidate( \43385_nG4fb4 , \43384 );
buf \U$42876 ( \43386 , \43385_nG4fb4 );
xor \U$42877 ( \43387 , \35516 , \42792 );
buf g50eb_GF_PartitionCandidate( \43388_nG50eb , \43387 );
buf \U$42878 ( \43389 , \43388_nG50eb );
and \U$42879 ( \43390 , \43386 , \43389 );
xor \U$42880 ( \43391 , \14511 , \21515 );
buf g4d41_GF_PartitionCandidate( \43392_nG4d41 , \43391 );
buf \U$42881 ( \43393 , \43392_nG4d41 );
xor \U$42882 ( \43394 , \35786 , \42790 );
buf g4e75_GF_PartitionCandidate( \43395_nG4e75 , \43394 );
buf \U$42883 ( \43396 , \43395_nG4e75 );
and \U$42884 ( \43397 , \43393 , \43396 );
xor \U$42885 ( \43398 , \14773 , \21513 );
buf g4ad8_GF_PartitionCandidate( \43399_nG4ad8 , \43398 );
buf \U$42886 ( \43400 , \43399_nG4ad8 );
xor \U$42887 ( \43401 , \36048 , \42788 );
buf g4c05_GF_PartitionCandidate( \43402_nG4c05 , \43401 );
buf \U$42888 ( \43403 , \43402_nG4c05 );
and \U$42889 ( \43404 , \43400 , \43403 );
xor \U$42890 ( \43405 , \15034 , \21511 );
buf g4879_GF_PartitionCandidate( \43406_nG4879 , \43405 );
buf \U$42891 ( \43407 , \43406_nG4879 );
xor \U$42892 ( \43408 , \36309 , \42786 );
buf g49a3_GF_PartitionCandidate( \43409_nG49a3 , \43408 );
buf \U$42893 ( \43410 , \43409_nG49a3 );
and \U$42894 ( \43411 , \43407 , \43410 );
xor \U$42895 ( \43412 , \15042 , \21509 );
buf g4624_GF_PartitionCandidate( \43413_nG4624 , \43412 );
buf \U$42896 ( \43414 , \43413_nG4624 );
xor \U$42897 ( \43415 , \36317 , \42784 );
buf g4747_GF_PartitionCandidate( \43416_nG4747 , \43415 );
buf \U$42898 ( \43417 , \43416_nG4747 );
and \U$42899 ( \43418 , \43414 , \43417 );
xor \U$42900 ( \43419 , \15288 , \21507 );
buf g43d9_GF_PartitionCandidate( \43420_nG43d9 , \43419 );
buf \U$42901 ( \43421 , \43420_nG43d9 );
xor \U$42902 ( \43422 , \36563 , \42782 );
buf g44f9_GF_PartitionCandidate( \43423_nG44f9 , \43422 );
buf \U$42903 ( \43424 , \43423_nG44f9 );
and \U$42904 ( \43425 , \43421 , \43424 );
xor \U$42905 ( \43426 , \15518 , \21505 );
buf g4198_GF_PartitionCandidate( \43427_nG4198 , \43426 );
buf \U$42906 ( \43428 , \43427_nG4198 );
xor \U$42907 ( \43429 , \36793 , \42780 );
buf g42b1_GF_PartitionCandidate( \43430_nG42b1 , \43429 );
buf \U$42908 ( \43431 , \43430_nG42b1 );
and \U$42909 ( \43432 , \43428 , \43431 );
xor \U$42910 ( \43433 , \15768 , \21503 );
buf g3f61_GF_PartitionCandidate( \43434_nG3f61 , \43433 );
buf \U$42911 ( \43435 , \43434_nG3f61 );
xor \U$42912 ( \43436 , \37043 , \42778 );
buf g4077_GF_PartitionCandidate( \43437_nG4077 , \43436 );
buf \U$42913 ( \43438 , \43437_nG4077 );
and \U$42914 ( \43439 , \43435 , \43438 );
xor \U$42915 ( \43440 , \15993 , \21501 );
buf g3d34_GF_PartitionCandidate( \43441_nG3d34 , \43440 );
buf \U$42916 ( \43442 , \43441_nG3d34 );
xor \U$42917 ( \43443 , \37268 , \42776 );
buf g3e43_GF_PartitionCandidate( \43444_nG3e43 , \43443 );
buf \U$42918 ( \43445 , \43444_nG3e43 );
and \U$42919 ( \43446 , \43442 , \43445 );
xor \U$42920 ( \43447 , \16212 , \21499 );
buf g3b11_GF_PartitionCandidate( \43448_nG3b11 , \43447 );
buf \U$42921 ( \43449 , \43448_nG3b11 );
xor \U$42922 ( \43450 , \37487 , \42774 );
buf g3c1d_GF_PartitionCandidate( \43451_nG3c1d , \43450 );
buf \U$42923 ( \43452 , \43451_nG3c1d );
and \U$42924 ( \43453 , \43449 , \43452 );
xor \U$42925 ( \43454 , \16442 , \21497 );
buf g38f8_GF_PartitionCandidate( \43455_nG38f8 , \43454 );
buf \U$42926 ( \43456 , \43455_nG38f8 );
xor \U$42927 ( \43457 , \37717 , \42772 );
buf g39fd_GF_PartitionCandidate( \43458_nG39fd , \43457 );
buf \U$42928 ( \43459 , \43458_nG39fd );
and \U$42929 ( \43460 , \43456 , \43459 );
xor \U$42930 ( \43461 , \16673 , \21495 );
buf g36e9_GF_PartitionCandidate( \43462_nG36e9 , \43461 );
buf \U$42931 ( \43463 , \43462_nG36e9 );
xor \U$42932 ( \43464 , \37948 , \42770 );
buf g37eb_GF_PartitionCandidate( \43465_nG37eb , \43464 );
buf \U$42933 ( \43466 , \43465_nG37eb );
and \U$42934 ( \43467 , \43463 , \43466 );
xor \U$42935 ( \43468 , \16884 , \21493 );
buf g34e4_GF_PartitionCandidate( \43469_nG34e4 , \43468 );
buf \U$42936 ( \43470 , \43469_nG34e4 );
xor \U$42937 ( \43471 , \38159 , \42768 );
buf g35df_GF_PartitionCandidate( \43472_nG35df , \43471 );
buf \U$42938 ( \43473 , \43472_nG35df );
and \U$42939 ( \43474 , \43470 , \43473 );
xor \U$42940 ( \43475 , \17097 , \21491 );
buf g32e9_GF_PartitionCandidate( \43476_nG32e9 , \43475 );
buf \U$42941 ( \43477 , \43476_nG32e9 );
xor \U$42942 ( \43478 , \38372 , \42766 );
buf g33e1_GF_PartitionCandidate( \43479_nG33e1 , \43478 );
buf \U$42943 ( \43480 , \43479_nG33e1 );
and \U$42944 ( \43481 , \43477 , \43480 );
xor \U$42945 ( \43482 , \17294 , \21489 );
buf g30f8_GF_PartitionCandidate( \43483_nG30f8 , \43482 );
buf \U$42946 ( \43484 , \43483_nG30f8 );
xor \U$42947 ( \43485 , \38569 , \42764 );
buf g31e9_GF_PartitionCandidate( \43486_nG31e9 , \43485 );
buf \U$42948 ( \43487 , \43486_nG31e9 );
and \U$42949 ( \43488 , \43484 , \43487 );
xor \U$42950 ( \43489 , \17490 , \21487 );
buf g2f11_GF_PartitionCandidate( \43490_nG2f11 , \43489 );
buf \U$42951 ( \43491 , \43490_nG2f11 );
xor \U$42952 ( \43492 , \38765 , \42762 );
buf g2fff_GF_PartitionCandidate( \43493_nG2fff , \43492 );
buf \U$42953 ( \43494 , \43493_nG2fff );
and \U$42954 ( \43495 , \43491 , \43494 );
xor \U$42955 ( \43496 , \17698 , \21485 );
buf g2d34_GF_PartitionCandidate( \43497_nG2d34 , \43496 );
buf \U$42956 ( \43498 , \43497_nG2d34 );
xor \U$42957 ( \43499 , \38973 , \42760 );
buf g2e1b_GF_PartitionCandidate( \43500_nG2e1b , \43499 );
buf \U$42958 ( \43501 , \43500_nG2e1b );
and \U$42959 ( \43502 , \43498 , \43501 );
xor \U$42960 ( \43503 , \17883 , \21483 );
buf g2b5e_GF_PartitionCandidate( \43504_nG2b5e , \43503 );
buf \U$42961 ( \43505 , \43504_nG2b5e );
xor \U$42962 ( \43506 , \39158 , \42758 );
buf g2c45_GF_PartitionCandidate( \43507_nG2c45 , \43506 );
buf \U$42963 ( \43508 , \43507_nG2c45 );
and \U$42964 ( \43509 , \43505 , \43508 );
xor \U$42965 ( \43510 , \18070 , \21481 );
buf g2993_GF_PartitionCandidate( \43511_nG2993 , \43510 );
buf \U$42966 ( \43512 , \43511_nG2993 );
xor \U$42967 ( \43513 , \39345 , \42756 );
buf g2a6f_GF_PartitionCandidate( \43514_nG2a6f , \43513 );
buf \U$42968 ( \43515 , \43514_nG2a6f );
and \U$42969 ( \43516 , \43512 , \43515 );
xor \U$42970 ( \43517 , \18260 , \21479 );
buf g27d5_GF_PartitionCandidate( \43518_nG27d5 , \43517 );
buf \U$42971 ( \43519 , \43518_nG27d5 );
xor \U$42972 ( \43520 , \39535 , \42754 );
buf g28af_GF_PartitionCandidate( \43521_nG28af , \43520 );
buf \U$42973 ( \43522 , \43521_nG28af );
and \U$42974 ( \43523 , \43519 , \43522 );
xor \U$42975 ( \43524 , \18436 , \21477 );
buf g2620_GF_PartitionCandidate( \43525_nG2620 , \43524 );
buf \U$42976 ( \43526 , \43525_nG2620 );
xor \U$42977 ( \43527 , \39711 , \42752 );
buf g26f3_GF_PartitionCandidate( \43528_nG26f3 , \43527 );
buf \U$42978 ( \43529 , \43528_nG26f3 );
and \U$42979 ( \43530 , \43526 , \43529 );
xor \U$42980 ( \43531 , \18607 , \21475 );
buf g2475_GF_PartitionCandidate( \43532_nG2475 , \43531 );
buf \U$42981 ( \43533 , \43532_nG2475 );
xor \U$42982 ( \43534 , \39882 , \42750 );
buf g2545_GF_PartitionCandidate( \43535_nG2545 , \43534 );
buf \U$42983 ( \43536 , \43535_nG2545 );
and \U$42984 ( \43537 , \43533 , \43536 );
xor \U$42985 ( \43538 , \18615 , \21473 );
buf g22d4_GF_PartitionCandidate( \43539_nG22d4 , \43538 );
buf \U$42986 ( \43540 , \43539_nG22d4 );
xor \U$42987 ( \43541 , \39890 , \42748 );
buf g239d_GF_PartitionCandidate( \43542_nG239d , \43541 );
buf \U$42988 ( \43543 , \43542_nG239d );
and \U$42989 ( \43544 , \43540 , \43543 );
xor \U$42990 ( \43545 , \18783 , \21471 );
buf g213d_GF_PartitionCandidate( \43546_nG213d , \43545 );
buf \U$42991 ( \43547 , \43546_nG213d );
xor \U$42992 ( \43548 , \40058 , \42746 );
buf g2203_GF_PartitionCandidate( \43549_nG2203 , \43548 );
buf \U$42993 ( \43550 , \43549_nG2203 );
and \U$42994 ( \43551 , \43547 , \43550 );
xor \U$42995 ( \43552 , \18923 , \21469 );
buf g1fb0_GF_PartitionCandidate( \43553_nG1fb0 , \43552 );
buf \U$42996 ( \43554 , \43553_nG1fb0 );
xor \U$42997 ( \43555 , \40198 , \42744 );
buf g206f_GF_PartitionCandidate( \43556_nG206f , \43555 );
buf \U$42998 ( \43557 , \43556_nG206f );
and \U$42999 ( \43558 , \43554 , \43557 );
xor \U$43000 ( \43559 , \19075 , \21467 );
buf g1e2d_GF_PartitionCandidate( \43560_nG1e2d , \43559 );
buf \U$43001 ( \43561 , \43560_nG1e2d );
xor \U$43002 ( \43562 , \40350 , \42742 );
buf g1ee9_GF_PartitionCandidate( \43563_nG1ee9 , \43562 );
buf \U$43003 ( \43564 , \43563_nG1ee9 );
and \U$43004 ( \43565 , \43561 , \43564 );
xor \U$43005 ( \43566 , \19239 , \21465 );
buf g1cb4_GF_PartitionCandidate( \43567_nG1cb4 , \43566 );
buf \U$43006 ( \43568 , \43567_nG1cb4 );
xor \U$43007 ( \43569 , \40514 , \42740 );
buf g1d69_GF_PartitionCandidate( \43570_nG1d69 , \43569 );
buf \U$43008 ( \43571 , \43570_nG1d69 );
and \U$43009 ( \43572 , \43568 , \43571 );
xor \U$43010 ( \43573 , \19378 , \21463 );
buf g1b45_GF_PartitionCandidate( \43574_nG1b45 , \43573 );
buf \U$43011 ( \43575 , \43574_nG1b45 );
xor \U$43012 ( \43576 , \40653 , \42738 );
buf g1bf7_GF_PartitionCandidate( \43577_nG1bf7 , \43576 );
buf \U$43013 ( \43578 , \43577_nG1bf7 );
and \U$43014 ( \43579 , \43575 , \43578 );
xor \U$43015 ( \43580 , \19503 , \21461 );
buf g19e0_GF_PartitionCandidate( \43581_nG19e0 , \43580 );
buf \U$43016 ( \43582 , \43581_nG19e0 );
xor \U$43017 ( \43583 , \40778 , \42736 );
buf g1a8b_GF_PartitionCandidate( \43584_nG1a8b , \43583 );
buf \U$43018 ( \43585 , \43584_nG1a8b );
and \U$43019 ( \43586 , \43582 , \43585 );
xor \U$43020 ( \43587 , \19647 , \21459 );
buf g1885_GF_PartitionCandidate( \43588_nG1885 , \43587 );
buf \U$43021 ( \43589 , \43588_nG1885 );
xor \U$43022 ( \43590 , \40922 , \42734 );
buf g192d_GF_PartitionCandidate( \43591_nG192d , \43590 );
buf \U$43023 ( \43592 , \43591_nG192d );
and \U$43024 ( \43593 , \43589 , \43592 );
xor \U$43025 ( \43594 , \19771 , \21457 );
buf g1734_GF_PartitionCandidate( \43595_nG1734 , \43594 );
buf \U$43026 ( \43596 , \43595_nG1734 );
xor \U$43027 ( \43597 , \41046 , \42732 );
buf g17d5_GF_PartitionCandidate( \43598_nG17d5 , \43597 );
buf \U$43028 ( \43599 , \43598_nG17d5 );
and \U$43029 ( \43600 , \43596 , \43599 );
xor \U$43030 ( \43601 , \19911 , \21455 );
buf g15ed_GF_PartitionCandidate( \43602_nG15ed , \43601 );
buf \U$43031 ( \43603 , \43602_nG15ed );
xor \U$43032 ( \43604 , \41186 , \42730 );
buf g168b_GF_PartitionCandidate( \43605_nG168b , \43604 );
buf \U$43033 ( \43606 , \43605_nG168b );
and \U$43034 ( \43607 , \43603 , \43606 );
xor \U$43035 ( \43608 , \20035 , \21453 );
buf g14b0_GF_PartitionCandidate( \43609_nG14b0 , \43608 );
buf \U$43036 ( \43610 , \43609_nG14b0 );
xor \U$43037 ( \43611 , \41310 , \42728 );
buf g1547_GF_PartitionCandidate( \43612_nG1547 , \43611 );
buf \U$43038 ( \43613 , \43612_nG1547 );
and \U$43039 ( \43614 , \43610 , \43613 );
xor \U$43040 ( \43615 , \20150 , \21451 );
buf g137d_GF_PartitionCandidate( \43616_nG137d , \43615 );
buf \U$43041 ( \43617 , \43616_nG137d );
xor \U$43042 ( \43618 , \41425 , \42726 );
buf g1411_GF_PartitionCandidate( \43619_nG1411 , \43618 );
buf \U$43043 ( \43620 , \43619_nG1411 );
and \U$43044 ( \43621 , \43617 , \43620 );
xor \U$43045 ( \43622 , \20158 , \21449 );
buf g1254_GF_PartitionCandidate( \43623_nG1254 , \43622 );
buf \U$43046 ( \43624 , \43623_nG1254 );
xor \U$43047 ( \43625 , \41433 , \42724 );
buf g12e1_GF_PartitionCandidate( \43626_nG12e1 , \43625 );
buf \U$43048 ( \43627 , \43626_nG12e1 );
and \U$43049 ( \43628 , \43624 , \43627 );
xor \U$43050 ( \43629 , \20254 , \21447 );
buf g1135_GF_PartitionCandidate( \43630_nG1135 , \43629 );
buf \U$43051 ( \43631 , \43630_nG1135 );
xor \U$43052 ( \43632 , \41529 , \42722 );
buf g11bf_GF_PartitionCandidate( \43633_nG11bf , \43632 );
buf \U$43053 ( \43634 , \43633_nG11bf );
and \U$43054 ( \43635 , \43631 , \43634 );
xor \U$43055 ( \43636 , \20369 , \21445 );
buf g1020_GF_PartitionCandidate( \43637_nG1020 , \43636 );
buf \U$43056 ( \43638 , \43637_nG1020 );
xor \U$43057 ( \43639 , \41644 , \42720 );
buf g10a3_GF_PartitionCandidate( \43640_nG10a3 , \43639 );
buf \U$43058 ( \43641 , \43640_nG10a3 );
and \U$43059 ( \43642 , \43638 , \43641 );
xor \U$43060 ( \43643 , \20457 , \21443 );
buf gf15_GF_PartitionCandidate( \43644_nGf15 , \43643 );
buf \U$43061 ( \43645 , \43644_nGf15 );
xor \U$43062 ( \43646 , \41732 , \42718 );
buf gf95_GF_PartitionCandidate( \43647_nGf95 , \43646 );
buf \U$43063 ( \43648 , \43647_nGf95 );
and \U$43064 ( \43649 , \43645 , \43648 );
xor \U$43065 ( \43650 , \20549 , \21441 );
buf ge14_GF_PartitionCandidate( \43651_nGe14 , \43650 );
buf \U$43066 ( \43652 , \43651_nGe14 );
xor \U$43067 ( \43653 , \41824 , \42716 );
buf ge8d_GF_PartitionCandidate( \43654_nGe8d , \43653 );
buf \U$43068 ( \43655 , \43654_nGe8d );
and \U$43069 ( \43656 , \43652 , \43655 );
xor \U$43070 ( \43657 , \20637 , \21439 );
buf gd1d_GF_PartitionCandidate( \43658_nGd1d , \43657 );
buf \U$43071 ( \43659 , \43658_nGd1d );
xor \U$43072 ( \43660 , \41912 , \42714 );
buf gd93_GF_PartitionCandidate( \43661_nGd93 , \43660 );
buf \U$43073 ( \43662 , \43661_nGd93 );
and \U$43074 ( \43663 , \43659 , \43662 );
xor \U$43075 ( \43664 , \20732 , \21437 );
buf gc30_GF_PartitionCandidate( \43665_nGc30 , \43664 );
buf \U$43076 ( \43666 , \43665_nGc30 );
xor \U$43077 ( \43667 , \42007 , \42712 );
buf gc9f_GF_PartitionCandidate( \43668_nGc9f , \43667 );
buf \U$43078 ( \43669 , \43668_nGc9f );
and \U$43079 ( \43670 , \43666 , \43669 );
xor \U$43080 ( \43671 , \20812 , \21435 );
buf gb4d_GF_PartitionCandidate( \43672_nGb4d , \43671 );
buf \U$43081 ( \43673 , \43672_nGb4d );
xor \U$43082 ( \43674 , \42087 , \42710 );
buf gbb9_GF_PartitionCandidate( \43675_nGbb9 , \43674 );
buf \U$43083 ( \43676 , \43675_nGbb9 );
and \U$43084 ( \43677 , \43673 , \43676 );
xor \U$43085 ( \43678 , \20891 , \21433 );
buf ga74_GF_PartitionCandidate( \43679_nGa74 , \43678 );
buf \U$43086 ( \43680 , \43679_nGa74 );
xor \U$43087 ( \43681 , \42166 , \42708 );
buf gad9_GF_PartitionCandidate( \43682_nGad9 , \43681 );
buf \U$43088 ( \43683 , \43682_nGad9 );
and \U$43089 ( \43684 , \43680 , \43683 );
xor \U$43090 ( \43685 , \20899 , \21431 );
buf g9a5_GF_PartitionCandidate( \43686_nG9a5 , \43685 );
buf \U$43091 ( \43687 , \43686_nG9a5 );
xor \U$43092 ( \43688 , \42174 , \42706 );
buf ga07_GF_PartitionCandidate( \43689_nGa07 , \43688 );
buf \U$43093 ( \43690 , \43689_nGa07 );
and \U$43094 ( \43691 , \43687 , \43690 );
xor \U$43095 ( \43692 , \20958 , \21429 );
buf g8e0_GF_PartitionCandidate( \43693_nG8e0 , \43692 );
buf \U$43096 ( \43694 , \43693_nG8e0 );
xor \U$43097 ( \43695 , \42233 , \42704 );
buf g93b_GF_PartitionCandidate( \43696_nG93b , \43695 );
buf \U$43098 ( \43697 , \43696_nG93b );
and \U$43099 ( \43698 , \43694 , \43697 );
xor \U$43100 ( \43699 , \21013 , \21427 );
buf g825_GF_PartitionCandidate( \43700_nG825 , \43699 );
buf \U$43101 ( \43701 , \43700_nG825 );
xor \U$43102 ( \43702 , \42288 , \42702 );
buf g87d_GF_PartitionCandidate( \43703_nG87d , \43702 );
buf \U$43103 ( \43704 , \43703_nG87d );
and \U$43104 ( \43705 , \43701 , \43704 );
xor \U$43105 ( \43706 , \21084 , \21425 );
buf g774_GF_PartitionCandidate( \43707_nG774 , \43706 );
buf \U$43106 ( \43708 , \43707_nG774 );
xor \U$43107 ( \43709 , \42359 , \42700 );
buf g7c5_GF_PartitionCandidate( \43710_nG7c5 , \43709 );
buf \U$43108 ( \43711 , \43710_nG7c5 );
and \U$43109 ( \43712 , \43708 , \43711 );
xor \U$43110 ( \43713 , \21137 , \21423 );
buf g6cd_GF_PartitionCandidate( \43714_nG6cd , \43713 );
buf \U$43111 ( \43715 , \43714_nG6cd );
xor \U$43112 ( \43716 , \42412 , \42698 );
buf g71b_GF_PartitionCandidate( \43717_nG71b , \43716 );
buf \U$43113 ( \43718 , \43717_nG71b );
and \U$43114 ( \43719 , \43715 , \43718 );
xor \U$43115 ( \43720 , \21176 , \21421 );
buf g630_GF_PartitionCandidate( \43721_nG630 , \43720 );
buf \U$43116 ( \43722 , \43721_nG630 );
xor \U$43117 ( \43723 , \42451 , \42696 );
buf g677_GF_PartitionCandidate( \43724_nG677 , \43723 );
buf \U$43118 ( \43725 , \43724_nG677 );
and \U$43119 ( \43726 , \43722 , \43725 );
xor \U$43120 ( \43727 , \21229 , \21419 );
buf g59d_GF_PartitionCandidate( \43728_nG59d , \43727 );
buf \U$43121 ( \43729 , \43728_nG59d );
xor \U$43122 ( \43730 , \42504 , \42694 );
buf g5e1_GF_PartitionCandidate( \43731_nG5e1 , \43730 );
buf \U$43123 ( \43732 , \43731_nG5e1 );
and \U$43124 ( \43733 , \43729 , \43732 );
xor \U$43125 ( \43734 , \21237 , \21417 );
buf g514_GF_PartitionCandidate( \43735_nG514 , \43734 );
buf \U$43126 ( \43736 , \43735_nG514 );
xor \U$43127 ( \43737 , \42512 , \42692 );
buf g551_GF_PartitionCandidate( \43738_nG551 , \43737 );
buf \U$43128 ( \43739 , \43738_nG551 );
and \U$43129 ( \43740 , \43736 , \43739 );
xor \U$43130 ( \43741 , \21271 , \21415 );
buf g495_GF_PartitionCandidate( \43742_nG495 , \43741 );
buf \U$43131 ( \43743 , \43742_nG495 );
xor \U$43132 ( \43744 , \42546 , \42690 );
buf g4cf_GF_PartitionCandidate( \43745_nG4cf , \43744 );
buf \U$43133 ( \43746 , \43745_nG4cf );
and \U$43134 ( \43747 , \43743 , \43746 );
xor \U$43135 ( \43748 , \21305 , \21413 );
buf g420_GF_PartitionCandidate( \43749_nG420 , \43748 );
buf \U$43136 ( \43750 , \43749_nG420 );
xor \U$43137 ( \43751 , \42580 , \42688 );
buf g453_GF_PartitionCandidate( \43752_nG453 , \43751 );
buf \U$43138 ( \43753 , \43752_nG453 );
and \U$43139 ( \43754 , \43750 , \43753 );
xor \U$43140 ( \43755 , \21313 , \21411 );
buf g3b5_GF_PartitionCandidate( \43756_nG3b5 , \43755 );
buf \U$43141 ( \43757 , \43756_nG3b5 );
xor \U$43142 ( \43758 , \42588 , \42686 );
buf g3e5_GF_PartitionCandidate( \43759_nG3e5 , \43758 );
buf \U$43143 ( \43760 , \43759_nG3e5 );
and \U$43144 ( \43761 , \43757 , \43760 );
xor \U$43145 ( \43762 , \21339 , \21409 );
buf g354_GF_PartitionCandidate( \43763_nG354 , \43762 );
buf \U$43146 ( \43764 , \43763_nG354 );
xor \U$43147 ( \43765 , \42614 , \42684 );
buf g37d_GF_PartitionCandidate( \43766_nG37d , \43765 );
buf \U$43148 ( \43767 , \43766_nG37d );
and \U$43149 ( \43768 , \43764 , \43767 );
xor \U$43150 ( \43769 , \21358 , \21407 );
buf g2fd_GF_PartitionCandidate( \43770_nG2fd , \43769 );
buf \U$43151 ( \43771 , \43770_nG2fd );
xor \U$43152 ( \43772 , \42633 , \42682 );
buf g323_GF_PartitionCandidate( \43773_nG323 , \43772 );
buf \U$43153 ( \43774 , \43773_nG323 );
and \U$43154 ( \43775 , \43771 , \43774 );
xor \U$43155 ( \43776 , \21366 , \21405 );
buf g2b0_GF_PartitionCandidate( \43777_nG2b0 , \43776 );
buf \U$43156 ( \43778 , \43777_nG2b0 );
xor \U$43157 ( \43779 , \42641 , \42680 );
buf g2cf_GF_PartitionCandidate( \43780_nG2cf , \43779 );
buf \U$43158 ( \43781 , \43780_nG2cf );
and \U$43159 ( \43782 , \43778 , \43781 );
xor \U$43160 ( \43783 , \21378 , \21403 );
buf g26d_GF_PartitionCandidate( \43784_nG26d , \43783 );
buf \U$43161 ( \43785 , \43784_nG26d );
xor \U$43162 ( \43786 , \42653 , \42678 );
buf g289_GF_PartitionCandidate( \43787_nG289 , \43786 );
buf \U$43163 ( \43788 , \43787_nG289 );
and \U$43164 ( \43789 , \43785 , \43788 );
xor \U$43165 ( \43790 , \21386 , \21401 );
buf g234_GF_PartitionCandidate( \43791_nG234 , \43790 );
buf \U$43166 ( \43792 , \43791_nG234 );
xor \U$43167 ( \43793 , \42661 , \42676 );
buf g249_GF_PartitionCandidate( \43794_nG249 , \43793 );
buf \U$43168 ( \43795 , \43794_nG249 );
and \U$43169 ( \43796 , \43792 , \43795 );
xor \U$43170 ( \43797 , \21391 , \21399 );
buf g204_GF_PartitionCandidate( \43798_nG204 , \43797 );
buf \U$43171 ( \43799 , \43798_nG204 );
xor \U$43172 ( \43800 , \42666 , \42674 );
buf g217_GF_PartitionCandidate( \43801_nG217 , \43800 );
buf \U$43173 ( \43802 , \43801_nG217 );
and \U$43174 ( \43803 , \43799 , \43802 );
xor \U$43175 ( \43804 , \21395 , \21398 );
buf g1e0_GF_PartitionCandidate( \43805_nG1e0 , \43804 );
buf \U$43176 ( \43806 , \43805_nG1e0 );
xor \U$43177 ( \43807 , \42670 , \42673 );
buf g1ec_GF_PartitionCandidate( \43808_nG1ec , \43807 );
buf \U$43178 ( \43809 , \43808_nG1ec );
and \U$43179 ( \43810 , \43806 , \43809 );
xor \U$43180 ( \43811 , \21397 , \9821 );
buf g189_GF_PartitionCandidate( \43812_nG189 , \43811 );
buf \U$43181 ( \43813 , \43812_nG189 );
xor \U$43182 ( \43814 , \42672 , \31096 );
buf g191_GF_PartitionCandidate( \43815_nG191 , \43814 );
buf \U$43183 ( \43816 , \43815_nG191 );
and \U$43184 ( \43817 , \43813 , \43816 );
and \U$43185 ( \43818 , \43809 , \43817 );
and \U$43186 ( \43819 , \43806 , \43817 );
or \U$43187 ( \43820 , \43810 , \43818 , \43819 );
and \U$43188 ( \43821 , \43802 , \43820 );
and \U$43189 ( \43822 , \43799 , \43820 );
or \U$43190 ( \43823 , \43803 , \43821 , \43822 );
and \U$43191 ( \43824 , \43795 , \43823 );
and \U$43192 ( \43825 , \43792 , \43823 );
or \U$43193 ( \43826 , \43796 , \43824 , \43825 );
and \U$43194 ( \43827 , \43788 , \43826 );
and \U$43195 ( \43828 , \43785 , \43826 );
or \U$43196 ( \43829 , \43789 , \43827 , \43828 );
and \U$43197 ( \43830 , \43781 , \43829 );
and \U$43198 ( \43831 , \43778 , \43829 );
or \U$43199 ( \43832 , \43782 , \43830 , \43831 );
and \U$43200 ( \43833 , \43774 , \43832 );
and \U$43201 ( \43834 , \43771 , \43832 );
or \U$43202 ( \43835 , \43775 , \43833 , \43834 );
and \U$43203 ( \43836 , \43767 , \43835 );
and \U$43204 ( \43837 , \43764 , \43835 );
or \U$43205 ( \43838 , \43768 , \43836 , \43837 );
and \U$43206 ( \43839 , \43760 , \43838 );
and \U$43207 ( \43840 , \43757 , \43838 );
or \U$43208 ( \43841 , \43761 , \43839 , \43840 );
and \U$43209 ( \43842 , \43753 , \43841 );
and \U$43210 ( \43843 , \43750 , \43841 );
or \U$43211 ( \43844 , \43754 , \43842 , \43843 );
and \U$43212 ( \43845 , \43746 , \43844 );
and \U$43213 ( \43846 , \43743 , \43844 );
or \U$43214 ( \43847 , \43747 , \43845 , \43846 );
and \U$43215 ( \43848 , \43739 , \43847 );
and \U$43216 ( \43849 , \43736 , \43847 );
or \U$43217 ( \43850 , \43740 , \43848 , \43849 );
and \U$43218 ( \43851 , \43732 , \43850 );
and \U$43219 ( \43852 , \43729 , \43850 );
or \U$43220 ( \43853 , \43733 , \43851 , \43852 );
and \U$43221 ( \43854 , \43725 , \43853 );
and \U$43222 ( \43855 , \43722 , \43853 );
or \U$43223 ( \43856 , \43726 , \43854 , \43855 );
and \U$43224 ( \43857 , \43718 , \43856 );
and \U$43225 ( \43858 , \43715 , \43856 );
or \U$43226 ( \43859 , \43719 , \43857 , \43858 );
and \U$43227 ( \43860 , \43711 , \43859 );
and \U$43228 ( \43861 , \43708 , \43859 );
or \U$43229 ( \43862 , \43712 , \43860 , \43861 );
and \U$43230 ( \43863 , \43704 , \43862 );
and \U$43231 ( \43864 , \43701 , \43862 );
or \U$43232 ( \43865 , \43705 , \43863 , \43864 );
and \U$43233 ( \43866 , \43697 , \43865 );
and \U$43234 ( \43867 , \43694 , \43865 );
or \U$43235 ( \43868 , \43698 , \43866 , \43867 );
and \U$43236 ( \43869 , \43690 , \43868 );
and \U$43237 ( \43870 , \43687 , \43868 );
or \U$43238 ( \43871 , \43691 , \43869 , \43870 );
and \U$43239 ( \43872 , \43683 , \43871 );
and \U$43240 ( \43873 , \43680 , \43871 );
or \U$43241 ( \43874 , \43684 , \43872 , \43873 );
and \U$43242 ( \43875 , \43676 , \43874 );
and \U$43243 ( \43876 , \43673 , \43874 );
or \U$43244 ( \43877 , \43677 , \43875 , \43876 );
and \U$43245 ( \43878 , \43669 , \43877 );
and \U$43246 ( \43879 , \43666 , \43877 );
or \U$43247 ( \43880 , \43670 , \43878 , \43879 );
and \U$43248 ( \43881 , \43662 , \43880 );
and \U$43249 ( \43882 , \43659 , \43880 );
or \U$43250 ( \43883 , \43663 , \43881 , \43882 );
and \U$43251 ( \43884 , \43655 , \43883 );
and \U$43252 ( \43885 , \43652 , \43883 );
or \U$43253 ( \43886 , \43656 , \43884 , \43885 );
and \U$43254 ( \43887 , \43648 , \43886 );
and \U$43255 ( \43888 , \43645 , \43886 );
or \U$43256 ( \43889 , \43649 , \43887 , \43888 );
and \U$43257 ( \43890 , \43641 , \43889 );
and \U$43258 ( \43891 , \43638 , \43889 );
or \U$43259 ( \43892 , \43642 , \43890 , \43891 );
and \U$43260 ( \43893 , \43634 , \43892 );
and \U$43261 ( \43894 , \43631 , \43892 );
or \U$43262 ( \43895 , \43635 , \43893 , \43894 );
and \U$43263 ( \43896 , \43627 , \43895 );
and \U$43264 ( \43897 , \43624 , \43895 );
or \U$43265 ( \43898 , \43628 , \43896 , \43897 );
and \U$43266 ( \43899 , \43620 , \43898 );
and \U$43267 ( \43900 , \43617 , \43898 );
or \U$43268 ( \43901 , \43621 , \43899 , \43900 );
and \U$43269 ( \43902 , \43613 , \43901 );
and \U$43270 ( \43903 , \43610 , \43901 );
or \U$43271 ( \43904 , \43614 , \43902 , \43903 );
and \U$43272 ( \43905 , \43606 , \43904 );
and \U$43273 ( \43906 , \43603 , \43904 );
or \U$43274 ( \43907 , \43607 , \43905 , \43906 );
and \U$43275 ( \43908 , \43599 , \43907 );
and \U$43276 ( \43909 , \43596 , \43907 );
or \U$43277 ( \43910 , \43600 , \43908 , \43909 );
and \U$43278 ( \43911 , \43592 , \43910 );
and \U$43279 ( \43912 , \43589 , \43910 );
or \U$43280 ( \43913 , \43593 , \43911 , \43912 );
and \U$43281 ( \43914 , \43585 , \43913 );
and \U$43282 ( \43915 , \43582 , \43913 );
or \U$43283 ( \43916 , \43586 , \43914 , \43915 );
and \U$43284 ( \43917 , \43578 , \43916 );
and \U$43285 ( \43918 , \43575 , \43916 );
or \U$43286 ( \43919 , \43579 , \43917 , \43918 );
and \U$43287 ( \43920 , \43571 , \43919 );
and \U$43288 ( \43921 , \43568 , \43919 );
or \U$43289 ( \43922 , \43572 , \43920 , \43921 );
and \U$43290 ( \43923 , \43564 , \43922 );
and \U$43291 ( \43924 , \43561 , \43922 );
or \U$43292 ( \43925 , \43565 , \43923 , \43924 );
and \U$43293 ( \43926 , \43557 , \43925 );
and \U$43294 ( \43927 , \43554 , \43925 );
or \U$43295 ( \43928 , \43558 , \43926 , \43927 );
and \U$43296 ( \43929 , \43550 , \43928 );
and \U$43297 ( \43930 , \43547 , \43928 );
or \U$43298 ( \43931 , \43551 , \43929 , \43930 );
and \U$43299 ( \43932 , \43543 , \43931 );
and \U$43300 ( \43933 , \43540 , \43931 );
or \U$43301 ( \43934 , \43544 , \43932 , \43933 );
and \U$43302 ( \43935 , \43536 , \43934 );
and \U$43303 ( \43936 , \43533 , \43934 );
or \U$43304 ( \43937 , \43537 , \43935 , \43936 );
and \U$43305 ( \43938 , \43529 , \43937 );
and \U$43306 ( \43939 , \43526 , \43937 );
or \U$43307 ( \43940 , \43530 , \43938 , \43939 );
and \U$43308 ( \43941 , \43522 , \43940 );
and \U$43309 ( \43942 , \43519 , \43940 );
or \U$43310 ( \43943 , \43523 , \43941 , \43942 );
and \U$43311 ( \43944 , \43515 , \43943 );
and \U$43312 ( \43945 , \43512 , \43943 );
or \U$43313 ( \43946 , \43516 , \43944 , \43945 );
and \U$43314 ( \43947 , \43508 , \43946 );
and \U$43315 ( \43948 , \43505 , \43946 );
or \U$43316 ( \43949 , \43509 , \43947 , \43948 );
and \U$43317 ( \43950 , \43501 , \43949 );
and \U$43318 ( \43951 , \43498 , \43949 );
or \U$43319 ( \43952 , \43502 , \43950 , \43951 );
and \U$43320 ( \43953 , \43494 , \43952 );
and \U$43321 ( \43954 , \43491 , \43952 );
or \U$43322 ( \43955 , \43495 , \43953 , \43954 );
and \U$43323 ( \43956 , \43487 , \43955 );
and \U$43324 ( \43957 , \43484 , \43955 );
or \U$43325 ( \43958 , \43488 , \43956 , \43957 );
and \U$43326 ( \43959 , \43480 , \43958 );
and \U$43327 ( \43960 , \43477 , \43958 );
or \U$43328 ( \43961 , \43481 , \43959 , \43960 );
and \U$43329 ( \43962 , \43473 , \43961 );
and \U$43330 ( \43963 , \43470 , \43961 );
or \U$43331 ( \43964 , \43474 , \43962 , \43963 );
and \U$43332 ( \43965 , \43466 , \43964 );
and \U$43333 ( \43966 , \43463 , \43964 );
or \U$43334 ( \43967 , \43467 , \43965 , \43966 );
and \U$43335 ( \43968 , \43459 , \43967 );
and \U$43336 ( \43969 , \43456 , \43967 );
or \U$43337 ( \43970 , \43460 , \43968 , \43969 );
and \U$43338 ( \43971 , \43452 , \43970 );
and \U$43339 ( \43972 , \43449 , \43970 );
or \U$43340 ( \43973 , \43453 , \43971 , \43972 );
and \U$43341 ( \43974 , \43445 , \43973 );
and \U$43342 ( \43975 , \43442 , \43973 );
or \U$43343 ( \43976 , \43446 , \43974 , \43975 );
and \U$43344 ( \43977 , \43438 , \43976 );
and \U$43345 ( \43978 , \43435 , \43976 );
or \U$43346 ( \43979 , \43439 , \43977 , \43978 );
and \U$43347 ( \43980 , \43431 , \43979 );
and \U$43348 ( \43981 , \43428 , \43979 );
or \U$43349 ( \43982 , \43432 , \43980 , \43981 );
and \U$43350 ( \43983 , \43424 , \43982 );
and \U$43351 ( \43984 , \43421 , \43982 );
or \U$43352 ( \43985 , \43425 , \43983 , \43984 );
and \U$43353 ( \43986 , \43417 , \43985 );
and \U$43354 ( \43987 , \43414 , \43985 );
or \U$43355 ( \43988 , \43418 , \43986 , \43987 );
and \U$43356 ( \43989 , \43410 , \43988 );
and \U$43357 ( \43990 , \43407 , \43988 );
or \U$43358 ( \43991 , \43411 , \43989 , \43990 );
and \U$43359 ( \43992 , \43403 , \43991 );
and \U$43360 ( \43993 , \43400 , \43991 );
or \U$43361 ( \43994 , \43404 , \43992 , \43993 );
and \U$43362 ( \43995 , \43396 , \43994 );
and \U$43363 ( \43996 , \43393 , \43994 );
or \U$43364 ( \43997 , \43397 , \43995 , \43996 );
and \U$43365 ( \43998 , \43389 , \43997 );
and \U$43366 ( \43999 , \43386 , \43997 );
or \U$43367 ( \44000 , \43390 , \43998 , \43999 );
and \U$43368 ( \44001 , \43382 , \44000 );
and \U$43369 ( \44002 , \43379 , \44000 );
or \U$43370 ( \44003 , \43383 , \44001 , \44002 );
and \U$43371 ( \44004 , \43375 , \44003 );
and \U$43372 ( \44005 , \43372 , \44003 );
or \U$43373 ( \44006 , \43376 , \44004 , \44005 );
and \U$43374 ( \44007 , \43368 , \44006 );
and \U$43375 ( \44008 , \43365 , \44006 );
or \U$43376 ( \44009 , \43369 , \44007 , \44008 );
and \U$43377 ( \44010 , \43361 , \44009 );
and \U$43378 ( \44011 , \43358 , \44009 );
or \U$43379 ( \44012 , \43362 , \44010 , \44011 );
and \U$43380 ( \44013 , \43354 , \44012 );
and \U$43381 ( \44014 , \43351 , \44012 );
or \U$43382 ( \44015 , \43355 , \44013 , \44014 );
and \U$43383 ( \44016 , \43347 , \44015 );
and \U$43384 ( \44017 , \43344 , \44015 );
or \U$43385 ( \44018 , \43348 , \44016 , \44017 );
and \U$43386 ( \44019 , \43340 , \44018 );
and \U$43387 ( \44020 , \43337 , \44018 );
or \U$43388 ( \44021 , \43341 , \44019 , \44020 );
and \U$43389 ( \44022 , \43333 , \44021 );
and \U$43390 ( \44023 , \43330 , \44021 );
or \U$43391 ( \44024 , \43334 , \44022 , \44023 );
and \U$43392 ( \44025 , \43326 , \44024 );
and \U$43393 ( \44026 , \43323 , \44024 );
or \U$43394 ( \44027 , \43327 , \44025 , \44026 );
and \U$43395 ( \44028 , \43319 , \44027 );
and \U$43396 ( \44029 , \43316 , \44027 );
or \U$43397 ( \44030 , \43320 , \44028 , \44029 );
and \U$43398 ( \44031 , \43312 , \44030 );
and \U$43399 ( \44032 , \43309 , \44030 );
or \U$43400 ( \44033 , \43313 , \44031 , \44032 );
and \U$43401 ( \44034 , \43305 , \44033 );
and \U$43402 ( \44035 , \43302 , \44033 );
or \U$43403 ( \44036 , \43306 , \44034 , \44035 );
and \U$43404 ( \44037 , \43298 , \44036 );
and \U$43405 ( \44038 , \43295 , \44036 );
or \U$43406 ( \44039 , \43299 , \44037 , \44038 );
and \U$43407 ( \44040 , \43291 , \44039 );
and \U$43408 ( \44041 , \43288 , \44039 );
or \U$43409 ( \44042 , \43292 , \44040 , \44041 );
and \U$43410 ( \44043 , \43284 , \44042 );
and \U$43411 ( \44044 , \43281 , \44042 );
or \U$43412 ( \44045 , \43285 , \44043 , \44044 );
and \U$43413 ( \44046 , \43277 , \44045 );
and \U$43414 ( \44047 , \43274 , \44045 );
or \U$43415 ( \44048 , \43278 , \44046 , \44047 );
and \U$43416 ( \44049 , \43270 , \44048 );
and \U$43417 ( \44050 , \43267 , \44048 );
or \U$43418 ( \44051 , \43271 , \44049 , \44050 );
and \U$43419 ( \44052 , \43263 , \44051 );
and \U$43420 ( \44053 , \43260 , \44051 );
or \U$43421 ( \44054 , \43264 , \44052 , \44053 );
and \U$43422 ( \44055 , \43256 , \44054 );
and \U$43423 ( \44056 , \43253 , \44054 );
or \U$43424 ( \44057 , \43257 , \44055 , \44056 );
and \U$43425 ( \44058 , \43249 , \44057 );
and \U$43426 ( \44059 , \43246 , \44057 );
or \U$43427 ( \44060 , \43250 , \44058 , \44059 );
and \U$43428 ( \44061 , \43242 , \44060 );
and \U$43429 ( \44062 , \43239 , \44060 );
or \U$43430 ( \44063 , \43243 , \44061 , \44062 );
and \U$43431 ( \44064 , \43235 , \44063 );
and \U$43432 ( \44065 , \43232 , \44063 );
or \U$43433 ( \44066 , \43236 , \44064 , \44065 );
and \U$43434 ( \44067 , \43228 , \44066 );
and \U$43435 ( \44068 , \43225 , \44066 );
or \U$43436 ( \44069 , \43229 , \44067 , \44068 );
and \U$43437 ( \44070 , \43221 , \44069 );
and \U$43438 ( \44071 , \43218 , \44069 );
or \U$43439 ( \44072 , \43222 , \44070 , \44071 );
and \U$43440 ( \44073 , \43214 , \44072 );
and \U$43441 ( \44074 , \43211 , \44072 );
or \U$43442 ( \44075 , \43215 , \44073 , \44074 );
and \U$43443 ( \44076 , \43207 , \44075 );
and \U$43444 ( \44077 , \43204 , \44075 );
or \U$43445 ( \44078 , \43208 , \44076 , \44077 );
and \U$43446 ( \44079 , \43200 , \44078 );
and \U$43447 ( \44080 , \43197 , \44078 );
or \U$43448 ( \44081 , \43201 , \44079 , \44080 );
and \U$43449 ( \44082 , \43193 , \44081 );
and \U$43450 ( \44083 , \43190 , \44081 );
or \U$43451 ( \44084 , \43194 , \44082 , \44083 );
and \U$43452 ( \44085 , \43186 , \44084 );
and \U$43453 ( \44086 , \43183 , \44084 );
or \U$43454 ( \44087 , \43187 , \44085 , \44086 );
and \U$43455 ( \44088 , \43179 , \44087 );
and \U$43456 ( \44089 , \43176 , \44087 );
or \U$43457 ( \44090 , \43180 , \44088 , \44089 );
and \U$43458 ( \44091 , \43172 , \44090 );
and \U$43459 ( \44092 , \43169 , \44090 );
or \U$43460 ( \44093 , \43173 , \44091 , \44092 );
and \U$43461 ( \44094 , \43165 , \44093 );
and \U$43462 ( \44095 , \43162 , \44093 );
or \U$43463 ( \44096 , \43166 , \44094 , \44095 );
and \U$43464 ( \44097 , \43158 , \44096 );
and \U$43465 ( \44098 , \43155 , \44096 );
or \U$43466 ( \44099 , \43159 , \44097 , \44098 );
and \U$43467 ( \44100 , \43151 , \44099 );
and \U$43468 ( \44101 , \43148 , \44099 );
or \U$43469 ( \44102 , \43152 , \44100 , \44101 );
and \U$43470 ( \44103 , \43144 , \44102 );
and \U$43471 ( \44104 , \43141 , \44102 );
or \U$43472 ( \44105 , \43145 , \44103 , \44104 );
and \U$43473 ( \44106 , \43137 , \44105 );
and \U$43474 ( \44107 , \43134 , \44105 );
or \U$43475 ( \44108 , \43138 , \44106 , \44107 );
and \U$43476 ( \44109 , \43130 , \44108 );
and \U$43477 ( \44110 , \43127 , \44108 );
or \U$43478 ( \44111 , \43131 , \44109 , \44110 );
and \U$43479 ( \44112 , \43123 , \44111 );
and \U$43480 ( \44113 , \43120 , \44111 );
or \U$43481 ( \44114 , \43124 , \44112 , \44113 );
and \U$43482 ( \44115 , \43116 , \44114 );
and \U$43483 ( \44116 , \43113 , \44114 );
or \U$43484 ( \44117 , \43117 , \44115 , \44116 );
and \U$43485 ( \44118 , \43109 , \44117 );
and \U$43486 ( \44119 , \43106 , \44117 );
or \U$43487 ( \44120 , \43110 , \44118 , \44119 );
and \U$43488 ( \44121 , \43102 , \44120 );
and \U$43489 ( \44122 , \43099 , \44120 );
or \U$43490 ( \44123 , \43103 , \44121 , \44122 );
and \U$43491 ( \44124 , \43095 , \44123 );
and \U$43492 ( \44125 , \43092 , \44123 );
or \U$43493 ( \44126 , \43096 , \44124 , \44125 );
and \U$43494 ( \44127 , \43088 , \44126 );
and \U$43495 ( \44128 , \43085 , \44126 );
or \U$43496 ( \44129 , \43089 , \44127 , \44128 );
and \U$43497 ( \44130 , \43081 , \44129 );
and \U$43498 ( \44131 , \43078 , \44129 );
or \U$43499 ( \44132 , \43082 , \44130 , \44131 );
and \U$43500 ( \44133 , \43074 , \44132 );
and \U$43501 ( \44134 , \43071 , \44132 );
or \U$43502 ( \44135 , \43075 , \44133 , \44134 );
and \U$43503 ( \44136 , \43067 , \44135 );
and \U$43504 ( \44137 , \43064 , \44135 );
or \U$43505 ( \44138 , \43068 , \44136 , \44137 );
and \U$43506 ( \44139 , \43060 , \44138 );
and \U$43507 ( \44140 , \43057 , \44138 );
or \U$43508 ( \44141 , \43061 , \44139 , \44140 );
and \U$43509 ( \44142 , \43053 , \44141 );
and \U$43510 ( \44143 , \43050 , \44141 );
or \U$43511 ( \44144 , \43054 , \44142 , \44143 );
and \U$43512 ( \44145 , \43046 , \44144 );
and \U$43513 ( \44146 , \43043 , \44144 );
or \U$43514 ( \44147 , \43047 , \44145 , \44146 );
and \U$43515 ( \44148 , \43039 , \44147 );
and \U$43516 ( \44149 , \43036 , \44147 );
or \U$43517 ( \44150 , \43040 , \44148 , \44149 );
and \U$43518 ( \44151 , \43032 , \44150 );
and \U$43519 ( \44152 , \43029 , \44150 );
or \U$43520 ( \44153 , \43033 , \44151 , \44152 );
and \U$43521 ( \44154 , \43025 , \44153 );
and \U$43522 ( \44155 , \43022 , \44153 );
or \U$43523 ( \44156 , \43026 , \44154 , \44155 );
and \U$43524 ( \44157 , \43018 , \44156 );
and \U$43525 ( \44158 , \43015 , \44156 );
or \U$43526 ( \44159 , \43019 , \44157 , \44158 );
and \U$43527 ( \44160 , \43011 , \44159 );
and \U$43528 ( \44161 , \43008 , \44159 );
or \U$43529 ( \44162 , \43012 , \44160 , \44161 );
and \U$43530 ( \44163 , \43004 , \44162 );
and \U$43531 ( \44164 , \43001 , \44162 );
or \U$43532 ( \44165 , \43005 , \44163 , \44164 );
and \U$43533 ( \44166 , \42997 , \44165 );
and \U$43534 ( \44167 , \42994 , \44165 );
or \U$43535 ( \44168 , \42998 , \44166 , \44167 );
and \U$43536 ( \44169 , \42990 , \44168 );
and \U$43537 ( \44170 , \42987 , \44168 );
or \U$43538 ( \44171 , \42991 , \44169 , \44170 );
and \U$43539 ( \44172 , \42983 , \44171 );
and \U$43540 ( \44173 , \42980 , \44171 );
or \U$43541 ( \44174 , \42984 , \44172 , \44173 );
and \U$43542 ( \44175 , \42976 , \44174 );
and \U$43543 ( \44176 , \42973 , \44174 );
or \U$43544 ( \44177 , \42977 , \44175 , \44176 );
and \U$43545 ( \44178 , \42969 , \44177 );
and \U$43546 ( \44179 , \42966 , \44177 );
or \U$43547 ( \44180 , \42970 , \44178 , \44179 );
and \U$43548 ( \44181 , \42962 , \44180 );
and \U$43549 ( \44182 , \42959 , \44180 );
or \U$43550 ( \44183 , \42963 , \44181 , \44182 );
and \U$43551 ( \44184 , \42955 , \44183 );
and \U$43552 ( \44185 , \42952 , \44183 );
or \U$43553 ( \44186 , \42956 , \44184 , \44185 );
and \U$43554 ( \44187 , \42948 , \44186 );
and \U$43555 ( \44188 , \42945 , \44186 );
or \U$43556 ( \44189 , \42949 , \44187 , \44188 );
and \U$43557 ( \44190 , \42941 , \44189 );
and \U$43558 ( \44191 , \42938 , \44189 );
or \U$43559 ( \44192 , \42942 , \44190 , \44191 );
and \U$43560 ( \44193 , \42934 , \44192 );
and \U$43561 ( \44194 , \42931 , \44192 );
or \U$43562 ( \44195 , \42935 , \44193 , \44194 );
xor \U$43563 ( \44196 , \42928 , \44195 );
buf gaee9_GF_PartitionCandidate( \44197_nGaee9 , \44196 );
xor \U$43564 ( \44198 , RIc22b390_193, RIc22b408_194);
xor \U$43565 ( \44199 , RIc22b480_195, RIc22b4f8_196);
xor \U$43566 ( \44200 , \44198 , \44199 );
xor \U$43567 ( \44201 , RIc22b570_197, RIc22b5e8_198);
xor \U$43568 ( \44202 , RIc22b660_199, RIc22b6d8_200);
xor \U$43569 ( \44203 , \44201 , \44202 );
xor \U$43570 ( \44204 , \44200 , \44203 );
xor \U$43571 ( \44205 , RIc22b750_201, RIc22b7c8_202);
xor \U$43572 ( \44206 , RIc22b840_203, RIc22b8b8_204);
xor \U$43573 ( \44207 , \44205 , \44206 );
xor \U$43574 ( \44208 , RIc22b930_205, RIc22b9a8_206);
xor \U$43575 ( \44209 , RIc22ba20_207, RIc22ba98_208);
xor \U$43576 ( \44210 , \44208 , \44209 );
xor \U$43577 ( \44211 , \44207 , \44210 );
xor \U$43578 ( \44212 , \44204 , \44211 );
xor \U$43579 ( \44213 , RIc22bb10_209, RIc22bb88_210);
xor \U$43580 ( \44214 , RIc22bc00_211, RIc22bc78_212);
xor \U$43581 ( \44215 , \44213 , \44214 );
xor \U$43582 ( \44216 , RIc22bcf0_213, RIc22bd68_214);
xor \U$43583 ( \44217 , RIc22bde0_215, RIc22be58_216);
xor \U$43584 ( \44218 , \44216 , \44217 );
xor \U$43585 ( \44219 , \44215 , \44218 );
xor \U$43586 ( \44220 , RIc22bed0_217, RIc22bf48_218);
xor \U$43587 ( \44221 , RIc22bfc0_219, RIc22c038_220);
xor \U$43588 ( \44222 , \44220 , \44221 );
xor \U$43589 ( \44223 , RIc22c0b0_221, RIc22c128_222);
xor \U$43590 ( \44224 , RIc22c1a0_223, RIc22c218_224);
xor \U$43591 ( \44225 , \44223 , \44224 );
xor \U$43592 ( \44226 , \44222 , \44225 );
xor \U$43593 ( \44227 , \44219 , \44226 );
xor \U$43594 ( \44228 , \44212 , \44227 );
xor \U$43595 ( \44229 , RIc22c290_225, RIc22c308_226);
xor \U$43596 ( \44230 , RIc22c380_227, RIc22c3f8_228);
xor \U$43597 ( \44231 , \44229 , \44230 );
xor \U$43598 ( \44232 , RIc22c470_229, RIc22c4e8_230);
xor \U$43599 ( \44233 , RIc22c560_231, RIc22c5d8_232);
xor \U$43600 ( \44234 , \44232 , \44233 );
xor \U$43601 ( \44235 , \44231 , \44234 );
xor \U$43602 ( \44236 , RIc22c650_233, RIc22c6c8_234);
xor \U$43603 ( \44237 , RIc22c740_235, RIc22c7b8_236);
xor \U$43604 ( \44238 , \44236 , \44237 );
xor \U$43605 ( \44239 , RIc22c830_237, RIc22c8a8_238);
xor \U$43606 ( \44240 , RIc22c920_239, RIc22c998_240);
xor \U$43607 ( \44241 , \44239 , \44240 );
xor \U$43608 ( \44242 , \44238 , \44241 );
xor \U$43609 ( \44243 , \44235 , \44242 );
xor \U$43610 ( \44244 , RIc22ca10_241, RIc22ca88_242);
xor \U$43611 ( \44245 , RIc22cb00_243, RIc22cb78_244);
xor \U$43612 ( \44246 , \44244 , \44245 );
xor \U$43613 ( \44247 , RIc22cbf0_245, RIc22cc68_246);
xor \U$43614 ( \44248 , RIc22cce0_247, RIc22cd58_248);
xor \U$43615 ( \44249 , \44247 , \44248 );
xor \U$43616 ( \44250 , \44246 , \44249 );
xor \U$43617 ( \44251 , RIc22cdd0_249, RIc22ce48_250);
xor \U$43618 ( \44252 , RIc22cec0_251, RIc22cf38_252);
xor \U$43619 ( \44253 , \44251 , \44252 );
xor \U$43620 ( \44254 , RIc22cfb0_253, RIc22d028_254);
xor \U$43621 ( \44255 , RIc22d0a0_255, RIc22d118_256);
xor \U$43622 ( \44256 , \44254 , \44255 );
xor \U$43623 ( \44257 , \44253 , \44256 );
xor \U$43624 ( \44258 , \44250 , \44257 );
xor \U$43625 ( \44259 , \44243 , \44258 );
xor \U$43626 ( \44260 , \44228 , \44259 );
not \U$43627 ( \44261 , \44260 );
_DC gaeea ( \44262_nGaeea , \44197_nGaee9 , \44261 );
buf \U$43628 ( \44263 , \44262_nGaeea );
xor \U$43629 ( \44264 , \42931 , \42934 );
xor \U$43630 ( \44265 , \44264 , \44192 );
buf gaec7_GF_PartitionCandidate( \44266_nGaec7 , \44265 );
_DC gaec8 ( \44267_nGaec8 , \44266_nGaec7 , \44261 );
buf \U$43631 ( \44268 , \44267_nGaec8 );
xor \U$43632 ( \44269 , \42938 , \42941 );
xor \U$43633 ( \44270 , \44269 , \44189 );
buf gae95_GF_PartitionCandidate( \44271_nGae95 , \44270 );
_DC gae96 ( \44272_nGae96 , \44271_nGae95 , \44261 );
buf \U$43634 ( \44273 , \44272_nGae96 );
xor \U$43635 ( \44274 , \42945 , \42948 );
xor \U$43636 ( \44275 , \44274 , \44186 );
buf gae59_GF_PartitionCandidate( \44276_nGae59 , \44275 );
_DC gae5a ( \44277_nGae5a , \44276_nGae59 , \44261 );
buf \U$43637 ( \44278 , \44277_nGae5a );
xor \U$43638 ( \44279 , \42952 , \42955 );
xor \U$43639 ( \44280 , \44279 , \44183 );
buf gae0f_GF_PartitionCandidate( \44281_nGae0f , \44280 );
_DC gae10 ( \44282_nGae10 , \44281_nGae0f , \44261 );
buf \U$43640 ( \44283 , \44282_nGae10 );
xor \U$43641 ( \44284 , \42959 , \42962 );
xor \U$43642 ( \44285 , \44284 , \44180 );
buf gadbb_GF_PartitionCandidate( \44286_nGadbb , \44285 );
_DC gadbc ( \44287_nGadbc , \44286_nGadbb , \44261 );
buf \U$43643 ( \44288 , \44287_nGadbc );
xor \U$43644 ( \44289 , \42966 , \42969 );
xor \U$43645 ( \44290 , \44289 , \44177 );
buf gad61_GF_PartitionCandidate( \44291_nGad61 , \44290 );
_DC gad62 ( \44292_nGad62 , \44291_nGad61 , \44261 );
buf \U$43646 ( \44293 , \44292_nGad62 );
xor \U$43647 ( \44294 , \42973 , \42976 );
xor \U$43648 ( \44295 , \44294 , \44174 );
buf gacfd_GF_PartitionCandidate( \44296_nGacfd , \44295 );
_DC gacfe ( \44297_nGacfe , \44296_nGacfd , \44261 );
buf \U$43649 ( \44298 , \44297_nGacfe );
xor \U$43650 ( \44299 , \42980 , \42983 );
xor \U$43651 ( \44300 , \44299 , \44171 );
buf gac8b_GF_PartitionCandidate( \44301_nGac8b , \44300 );
_DC gac8c ( \44302_nGac8c , \44301_nGac8b , \44261 );
buf \U$43652 ( \44303 , \44302_nGac8c );
xor \U$43653 ( \44304 , \42987 , \42990 );
xor \U$43654 ( \44305 , \44304 , \44168 );
buf gac15_GF_PartitionCandidate( \44306_nGac15 , \44305 );
_DC gac16 ( \44307_nGac16 , \44306_nGac15 , \44261 );
buf \U$43655 ( \44308 , \44307_nGac16 );
xor \U$43656 ( \44309 , \42994 , \42997 );
xor \U$43657 ( \44310 , \44309 , \44165 );
buf gab8f_GF_PartitionCandidate( \44311_nGab8f , \44310 );
_DC gab90 ( \44312_nGab90 , \44311_nGab8f , \44261 );
buf \U$43658 ( \44313 , \44312_nGab90 );
xor \U$43659 ( \44314 , \43001 , \43004 );
xor \U$43660 ( \44315 , \44314 , \44162 );
buf gaaff_GF_PartitionCandidate( \44316_nGaaff , \44315 );
_DC gab00 ( \44317_nGab00 , \44316_nGaaff , \44261 );
buf \U$43661 ( \44318 , \44317_nGab00 );
xor \U$43662 ( \44319 , \43008 , \43011 );
xor \U$43663 ( \44320 , \44319 , \44159 );
buf gaa69_GF_PartitionCandidate( \44321_nGaa69 , \44320 );
_DC gaa6a ( \44322_nGaa6a , \44321_nGaa69 , \44261 );
buf \U$43664 ( \44323 , \44322_nGaa6a );
xor \U$43665 ( \44324 , \43015 , \43018 );
xor \U$43666 ( \44325 , \44324 , \44156 );
buf ga9c9_GF_PartitionCandidate( \44326_nGa9c9 , \44325 );
_DC ga9ca ( \44327_nGa9ca , \44326_nGa9c9 , \44261 );
buf \U$43667 ( \44328 , \44327_nGa9ca );
xor \U$43668 ( \44329 , \43022 , \43025 );
xor \U$43669 ( \44330 , \44329 , \44153 );
buf ga91b_GF_PartitionCandidate( \44331_nGa91b , \44330 );
_DC ga91c ( \44332_nGa91c , \44331_nGa91b , \44261 );
buf \U$43670 ( \44333 , \44332_nGa91c );
xor \U$43671 ( \44334 , \43029 , \43032 );
xor \U$43672 ( \44335 , \44334 , \44150 );
buf ga869_GF_PartitionCandidate( \44336_nGa869 , \44335 );
_DC ga86a ( \44337_nGa86a , \44336_nGa869 , \44261 );
buf \U$43673 ( \44338 , \44337_nGa86a );
xor \U$43674 ( \44339 , \43036 , \43039 );
xor \U$43675 ( \44340 , \44339 , \44147 );
buf ga7a7_GF_PartitionCandidate( \44341_nGa7a7 , \44340 );
_DC ga7a8 ( \44342_nGa7a8 , \44341_nGa7a7 , \44261 );
buf \U$43676 ( \44343 , \44342_nGa7a8 );
xor \U$43677 ( \44344 , \43043 , \43046 );
xor \U$43678 ( \44345 , \44344 , \44144 );
buf ga6e1_GF_PartitionCandidate( \44346_nGa6e1 , \44345 );
_DC ga6e2 ( \44347_nGa6e2 , \44346_nGa6e1 , \44261 );
buf \U$43679 ( \44348 , \44347_nGa6e2 );
xor \U$43680 ( \44349 , \43050 , \43053 );
xor \U$43681 ( \44350 , \44349 , \44141 );
buf ga60b_GF_PartitionCandidate( \44351_nGa60b , \44350 );
_DC ga60c ( \44352_nGa60c , \44351_nGa60b , \44261 );
buf \U$43682 ( \44353 , \44352_nGa60c );
xor \U$43683 ( \44354 , \43057 , \43060 );
xor \U$43684 ( \44355 , \44354 , \44138 );
buf ga531_GF_PartitionCandidate( \44356_nGa531 , \44355 );
_DC ga532 ( \44357_nGa532 , \44356_nGa531 , \44261 );
buf \U$43685 ( \44358 , \44357_nGa532 );
xor \U$43686 ( \44359 , \43064 , \43067 );
xor \U$43687 ( \44360 , \44359 , \44135 );
buf ga44d_GF_PartitionCandidate( \44361_nGa44d , \44360 );
_DC ga44e ( \44362_nGa44e , \44361_nGa44d , \44261 );
buf \U$43688 ( \44363 , \44362_nGa44e );
xor \U$43689 ( \44364 , \43071 , \43074 );
xor \U$43690 ( \44365 , \44364 , \44132 );
buf ga35d_GF_PartitionCandidate( \44366_nGa35d , \44365 );
_DC ga35e ( \44367_nGa35e , \44366_nGa35d , \44261 );
buf \U$43691 ( \44368 , \44367_nGa35e );
xor \U$43692 ( \44369 , \43078 , \43081 );
xor \U$43693 ( \44370 , \44369 , \44129 );
buf ga25f_GF_PartitionCandidate( \44371_nGa25f , \44370 );
_DC ga260 ( \44372_nGa260 , \44371_nGa25f , \44261 );
buf \U$43694 ( \44373 , \44372_nGa260 );
xor \U$43695 ( \44374 , \43085 , \43088 );
xor \U$43696 ( \44375 , \44374 , \44126 );
buf ga157_GF_PartitionCandidate( \44376_nGa157 , \44375 );
_DC ga158 ( \44377_nGa158 , \44376_nGa157 , \44261 );
buf \U$43697 ( \44378 , \44377_nGa158 );
xor \U$43698 ( \44379 , \43092 , \43095 );
xor \U$43699 ( \44380 , \44379 , \44123 );
buf ga043_GF_PartitionCandidate( \44381_nGa043 , \44380 );
_DC ga044 ( \44382_nGa044 , \44381_nGa043 , \44261 );
buf \U$43700 ( \44383 , \44382_nGa044 );
xor \U$43701 ( \44384 , \43099 , \43102 );
xor \U$43702 ( \44385 , \44384 , \44120 );
buf g9f2d_GF_PartitionCandidate( \44386_nG9f2d , \44385 );
_DC g9f2e ( \44387_nG9f2e , \44386_nG9f2d , \44261 );
buf \U$43703 ( \44388 , \44387_nG9f2e );
xor \U$43704 ( \44389 , \43106 , \43109 );
xor \U$43705 ( \44390 , \44389 , \44117 );
buf g9e07_GF_PartitionCandidate( \44391_nG9e07 , \44390 );
_DC g9e08 ( \44392_nG9e08 , \44391_nG9e07 , \44261 );
buf \U$43706 ( \44393 , \44392_nG9e08 );
xor \U$43707 ( \44394 , \43113 , \43116 );
xor \U$43708 ( \44395 , \44394 , \44114 );
buf g9cd7_GF_PartitionCandidate( \44396_nG9cd7 , \44395 );
_DC g9cd8 ( \44397_nG9cd8 , \44396_nG9cd7 , \44261 );
buf \U$43709 ( \44398 , \44397_nG9cd8 );
xor \U$43710 ( \44399 , \43120 , \43123 );
xor \U$43711 ( \44400 , \44399 , \44111 );
buf g9b99_GF_PartitionCandidate( \44401_nG9b99 , \44400 );
_DC g9b9a ( \44402_nG9b9a , \44401_nG9b99 , \44261 );
buf \U$43712 ( \44403 , \44402_nG9b9a );
xor \U$43713 ( \44404 , \43127 , \43130 );
xor \U$43714 ( \44405 , \44404 , \44108 );
buf g9a51_GF_PartitionCandidate( \44406_nG9a51 , \44405 );
_DC g9a52 ( \44407_nG9a52 , \44406_nG9a51 , \44261 );
buf \U$43715 ( \44408 , \44407_nG9a52 );
xor \U$43716 ( \44409 , \43134 , \43137 );
xor \U$43717 ( \44410 , \44409 , \44105 );
buf g9903_GF_PartitionCandidate( \44411_nG9903 , \44410 );
_DC g9904 ( \44412_nG9904 , \44411_nG9903 , \44261 );
buf \U$43718 ( \44413 , \44412_nG9904 );
xor \U$43719 ( \44414 , \43141 , \43144 );
xor \U$43720 ( \44415 , \44414 , \44102 );
buf g97b1_GF_PartitionCandidate( \44416_nG97b1 , \44415 );
_DC g97b2 ( \44417_nG97b2 , \44416_nG97b1 , \44261 );
buf \U$43721 ( \44418 , \44417_nG97b2 );
xor \U$43722 ( \44419 , \43148 , \43151 );
xor \U$43723 ( \44420 , \44419 , \44099 );
buf g9655_GF_PartitionCandidate( \44421_nG9655 , \44420 );
_DC g9656 ( \44422_nG9656 , \44421_nG9655 , \44261 );
buf \U$43724 ( \44423 , \44422_nG9656 );
xor \U$43725 ( \44424 , \43155 , \43158 );
xor \U$43726 ( \44425 , \44424 , \44096 );
buf g94f3_GF_PartitionCandidate( \44426_nG94f3 , \44425 );
_DC g94f4 ( \44427_nG94f4 , \44426_nG94f3 , \44261 );
buf \U$43727 ( \44428 , \44427_nG94f4 );
xor \U$43728 ( \44429 , \43162 , \43165 );
xor \U$43729 ( \44430 , \44429 , \44093 );
buf g9381_GF_PartitionCandidate( \44431_nG9381 , \44430 );
_DC g9382 ( \44432_nG9382 , \44431_nG9381 , \44261 );
buf \U$43730 ( \44433 , \44432_nG9382 );
xor \U$43731 ( \44434 , \43169 , \43172 );
xor \U$43732 ( \44435 , \44434 , \44090 );
buf g9205_GF_PartitionCandidate( \44436_nG9205 , \44435 );
_DC g9206 ( \44437_nG9206 , \44436_nG9205 , \44261 );
buf \U$43733 ( \44438 , \44437_nG9206 );
xor \U$43734 ( \44439 , \43176 , \43179 );
xor \U$43735 ( \44440 , \44439 , \44087 );
buf g907b_GF_PartitionCandidate( \44441_nG907b , \44440 );
_DC g907c ( \44442_nG907c , \44441_nG907b , \44261 );
buf \U$43736 ( \44443 , \44442_nG907c );
xor \U$43737 ( \44444 , \43183 , \43186 );
xor \U$43738 ( \44445 , \44444 , \44084 );
buf g8eed_GF_PartitionCandidate( \44446_nG8eed , \44445 );
_DC g8eee ( \44447_nG8eee , \44446_nG8eed , \44261 );
buf \U$43739 ( \44448 , \44447_nG8eee );
xor \U$43740 ( \44449 , \43190 , \43193 );
xor \U$43741 ( \44450 , \44449 , \44081 );
buf g8d4f_GF_PartitionCandidate( \44451_nG8d4f , \44450 );
_DC g8d50 ( \44452_nG8d50 , \44451_nG8d4f , \44261 );
buf \U$43742 ( \44453 , \44452_nG8d50 );
xor \U$43743 ( \44454 , \43197 , \43200 );
xor \U$43744 ( \44455 , \44454 , \44078 );
buf g8bad_GF_PartitionCandidate( \44456_nG8bad , \44455 );
_DC g8bae ( \44457_nG8bae , \44456_nG8bad , \44261 );
buf \U$43745 ( \44458 , \44457_nG8bae );
xor \U$43746 ( \44459 , \43204 , \43207 );
xor \U$43747 ( \44460 , \44459 , \44075 );
buf g89fb_GF_PartitionCandidate( \44461_nG89fb , \44460 );
_DC g89fc ( \44462_nG89fc , \44461_nG89fb , \44261 );
buf \U$43748 ( \44463 , \44462_nG89fc );
xor \U$43749 ( \44464 , \43211 , \43214 );
xor \U$43750 ( \44465 , \44464 , \44072 );
buf g883f_GF_PartitionCandidate( \44466_nG883f , \44465 );
_DC g8840 ( \44467_nG8840 , \44466_nG883f , \44261 );
buf \U$43751 ( \44468 , \44467_nG8840 );
xor \U$43752 ( \44469 , \43218 , \43221 );
xor \U$43753 ( \44470 , \44469 , \44069 );
buf g8677_GF_PartitionCandidate( \44471_nG8677 , \44470 );
_DC g8678 ( \44472_nG8678 , \44471_nG8677 , \44261 );
buf \U$43754 ( \44473 , \44472_nG8678 );
xor \U$43755 ( \44474 , \43225 , \43228 );
xor \U$43756 ( \44475 , \44474 , \44066 );
buf g84a7_GF_PartitionCandidate( \44476_nG84a7 , \44475 );
_DC g84a8 ( \44477_nG84a8 , \44476_nG84a7 , \44261 );
buf \U$43757 ( \44478 , \44477_nG84a8 );
xor \U$43758 ( \44479 , \43232 , \43235 );
xor \U$43759 ( \44480 , \44479 , \44063 );
buf g82c9_GF_PartitionCandidate( \44481_nG82c9 , \44480 );
_DC g82ca ( \44482_nG82ca , \44481_nG82c9 , \44261 );
buf \U$43760 ( \44483 , \44482_nG82ca );
xor \U$43761 ( \44484 , \43239 , \43242 );
xor \U$43762 ( \44485 , \44484 , \44060 );
buf g80e7_GF_PartitionCandidate( \44486_nG80e7 , \44485 );
_DC g80e8 ( \44487_nG80e8 , \44486_nG80e7 , \44261 );
buf \U$43763 ( \44488 , \44487_nG80e8 );
xor \U$43764 ( \44489 , \43246 , \43249 );
xor \U$43765 ( \44490 , \44489 , \44057 );
buf g7ef5_GF_PartitionCandidate( \44491_nG7ef5 , \44490 );
_DC g7ef6 ( \44492_nG7ef6 , \44491_nG7ef5 , \44261 );
buf \U$43766 ( \44493 , \44492_nG7ef6 );
xor \U$43767 ( \44494 , \43253 , \43256 );
xor \U$43768 ( \44495 , \44494 , \44054 );
buf g7cf9_GF_PartitionCandidate( \44496_nG7cf9 , \44495 );
_DC g7cfa ( \44497_nG7cfa , \44496_nG7cf9 , \44261 );
buf \U$43769 ( \44498 , \44497_nG7cfa );
xor \U$43770 ( \44499 , \43260 , \43263 );
xor \U$43771 ( \44500 , \44499 , \44051 );
buf g7af7_GF_PartitionCandidate( \44501_nG7af7 , \44500 );
_DC g7af8 ( \44502_nG7af8 , \44501_nG7af7 , \44261 );
buf \U$43772 ( \44503 , \44502_nG7af8 );
xor \U$43773 ( \44504 , \43267 , \43270 );
xor \U$43774 ( \44505 , \44504 , \44048 );
buf g78f1_GF_PartitionCandidate( \44506_nG78f1 , \44505 );
_DC g78f2 ( \44507_nG78f2 , \44506_nG78f1 , \44261 );
buf \U$43775 ( \44508 , \44507_nG78f2 );
xor \U$43776 ( \44509 , \43274 , \43277 );
xor \U$43777 ( \44510 , \44509 , \44045 );
buf g76e1_GF_PartitionCandidate( \44511_nG76e1 , \44510 );
_DC g76e2 ( \44512_nG76e2 , \44511_nG76e1 , \44261 );
buf \U$43778 ( \44513 , \44512_nG76e2 );
xor \U$43779 ( \44514 , \43281 , \43284 );
xor \U$43780 ( \44515 , \44514 , \44042 );
buf g74c5_GF_PartitionCandidate( \44516_nG74c5 , \44515 );
_DC g74c6 ( \44517_nG74c6 , \44516_nG74c5 , \44261 );
buf \U$43781 ( \44518 , \44517_nG74c6 );
xor \U$43782 ( \44519 , \43288 , \43291 );
xor \U$43783 ( \44520 , \44519 , \44039 );
buf g72a1_GF_PartitionCandidate( \44521_nG72a1 , \44520 );
_DC g72a2 ( \44522_nG72a2 , \44521_nG72a1 , \44261 );
buf \U$43784 ( \44523 , \44522_nG72a2 );
xor \U$43785 ( \44524 , \43295 , \43298 );
xor \U$43786 ( \44525 , \44524 , \44036 );
buf g7077_GF_PartitionCandidate( \44526_nG7077 , \44525 );
_DC g7078 ( \44527_nG7078 , \44526_nG7077 , \44261 );
buf \U$43787 ( \44528 , \44527_nG7078 );
xor \U$43788 ( \44529 , \43302 , \43305 );
xor \U$43789 ( \44530 , \44529 , \44033 );
buf g6e3d_GF_PartitionCandidate( \44531_nG6e3d , \44530 );
_DC g6e3e ( \44532_nG6e3e , \44531_nG6e3d , \44261 );
buf \U$43790 ( \44533 , \44532_nG6e3e );
xor \U$43791 ( \44534 , \43309 , \43312 );
xor \U$43792 ( \44535 , \44534 , \44030 );
buf g6bff_GF_PartitionCandidate( \44536_nG6bff , \44535 );
_DC g6c00 ( \44537_nG6c00 , \44536_nG6bff , \44261 );
buf \U$43793 ( \44538 , \44537_nG6c00 );
xor \U$43794 ( \44539 , \43316 , \43319 );
xor \U$43795 ( \44540 , \44539 , \44027 );
buf g69b1_GF_PartitionCandidate( \44541_nG69b1 , \44540 );
_DC g69b2 ( \44542_nG69b2 , \44541_nG69b1 , \44261 );
buf \U$43796 ( \44543 , \44542_nG69b2 );
xor \U$43797 ( \44544 , \43323 , \43326 );
xor \U$43798 ( \44545 , \44544 , \44024 );
buf g6759_GF_PartitionCandidate( \44546_nG6759 , \44545 );
_DC g675a ( \44547_nG675a , \44546_nG6759 , \44261 );
buf \U$43799 ( \44548 , \44547_nG675a );
xor \U$43800 ( \44549 , \43330 , \43333 );
xor \U$43801 ( \44550 , \44549 , \44021 );
buf g64f3_GF_PartitionCandidate( \44551_nG64f3 , \44550 );
_DC g64f4 ( \44552_nG64f4 , \44551_nG64f3 , \44261 );
buf \U$43802 ( \44553 , \44552_nG64f4 );
xor \U$43803 ( \44554 , \43337 , \43340 );
xor \U$43804 ( \44555 , \44554 , \44018 );
buf g6283_GF_PartitionCandidate( \44556_nG6283 , \44555 );
_DC g6284 ( \44557_nG6284 , \44556_nG6283 , \44261 );
buf \U$43805 ( \44558 , \44557_nG6284 );
xor \U$43806 ( \44559 , \43344 , \43347 );
xor \U$43807 ( \44560 , \44559 , \44015 );
buf g600d_GF_PartitionCandidate( \44561_nG600d , \44560 );
_DC g600e ( \44562_nG600e , \44561_nG600d , \44261 );
buf \U$43808 ( \44563 , \44562_nG600e );
xor \U$43809 ( \44564 , \43351 , \43354 );
xor \U$43810 ( \44565 , \44564 , \44012 );
buf g5d8d_GF_PartitionCandidate( \44566_nG5d8d , \44565 );
_DC g5d8e ( \44567_nG5d8e , \44566_nG5d8d , \44261 );
buf \U$43811 ( \44568 , \44567_nG5d8e );
xor \U$43812 ( \44569 , \43358 , \43361 );
xor \U$43813 ( \44570 , \44569 , \44009 );
buf g5b0b_GF_PartitionCandidate( \44571_nG5b0b , \44570 );
_DC g5b0c ( \44572_nG5b0c , \44571_nG5b0b , \44261 );
buf \U$43814 ( \44573 , \44572_nG5b0c );
xor \U$43815 ( \44574 , \43365 , \43368 );
xor \U$43816 ( \44575 , \44574 , \44006 );
buf g5887_GF_PartitionCandidate( \44576_nG5887 , \44575 );
_DC g5888 ( \44577_nG5888 , \44576_nG5887 , \44261 );
buf \U$43817 ( \44578 , \44577_nG5888 );
xor \U$43818 ( \44579 , \43372 , \43375 );
xor \U$43819 ( \44580 , \44579 , \44003 );
buf g5601_GF_PartitionCandidate( \44581_nG5601 , \44580 );
_DC g5602 ( \44582_nG5602 , \44581_nG5601 , \44261 );
buf \U$43820 ( \44583 , \44582_nG5602 );
xor \U$43821 ( \44584 , \43379 , \43382 );
xor \U$43822 ( \44585 , \44584 , \44000 );
buf g5377_GF_PartitionCandidate( \44586_nG5377 , \44585 );
_DC g5378 ( \44587_nG5378 , \44586_nG5377 , \44261 );
buf \U$43823 ( \44588 , \44587_nG5378 );
xor \U$43824 ( \44589 , \43386 , \43389 );
xor \U$43825 ( \44590 , \44589 , \43997 );
buf g50f3_GF_PartitionCandidate( \44591_nG50f3 , \44590 );
_DC g50f4 ( \44592_nG50f4 , \44591_nG50f3 , \44261 );
buf \U$43826 ( \44593 , \44592_nG50f4 );
xor \U$43827 ( \44594 , \43393 , \43396 );
xor \U$43828 ( \44595 , \44594 , \43994 );
buf g4e7d_GF_PartitionCandidate( \44596_nG4e7d , \44595 );
_DC g4e7e ( \44597_nG4e7e , \44596_nG4e7d , \44261 );
buf \U$43829 ( \44598 , \44597_nG4e7e );
xor \U$43830 ( \44599 , \43400 , \43403 );
xor \U$43831 ( \44600 , \44599 , \43991 );
buf g4c0d_GF_PartitionCandidate( \44601_nG4c0d , \44600 );
_DC g4c0e ( \44602_nG4c0e , \44601_nG4c0d , \44261 );
buf \U$43832 ( \44603 , \44602_nG4c0e );
xor \U$43833 ( \44604 , \43407 , \43410 );
xor \U$43834 ( \44605 , \44604 , \43988 );
buf g49ab_GF_PartitionCandidate( \44606_nG49ab , \44605 );
_DC g49ac ( \44607_nG49ac , \44606_nG49ab , \44261 );
buf \U$43835 ( \44608 , \44607_nG49ac );
xor \U$43836 ( \44609 , \43414 , \43417 );
xor \U$43837 ( \44610 , \44609 , \43985 );
buf g474f_GF_PartitionCandidate( \44611_nG474f , \44610 );
_DC g4750 ( \44612_nG4750 , \44611_nG474f , \44261 );
buf \U$43838 ( \44613 , \44612_nG4750 );
xor \U$43839 ( \44614 , \43421 , \43424 );
xor \U$43840 ( \44615 , \44614 , \43982 );
buf g4501_GF_PartitionCandidate( \44616_nG4501 , \44615 );
_DC g4502 ( \44617_nG4502 , \44616_nG4501 , \44261 );
buf \U$43841 ( \44618 , \44617_nG4502 );
xor \U$43842 ( \44619 , \43428 , \43431 );
xor \U$43843 ( \44620 , \44619 , \43979 );
buf g42b9_GF_PartitionCandidate( \44621_nG42b9 , \44620 );
_DC g42ba ( \44622_nG42ba , \44621_nG42b9 , \44261 );
buf \U$43844 ( \44623 , \44622_nG42ba );
xor \U$43845 ( \44624 , \43435 , \43438 );
xor \U$43846 ( \44625 , \44624 , \43976 );
buf g407f_GF_PartitionCandidate( \44626_nG407f , \44625 );
_DC g4080 ( \44627_nG4080 , \44626_nG407f , \44261 );
buf \U$43847 ( \44628 , \44627_nG4080 );
xor \U$43848 ( \44629 , \43442 , \43445 );
xor \U$43849 ( \44630 , \44629 , \43973 );
buf g3e4b_GF_PartitionCandidate( \44631_nG3e4b , \44630 );
_DC g3e4c ( \44632_nG3e4c , \44631_nG3e4b , \44261 );
buf \U$43850 ( \44633 , \44632_nG3e4c );
xor \U$43851 ( \44634 , \43449 , \43452 );
xor \U$43852 ( \44635 , \44634 , \43970 );
buf g3c25_GF_PartitionCandidate( \44636_nG3c25 , \44635 );
_DC g3c26 ( \44637_nG3c26 , \44636_nG3c25 , \44261 );
buf \U$43853 ( \44638 , \44637_nG3c26 );
xor \U$43854 ( \44639 , \43456 , \43459 );
xor \U$43855 ( \44640 , \44639 , \43967 );
buf g3a05_GF_PartitionCandidate( \44641_nG3a05 , \44640 );
_DC g3a06 ( \44642_nG3a06 , \44641_nG3a05 , \44261 );
buf \U$43856 ( \44643 , \44642_nG3a06 );
xor \U$43857 ( \44644 , \43463 , \43466 );
xor \U$43858 ( \44645 , \44644 , \43964 );
buf g37f3_GF_PartitionCandidate( \44646_nG37f3 , \44645 );
_DC g37f4 ( \44647_nG37f4 , \44646_nG37f3 , \44261 );
buf \U$43859 ( \44648 , \44647_nG37f4 );
xor \U$43860 ( \44649 , \43470 , \43473 );
xor \U$43861 ( \44650 , \44649 , \43961 );
buf g35e7_GF_PartitionCandidate( \44651_nG35e7 , \44650 );
_DC g35e8 ( \44652_nG35e8 , \44651_nG35e7 , \44261 );
buf \U$43862 ( \44653 , \44652_nG35e8 );
xor \U$43863 ( \44654 , \43477 , \43480 );
xor \U$43864 ( \44655 , \44654 , \43958 );
buf g33e9_GF_PartitionCandidate( \44656_nG33e9 , \44655 );
_DC g33ea ( \44657_nG33ea , \44656_nG33e9 , \44261 );
buf \U$43865 ( \44658 , \44657_nG33ea );
xor \U$43866 ( \44659 , \43484 , \43487 );
xor \U$43867 ( \44660 , \44659 , \43955 );
buf g31f1_GF_PartitionCandidate( \44661_nG31f1 , \44660 );
_DC g31f2 ( \44662_nG31f2 , \44661_nG31f1 , \44261 );
buf \U$43868 ( \44663 , \44662_nG31f2 );
xor \U$43869 ( \44664 , \43491 , \43494 );
xor \U$43870 ( \44665 , \44664 , \43952 );
buf g3007_GF_PartitionCandidate( \44666_nG3007 , \44665 );
_DC g3008 ( \44667_nG3008 , \44666_nG3007 , \44261 );
buf \U$43871 ( \44668 , \44667_nG3008 );
xor \U$43872 ( \44669 , \43498 , \43501 );
xor \U$43873 ( \44670 , \44669 , \43949 );
buf g2e23_GF_PartitionCandidate( \44671_nG2e23 , \44670 );
_DC g2e24 ( \44672_nG2e24 , \44671_nG2e23 , \44261 );
buf \U$43874 ( \44673 , \44672_nG2e24 );
xor \U$43875 ( \44674 , \43505 , \43508 );
xor \U$43876 ( \44675 , \44674 , \43946 );
buf g2c4d_GF_PartitionCandidate( \44676_nG2c4d , \44675 );
_DC g2c4e ( \44677_nG2c4e , \44676_nG2c4d , \44261 );
buf \U$43877 ( \44678 , \44677_nG2c4e );
xor \U$43878 ( \44679 , \43512 , \43515 );
xor \U$43879 ( \44680 , \44679 , \43943 );
buf g2a77_GF_PartitionCandidate( \44681_nG2a77 , \44680 );
_DC g2a78 ( \44682_nG2a78 , \44681_nG2a77 , \44261 );
buf \U$43880 ( \44683 , \44682_nG2a78 );
xor \U$43881 ( \44684 , \43519 , \43522 );
xor \U$43882 ( \44685 , \44684 , \43940 );
buf g28b7_GF_PartitionCandidate( \44686_nG28b7 , \44685 );
_DC g28b8 ( \44687_nG28b8 , \44686_nG28b7 , \44261 );
buf \U$43883 ( \44688 , \44687_nG28b8 );
xor \U$43884 ( \44689 , \43526 , \43529 );
xor \U$43885 ( \44690 , \44689 , \43937 );
buf g26fb_GF_PartitionCandidate( \44691_nG26fb , \44690 );
_DC g26fc ( \44692_nG26fc , \44691_nG26fb , \44261 );
buf \U$43886 ( \44693 , \44692_nG26fc );
xor \U$43887 ( \44694 , \43533 , \43536 );
xor \U$43888 ( \44695 , \44694 , \43934 );
buf g254d_GF_PartitionCandidate( \44696_nG254d , \44695 );
_DC g254e ( \44697_nG254e , \44696_nG254d , \44261 );
buf \U$43889 ( \44698 , \44697_nG254e );
xor \U$43890 ( \44699 , \43540 , \43543 );
xor \U$43891 ( \44700 , \44699 , \43931 );
buf g23a5_GF_PartitionCandidate( \44701_nG23a5 , \44700 );
_DC g23a6 ( \44702_nG23a6 , \44701_nG23a5 , \44261 );
buf \U$43892 ( \44703 , \44702_nG23a6 );
xor \U$43893 ( \44704 , \43547 , \43550 );
xor \U$43894 ( \44705 , \44704 , \43928 );
buf g220b_GF_PartitionCandidate( \44706_nG220b , \44705 );
_DC g220c ( \44707_nG220c , \44706_nG220b , \44261 );
buf \U$43895 ( \44708 , \44707_nG220c );
xor \U$43896 ( \44709 , \43554 , \43557 );
xor \U$43897 ( \44710 , \44709 , \43925 );
buf g2077_GF_PartitionCandidate( \44711_nG2077 , \44710 );
_DC g2078 ( \44712_nG2078 , \44711_nG2077 , \44261 );
buf \U$43898 ( \44713 , \44712_nG2078 );
xor \U$43899 ( \44714 , \43561 , \43564 );
xor \U$43900 ( \44715 , \44714 , \43922 );
buf g1ef1_GF_PartitionCandidate( \44716_nG1ef1 , \44715 );
_DC g1ef2 ( \44717_nG1ef2 , \44716_nG1ef1 , \44261 );
buf \U$43901 ( \44718 , \44717_nG1ef2 );
xor \U$43902 ( \44719 , \43568 , \43571 );
xor \U$43903 ( \44720 , \44719 , \43919 );
buf g1d71_GF_PartitionCandidate( \44721_nG1d71 , \44720 );
_DC g1d72 ( \44722_nG1d72 , \44721_nG1d71 , \44261 );
buf \U$43904 ( \44723 , \44722_nG1d72 );
xor \U$43905 ( \44724 , \43575 , \43578 );
xor \U$43906 ( \44725 , \44724 , \43916 );
buf g1bff_GF_PartitionCandidate( \44726_nG1bff , \44725 );
_DC g1c00 ( \44727_nG1c00 , \44726_nG1bff , \44261 );
buf \U$43907 ( \44728 , \44727_nG1c00 );
xor \U$43908 ( \44729 , \43582 , \43585 );
xor \U$43909 ( \44730 , \44729 , \43913 );
buf g1a93_GF_PartitionCandidate( \44731_nG1a93 , \44730 );
_DC g1a94 ( \44732_nG1a94 , \44731_nG1a93 , \44261 );
buf \U$43910 ( \44733 , \44732_nG1a94 );
xor \U$43911 ( \44734 , \43589 , \43592 );
xor \U$43912 ( \44735 , \44734 , \43910 );
buf g1935_GF_PartitionCandidate( \44736_nG1935 , \44735 );
_DC g1936 ( \44737_nG1936 , \44736_nG1935 , \44261 );
buf \U$43913 ( \44738 , \44737_nG1936 );
xor \U$43914 ( \44739 , \43596 , \43599 );
xor \U$43915 ( \44740 , \44739 , \43907 );
buf g17dd_GF_PartitionCandidate( \44741_nG17dd , \44740 );
_DC g17de ( \44742_nG17de , \44741_nG17dd , \44261 );
buf \U$43916 ( \44743 , \44742_nG17de );
xor \U$43917 ( \44744 , \43603 , \43606 );
xor \U$43918 ( \44745 , \44744 , \43904 );
buf g1693_GF_PartitionCandidate( \44746_nG1693 , \44745 );
_DC g1694 ( \44747_nG1694 , \44746_nG1693 , \44261 );
buf \U$43919 ( \44748 , \44747_nG1694 );
xor \U$43920 ( \44749 , \43610 , \43613 );
xor \U$43921 ( \44750 , \44749 , \43901 );
buf g154f_GF_PartitionCandidate( \44751_nG154f , \44750 );
_DC g1550 ( \44752_nG1550 , \44751_nG154f , \44261 );
buf \U$43922 ( \44753 , \44752_nG1550 );
xor \U$43923 ( \44754 , \43617 , \43620 );
xor \U$43924 ( \44755 , \44754 , \43898 );
buf g1419_GF_PartitionCandidate( \44756_nG1419 , \44755 );
_DC g141a ( \44757_nG141a , \44756_nG1419 , \44261 );
buf \U$43925 ( \44758 , \44757_nG141a );
xor \U$43926 ( \44759 , \43624 , \43627 );
xor \U$43927 ( \44760 , \44759 , \43895 );
buf g12e9_GF_PartitionCandidate( \44761_nG12e9 , \44760 );
_DC g12ea ( \44762_nG12ea , \44761_nG12e9 , \44261 );
buf \U$43928 ( \44763 , \44762_nG12ea );
xor \U$43929 ( \44764 , \43631 , \43634 );
xor \U$43930 ( \44765 , \44764 , \43892 );
buf g11c7_GF_PartitionCandidate( \44766_nG11c7 , \44765 );
_DC g11c8 ( \44767_nG11c8 , \44766_nG11c7 , \44261 );
buf \U$43931 ( \44768 , \44767_nG11c8 );
xor \U$43932 ( \44769 , \43638 , \43641 );
xor \U$43933 ( \44770 , \44769 , \43889 );
buf g10ab_GF_PartitionCandidate( \44771_nG10ab , \44770 );
_DC g10ac ( \44772_nG10ac , \44771_nG10ab , \44261 );
buf \U$43934 ( \44773 , \44772_nG10ac );
xor \U$43935 ( \44774 , \43645 , \43648 );
xor \U$43936 ( \44775 , \44774 , \43886 );
buf gf9d_GF_PartitionCandidate( \44776_nGf9d , \44775 );
_DC gf9e ( \44777_nGf9e , \44776_nGf9d , \44261 );
buf \U$43937 ( \44778 , \44777_nGf9e );
xor \U$43938 ( \44779 , \43652 , \43655 );
xor \U$43939 ( \44780 , \44779 , \43883 );
buf ge95_GF_PartitionCandidate( \44781_nGe95 , \44780 );
_DC ge96 ( \44782_nGe96 , \44781_nGe95 , \44261 );
buf \U$43940 ( \44783 , \44782_nGe96 );
xor \U$43941 ( \44784 , \43659 , \43662 );
xor \U$43942 ( \44785 , \44784 , \43880 );
buf gd9b_GF_PartitionCandidate( \44786_nGd9b , \44785 );
_DC gd9c ( \44787_nGd9c , \44786_nGd9b , \44261 );
buf \U$43943 ( \44788 , \44787_nGd9c );
xor \U$43944 ( \44789 , \43666 , \43669 );
xor \U$43945 ( \44790 , \44789 , \43877 );
buf gca7_GF_PartitionCandidate( \44791_nGca7 , \44790 );
_DC gca8 ( \44792_nGca8 , \44791_nGca7 , \44261 );
buf \U$43946 ( \44793 , \44792_nGca8 );
xor \U$43947 ( \44794 , \43673 , \43676 );
xor \U$43948 ( \44795 , \44794 , \43874 );
buf gbc1_GF_PartitionCandidate( \44796_nGbc1 , \44795 );
_DC gbc2 ( \44797_nGbc2 , \44796_nGbc1 , \44261 );
buf \U$43949 ( \44798 , \44797_nGbc2 );
xor \U$43950 ( \44799 , \43680 , \43683 );
xor \U$43951 ( \44800 , \44799 , \43871 );
buf gae1_GF_PartitionCandidate( \44801_nGae1 , \44800 );
_DC gae2 ( \44802_nGae2 , \44801_nGae1 , \44261 );
buf \U$43952 ( \44803 , \44802_nGae2 );
xor \U$43953 ( \44804 , \43687 , \43690 );
xor \U$43954 ( \44805 , \44804 , \43868 );
buf ga0f_GF_PartitionCandidate( \44806_nGa0f , \44805 );
_DC ga10 ( \44807_nGa10 , \44806_nGa0f , \44261 );
buf \U$43955 ( \44808 , \44807_nGa10 );
xor \U$43956 ( \44809 , \43694 , \43697 );
xor \U$43957 ( \44810 , \44809 , \43865 );
buf g943_GF_PartitionCandidate( \44811_nG943 , \44810 );
_DC g944 ( \44812_nG944 , \44811_nG943 , \44261 );
buf \U$43958 ( \44813 , \44812_nG944 );
xor \U$43959 ( \44814 , \43701 , \43704 );
xor \U$43960 ( \44815 , \44814 , \43862 );
buf g885_GF_PartitionCandidate( \44816_nG885 , \44815 );
_DC g886 ( \44817_nG886 , \44816_nG885 , \44261 );
buf \U$43961 ( \44818 , \44817_nG886 );
xor \U$43962 ( \44819 , \43708 , \43711 );
xor \U$43963 ( \44820 , \44819 , \43859 );
buf g7cd_GF_PartitionCandidate( \44821_nG7cd , \44820 );
_DC g7ce ( \44822_nG7ce , \44821_nG7cd , \44261 );
buf \U$43964 ( \44823 , \44822_nG7ce );
xor \U$43965 ( \44824 , \43715 , \43718 );
xor \U$43966 ( \44825 , \44824 , \43856 );
buf g723_GF_PartitionCandidate( \44826_nG723 , \44825 );
_DC g724 ( \44827_nG724 , \44826_nG723 , \44261 );
buf \U$43967 ( \44828 , \44827_nG724 );
xor \U$43968 ( \44829 , \43722 , \43725 );
xor \U$43969 ( \44830 , \44829 , \43853 );
buf g67f_GF_PartitionCandidate( \44831_nG67f , \44830 );
_DC g680 ( \44832_nG680 , \44831_nG67f , \44261 );
buf \U$43970 ( \44833 , \44832_nG680 );
xor \U$43971 ( \44834 , \43729 , \43732 );
xor \U$43972 ( \44835 , \44834 , \43850 );
buf g5e9_GF_PartitionCandidate( \44836_nG5e9 , \44835 );
_DC g5ea ( \44837_nG5ea , \44836_nG5e9 , \44261 );
buf \U$43973 ( \44838 , \44837_nG5ea );
xor \U$43974 ( \44839 , \43736 , \43739 );
xor \U$43975 ( \44840 , \44839 , \43847 );
buf g559_GF_PartitionCandidate( \44841_nG559 , \44840 );
_DC g55a ( \44842_nG55a , \44841_nG559 , \44261 );
buf \U$43976 ( \44843 , \44842_nG55a );
xor \U$43977 ( \44844 , \43743 , \43746 );
xor \U$43978 ( \44845 , \44844 , \43844 );
buf g4d7_GF_PartitionCandidate( \44846_nG4d7 , \44845 );
_DC g4d8 ( \44847_nG4d8 , \44846_nG4d7 , \44261 );
buf \U$43979 ( \44848 , \44847_nG4d8 );
xor \U$43980 ( \44849 , \43750 , \43753 );
xor \U$43981 ( \44850 , \44849 , \43841 );
buf g45b_GF_PartitionCandidate( \44851_nG45b , \44850 );
_DC g45c ( \44852_nG45c , \44851_nG45b , \44261 );
buf \U$43982 ( \44853 , \44852_nG45c );
endmodule

