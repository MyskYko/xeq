//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RI994e460_14,RI994e028_23,RI994dfb0_24,RI994df38_25,RI994e0a0_22,RI994e118_21,RI994e190_20,RI994e208_19,RI994e3e8_15,
        RI994e370_16,RI994e2f8_17,RI994e280_18,RI9921898_610,RI9921820_611,RI99217a8_612,RI9921910_609,RI9921730_613,RI994de48_27,RI98bc948_40,
        RI995e4c8_235,RI98abcb0_53,RI98197a8_66,RI890f600_209,RI99670f0_222,RI89ec0a0_131,RI8946038_144,RI8924e10_183,RI89185e8_196,RI8939810_157,
        RI8930828_170,RI9776ff8_105,RI98084f8_92,RI9808b10_79,RI89ec6b8_118,RI98bc8d0_41,RI994ddd0_28,RI995e450_236,RI9967690_210,RI9967078_223,
        RI98abc38_54,RI9819730_67,RI89465d8_132,RI8939db0_145,RI890fba0_197,RI9808a98_80,RI8930dc8_158,RI89253b0_171,RI8918b88_184,RI89ec640_119,
        RI9776f80_106,RI9808480_93,RI98bc768_44,RI994dc68_31,RI9959f68_239,RI9967528_213,RI995e900_226,RI890fa38_200,RI9808930_83,RI8930c60_161,
        RI8925248_174,RI98195c8_70,RI98abad0_57,RI8946470_135,RI8939c48_148,RI8918a20_187,RI89ec4d8_122,RI9808318_96,RI9776e18_109,RI98082a0_97,
        RI9776da0_110,RI8930be8_162,RI89251d0_175,RI98bc6f0_45,RI994dbf0_32,RI9959860_240,RI99674b0_214,RI995e888_227,RI9819550_71,RI98aba58_58,
        RI89463f8_136,RI8939bd0_149,RI890f9c0_201,RI89189a8_188,RI98088b8_84,RI89ec460_123,RI98abff8_46,RI994d998_241,RI9967438_215,RI98bcc90_33,
        RI995e810_228,RI8946380_137,RI98194d8_72,RI98ab9e0_59,RI8939b58_150,RI9808840_85,RI890f948_202,RI9808228_98,RI9776d28_111,RI8918930_189,
        RI8930b70_163,RI8925158_176,RI89ec3e8_124,RI98abf80_47,RI98bcc18_34,RI994d920_242,RI99673c0_216,RI995e798_229,RI98087c8_86,RI890f8d0_203,
        RI97772c8_99,RI89ec988_112,RI89188b8_190,RI89250e0_177,RI8930af8_164,RI89ec370_125,RI98ab968_60,RI9819460_73,RI8946308_138,RI8939ae0_151,
        RI98abe90_49,RI98bcb28_36,RI994d830_244,RI99672d0_218,RI995e6a8_231,RI98086d8_88,RI890f7e0_205,RI97771d8_101,RI89ec898_114,RI89187c8_192,
        RI8924ff0_179,RI8930a08_166,RI89ec280_127,RI8946218_140,RI89399f0_153,RI9819370_75,RI98ab878_62,RI890f768_206,RI9808660_89,RI9777160_102,
        RI89ec820_115,RI98abe18_50,RI98bcab0_37,RI994d7b8_245,RI9967258_219,RI995e630_232,RI8918750_193,RI8924f78_180,RI8930990_167,RI89ec208_128,
        RI98192f8_76,RI98ab800_63,RI89461a0_141,RI8939978_154,RI89186d8_194,RI89ec190_129,RI98ab788_64,RI9819280_77,RI98abda0_51,RI98bca38_38,
        RI994d740_246,RI995e5b8_233,RI99671e0_220,RI97770e8_103,RI98085e8_90,RI8930918_168,RI8924f00_181,RI8946128_142,RI8939900_155,RI89ec7a8_116,
        RI890f6f0_207,RI9967168_221,RI98abd28_52,RI994d6c8_247,RI98bc9c0_39,RI995e540_234,RI890f678_208,RI89ec730_117,RI9819208_78,RI89308a0_169,
        RI89460b0_143,RI98ab710_65,RI8939888_156,RI8924e88_182,RI9777070_104,RI9808570_91,RI8918660_195,RI89ec118_130,RI994dec0_26,RI994d8a8_243,
        RI9967348_217,RI995e720_230,RI98abf08_48,RI98bcba0_35,RI890f858_204,RI9808750_87,RI9777250_100,RI89ec910_113,RI8918840_191,RI8925068_178,
        RI8930a80_165,RI89ec2f8_126,RI98193e8_74,RI98ab8f0_61,RI8946290_139,RI8939a68_152,RI8918a98_186,RI890fab0_199,RI98089a8_82,RI89ec550_121,
        RI8930cd8_160,RI89252c0_173,RI9776e90_108,RI9808390_95,RI98bc7e0_43,RI994dce0_30,RI9959fe0_238,RI98abb48_56,RI9819640_69,RI89464e8_134,
        RI8939cc0_147,RI99675a0_212,RI995e978_225,RI98bc858_42,RI994dd58_29,RI995e3d8_237,RI98abbc0_55,RI98196b8_68,RI9967618_211,RI99669e8_224,
        RI8946560_133,RI8939d38_146,RI8918b10_185,RI890fb28_198,RI8930d50_159,RI8925338_172,RI9776f08_107,RI9808408_94,RI9808a20_81,RI89ec5c8_120,
        RI9921a00_607,RI9921988_608,RI9921a78_606,RI9921cd0_601,RI9921b68_604,RI9921c58_602,RI9921af0_605,RI9921be0_603,RI994d650_248,RI9931b58_268,
        RI9923878_548,RI9922f18_568,RI992a268_388,RI992f8a8_288,RI9928198_428,RI992c6f8_348,RI992ef48_308,RI9926de8_448,RI9926488_468,RI992abc8_368,
        RI99241d8_528,RI9925b28_488,RI9928af8_408,RI992d058_328,RI9924b38_508,RI994d5d8_249,RI992a1f0_389,RI992f830_289,RI9928120_429,RI992eed0_309,
        RI992b4b0_349,RI9931ae0_269,RI9922bd0_569,RI9923800_549,RI9926d70_449,RI9926410_469,RI9928a80_409,RI9925ab0_489,RI992cfe0_329,RI9924ac0_509,
        RI992ab50_369,RI9924160_529,RI992cf68_330,RI9924a48_510,RI994d560_250,RI9931a68_270,RI9922b58_570,RI9923788_550,RI992aad8_370,RI99240e8_530,
        RI992ee58_310,RI9928a08_410,RI9925a38_490,RI9926cf8_450,RI9926398_470,RI99280a8_430,RI992b438_350,RI992f7b8_290,RI992a178_390,RI9928990_411,
        RI99259c0_491,RI992aa60_371,RI9924070_531,RI992ede0_311,RI9928030_431,RI992b3c0_351,RI9926c80_451,RI9926320_471,RI992f740_291,RI992a100_391,
        RI99319f0_271,RI9922ae0_571,RI9923710_551,RI99249d0_511,RI992cef0_331,RI994d4e8_251,RI9927fb8_432,RI992b348_352,RI9926c08_452,RI99262a8_472,
        RI992f6c8_292,RI9929278_392,RI9928918_412,RI9925948_492,RI992a9e8_372,RI9923ff8_532,RI992ed68_312,RI9931978_272,RI9922a68_572,RI9923698_552,
        RI9924958_512,RI992ce78_332,RI994d470_252,RI9935fc8_254,RI9931888_274,RI9922978_574,RI99235a8_554,RI9929188_394,RI992f5d8_294,RI9927ec8_434,
        RI992d6e8_314,RI992b258_354,RI9926b18_454,RI99261b8_474,RI992a8f8_374,RI9923f08_534,RI9928828_414,RI9925858_494,RI992cd88_334,RI9924868_514,
        RI994d3f8_253,RI9931900_273,RI99229f0_573,RI9923620_553,RI9929200_393,RI992f650_293,RI9927f40_433,RI992ecf0_313,RI992b2d0_353,RI9926b90_453,
        RI9926230_473,RI992a970_373,RI9923f80_533,RI99288a0_413,RI99258d0_493,RI992ce00_333,RI99248e0_513,RI9923e18_536,RI992a808_376,RI9928738_416,
        RI9925768_496,RI992d5f8_316,RI9926a28_456,RI99260c8_476,RI9927dd8_436,RI992b168_356,RI992f4e8_296,RI9929098_396,RI992cc98_336,RI9924778_516,
        RI9931798_276,RI9922888_576,RI99234b8_556,RI9935ed8_256,RI9926140_475,RI9926aa0_455,RI992b1e0_355,RI9927e50_435,RI9929110_395,RI992f560_295,
        RI99257e0_495,RI99287b0_415,RI9923e90_535,RI992a880_375,RI992d670_315,RI99247f0_515,RI992cd10_335,RI9931810_275,RI9923530_555,RI9922900_575,
        RI9935f50_255,RI9933d18_258,RI9928fa8_398,RI9927ce8_438,RI992f3f8_298,RI992d508_318,RI992b078_358,RI99316a8_278,RI9922798_578,RI99233c8_558,
        RI992cba8_338,RI9924688_518,RI9928648_418,RI9925678_498,RI9926938_458,RI9925fd8_478,RI992a718_378,RI9923d28_538,RI99269b0_457,RI9926050_477,
        RI99286c0_417,RI99256f0_497,RI992cc20_337,RI9924700_517,RI992a790_377,RI9923da0_537,RI9933d90_257,RI9929020_397,RI9927d60_437,RI992f470_297,
        RI992d580_317,RI992b0f0_357,RI9931720_277,RI9922810_577,RI9923440_557,RI9933ca0_259,RI9931630_279,RI9922720_579,RI9923350_559,RI9928f30_399,
        RI992f380_299,RI9927c70_439,RI992d490_319,RI992b000_359,RI99268c0_459,RI9925f60_479,RI992a6a0_379,RI9923cb0_539,RI99285d0_419,RI9925600_499,
        RI992cb30_339,RI9924610_519,RI992c9c8_342,RI99244a8_522,RI9933b38_262,RI99314c8_282,RI99225b8_582,RI99231e8_562,RI9923b48_542,RI992a538_382,
        RI992d328_322,RI9925df8_482,RI9926758_462,RI992ae98_362,RI9927b08_442,RI9928dc8_402,RI992f218_302,RI9928468_422,RI9924e08_502,RI9933bb0_261,
        RI9928e40_401,RI9927b80_441,RI992f290_301,RI992d3a0_321,RI992af10_361,RI9931540_281,RI9923260_561,RI9922630_581,RI99267d0_461,RI9925e70_481,
        RI99284e0_421,RI9925510_501,RI992ca40_341,RI9924520_521,RI9923bc0_541,RI992a5b0_381,RI99266e0_463,RI9925d80_483,RI992ae20_363,RI9927040_443,
        RI9928d50_403,RI992f1a0_303,RI992c950_343,RI9924430_523,RI9933ac0_263,RI9931450_283,RI9922540_583,RI9923170_563,RI9923ad0_543,RI992a4c0_383,
        RI992d2b0_323,RI99283f0_423,RI9924d90_503,RI9933c28_260,RI99315b8_280,RI99226a8_580,RI99232d8_560,RI9928eb8_400,RI992f308_300,RI9927bf8_440,
        RI992af88_360,RI992d418_320,RI9925588_500,RI9928558_420,RI992cab8_340,RI9924598_520,RI9925ee8_480,RI9926848_460,RI992a628_380,RI9923c38_540,
        RI9926fc8_444,RI992ada8_364,RI9925d08_484,RI9926668_464,RI992f128_304,RI9928cd8_404,RI992a448_384,RI9923a58_544,RI9928378_424,RI9924d18_504,
        RI992d238_324,RI992c8d8_344,RI99243b8_524,RI99313d8_284,RI99224c8_584,RI99230f8_564,RI9933a48_264,RI99339d0_265,RI9931360_285,RI9922450_585,
        RI9923080_565,RI9928c60_405,RI992f0b0_305,RI9926f50_445,RI992d1c0_325,RI992ad30_365,RI99265f0_465,RI9925c90_485,RI992a3d0_385,RI99239e0_545,
        RI9928300_425,RI9924ca0_505,RI992c860_345,RI9924340_525,RI9926500_467,RI9925ba0_487,RI9926e60_447,RI992ac40_367,RI9928b70_407,RI992efc0_307,
        RI9924250_527,RI992c770_347,RI992f920_287,RI9922f90_567,RI9922360_587,RI99338e0_267,RI992a2e0_387,RI99238f0_547,RI992d0d0_327,RI9928210_427,
        RI9924bb0_507,RI9933958_266,RI99312e8_286,RI99223d8_586,RI9923008_566,RI9928be8_406,RI9926ed8_446,RI992f038_306,RI992d148_326,RI992acb8_366,
        RI9926578_466,RI9925c18_486,RI992a358_386,RI9923968_546,RI9928288_426,RI9924c28_506,RI992c7e8_346,RI99242c8_526,RI99216b8_614,RI9921f28_596,
        RI99222e8_588,RI9922090_593,RI99221f8_590,RI9922180_591,RI9922018_594,RI9921fa0_595,RI9922270_589,RI9922108_592,RI9921eb0_597,RI9921e38_598,
        RI9921dc0_599,RI9921d48_600,RI995ef90_4,RI995ecc0_10,RI995ec48_11,RI995ebd0_12,RI995ed38_9,RI995edb0_8,RI995ee28_7,RI995eea0_6,
        RI995ef18_5,RI995f008_3,RI995f080_2,RI994e4d8_13,RI995f0f8_1,R_289_8400778,R_28a_8401e70,R_28b_8401f18,R_28c_8401fc0,R_28d_8402068,
        R_28e_8402110,R_28f_84021b8,R_290_8402260,R_291_8402308,R_292_84023b0,R_293_8402458,R_294_8402500,R_295_84025a8,R_296_8402650,R_297_84026f8,
        R_298_84027a0,R_299_8402848,R_29a_84028f0,R_29b_8402998,R_29c_8402a40,R_29d_8402ae8,R_29e_8402b90,R_29f_8402c38,R_2a0_8402ce0,R_2a1_8402d88,
        R_2a2_8402e30,R_2a3_8402ed8,R_267_8403418,R_268_8400820,R_269_84008c8,R_26a_8400970,R_26b_8400a18,R_26c_8400ac0,R_26d_8400b68,R_26e_8400c10,
        R_26f_8400cb8,R_270_8400d60,R_271_8400e08,R_272_8400eb0,R_273_8400f58,R_274_8401000,R_275_84010a8,R_276_8401150,R_277_84011f8,R_278_84012a0,
        R_279_8401348,R_27a_84013f0,R_27b_8401498,R_27c_8401540,R_27d_84015e8,R_27e_8401690,R_27f_8401738,R_280_84017e0,R_281_8401888);
input RI994e460_14,RI994e028_23,RI994dfb0_24,RI994df38_25,RI994e0a0_22,RI994e118_21,RI994e190_20,RI994e208_19,RI994e3e8_15,
        RI994e370_16,RI994e2f8_17,RI994e280_18,RI9921898_610,RI9921820_611,RI99217a8_612,RI9921910_609,RI9921730_613,RI994de48_27,RI98bc948_40,
        RI995e4c8_235,RI98abcb0_53,RI98197a8_66,RI890f600_209,RI99670f0_222,RI89ec0a0_131,RI8946038_144,RI8924e10_183,RI89185e8_196,RI8939810_157,
        RI8930828_170,RI9776ff8_105,RI98084f8_92,RI9808b10_79,RI89ec6b8_118,RI98bc8d0_41,RI994ddd0_28,RI995e450_236,RI9967690_210,RI9967078_223,
        RI98abc38_54,RI9819730_67,RI89465d8_132,RI8939db0_145,RI890fba0_197,RI9808a98_80,RI8930dc8_158,RI89253b0_171,RI8918b88_184,RI89ec640_119,
        RI9776f80_106,RI9808480_93,RI98bc768_44,RI994dc68_31,RI9959f68_239,RI9967528_213,RI995e900_226,RI890fa38_200,RI9808930_83,RI8930c60_161,
        RI8925248_174,RI98195c8_70,RI98abad0_57,RI8946470_135,RI8939c48_148,RI8918a20_187,RI89ec4d8_122,RI9808318_96,RI9776e18_109,RI98082a0_97,
        RI9776da0_110,RI8930be8_162,RI89251d0_175,RI98bc6f0_45,RI994dbf0_32,RI9959860_240,RI99674b0_214,RI995e888_227,RI9819550_71,RI98aba58_58,
        RI89463f8_136,RI8939bd0_149,RI890f9c0_201,RI89189a8_188,RI98088b8_84,RI89ec460_123,RI98abff8_46,RI994d998_241,RI9967438_215,RI98bcc90_33,
        RI995e810_228,RI8946380_137,RI98194d8_72,RI98ab9e0_59,RI8939b58_150,RI9808840_85,RI890f948_202,RI9808228_98,RI9776d28_111,RI8918930_189,
        RI8930b70_163,RI8925158_176,RI89ec3e8_124,RI98abf80_47,RI98bcc18_34,RI994d920_242,RI99673c0_216,RI995e798_229,RI98087c8_86,RI890f8d0_203,
        RI97772c8_99,RI89ec988_112,RI89188b8_190,RI89250e0_177,RI8930af8_164,RI89ec370_125,RI98ab968_60,RI9819460_73,RI8946308_138,RI8939ae0_151,
        RI98abe90_49,RI98bcb28_36,RI994d830_244,RI99672d0_218,RI995e6a8_231,RI98086d8_88,RI890f7e0_205,RI97771d8_101,RI89ec898_114,RI89187c8_192,
        RI8924ff0_179,RI8930a08_166,RI89ec280_127,RI8946218_140,RI89399f0_153,RI9819370_75,RI98ab878_62,RI890f768_206,RI9808660_89,RI9777160_102,
        RI89ec820_115,RI98abe18_50,RI98bcab0_37,RI994d7b8_245,RI9967258_219,RI995e630_232,RI8918750_193,RI8924f78_180,RI8930990_167,RI89ec208_128,
        RI98192f8_76,RI98ab800_63,RI89461a0_141,RI8939978_154,RI89186d8_194,RI89ec190_129,RI98ab788_64,RI9819280_77,RI98abda0_51,RI98bca38_38,
        RI994d740_246,RI995e5b8_233,RI99671e0_220,RI97770e8_103,RI98085e8_90,RI8930918_168,RI8924f00_181,RI8946128_142,RI8939900_155,RI89ec7a8_116,
        RI890f6f0_207,RI9967168_221,RI98abd28_52,RI994d6c8_247,RI98bc9c0_39,RI995e540_234,RI890f678_208,RI89ec730_117,RI9819208_78,RI89308a0_169,
        RI89460b0_143,RI98ab710_65,RI8939888_156,RI8924e88_182,RI9777070_104,RI9808570_91,RI8918660_195,RI89ec118_130,RI994dec0_26,RI994d8a8_243,
        RI9967348_217,RI995e720_230,RI98abf08_48,RI98bcba0_35,RI890f858_204,RI9808750_87,RI9777250_100,RI89ec910_113,RI8918840_191,RI8925068_178,
        RI8930a80_165,RI89ec2f8_126,RI98193e8_74,RI98ab8f0_61,RI8946290_139,RI8939a68_152,RI8918a98_186,RI890fab0_199,RI98089a8_82,RI89ec550_121,
        RI8930cd8_160,RI89252c0_173,RI9776e90_108,RI9808390_95,RI98bc7e0_43,RI994dce0_30,RI9959fe0_238,RI98abb48_56,RI9819640_69,RI89464e8_134,
        RI8939cc0_147,RI99675a0_212,RI995e978_225,RI98bc858_42,RI994dd58_29,RI995e3d8_237,RI98abbc0_55,RI98196b8_68,RI9967618_211,RI99669e8_224,
        RI8946560_133,RI8939d38_146,RI8918b10_185,RI890fb28_198,RI8930d50_159,RI8925338_172,RI9776f08_107,RI9808408_94,RI9808a20_81,RI89ec5c8_120,
        RI9921a00_607,RI9921988_608,RI9921a78_606,RI9921cd0_601,RI9921b68_604,RI9921c58_602,RI9921af0_605,RI9921be0_603,RI994d650_248,RI9931b58_268,
        RI9923878_548,RI9922f18_568,RI992a268_388,RI992f8a8_288,RI9928198_428,RI992c6f8_348,RI992ef48_308,RI9926de8_448,RI9926488_468,RI992abc8_368,
        RI99241d8_528,RI9925b28_488,RI9928af8_408,RI992d058_328,RI9924b38_508,RI994d5d8_249,RI992a1f0_389,RI992f830_289,RI9928120_429,RI992eed0_309,
        RI992b4b0_349,RI9931ae0_269,RI9922bd0_569,RI9923800_549,RI9926d70_449,RI9926410_469,RI9928a80_409,RI9925ab0_489,RI992cfe0_329,RI9924ac0_509,
        RI992ab50_369,RI9924160_529,RI992cf68_330,RI9924a48_510,RI994d560_250,RI9931a68_270,RI9922b58_570,RI9923788_550,RI992aad8_370,RI99240e8_530,
        RI992ee58_310,RI9928a08_410,RI9925a38_490,RI9926cf8_450,RI9926398_470,RI99280a8_430,RI992b438_350,RI992f7b8_290,RI992a178_390,RI9928990_411,
        RI99259c0_491,RI992aa60_371,RI9924070_531,RI992ede0_311,RI9928030_431,RI992b3c0_351,RI9926c80_451,RI9926320_471,RI992f740_291,RI992a100_391,
        RI99319f0_271,RI9922ae0_571,RI9923710_551,RI99249d0_511,RI992cef0_331,RI994d4e8_251,RI9927fb8_432,RI992b348_352,RI9926c08_452,RI99262a8_472,
        RI992f6c8_292,RI9929278_392,RI9928918_412,RI9925948_492,RI992a9e8_372,RI9923ff8_532,RI992ed68_312,RI9931978_272,RI9922a68_572,RI9923698_552,
        RI9924958_512,RI992ce78_332,RI994d470_252,RI9935fc8_254,RI9931888_274,RI9922978_574,RI99235a8_554,RI9929188_394,RI992f5d8_294,RI9927ec8_434,
        RI992d6e8_314,RI992b258_354,RI9926b18_454,RI99261b8_474,RI992a8f8_374,RI9923f08_534,RI9928828_414,RI9925858_494,RI992cd88_334,RI9924868_514,
        RI994d3f8_253,RI9931900_273,RI99229f0_573,RI9923620_553,RI9929200_393,RI992f650_293,RI9927f40_433,RI992ecf0_313,RI992b2d0_353,RI9926b90_453,
        RI9926230_473,RI992a970_373,RI9923f80_533,RI99288a0_413,RI99258d0_493,RI992ce00_333,RI99248e0_513,RI9923e18_536,RI992a808_376,RI9928738_416,
        RI9925768_496,RI992d5f8_316,RI9926a28_456,RI99260c8_476,RI9927dd8_436,RI992b168_356,RI992f4e8_296,RI9929098_396,RI992cc98_336,RI9924778_516,
        RI9931798_276,RI9922888_576,RI99234b8_556,RI9935ed8_256,RI9926140_475,RI9926aa0_455,RI992b1e0_355,RI9927e50_435,RI9929110_395,RI992f560_295,
        RI99257e0_495,RI99287b0_415,RI9923e90_535,RI992a880_375,RI992d670_315,RI99247f0_515,RI992cd10_335,RI9931810_275,RI9923530_555,RI9922900_575,
        RI9935f50_255,RI9933d18_258,RI9928fa8_398,RI9927ce8_438,RI992f3f8_298,RI992d508_318,RI992b078_358,RI99316a8_278,RI9922798_578,RI99233c8_558,
        RI992cba8_338,RI9924688_518,RI9928648_418,RI9925678_498,RI9926938_458,RI9925fd8_478,RI992a718_378,RI9923d28_538,RI99269b0_457,RI9926050_477,
        RI99286c0_417,RI99256f0_497,RI992cc20_337,RI9924700_517,RI992a790_377,RI9923da0_537,RI9933d90_257,RI9929020_397,RI9927d60_437,RI992f470_297,
        RI992d580_317,RI992b0f0_357,RI9931720_277,RI9922810_577,RI9923440_557,RI9933ca0_259,RI9931630_279,RI9922720_579,RI9923350_559,RI9928f30_399,
        RI992f380_299,RI9927c70_439,RI992d490_319,RI992b000_359,RI99268c0_459,RI9925f60_479,RI992a6a0_379,RI9923cb0_539,RI99285d0_419,RI9925600_499,
        RI992cb30_339,RI9924610_519,RI992c9c8_342,RI99244a8_522,RI9933b38_262,RI99314c8_282,RI99225b8_582,RI99231e8_562,RI9923b48_542,RI992a538_382,
        RI992d328_322,RI9925df8_482,RI9926758_462,RI992ae98_362,RI9927b08_442,RI9928dc8_402,RI992f218_302,RI9928468_422,RI9924e08_502,RI9933bb0_261,
        RI9928e40_401,RI9927b80_441,RI992f290_301,RI992d3a0_321,RI992af10_361,RI9931540_281,RI9923260_561,RI9922630_581,RI99267d0_461,RI9925e70_481,
        RI99284e0_421,RI9925510_501,RI992ca40_341,RI9924520_521,RI9923bc0_541,RI992a5b0_381,RI99266e0_463,RI9925d80_483,RI992ae20_363,RI9927040_443,
        RI9928d50_403,RI992f1a0_303,RI992c950_343,RI9924430_523,RI9933ac0_263,RI9931450_283,RI9922540_583,RI9923170_563,RI9923ad0_543,RI992a4c0_383,
        RI992d2b0_323,RI99283f0_423,RI9924d90_503,RI9933c28_260,RI99315b8_280,RI99226a8_580,RI99232d8_560,RI9928eb8_400,RI992f308_300,RI9927bf8_440,
        RI992af88_360,RI992d418_320,RI9925588_500,RI9928558_420,RI992cab8_340,RI9924598_520,RI9925ee8_480,RI9926848_460,RI992a628_380,RI9923c38_540,
        RI9926fc8_444,RI992ada8_364,RI9925d08_484,RI9926668_464,RI992f128_304,RI9928cd8_404,RI992a448_384,RI9923a58_544,RI9928378_424,RI9924d18_504,
        RI992d238_324,RI992c8d8_344,RI99243b8_524,RI99313d8_284,RI99224c8_584,RI99230f8_564,RI9933a48_264,RI99339d0_265,RI9931360_285,RI9922450_585,
        RI9923080_565,RI9928c60_405,RI992f0b0_305,RI9926f50_445,RI992d1c0_325,RI992ad30_365,RI99265f0_465,RI9925c90_485,RI992a3d0_385,RI99239e0_545,
        RI9928300_425,RI9924ca0_505,RI992c860_345,RI9924340_525,RI9926500_467,RI9925ba0_487,RI9926e60_447,RI992ac40_367,RI9928b70_407,RI992efc0_307,
        RI9924250_527,RI992c770_347,RI992f920_287,RI9922f90_567,RI9922360_587,RI99338e0_267,RI992a2e0_387,RI99238f0_547,RI992d0d0_327,RI9928210_427,
        RI9924bb0_507,RI9933958_266,RI99312e8_286,RI99223d8_586,RI9923008_566,RI9928be8_406,RI9926ed8_446,RI992f038_306,RI992d148_326,RI992acb8_366,
        RI9926578_466,RI9925c18_486,RI992a358_386,RI9923968_546,RI9928288_426,RI9924c28_506,RI992c7e8_346,RI99242c8_526,RI99216b8_614,RI9921f28_596,
        RI99222e8_588,RI9922090_593,RI99221f8_590,RI9922180_591,RI9922018_594,RI9921fa0_595,RI9922270_589,RI9922108_592,RI9921eb0_597,RI9921e38_598,
        RI9921dc0_599,RI9921d48_600,RI995ef90_4,RI995ecc0_10,RI995ec48_11,RI995ebd0_12,RI995ed38_9,RI995edb0_8,RI995ee28_7,RI995eea0_6,
        RI995ef18_5,RI995f008_3,RI995f080_2,RI994e4d8_13,RI995f0f8_1;
output R_289_8400778,R_28a_8401e70,R_28b_8401f18,R_28c_8401fc0,R_28d_8402068,R_28e_8402110,R_28f_84021b8,R_290_8402260,R_291_8402308,
        R_292_84023b0,R_293_8402458,R_294_8402500,R_295_84025a8,R_296_8402650,R_297_84026f8,R_298_84027a0,R_299_8402848,R_29a_84028f0,R_29b_8402998,
        R_29c_8402a40,R_29d_8402ae8,R_29e_8402b90,R_29f_8402c38,R_2a0_8402ce0,R_2a1_8402d88,R_2a2_8402e30,R_2a3_8402ed8,R_267_8403418,R_268_8400820,
        R_269_84008c8,R_26a_8400970,R_26b_8400a18,R_26c_8400ac0,R_26d_8400b68,R_26e_8400c10,R_26f_8400cb8,R_270_8400d60,R_271_8400e08,R_272_8400eb0,
        R_273_8400f58,R_274_8401000,R_275_84010a8,R_276_8401150,R_277_84011f8,R_278_84012a0,R_279_8401348,R_27a_84013f0,R_27b_8401498,R_27c_8401540,
        R_27d_84015e8,R_27e_8401690,R_27f_8401738,R_280_84017e0,R_281_8401888;

wire \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677_N$1 ,
         \678_N$2 , \679_N$4 , \680_N$5 , \681_N$6 , \682_N$7 , \683_N$9 , \684_N$10 , \685_ZERO , \686 , \687 ,
         \688 , \689_N$3 , \690_N$8 , \691_N$11 , \692_ONE , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 ,
         \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 ,
         \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 ,
         \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 ,
         \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 ,
         \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 ,
         \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 ,
         \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 ,
         \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 ,
         \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 ,
         \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 ,
         \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 ,
         \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 ,
         \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 ,
         \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 ,
         \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 ,
         \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 ,
         \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 ,
         \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 ,
         \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 ,
         \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 ,
         \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 ,
         \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 ,
         \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 ,
         \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 ,
         \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 ,
         \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 ,
         \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 ,
         \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 ,
         \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 ,
         \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 ,
         \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 ,
         \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 ,
         \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 ,
         \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 ,
         \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 ,
         \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 ,
         \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 ,
         \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 ,
         \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 ,
         \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 ,
         \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 ,
         \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 ,
         \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 ,
         \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 ,
         \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 ,
         \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 ,
         \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 ,
         \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 ,
         \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 ,
         \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 ,
         \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 ,
         \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 ,
         \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 ,
         \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 ,
         \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 ,
         \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 ,
         \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 ,
         \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 ,
         \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 ,
         \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 ,
         \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 ,
         \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 ,
         \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 ,
         \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 ,
         \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 ,
         \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 ,
         \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 ,
         \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 ,
         \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 ,
         \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 ,
         \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 ,
         \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 ,
         \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 ,
         \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 ,
         \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 ,
         \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 ,
         \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 ,
         \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 ,
         \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 ,
         \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 ,
         \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 ,
         \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 ,
         \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 ,
         \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 ,
         \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 ,
         \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 ,
         \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 ,
         \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 ,
         \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 ,
         \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 ,
         \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 ,
         \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 ,
         \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 ,
         \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 ,
         \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 ,
         \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 ,
         \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 ,
         \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 ,
         \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 ,
         \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 ,
         \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 ,
         \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 ,
         \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 ,
         \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 ,
         \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 ,
         \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 ,
         \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 ,
         \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 ,
         \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 ,
         \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 ,
         \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 ,
         \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 ,
         \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 ,
         \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 ,
         \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 ,
         \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 ,
         \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 ,
         \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 ,
         \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 ,
         \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 ,
         \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 ,
         \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 ,
         \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 ,
         \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 ,
         \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 ,
         \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 ,
         \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 ,
         \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 ,
         \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 ,
         \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 ,
         \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 ,
         \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 ,
         \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 ,
         \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 ,
         \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 ,
         \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 ,
         \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 ,
         \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 ,
         \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 ,
         \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 ,
         \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 ,
         \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 ,
         \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 ,
         \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 ,
         \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 ,
         \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 ,
         \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 ,
         \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 ,
         \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 ,
         \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 ,
         \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 ,
         \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 ,
         \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 ,
         \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 ,
         \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 ,
         \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 ,
         \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 ,
         \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 ,
         \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 ,
         \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 ,
         \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 ,
         \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 ,
         \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 ,
         \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 ,
         \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 ,
         \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 ,
         \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 ,
         \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 ,
         \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 ,
         \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 ,
         \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 ,
         \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 ,
         \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 ,
         \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 ,
         \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 ,
         \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 ,
         \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 ,
         \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 ,
         \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 ,
         \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 ,
         \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 ,
         \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 ,
         \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 ,
         \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 ,
         \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 ,
         \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 ,
         \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 ,
         \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 ,
         \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 ,
         \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 ,
         \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 ,
         \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 ,
         \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 ,
         \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 ,
         \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 ,
         \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 ,
         \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 ,
         \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 ,
         \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 ,
         \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 ,
         \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 ,
         \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 ,
         \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 ,
         \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 ,
         \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 ,
         \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 ,
         \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 ,
         \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 ,
         \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 ,
         \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 ,
         \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 ,
         \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 ,
         \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 ,
         \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 ,
         \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 ,
         \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 ,
         \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 ,
         \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 ,
         \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 ,
         \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 ,
         \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 ,
         \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 ,
         \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 ,
         \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 ,
         \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 ,
         \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 ,
         \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 ,
         \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 ,
         \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 ,
         \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 ,
         \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 ,
         \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 ,
         \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 ,
         \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 ,
         \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 ,
         \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 ,
         \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 ,
         \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 ,
         \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 ,
         \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 ,
         \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 ,
         \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 ,
         \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 ,
         \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 ,
         \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 ,
         \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 ,
         \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 ,
         \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 ,
         \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 ,
         \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 ,
         \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 ,
         \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 ,
         \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 ,
         \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 ,
         \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 ,
         \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 ,
         \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 ,
         \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 ,
         \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 ,
         \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 ,
         \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 ,
         \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 ,
         \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 ,
         \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 ,
         \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 ,
         \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 ,
         \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 ,
         \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 ,
         \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 ,
         \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 ,
         \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 ,
         \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 ,
         \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 ,
         \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 ,
         \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 ,
         \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 ,
         \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 ,
         \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 ,
         \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 ,
         \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 ,
         \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 ,
         \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 ,
         \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 ,
         \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 ,
         \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 ,
         \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 ,
         \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 ,
         \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 ,
         \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 ,
         \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 ,
         \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 ,
         \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 ,
         \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 ,
         \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 ,
         \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 ,
         \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 ,
         \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 ,
         \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 ,
         \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 ,
         \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 ,
         \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 ,
         \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 ,
         \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 ,
         \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 ,
         \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 ,
         \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 ,
         \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 ,
         \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 ,
         \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 ,
         \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 ,
         \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 ,
         \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 ,
         \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 ,
         \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 ,
         \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 ,
         \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 ,
         \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 ,
         \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 ,
         \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 ,
         \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 ,
         \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 ,
         \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 ,
         \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 ,
         \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 ,
         \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 ,
         \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 ,
         \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 ,
         \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 ,
         \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 ,
         \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 ,
         \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 ,
         \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 ,
         \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 ,
         \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 ,
         \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 ,
         \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 ,
         \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 ,
         \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 ,
         \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 ,
         \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 ,
         \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 ,
         \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 ,
         \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 ,
         \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 ,
         \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 ,
         \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 ,
         \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 ,
         \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 ,
         \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 ,
         \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 ,
         \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 ,
         \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 ,
         \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 ,
         \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 ,
         \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 ,
         \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 ,
         \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 ,
         \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 ,
         \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 ,
         \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 ,
         \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 ,
         \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 ,
         \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 ,
         \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 ,
         \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 ,
         \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 ,
         \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 ,
         \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 ,
         \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 ,
         \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 ,
         \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 ,
         \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 ,
         \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 ,
         \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 ,
         \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 ,
         \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 ,
         \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 ,
         \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 ,
         \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 ,
         \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 ,
         \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 ,
         \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 ,
         \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 ,
         \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 ,
         \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 ,
         \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 ,
         \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 ,
         \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 ,
         \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 ,
         \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 ,
         \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 ,
         \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 ,
         \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 ,
         \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 ,
         \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 ,
         \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 ,
         \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 ,
         \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 ,
         \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 ,
         \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 ,
         \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 ,
         \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 ,
         \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 ,
         \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 ,
         \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 ,
         \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 ,
         \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 ,
         \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 ,
         \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 ,
         \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 ,
         \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 ,
         \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 ,
         \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 ,
         \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 ,
         \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 ,
         \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 ,
         \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 ,
         \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 ,
         \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 ,
         \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 ,
         \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 ,
         \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 ,
         \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 ,
         \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 ,
         \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 ,
         \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 ,
         \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 ,
         \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 ,
         \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 ,
         \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 ,
         \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 ,
         \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 ,
         \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 ,
         \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 ,
         \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 ,
         \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 ,
         \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 ,
         \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 ,
         \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 ,
         \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 ,
         \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 ,
         \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 ,
         \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 ,
         \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 ,
         \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 ,
         \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 ,
         \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 ,
         \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 ,
         \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 ,
         \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 ,
         \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 ,
         \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 ,
         \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 ,
         \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 ,
         \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 ,
         \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 ,
         \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 ,
         \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 ,
         \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 ,
         \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 ,
         \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 ,
         \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 ,
         \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 ,
         \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 ,
         \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 ,
         \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 ,
         \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 ,
         \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 ,
         \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 ,
         \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 ,
         \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 ,
         \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 ,
         \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 ,
         \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 ,
         \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 ,
         \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 ,
         \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 ,
         \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 ,
         \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 ,
         \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 ,
         \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 ,
         \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 ,
         \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 ,
         \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 ,
         \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 ,
         \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 ,
         \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 ,
         \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 ,
         \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 ,
         \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 ,
         \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 ,
         \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 ,
         \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 ,
         \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 ,
         \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 ,
         \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 ,
         \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 ,
         \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 ,
         \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 ,
         \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 ,
         \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 ,
         \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 ,
         \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 ,
         \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 ,
         \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 ,
         \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 ,
         \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 ,
         \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 ,
         \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 ,
         \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 ,
         \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 ,
         \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 ,
         \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 ,
         \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 ,
         \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 ,
         \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 ,
         \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 ,
         \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 ,
         \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 ,
         \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 ,
         \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 ,
         \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 ,
         \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 ,
         \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 ,
         \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 ,
         \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 ,
         \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 ,
         \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 ,
         \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 ,
         \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 ,
         \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 ,
         \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 ,
         \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 ,
         \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 ,
         \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 ,
         \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 ,
         \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 ,
         \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 ,
         \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 ,
         \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 ,
         \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 ,
         \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 ,
         \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 ,
         \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 ,
         \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 ,
         \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 ,
         \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 ,
         \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 ,
         \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 ,
         \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 ,
         \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 ,
         \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 ,
         \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 ,
         \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 ,
         \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 ,
         \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 ,
         \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 ,
         \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 ,
         \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 ,
         \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 ,
         \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 ,
         \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 ,
         \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 ,
         \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 ,
         \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 ,
         \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 ,
         \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 ,
         \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 ,
         \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 ,
         \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 ,
         \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 ,
         \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 ,
         \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 ,
         \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 ,
         \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 ,
         \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 ,
         \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 ,
         \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 ,
         \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 ,
         \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 ,
         \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 ,
         \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 ,
         \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 ,
         \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 ,
         \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 ,
         \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 ,
         \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 ,
         \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 ,
         \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 ,
         \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 ,
         \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 ,
         \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 ,
         \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 ,
         \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 ,
         \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 ,
         \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 ,
         \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 ,
         \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 ,
         \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 ,
         \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 ,
         \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 ,
         \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 ,
         \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 ,
         \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 ,
         \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 ,
         \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 ,
         \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 ,
         \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 ,
         \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 ,
         \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 ,
         \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 ,
         \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 ,
         \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 ,
         \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 ,
         \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 ,
         \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 ,
         \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 ,
         \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 ,
         \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 ,
         \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 ,
         \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 ,
         \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 ,
         \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 ,
         \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 ,
         \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 ,
         \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 ,
         \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 ,
         \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 ,
         \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 ,
         \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 ,
         \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 ,
         \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 ,
         \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 ,
         \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 ,
         \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 ,
         \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
         \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 ,
         \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 ,
         \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 ,
         \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 ,
         \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 ,
         \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 ,
         \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 ,
         \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 ,
         \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 ,
         \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 ,
         \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 ,
         \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 ,
         \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 ,
         \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 ,
         \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 ,
         \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 ,
         \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 ,
         \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 ,
         \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 ,
         \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 ,
         \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 ,
         \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 ,
         \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 ,
         \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 ,
         \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 ,
         \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 ,
         \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 ,
         \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 ,
         \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 ,
         \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 ,
         \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 ,
         \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 ,
         \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 ,
         \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 ,
         \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 ,
         \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 ,
         \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 ,
         \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 ,
         \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 ,
         \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 ,
         \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 ,
         \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 ,
         \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 ,
         \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 ,
         \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 ,
         \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 ,
         \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 ,
         \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 ,
         \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 ,
         \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 ,
         \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 ,
         \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 ,
         \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 ,
         \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 ,
         \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 ,
         \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 ,
         \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 ,
         \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 ,
         \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 ,
         \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 ,
         \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 ,
         \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 ,
         \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 ,
         \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 ,
         \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 ,
         \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 ,
         \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 ,
         \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 ,
         \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 ,
         \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 ,
         \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 ,
         \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 ,
         \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 ,
         \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 ,
         \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 ,
         \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 ,
         \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 ,
         \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 ,
         \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 ,
         \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 ,
         \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 ,
         \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 ,
         \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 ,
         \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 ,
         \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 ,
         \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 ,
         \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 ,
         \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 ,
         \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 ,
         \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 ,
         \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 ,
         \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 ,
         \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 ,
         \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 ,
         \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 ,
         \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 ,
         \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 ,
         \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 ,
         \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 ,
         \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 ,
         \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 ,
         \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 ,
         \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 ,
         \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 ,
         \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 ,
         \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 ,
         \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 ,
         \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 ,
         \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 ,
         \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 ,
         \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 ,
         \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 ,
         \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 ,
         \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 ,
         \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 ,
         \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 ,
         \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 ,
         \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 ,
         \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 ,
         \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 ,
         \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 ,
         \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 ,
         \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 ,
         \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 ,
         \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 ,
         \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 ,
         \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 ,
         \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 ,
         \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 ,
         \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 ,
         \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 ,
         \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 ,
         \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 ,
         \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 ,
         \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 ,
         \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 ,
         \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 ,
         \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 ,
         \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 ,
         \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 ,
         \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 ,
         \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 ,
         \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 ,
         \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 ,
         \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 ,
         \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 ,
         \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 ,
         \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 ,
         \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 ,
         \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 ,
         \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 ,
         \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 ,
         \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 ,
         \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 ,
         \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 ,
         \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 ,
         \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 ,
         \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 ,
         \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 ,
         \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 ,
         \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 ,
         \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 ,
         \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 ,
         \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 ,
         \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 ,
         \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 ,
         \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 ,
         \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 ,
         \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 ,
         \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 ,
         \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 ,
         \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 ,
         \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 ,
         \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 ,
         \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 ,
         \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 ,
         \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 ,
         \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 ,
         \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 ,
         \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 ,
         \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 ,
         \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 ,
         \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 ,
         \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 ,
         \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 ,
         \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 ,
         \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 ,
         \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 ,
         \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 ,
         \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 ,
         \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 ,
         \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 ,
         \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 ,
         \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 ,
         \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 ,
         \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 ,
         \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 ,
         \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 ,
         \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 ,
         \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 ,
         \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 ,
         \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 ,
         \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 ,
         \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 ,
         \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 ,
         \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 ,
         \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 ,
         \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 ,
         \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 ,
         \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 ,
         \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 ,
         \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 ,
         \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 ,
         \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 ,
         \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 ,
         \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 ,
         \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 ,
         \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 ,
         \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 ,
         \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 ,
         \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 ,
         \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 ,
         \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 ,
         \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 ,
         \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 ,
         \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 ,
         \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 ,
         \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 ,
         \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 ,
         \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 ,
         \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 ,
         \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 ,
         \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 ,
         \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 ,
         \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 ,
         \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 ,
         \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 ,
         \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 ,
         \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 ,
         \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 ,
         \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 ,
         \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 ,
         \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 ,
         \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 ,
         \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 ,
         \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 ,
         \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 ,
         \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 ,
         \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 ,
         \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 ,
         \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 ,
         \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 ,
         \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 ,
         \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 ,
         \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 ,
         \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 ,
         \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 ,
         \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 ,
         \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 ,
         \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 ,
         \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 ,
         \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 ,
         \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 ,
         \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 ,
         \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 ,
         \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 ,
         \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 ,
         \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 ,
         \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 ,
         \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 ,
         \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 ,
         \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 ,
         \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 ,
         \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 ,
         \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 ,
         \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 ,
         \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 ,
         \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 ,
         \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 ,
         \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 ,
         \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 ,
         \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 ,
         \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 ,
         \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 ,
         \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 ,
         \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 ,
         \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 ,
         \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 ,
         \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 ,
         \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 ,
         \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 ,
         \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 ,
         \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 ,
         \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 ,
         \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 ,
         \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 ,
         \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 ,
         \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 ,
         \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 ,
         \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 ,
         \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 ,
         \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 ,
         \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 ,
         \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 ,
         \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 ,
         \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 ,
         \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 ,
         \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 ,
         \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 ,
         \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 ,
         \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 ,
         \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 ,
         \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 ,
         \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 ,
         \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 ,
         \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 ,
         \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 ,
         \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 ,
         \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 ,
         \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 ,
         \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 ,
         \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 ,
         \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 ,
         \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 ,
         \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 ,
         \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 ,
         \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 ,
         \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 ,
         \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 ,
         \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 ,
         \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 ,
         \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 ,
         \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 ,
         \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 ,
         \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 ,
         \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 ,
         \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 ,
         \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 ,
         \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 ,
         \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 ,
         \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 ,
         \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 ,
         \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 ,
         \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 ,
         \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 ,
         \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 ,
         \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 ,
         \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 ,
         \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 ,
         \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 ,
         \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 ,
         \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 ,
         \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 ,
         \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 ,
         \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 ,
         \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 ,
         \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 ,
         \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 ,
         \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 ,
         \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 ,
         \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 ,
         \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 ,
         \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 ,
         \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 ,
         \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 ,
         \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 ,
         \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 ,
         \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 ,
         \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 ,
         \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 ,
         \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 ,
         \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 ,
         \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 ,
         \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 ,
         \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 ,
         \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 ,
         \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 ,
         \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 ,
         \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 ,
         \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 ,
         \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 ,
         \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 ,
         \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 ,
         \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 ,
         \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 ,
         \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 ,
         \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 ,
         \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 ,
         \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 ,
         \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 ,
         \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 ,
         \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 ,
         \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 ,
         \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 ,
         \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 ,
         \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 ,
         \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 ,
         \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 ,
         \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 ,
         \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 ,
         \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 ,
         \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 ,
         \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 ,
         \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 ,
         \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 ,
         \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 ,
         \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 ,
         \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 ,
         \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 ,
         \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 ,
         \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 ,
         \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 ,
         \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 ,
         \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 ,
         \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 ,
         \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 ,
         \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 ,
         \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 ,
         \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 ,
         \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 ,
         \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 ,
         \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 ,
         \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 ,
         \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 ,
         \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 ,
         \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 ,
         \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 ,
         \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 ,
         \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 ,
         \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 ,
         \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 ,
         \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 ,
         \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 ,
         \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 ,
         \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 ,
         \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 ,
         \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 ,
         \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 ,
         \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 ,
         \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 ,
         \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 ,
         \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 ,
         \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 ,
         \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 ,
         \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 ,
         \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 ,
         \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 ,
         \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 ,
         \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 ,
         \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 ,
         \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 ,
         \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 ,
         \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 ,
         \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 ,
         \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 ,
         \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 ,
         \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 ,
         \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 ,
         \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 ,
         \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 ,
         \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 ,
         \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 ,
         \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 ,
         \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 ,
         \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 ,
         \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 ,
         \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 ,
         \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 ,
         \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 ,
         \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 ,
         \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 ,
         \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 ,
         \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 ,
         \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 ,
         \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 ,
         \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 ,
         \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 ,
         \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 ,
         \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 ,
         \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 ,
         \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 ,
         \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 ,
         \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 ,
         \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 ,
         \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 ,
         \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 ,
         \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 ,
         \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 ,
         \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 ,
         \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 ,
         \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 ,
         \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 ,
         \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 ,
         \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 ,
         \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 ,
         \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 ,
         \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 ,
         \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 ,
         \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 ,
         \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 ,
         \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 ,
         \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 ,
         \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 ,
         \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 ,
         \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 ,
         \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 ,
         \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 ,
         \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 ,
         \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 ,
         \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 ,
         \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 ,
         \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 ,
         \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 ,
         \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 ,
         \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 ,
         \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 ,
         \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 ,
         \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 ,
         \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 ,
         \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 ,
         \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 ,
         \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 ,
         \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 ,
         \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 ,
         \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 ,
         \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 ,
         \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 ,
         \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 ,
         \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 ,
         \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 ,
         \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 ,
         \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 ,
         \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 ,
         \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 ,
         \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 ,
         \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 ,
         \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 ,
         \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 ,
         \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 ,
         \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 ,
         \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 ,
         \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 ,
         \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 ,
         \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 ,
         \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 ,
         \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 ,
         \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 ,
         \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 ,
         \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 ,
         \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 ,
         \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 ,
         \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 ,
         \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 ,
         \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 ,
         \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 ,
         \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 ,
         \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 ,
         \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 ,
         \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 ,
         \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 ,
         \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 ,
         \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 ,
         \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 ,
         \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 ,
         \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 ,
         \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 ,
         \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 ,
         \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 ,
         \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 ,
         \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 ,
         \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 ,
         \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 ,
         \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 ,
         \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 ,
         \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 ,
         \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 ,
         \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 ,
         \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 ,
         \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 ,
         \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 ,
         \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 ,
         \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 ,
         \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 ,
         \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 ,
         \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 ,
         \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 ,
         \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 ,
         \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 ,
         \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 ,
         \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 ,
         \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 ,
         \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 ,
         \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 ,
         \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 ,
         \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 ,
         \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 ,
         \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 ,
         \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 ,
         \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 ,
         \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 ,
         \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 ,
         \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 ,
         \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 ,
         \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 ,
         \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 ,
         \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 ,
         \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 ,
         \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 ,
         \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 ,
         \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 ,
         \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 ,
         \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 ,
         \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 ,
         \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 ,
         \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 ,
         \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 ,
         \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 ,
         \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 ,
         \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 ,
         \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 ,
         \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 ,
         \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 ,
         \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 ,
         \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 ,
         \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 ,
         \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 ,
         \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 ,
         \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 ,
         \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 ,
         \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 ,
         \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 ,
         \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 ,
         \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 ,
         \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 ,
         \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 ,
         \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 ,
         \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 ,
         \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 ,
         \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 ,
         \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 ,
         \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 ,
         \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 ,
         \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 ,
         \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 ,
         \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 ,
         \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 ,
         \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 ,
         \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 ,
         \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 ,
         \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 ,
         \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 ,
         \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 ,
         \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 ,
         \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 ,
         \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 ,
         \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 ,
         \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 ,
         \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 ,
         \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 ,
         \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 ,
         \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 ,
         \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 ,
         \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 ,
         \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 ,
         \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 ,
         \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 ,
         \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 ,
         \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 ,
         \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 ,
         \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 ,
         \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 ,
         \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 ,
         \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 ,
         \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 ,
         \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 ,
         \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 ,
         \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 ,
         \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 ,
         \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 ,
         \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 ,
         \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 ,
         \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 ,
         \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 ,
         \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 ,
         \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 ,
         \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 ,
         \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 ,
         \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 ,
         \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 ,
         \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 ,
         \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 ,
         \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 ,
         \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 ,
         \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 ,
         \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 ,
         \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 ,
         \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 ,
         \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 ,
         \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 ,
         \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 ,
         \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 ,
         \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 ,
         \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 ,
         \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 ,
         \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 ,
         \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 ,
         \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 ,
         \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 ,
         \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 ,
         \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 ,
         \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 ,
         \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 ,
         \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 ,
         \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 ,
         \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 ,
         \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 ,
         \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 ,
         \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 ,
         \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 ,
         \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 ,
         \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 ,
         \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 ,
         \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 ,
         \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 ,
         \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 ,
         \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 ,
         \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 ,
         \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 ,
         \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 ,
         \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 ,
         \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 ,
         \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 ,
         \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 ,
         \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 ,
         \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 ,
         \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 ,
         \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 ,
         \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 ,
         \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 ,
         \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 ,
         \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 ,
         \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 ,
         \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 ,
         \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 ,
         \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 ,
         \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 ,
         \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 ,
         \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 ,
         \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 ,
         \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 ,
         \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 ,
         \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 ,
         \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 ,
         \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 ,
         \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 ,
         \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 ,
         \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 ,
         \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 ,
         \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 ,
         \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 ,
         \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 ,
         \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 ,
         \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 ,
         \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 ,
         \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 ,
         \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 ,
         \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 ,
         \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 ,
         \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 ,
         \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 ,
         \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 ,
         \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 ,
         \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 ,
         \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 ,
         \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 ,
         \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 ,
         \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 ,
         \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 ,
         \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 ,
         \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 ,
         \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 ,
         \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 ,
         \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 ,
         \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 ,
         \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 ,
         \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 ,
         \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 ,
         \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 ,
         \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 ,
         \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 ,
         \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 ,
         \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 ,
         \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 ,
         \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 ,
         \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 ,
         \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 ,
         \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 ,
         \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 ,
         \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 ,
         \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 ,
         \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 ,
         \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 ,
         \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 ,
         \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 ,
         \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 ,
         \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 ,
         \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 ,
         \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 ,
         \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 ,
         \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 ,
         \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 ,
         \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 ,
         \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 ,
         \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 ,
         \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 ,
         \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 ,
         \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 ,
         \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 ,
         \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 ,
         \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 ,
         \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 ,
         \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 ,
         \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 ,
         \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 ,
         \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 ,
         \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 ,
         \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 ,
         \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 ,
         \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 ,
         \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 ,
         \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 ,
         \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 ,
         \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 ,
         \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 ,
         \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 ,
         \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 ,
         \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 ,
         \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 ,
         \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 ,
         \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 ,
         \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 ,
         \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 ,
         \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 ,
         \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 ,
         \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 ,
         \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 ,
         \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 ,
         \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 ,
         \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 ,
         \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 ,
         \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 ,
         \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 ,
         \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 ,
         \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 ,
         \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 ,
         \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 ,
         \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 ,
         \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 ,
         \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 ,
         \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 ,
         \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 ,
         \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 ,
         \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 ,
         \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 ,
         \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 ,
         \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 ,
         \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 ,
         \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 ,
         \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 ,
         \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 ,
         \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 ,
         \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 ,
         \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 ,
         \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 ,
         \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 ,
         \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 ,
         \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 ,
         \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 ,
         \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 ,
         \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 ,
         \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 ,
         \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 ,
         \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 ,
         \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 ,
         \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 ,
         \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 ,
         \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 ,
         \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 ,
         \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 ,
         \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 ,
         \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 ,
         \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 ,
         \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 ,
         \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 ,
         \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 ,
         \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 ,
         \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 ,
         \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 ,
         \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 ,
         \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 ,
         \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 ,
         \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 ,
         \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 ,
         \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 ,
         \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 ,
         \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 ,
         \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 ,
         \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 ,
         \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 ,
         \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 ,
         \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 ,
         \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 ,
         \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 ,
         \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 ,
         \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 ,
         \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 ,
         \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 ,
         \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 ,
         \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 ,
         \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 ,
         \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 ,
         \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 ,
         \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 ,
         \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 ,
         \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 ,
         \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 ,
         \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 ,
         \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 ,
         \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 ,
         \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 ,
         \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 ,
         \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 ,
         \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 ,
         \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 ,
         \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 ,
         \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 ,
         \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 ,
         \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 ,
         \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 ,
         \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 ,
         \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 ,
         \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 ,
         \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 ,
         \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 ,
         \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 ,
         \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 ,
         \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 ,
         \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 ,
         \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 ,
         \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 ,
         \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 ,
         \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 ,
         \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 ,
         \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 ,
         \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 ,
         \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 ,
         \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 ,
         \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 ,
         \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 ,
         \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 ,
         \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 ,
         \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 ,
         \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 ,
         \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 ,
         \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 ,
         \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 ,
         \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 ,
         \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 ,
         \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 ,
         \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 ,
         \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 ,
         \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 ,
         \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 ,
         \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 ,
         \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 ,
         \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 ,
         \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 ,
         \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 ,
         \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 ,
         \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 ,
         \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 ,
         \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 ,
         \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 ,
         \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 ,
         \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 ,
         \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 ,
         \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 ,
         \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 ,
         \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 ,
         \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 ,
         \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 ,
         \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 ,
         \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 ,
         \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 ,
         \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 ,
         \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 ,
         \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 ,
         \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 ,
         \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 ,
         \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 ,
         \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 ,
         \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 ,
         \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 ,
         \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 ,
         \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 ,
         \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 ,
         \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 ,
         \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 ,
         \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 ,
         \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 ,
         \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 ,
         \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 ,
         \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 ,
         \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 ,
         \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 ,
         \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 ,
         \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 ,
         \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 ,
         \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 ,
         \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 ,
         \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 ,
         \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 ,
         \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 ,
         \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 ,
         \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 ,
         \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 ,
         \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 ,
         \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 ,
         \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 ,
         \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 ,
         \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 ,
         \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 ,
         \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 ,
         \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 ,
         \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 ,
         \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 ,
         \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 ,
         \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 ,
         \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 ,
         \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 ,
         \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 ,
         \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 ,
         \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 ,
         \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 ,
         \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 ,
         \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 ,
         \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 ,
         \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 ,
         \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 ,
         \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 ,
         \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 ,
         \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 ,
         \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 ,
         \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 ,
         \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 ,
         \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 ,
         \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 ,
         \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 ,
         \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 ,
         \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 ,
         \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 ,
         \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 ,
         \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 ,
         \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 ,
         \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 ,
         \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 ,
         \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 ,
         \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 ,
         \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 ,
         \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 ,
         \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 ,
         \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 ,
         \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 ,
         \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 ,
         \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 ,
         \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 ,
         \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 ,
         \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 ,
         \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 ,
         \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 ,
         \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 ,
         \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 ,
         \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 ,
         \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 ,
         \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 ,
         \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 ,
         \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 ,
         \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 ,
         \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 ,
         \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 ,
         \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 ,
         \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 ,
         \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 ,
         \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 ,
         \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 ,
         \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 ,
         \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 ,
         \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 ,
         \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 ,
         \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 ,
         \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 ,
         \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 ,
         \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 ,
         \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 ,
         \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 ,
         \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 ,
         \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 ,
         \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 ,
         \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 ,
         \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 ,
         \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 ,
         \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 ,
         \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 ,
         \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 ,
         \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 ,
         \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 ,
         \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 ,
         \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 ,
         \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 ,
         \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 ,
         \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 ,
         \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 ,
         \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 ,
         \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 ,
         \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 ,
         \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 ,
         \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 ,
         \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 ,
         \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 ,
         \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 ,
         \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 ,
         \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 ,
         \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 ,
         \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 ,
         \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 ,
         \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 ,
         \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 ,
         \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 ,
         \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 ,
         \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 ,
         \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 ,
         \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 ,
         \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 ,
         \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 ,
         \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 ,
         \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 ,
         \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 ,
         \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 ,
         \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 ,
         \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 ,
         \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 ,
         \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 ,
         \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 ,
         \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 ,
         \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 ,
         \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 ,
         \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 ,
         \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 ,
         \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 ,
         \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 ,
         \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 ,
         \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 ,
         \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 ,
         \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 ,
         \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 ,
         \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 ,
         \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 ,
         \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 ,
         \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 ,
         \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 ,
         \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 ,
         \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 ,
         \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 ,
         \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 ,
         \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 ,
         \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 ,
         \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 ,
         \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 ,
         \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 ,
         \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 ,
         \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 ,
         \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 ,
         \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 ,
         \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 ,
         \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 ,
         \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 ,
         \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 ,
         \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 ,
         \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 ,
         \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 ,
         \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 ,
         \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 ,
         \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 ,
         \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 ,
         \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 ,
         \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 ,
         \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 ,
         \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 ,
         \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 ,
         \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 ,
         \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 ,
         \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 ,
         \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 ,
         \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 ,
         \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 ,
         \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 ,
         \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 ,
         \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 ,
         \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 ,
         \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 ,
         \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 ,
         \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 ,
         \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 ,
         \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 ,
         \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 ,
         \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 ,
         \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 ,
         \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 ,
         \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 ,
         \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 ,
         \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 ,
         \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 ,
         \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 ,
         \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 ,
         \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 ,
         \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 ,
         \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 ,
         \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 ,
         \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 ,
         \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 ,
         \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 ,
         \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 ,
         \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 ,
         \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 ,
         \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 ,
         \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 ,
         \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 ,
         \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 ,
         \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 ,
         \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 ,
         \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 ,
         \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 ,
         \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 ,
         \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 ,
         \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 ,
         \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 ,
         \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 ,
         \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 ,
         \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 ,
         \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 ,
         \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 ,
         \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 ,
         \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 ,
         \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 ,
         \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 ,
         \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 ,
         \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 ,
         \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 ,
         \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 ,
         \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 ,
         \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 ,
         \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 ,
         \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 ,
         \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 ,
         \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 ,
         \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 ,
         \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 ,
         \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 ,
         \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 ,
         \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 ,
         \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 ,
         \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 ,
         \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 ,
         \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 ,
         \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 ,
         \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 ,
         \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 ,
         \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 ,
         \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 ,
         \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 ,
         \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 ,
         \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 ,
         \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 ,
         \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 ,
         \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 ,
         \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 ,
         \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 ,
         \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 ,
         \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 ,
         \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 ,
         \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 ,
         \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 ,
         \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 ,
         \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 ,
         \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 ,
         \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 ,
         \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 ,
         \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 ,
         \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 ,
         \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 ,
         \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 ,
         \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 ,
         \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 ,
         \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 ,
         \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 ,
         \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 ,
         \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 ,
         \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 ,
         \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 ,
         \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 ,
         \20708 , \20709 , \20710 , \20711 , \20712 , \20713 ;
buf \U$labaj2145 ( R_289_8400778, \10196 );
buf \U$labaj2146 ( R_28a_8401e70, \10205 );
buf \U$labaj2147 ( R_28b_8401f18, \10255 );
buf \U$labaj2148 ( R_28c_8401fc0, \10315 );
buf \U$labaj2149 ( R_28d_8402068, \10333 );
buf \U$labaj2150 ( R_28e_8402110, \10347 );
buf \U$labaj2151 ( R_28f_84021b8, \10377 );
buf \U$labaj2152 ( R_290_8402260, \10386 );
buf \U$labaj2153 ( R_291_8402308, \10404 );
buf \U$labaj2154 ( R_292_84023b0, \10419 );
buf \U$labaj2155 ( R_293_8402458, \10456 );
buf \U$labaj2156 ( R_294_8402500, \10465 );
buf \U$labaj2157 ( R_295_84025a8, \10490 );
buf \U$labaj2158 ( R_296_8402650, \10500 );
buf \U$labaj2159 ( R_297_84026f8, \10529 );
buf \U$labaj2160 ( R_298_84027a0, \10543 );
buf \U$labaj2161 ( R_299_8402848, \10559 );
buf \U$labaj2162 ( R_29a_84028f0, \10578 );
buf \U$labaj2163 ( R_29b_8402998, \10612 );
buf \U$labaj2164 ( R_29c_8402a40, \10625 );
buf \U$labaj2165 ( R_29d_8402ae8, \10651 );
buf \U$labaj2166 ( R_29e_8402b90, \10665 );
buf \U$labaj2167 ( R_29f_8402c38, \10684 );
buf \U$labaj2168 ( R_2a0_8402ce0, \10695 );
buf \U$labaj2169 ( R_2a1_8402d88, \10704 );
buf \U$labaj2170 ( R_2a2_8402e30, \10719 );
buf \U$labaj2171 ( R_2a3_8402ed8, \10734 );
buf \U$labaj2172 ( R_267_8403418, \20170 );
buf \U$labaj2173 ( R_268_8400820, \20181 );
buf \U$labaj2174 ( R_269_84008c8, \20232 );
buf \U$labaj2175 ( R_26a_8400970, \20288 );
buf \U$labaj2176 ( R_26b_8400a18, \20307 );
buf \U$labaj2177 ( R_26c_8400ac0, \20325 );
buf \U$labaj2178 ( R_26d_8400b68, \20360 );
buf \U$labaj2179 ( R_26e_8400c10, \20369 );
buf \U$labaj2180 ( R_26f_8400cb8, \20387 );
buf \U$labaj2181 ( R_270_8400d60, \20398 );
buf \U$labaj2182 ( R_271_8400e08, \20441 );
buf \U$labaj2183 ( R_272_8400eb0, \20450 );
buf \U$labaj2184 ( R_273_8400f58, \20476 );
buf \U$labaj2185 ( R_274_8401000, \20486 );
buf \U$labaj2186 ( R_275_84010a8, \20515 );
buf \U$labaj2187 ( R_276_8401150, \20524 );
buf \U$labaj2188 ( R_277_84011f8, \20539 );
buf \U$labaj2189 ( R_278_84012a0, \20558 );
buf \U$labaj2190 ( R_279_8401348, \20592 );
buf \U$labaj2191 ( R_27a_84013f0, \20605 );
buf \U$labaj2192 ( R_27b_8401498, \20630 );
buf \U$labaj2193 ( R_27c_8401540, \20644 );
buf \U$labaj2194 ( R_27d_84015e8, \20664 );
buf \U$labaj2195 ( R_27e_8401690, \20674 );
buf \U$labaj2196 ( R_27f_8401738, \20683 );
buf \U$labaj2197 ( R_280_84017e0, \20699 );
buf \U$labaj2198 ( R_281_8401888, \20713 );
not \U$1 ( \693 , RI994e028_23);
nand \U$2 ( \694 , RI994dfb0_24, RI994df38_25);
nor \U$3 ( \695 , \693 , \694 );
nand \U$4 ( \696 , \695 , RI994e0a0_22);
not \U$5 ( \697 , RI994e118_21);
nor \U$6 ( \698 , \696 , \697 );
nand \U$7 ( \699 , \698 , RI994e190_20);
not \U$8 ( \700 , \699 );
nand \U$9 ( \701 , \700 , RI994e208_19);
nand \U$10 ( \702 , RI994e3e8_15, RI994e370_16, RI994e2f8_17, RI994e280_18);
nor \U$11 ( \703 , \701 , \702 );
xor \U$12 ( \704 , RI994e460_14, \703 );
nor \U$13 ( \705 , RI9921898_610, RI9921820_611);
nor \U$14 ( \706 , RI99217a8_612, RI9921910_609, RI9921730_613);
and \U$15 ( \707 , \705 , \706 );
buf \U$16 ( \708 , \707 );
and \U$17 ( \709 , \708 , RI994de48_27);
not \U$18 ( \710 , RI99217a8_612);
nand \U$19 ( \711 , \710 , \705 , RI9921730_613);
not \U$20 ( \712 , \711 );
not \U$21 ( \713 , \712 );
not \U$22 ( \714 , RI98bc948_40);
or \U$23 ( \715 , \713 , \714 );
nand \U$24 ( \716 , RI995e4c8_235, RI9921910_609);
nand \U$25 ( \717 , \715 , \716 );
nor \U$26 ( \718 , \709 , \717 );
not \U$27 ( \719 , RI99217a8_612);
nor \U$28 ( \720 , \719 , RI9921730_613);
and \U$29 ( \721 , \705 , \720 );
buf \U$30 ( \722 , \721 );
and \U$31 ( \723 , \722 , RI98abcb0_53);
nand \U$32 ( \724 , RI99217a8_612, RI9921730_613);
not \U$33 ( \725 , \724 );
nand \U$34 ( \726 , \725 , \705 );
not \U$35 ( \727 , \726 );
and \U$36 ( \728 , \727 , RI98197a8_66);
nor \U$37 ( \729 , \723 , \728 );
nand \U$38 ( \730 , RI9921820_611, RI99217a8_612);
not \U$39 ( \731 , \730 );
not \U$40 ( \732 , RI9921898_610);
nor \U$41 ( \733 , \732 , RI9921730_613);
nand \U$42 ( \734 , \731 , \733 );
not \U$43 ( \735 , \734 );
and \U$44 ( \736 , \735 , RI890f600_209);
nand \U$45 ( \737 , RI9921898_610, RI9921730_613);
nor \U$46 ( \738 , \730 , \737 );
buf \U$47 ( \739 , \738 );
and \U$48 ( \740 , \739 , RI99670f0_222);
nor \U$49 ( \741 , \736 , \740 );
nor \U$50 ( \742 , RI9921820_611, RI99217a8_612);
and \U$51 ( \743 , \733 , \742 );
buf \U$52 ( \744 , \743 );
and \U$53 ( \745 , \744 , RI89ec0a0_131);
not \U$54 ( \746 , \742 );
nor \U$55 ( \747 , \746 , \737 );
buf \U$56 ( \748 , \747 );
and \U$57 ( \749 , \748 , RI8946038_144);
nor \U$58 ( \750 , \745 , \749 );
nand \U$59 ( \751 , \718 , \729 , \741 , \750 );
not \U$60 ( \752 , RI9921820_611);
nor \U$61 ( \753 , \752 , RI99217a8_612);
and \U$62 ( \754 , \753 , \733 );
buf \U$63 ( \755 , \754 );
and \U$64 ( \756 , \755 , RI8924e10_183);
not \U$65 ( \757 , RI9921730_613);
not \U$66 ( \758 , RI9921898_610);
nor \U$67 ( \759 , \757 , \758 );
nand \U$68 ( \760 , \759 , \753 );
not \U$69 ( \761 , \760 );
and \U$70 ( \762 , \761 , RI89185e8_196);
nor \U$71 ( \763 , \756 , \762 );
not \U$72 ( \764 , RI9921820_611);
nand \U$73 ( \765 , \764 , RI99217a8_612);
not \U$74 ( \766 , \765 );
nand \U$75 ( \767 , \766 , \733 );
not \U$76 ( \768 , \767 );
buf \U$77 ( \769 , \768 );
and \U$78 ( \770 , \769 , RI8939810_157);
not \U$79 ( \771 , RI99217a8_612);
nor \U$80 ( \772 , \771 , \737 , RI9921820_611);
buf \U$81 ( \773 , \772 );
and \U$82 ( \774 , \773 , RI8930828_170);
nor \U$83 ( \775 , \770 , \774 );
nor \U$84 ( \776 , RI9921898_610, RI9921730_613);
not \U$85 ( \777 , \776 );
nor \U$86 ( \778 , \777 , \730 );
buf \U$87 ( \779 , \778 );
and \U$88 ( \780 , \779 , RI9776ff8_105);
not \U$89 ( \781 , RI9921730_613);
nor \U$90 ( \782 , \781 , RI9921898_610);
and \U$91 ( \783 , \753 , \782 );
buf \U$92 ( \784 , \783 );
and \U$93 ( \785 , \784 , RI98084f8_92);
nor \U$94 ( \786 , \780 , \785 );
and \U$95 ( \787 , \753 , \776 );
buf \U$96 ( \788 , \787 );
and \U$97 ( \789 , \788 , RI9808b10_79);
not \U$98 ( \790 , \782 );
nor \U$99 ( \791 , \790 , \730 );
buf \U$100 ( \792 , \791 );
and \U$101 ( \793 , \792 , RI89ec6b8_118);
nor \U$102 ( \794 , \789 , \793 );
nand \U$103 ( \795 , \763 , \775 , \786 , \794 );
nor \U$104 ( \796 , \751 , \795 );
or \U$105 ( \797 , \704 , \796 );
not \U$106 ( \798 , \797 );
not \U$107 ( \799 , \713 );
nand \U$108 ( \800 , \799 , RI98bc8d0_41);
nand \U$109 ( \801 , \708 , RI994ddd0_28);
nand \U$110 ( \802 , RI995e450_236, RI9921910_609);
and \U$111 ( \803 , \800 , \801 , \802 );
and \U$112 ( \804 , \735 , RI9967690_210);
and \U$113 ( \805 , \739 , RI9967078_223);
nor \U$114 ( \806 , \804 , \805 );
and \U$115 ( \807 , \722 , RI98abc38_54);
and \U$116 ( \808 , \727 , RI9819730_67);
nor \U$117 ( \809 , \807 , \808 );
and \U$118 ( \810 , \744 , RI89465d8_132);
and \U$119 ( \811 , \748 , RI8939db0_145);
nor \U$120 ( \812 , \810 , \811 );
nand \U$121 ( \813 , \803 , \806 , \809 , \812 );
not \U$122 ( \814 , \760 );
not \U$123 ( \815 , RI890fba0_197);
not \U$124 ( \816 , \815 );
and \U$125 ( \817 , \814 , \816 );
and \U$126 ( \818 , \788 , RI9808a98_80);
nor \U$127 ( \819 , \817 , \818 );
and \U$128 ( \820 , \769 , RI8930dc8_158);
and \U$129 ( \821 , \773 , RI89253b0_171);
nor \U$130 ( \822 , \820 , \821 );
and \U$131 ( \823 , \755 , RI8918b88_184);
and \U$132 ( \824 , \792 , RI89ec640_119);
nor \U$133 ( \825 , \823 , \824 );
not \U$134 ( \826 , \730 );
nand \U$135 ( \827 , \826 , \776 );
not \U$136 ( \828 , \827 );
not \U$137 ( \829 , RI9776f80_106);
not \U$138 ( \830 , \829 );
and \U$139 ( \831 , \828 , \830 );
and \U$140 ( \832 , \784 , RI9808480_93);
nor \U$141 ( \833 , \831 , \832 );
nand \U$142 ( \834 , \819 , \822 , \825 , \833 );
nor \U$143 ( \835 , \813 , \834 );
not \U$144 ( \836 , \835 );
not \U$145 ( \837 , RI994e280_18);
nor \U$146 ( \838 , \837 , \701 );
nand \U$147 ( \839 , \838 , RI994e2f8_17);
not \U$148 ( \840 , \839 );
nand \U$149 ( \841 , \840 , RI994e370_16);
xor \U$150 ( \842 , \841 , RI994e3e8_15);
nand \U$151 ( \843 , \836 , \842 );
not \U$152 ( \844 , \843 );
xor \U$153 ( \845 , \701 , RI994e280_18);
nand \U$154 ( \846 , \799 , RI98bc768_44);
nand \U$155 ( \847 , \708 , RI994dc68_31);
nand \U$156 ( \848 , RI9959f68_239, RI9921910_609);
nand \U$157 ( \849 , \846 , \847 , \848 );
not \U$158 ( \850 , RI9967528_213);
not \U$159 ( \851 , \735 );
or \U$160 ( \852 , \850 , \851 );
nand \U$161 ( \853 , \739 , RI995e900_226);
nand \U$162 ( \854 , \852 , \853 );
nor \U$163 ( \855 , \849 , \854 );
not \U$164 ( \856 , RI890fa38_200);
not \U$165 ( \857 , \761 );
or \U$166 ( \858 , \856 , \857 );
nand \U$167 ( \859 , \788 , RI9808930_83);
nand \U$168 ( \860 , \858 , \859 );
not \U$169 ( \861 , RI8930c60_161);
not \U$170 ( \862 , \769 );
or \U$171 ( \863 , \861 , \862 );
nand \U$172 ( \864 , \773 , RI8925248_174);
nand \U$173 ( \865 , \863 , \864 );
nor \U$174 ( \866 , \860 , \865 );
not \U$175 ( \867 , RI98195c8_70);
not \U$176 ( \868 , \727 );
or \U$177 ( \869 , \867 , \868 );
nand \U$178 ( \870 , \722 , RI98abad0_57);
nand \U$179 ( \871 , \869 , \870 );
not \U$180 ( \872 , RI8946470_135);
not \U$181 ( \873 , \744 );
or \U$182 ( \874 , \872 , \873 );
nand \U$183 ( \875 , \748 , RI8939c48_148);
nand \U$184 ( \876 , \874 , \875 );
nor \U$185 ( \877 , \871 , \876 );
not \U$186 ( \878 , RI8918a20_187);
not \U$187 ( \879 , \755 );
or \U$188 ( \880 , \878 , \879 );
nand \U$189 ( \881 , \792 , RI89ec4d8_122);
nand \U$190 ( \882 , \880 , \881 );
not \U$191 ( \883 , RI9808318_96);
not \U$192 ( \884 , \784 );
or \U$193 ( \885 , \883 , \884 );
nand \U$194 ( \886 , \779 , RI9776e18_109);
nand \U$195 ( \887 , \885 , \886 );
nor \U$196 ( \888 , \882 , \887 );
nand \U$197 ( \889 , \855 , \866 , \877 , \888 );
nand \U$198 ( \890 , \845 , \889 );
and \U$199 ( \891 , RI98082a0_97, \784 );
and \U$200 ( \892 , \779 , RI9776da0_110);
not \U$201 ( \893 , RI8930be8_162);
not \U$202 ( \894 , \769 );
or \U$203 ( \895 , \893 , \894 );
nand \U$204 ( \896 , \773 , RI89251d0_175);
nand \U$205 ( \897 , \895 , \896 );
nor \U$206 ( \898 , \891 , \892 , \897 );
nand \U$207 ( \899 , \799 , RI98bc6f0_45);
nand \U$208 ( \900 , \708 , RI994dbf0_32);
nand \U$209 ( \901 , RI9959860_240, RI9921910_609);
nand \U$210 ( \902 , \899 , \900 , \901 );
not \U$211 ( \903 , RI99674b0_214);
not \U$212 ( \904 , \735 );
or \U$213 ( \905 , \903 , \904 );
nand \U$214 ( \906 , \739 , RI995e888_227);
nand \U$215 ( \907 , \905 , \906 );
nor \U$216 ( \908 , \902 , \907 );
not \U$217 ( \909 , RI9819550_71);
not \U$218 ( \910 , \727 );
or \U$219 ( \911 , \909 , \910 );
nand \U$220 ( \912 , \722 , RI98aba58_58);
nand \U$221 ( \913 , \911 , \912 );
not \U$222 ( \914 , RI89463f8_136);
not \U$223 ( \915 , \744 );
or \U$224 ( \916 , \914 , \915 );
nand \U$225 ( \917 , \748 , RI8939bd0_149);
nand \U$226 ( \918 , \916 , \917 );
nor \U$227 ( \919 , \913 , \918 );
not \U$228 ( \920 , RI890f9c0_201);
not \U$229 ( \921 , \761 );
or \U$230 ( \922 , \920 , \921 );
nand \U$231 ( \923 , \755 , RI89189a8_188);
nand \U$232 ( \924 , \922 , \923 );
not \U$233 ( \925 , RI98088b8_84);
not \U$234 ( \926 , \788 );
or \U$235 ( \927 , \925 , \926 );
nand \U$236 ( \928 , \792 , RI89ec460_123);
nand \U$237 ( \929 , \927 , \928 );
nor \U$238 ( \930 , \924 , \929 );
nand \U$239 ( \931 , \898 , \908 , \919 , \930 );
and \U$240 ( \932 , \699 , RI994e208_19);
not \U$241 ( \933 , \699 );
not \U$242 ( \934 , RI994e208_19);
and \U$243 ( \935 , \933 , \934 );
nor \U$244 ( \936 , \932 , \935 );
nand \U$245 ( \937 , \931 , \936 );
nand \U$246 ( \938 , \890 , \937 );
and \U$247 ( \939 , \799 , RI98abff8_46);
nand \U$248 ( \940 , RI994d998_241, RI9921910_609);
not \U$249 ( \941 , \940 );
nor \U$250 ( \942 , \939 , \941 );
nand \U$251 ( \943 , \735 , RI9967438_215);
nand \U$252 ( \944 , \708 , RI98bcc90_33);
nand \U$253 ( \945 , \739 , RI995e810_228);
nand \U$254 ( \946 , \942 , \943 , \944 , \945 );
nand \U$255 ( \947 , \744 , RI8946380_137);
nand \U$256 ( \948 , \727 , RI98194d8_72);
nand \U$257 ( \949 , \722 , RI98ab9e0_59);
nand \U$258 ( \950 , \748 , RI8939b58_150);
nand \U$259 ( \951 , \947 , \948 , \949 , \950 );
nor \U$260 ( \952 , \946 , \951 );
nand \U$261 ( \953 , \788 , RI9808840_85);
nand \U$262 ( \954 , \761 , RI890f948_202);
nand \U$263 ( \955 , \784 , RI9808228_98);
nand \U$264 ( \956 , \779 , RI9776d28_111);
nand \U$265 ( \957 , \953 , \954 , \955 , \956 );
nand \U$266 ( \958 , \755 , RI8918930_189);
nand \U$267 ( \959 , \769 , RI8930b70_163);
nand \U$268 ( \960 , \773 , RI8925158_176);
nand \U$269 ( \961 , \792 , RI89ec3e8_124);
nand \U$270 ( \962 , \958 , \959 , \960 , \961 );
nor \U$271 ( \963 , \957 , \962 );
nand \U$272 ( \964 , \952 , \963 );
xnor \U$273 ( \965 , \698 , RI994e190_20);
nand \U$274 ( \966 , \964 , \965 );
nand \U$275 ( \967 , \799 , RI98abf80_47);
nand \U$276 ( \968 , \708 , RI98bcc18_34);
nand \U$277 ( \969 , RI994d920_242, RI9921910_609);
nand \U$278 ( \970 , \967 , \968 , \969 );
not \U$279 ( \971 , RI99673c0_216);
not \U$280 ( \972 , \735 );
or \U$281 ( \973 , \971 , \972 );
nand \U$282 ( \974 , \739 , RI995e798_229);
nand \U$283 ( \975 , \973 , \974 );
nor \U$284 ( \976 , \970 , \975 );
not \U$285 ( \977 , RI98087c8_86);
not \U$286 ( \978 , \788 );
or \U$287 ( \979 , \977 , \978 );
nand \U$288 ( \980 , \761 , RI890f8d0_203);
nand \U$289 ( \981 , \979 , \980 );
not \U$290 ( \982 , RI97772c8_99);
not \U$291 ( \983 , \784 );
or \U$292 ( \984 , \982 , \983 );
nand \U$293 ( \985 , \779 , RI89ec988_112);
nand \U$294 ( \986 , \984 , \985 );
nor \U$295 ( \987 , \981 , \986 );
not \U$296 ( \988 , RI89188b8_190);
not \U$297 ( \989 , \755 );
or \U$298 ( \990 , \988 , \989 );
nand \U$299 ( \991 , \773 , RI89250e0_177);
nand \U$300 ( \992 , \990 , \991 );
not \U$301 ( \993 , RI8930af8_164);
not \U$302 ( \994 , \769 );
or \U$303 ( \995 , \993 , \994 );
nand \U$304 ( \996 , \792 , RI89ec370_125);
nand \U$305 ( \997 , \995 , \996 );
nor \U$306 ( \998 , \992 , \997 );
not \U$307 ( \999 , RI98ab968_60);
not \U$308 ( \1000 , \722 );
or \U$309 ( \1001 , \999 , \1000 );
nand \U$310 ( \1002 , \727 , RI9819460_73);
nand \U$311 ( \1003 , \1001 , \1002 );
not \U$312 ( \1004 , RI8946308_138);
not \U$313 ( \1005 , \744 );
or \U$314 ( \1006 , \1004 , \1005 );
nand \U$315 ( \1007 , \748 , RI8939ae0_151);
nand \U$316 ( \1008 , \1006 , \1007 );
nor \U$317 ( \1009 , \1003 , \1008 );
nand \U$318 ( \1010 , \976 , \987 , \998 , \1009 );
and \U$319 ( \1011 , \696 , \697 );
not \U$320 ( \1012 , \696 );
and \U$321 ( \1013 , \1012 , RI994e118_21);
or \U$322 ( \1014 , \1011 , \1013 );
nand \U$323 ( \1015 , \1010 , \1014 );
nand \U$324 ( \1016 , \966 , \1015 );
nor \U$325 ( \1017 , \938 , \1016 );
not \U$326 ( \1018 , \1017 );
xnor \U$327 ( \1019 , \694 , RI994e028_23);
nand \U$328 ( \1020 , \799 , RI98abe90_49);
nand \U$329 ( \1021 , \708 , RI98bcb28_36);
nand \U$330 ( \1022 , RI994d830_244, RI9921910_609);
nand \U$331 ( \1023 , \1020 , \1021 , \1022 );
not \U$332 ( \1024 , RI99672d0_218);
not \U$333 ( \1025 , \735 );
or \U$334 ( \1026 , \1024 , \1025 );
nand \U$335 ( \1027 , \739 , RI995e6a8_231);
nand \U$336 ( \1028 , \1026 , \1027 );
nor \U$337 ( \1029 , \1023 , \1028 );
not \U$338 ( \1030 , RI98086d8_88);
not \U$339 ( \1031 , \788 );
or \U$340 ( \1032 , \1030 , \1031 );
nand \U$341 ( \1033 , \761 , RI890f7e0_205);
nand \U$342 ( \1034 , \1032 , \1033 );
not \U$343 ( \1035 , RI97771d8_101);
not \U$344 ( \1036 , \784 );
or \U$345 ( \1037 , \1035 , \1036 );
nand \U$346 ( \1038 , \779 , RI89ec898_114);
nand \U$347 ( \1039 , \1037 , \1038 );
nor \U$348 ( \1040 , \1034 , \1039 );
not \U$349 ( \1041 , RI89187c8_192);
not \U$350 ( \1042 , \755 );
or \U$351 ( \1043 , \1041 , \1042 );
nand \U$352 ( \1044 , \773 , RI8924ff0_179);
nand \U$353 ( \1045 , \1043 , \1044 );
not \U$354 ( \1046 , RI8930a08_166);
not \U$355 ( \1047 , \769 );
or \U$356 ( \1048 , \1046 , \1047 );
nand \U$357 ( \1049 , \792 , RI89ec280_127);
nand \U$358 ( \1050 , \1048 , \1049 );
nor \U$359 ( \1051 , \1045 , \1050 );
not \U$360 ( \1052 , RI8946218_140);
not \U$361 ( \1053 , \744 );
or \U$362 ( \1054 , \1052 , \1053 );
nand \U$363 ( \1055 , \748 , RI89399f0_153);
nand \U$364 ( \1056 , \1054 , \1055 );
not \U$365 ( \1057 , RI9819370_75);
not \U$366 ( \1058 , \727 );
or \U$367 ( \1059 , \1057 , \1058 );
nand \U$368 ( \1060 , \722 , RI98ab878_62);
nand \U$369 ( \1061 , \1059 , \1060 );
nor \U$370 ( \1062 , \1056 , \1061 );
nand \U$371 ( \1063 , \1029 , \1040 , \1051 , \1062 );
not \U$372 ( \1064 , \1063 );
xor \U$373 ( \1065 , \1019 , \1064 );
not \U$374 ( \1066 , RI890f768_206);
not \U$375 ( \1067 , \761 );
or \U$376 ( \1068 , \1066 , \1067 );
nand \U$377 ( \1069 , \788 , RI9808660_89);
nand \U$378 ( \1070 , \1068 , \1069 );
not \U$379 ( \1071 , RI9777160_102);
not \U$380 ( \1072 , \784 );
or \U$381 ( \1073 , \1071 , \1072 );
nand \U$382 ( \1074 , \778 , RI89ec820_115);
nand \U$383 ( \1075 , \1073 , \1074 );
nor \U$384 ( \1076 , \1070 , \1075 );
nand \U$385 ( \1077 , \712 , RI98abe18_50);
nand \U$386 ( \1078 , \707 , RI98bcab0_37);
nand \U$387 ( \1079 , RI994d7b8_245, RI9921910_609);
nand \U$388 ( \1080 , \1077 , \1078 , \1079 );
not \U$389 ( \1081 , RI9967258_219);
not \U$390 ( \1082 , \735 );
or \U$391 ( \1083 , \1081 , \1082 );
nand \U$392 ( \1084 , \738 , RI995e630_232);
nand \U$393 ( \1085 , \1083 , \1084 );
nor \U$394 ( \1086 , \1080 , \1085 );
not \U$395 ( \1087 , RI8918750_193);
not \U$396 ( \1088 , \755 );
or \U$397 ( \1089 , \1087 , \1088 );
nand \U$398 ( \1090 , \773 , RI8924f78_180);
nand \U$399 ( \1091 , \1089 , \1090 );
not \U$400 ( \1092 , RI8930990_167);
not \U$401 ( \1093 , \769 );
or \U$402 ( \1094 , \1092 , \1093 );
nand \U$403 ( \1095 , \792 , RI89ec208_128);
nand \U$404 ( \1096 , \1094 , \1095 );
nor \U$405 ( \1097 , \1091 , \1096 );
not \U$406 ( \1098 , RI98192f8_76);
not \U$407 ( \1099 , \727 );
or \U$408 ( \1100 , \1098 , \1099 );
nand \U$409 ( \1101 , \722 , RI98ab800_63);
nand \U$410 ( \1102 , \1100 , \1101 );
not \U$411 ( \1103 , RI89461a0_141);
not \U$412 ( \1104 , \743 );
or \U$413 ( \1105 , \1103 , \1104 );
nand \U$414 ( \1106 , \747 , RI8939978_154);
nand \U$415 ( \1107 , \1105 , \1106 );
nor \U$416 ( \1108 , \1102 , \1107 );
nand \U$417 ( \1109 , \1076 , \1086 , \1097 , \1108 );
and \U$418 ( \1110 , RI994dfb0_24, RI994df38_25);
not \U$419 ( \1111 , RI994dfb0_24);
not \U$420 ( \1112 , RI994df38_25);
and \U$421 ( \1113 , \1111 , \1112 );
nor \U$422 ( \1114 , \1110 , \1113 );
not \U$423 ( \1115 , \1114 );
nand \U$424 ( \1116 , \1109 , \1115 );
not \U$425 ( \1117 , \1116 );
not \U$426 ( \1118 , RI89186d8_194);
not \U$427 ( \1119 , \754 );
or \U$428 ( \1120 , \1118 , \1119 );
nand \U$429 ( \1121 , \791 , RI89ec190_129);
nand \U$430 ( \1122 , \1120 , \1121 );
not \U$431 ( \1123 , RI98ab788_64);
not \U$432 ( \1124 , \721 );
or \U$433 ( \1125 , \1123 , \1124 );
not \U$434 ( \1126 , \726 );
nand \U$435 ( \1127 , \1126 , RI9819280_77);
nand \U$436 ( \1128 , \1125 , \1127 );
nor \U$437 ( \1129 , \1122 , \1128 );
not \U$438 ( \1130 , RI98abda0_51);
nor \U$439 ( \1131 , \1130 , \711 );
not \U$440 ( \1132 , \1131 );
nand \U$441 ( \1133 , \707 , RI98bca38_38);
nand \U$442 ( \1134 , RI994d740_246, RI9921910_609);
nand \U$443 ( \1135 , \1132 , \1133 , \1134 );
nor \U$444 ( \1136 , \737 , \730 );
not \U$445 ( \1137 , \1136 );
not \U$446 ( \1138 , RI995e5b8_233);
or \U$447 ( \1139 , \1137 , \1138 );
not \U$448 ( \1140 , RI99671e0_220);
or \U$449 ( \1141 , \734 , \1140 );
nand \U$450 ( \1142 , \1139 , \1141 );
nor \U$451 ( \1143 , \1135 , \1142 );
not \U$452 ( \1144 , RI97770e8_103);
not \U$453 ( \1145 , \783 );
or \U$454 ( \1146 , \1144 , \1145 );
nand \U$455 ( \1147 , \787 , RI98085e8_90);
nand \U$456 ( \1148 , \1146 , \1147 );
not \U$457 ( \1149 , RI8930918_168);
not \U$458 ( \1150 , \768 );
or \U$459 ( \1151 , \1149 , \1150 );
nand \U$460 ( \1152 , \772 , RI8924f00_181);
nand \U$461 ( \1153 , \1151 , \1152 );
nor \U$462 ( \1154 , \1148 , \1153 );
not \U$463 ( \1155 , RI8946128_142);
not \U$464 ( \1156 , \743 );
or \U$465 ( \1157 , \1155 , \1156 );
nand \U$466 ( \1158 , \747 , RI8939900_155);
nand \U$467 ( \1159 , \1157 , \1158 );
not \U$468 ( \1160 , \778 );
not \U$469 ( \1161 , RI89ec7a8_116);
or \U$470 ( \1162 , \1160 , \1161 );
not \U$471 ( \1163 , \760 );
nand \U$472 ( \1164 , \1163 , RI890f6f0_207);
nand \U$473 ( \1165 , \1162 , \1164 );
nor \U$474 ( \1166 , \1159 , \1165 );
nand \U$475 ( \1167 , \1129 , \1143 , \1154 , \1166 );
nand \U$476 ( \1168 , \1167 , RI994df38_25);
not \U$477 ( \1169 , \1168 );
nand \U$478 ( \1170 , \735 , RI9967168_221);
and \U$479 ( \1171 , \712 , RI98abd28_52);
nand \U$480 ( \1172 , RI994d6c8_247, RI9921910_609);
not \U$481 ( \1173 , \1172 );
nor \U$482 ( \1174 , \1171 , \1173 );
nand \U$483 ( \1175 , \707 , RI98bc9c0_39);
nand \U$484 ( \1176 , \738 , RI995e540_234);
nand \U$485 ( \1177 , \1170 , \1174 , \1175 , \1176 );
and \U$486 ( \1178 , RI890f678_208, \761 );
not \U$487 ( \1179 , RI89ec730_117);
nor \U$488 ( \1180 , \1179 , \827 );
nor \U$489 ( \1181 , \1178 , \1180 );
and \U$490 ( \1182 , \727 , RI9819208_78);
and \U$491 ( \1183 , \768 , RI89308a0_169);
nor \U$492 ( \1184 , \1182 , \1183 );
nand \U$493 ( \1185 , \1181 , \1184 );
nor \U$494 ( \1186 , \1177 , \1185 );
nand \U$495 ( \1187 , \743 , RI89460b0_143);
nand \U$496 ( \1188 , \721 , RI98ab710_65);
nand \U$497 ( \1189 , \747 , RI8939888_156);
nand \U$498 ( \1190 , \772 , RI8924e88_182);
nand \U$499 ( \1191 , \1187 , \1188 , \1189 , \1190 );
not \U$500 ( \1192 , RI9777070_104);
not \U$501 ( \1193 , \783 );
or \U$502 ( \1194 , \1192 , \1193 );
nand \U$503 ( \1195 , \787 , RI9808570_91);
nand \U$504 ( \1196 , \1194 , \1195 );
not \U$505 ( \1197 , RI8918660_195);
not \U$506 ( \1198 , \754 );
or \U$507 ( \1199 , \1197 , \1198 );
nand \U$508 ( \1200 , \791 , RI89ec118_130);
nand \U$509 ( \1201 , \1199 , \1200 );
nor \U$510 ( \1202 , \1191 , \1196 , \1201 );
nand \U$511 ( \1203 , \1186 , \1202 );
not \U$512 ( \1204 , RI994dec0_26);
nand \U$513 ( \1205 , \1203 , \1204 );
not \U$514 ( \1206 , \1205 );
or \U$515 ( \1207 , \1169 , \1206 );
not \U$516 ( \1208 , \1167 );
nand \U$517 ( \1209 , \1208 , \1112 );
nand \U$518 ( \1210 , \1207 , \1209 );
not \U$519 ( \1211 , \1210 );
or \U$520 ( \1212 , \1117 , \1211 );
not \U$521 ( \1213 , \1109 );
nand \U$522 ( \1214 , \1213 , \1114 );
nand \U$523 ( \1215 , \1212 , \1214 );
and \U$524 ( \1216 , \1065 , \1215 );
and \U$525 ( \1217 , \1019 , \1064 );
or \U$526 ( \1218 , \1216 , \1217 );
not \U$527 ( \1219 , \1218 );
nand \U$528 ( \1220 , RI994d8a8_243, RI9921910_609);
not \U$529 ( \1221 , \1220 );
not \U$530 ( \1222 , RI9967348_217);
not \U$531 ( \1223 , \735 );
or \U$532 ( \1224 , \1222 , \1223 );
nand \U$533 ( \1225 , \739 , RI995e720_230);
nand \U$534 ( \1226 , \1224 , \1225 );
not \U$535 ( \1227 , \799 );
not \U$536 ( \1228 , RI98abf08_48);
or \U$537 ( \1229 , \1227 , \1228 );
nand \U$538 ( \1230 , \708 , RI98bcba0_35);
nand \U$539 ( \1231 , \1229 , \1230 );
nor \U$540 ( \1232 , \1221 , \1226 , \1231 );
not \U$541 ( \1233 , RI890f858_204);
not \U$542 ( \1234 , \761 );
or \U$543 ( \1235 , \1233 , \1234 );
nand \U$544 ( \1236 , \788 , RI9808750_87);
nand \U$545 ( \1237 , \1235 , \1236 );
not \U$546 ( \1238 , RI9777250_100);
not \U$547 ( \1239 , \784 );
or \U$548 ( \1240 , \1238 , \1239 );
nand \U$549 ( \1241 , \779 , RI89ec910_113);
nand \U$550 ( \1242 , \1240 , \1241 );
nor \U$551 ( \1243 , \1237 , \1242 );
not \U$552 ( \1244 , RI8918840_191);
not \U$553 ( \1245 , \755 );
or \U$554 ( \1246 , \1244 , \1245 );
nand \U$555 ( \1247 , \773 , RI8925068_178);
nand \U$556 ( \1248 , \1246 , \1247 );
not \U$557 ( \1249 , RI8930a80_165);
not \U$558 ( \1250 , \769 );
or \U$559 ( \1251 , \1249 , \1250 );
nand \U$560 ( \1252 , \792 , RI89ec2f8_126);
nand \U$561 ( \1253 , \1251 , \1252 );
nor \U$562 ( \1254 , \1248 , \1253 );
not \U$563 ( \1255 , RI98193e8_74);
not \U$564 ( \1256 , \727 );
or \U$565 ( \1257 , \1255 , \1256 );
nand \U$566 ( \1258 , \722 , RI98ab8f0_61);
nand \U$567 ( \1259 , \1257 , \1258 );
not \U$568 ( \1260 , RI8946290_139);
not \U$569 ( \1261 , \744 );
or \U$570 ( \1262 , \1260 , \1261 );
nand \U$571 ( \1263 , \748 , RI8939a68_152);
nand \U$572 ( \1264 , \1262 , \1263 );
nor \U$573 ( \1265 , \1259 , \1264 );
nand \U$574 ( \1266 , \1232 , \1243 , \1254 , \1265 );
not \U$575 ( \1267 , RI994e0a0_22);
and \U$576 ( \1268 , \695 , \1267 );
not \U$577 ( \1269 , \695 );
and \U$578 ( \1270 , \1269 , RI994e0a0_22);
nor \U$579 ( \1271 , \1268 , \1270 );
nand \U$580 ( \1272 , \1266 , \1271 );
not \U$581 ( \1273 , \1272 );
nor \U$582 ( \1274 , \1219 , \1273 );
not \U$583 ( \1275 , \1274 );
or \U$584 ( \1276 , \1018 , \1275 );
not \U$585 ( \1277 , \1010 );
not \U$586 ( \1278 , \1014 );
nand \U$587 ( \1279 , \1277 , \1278 );
nor \U$588 ( \1280 , \1266 , \1271 );
nand \U$589 ( \1281 , \1280 , \1015 );
nand \U$590 ( \1282 , \1279 , \1281 );
and \U$591 ( \1283 , \1282 , \966 );
nor \U$592 ( \1284 , \964 , \965 );
nor \U$593 ( \1285 , \1283 , \1284 );
nor \U$594 ( \1286 , \1285 , \938 );
not \U$595 ( \1287 , \890 );
or \U$596 ( \1288 , \931 , \936 );
or \U$597 ( \1289 , \1287 , \1288 );
not \U$598 ( \1290 , \845 );
not \U$599 ( \1291 , \889 );
nand \U$600 ( \1292 , \1290 , \1291 );
nand \U$601 ( \1293 , \1289 , \1292 );
nor \U$602 ( \1294 , \1286 , \1293 );
nand \U$603 ( \1295 , \1276 , \1294 );
xnor \U$604 ( \1296 , \838 , RI994e2f8_17);
and \U$605 ( \1297 , \755 , RI8918a98_186);
and \U$606 ( \1298 , \761 , RI890fab0_199);
nor \U$607 ( \1299 , \1297 , \1298 );
and \U$608 ( \1300 , \788 , RI98089a8_82);
and \U$609 ( \1301 , \792 , RI89ec550_121);
nor \U$610 ( \1302 , \1300 , \1301 );
and \U$611 ( \1303 , \769 , RI8930cd8_160);
and \U$612 ( \1304 , \773 , RI89252c0_173);
nor \U$613 ( \1305 , \1303 , \1304 );
and \U$614 ( \1306 , \779 , RI9776e90_108);
and \U$615 ( \1307 , \784 , RI9808390_95);
nor \U$616 ( \1308 , \1306 , \1307 );
nand \U$617 ( \1309 , \1299 , \1302 , \1305 , \1308 );
nand \U$618 ( \1310 , \799 , RI98bc7e0_43);
nand \U$619 ( \1311 , \708 , RI994dce0_30);
nand \U$620 ( \1312 , RI9959fe0_238, RI9921910_609);
and \U$621 ( \1313 , \1310 , \1311 , \1312 );
and \U$622 ( \1314 , \722 , RI98abb48_56);
and \U$623 ( \1315 , \727 , RI9819640_69);
nor \U$624 ( \1316 , \1314 , \1315 );
and \U$625 ( \1317 , \744 , RI89464e8_134);
and \U$626 ( \1318 , \748 , RI8939cc0_147);
nor \U$627 ( \1319 , \1317 , \1318 );
and \U$628 ( \1320 , \735 , RI99675a0_212);
and \U$629 ( \1321 , \739 , RI995e978_225);
nor \U$630 ( \1322 , \1320 , \1321 );
nand \U$631 ( \1323 , \1313 , \1316 , \1319 , \1322 );
or \U$632 ( \1324 , \1309 , \1323 );
nand \U$633 ( \1325 , \1296 , \1324 );
and \U$634 ( \1326 , \1295 , \1325 );
nor \U$635 ( \1327 , \1296 , \1324 );
nor \U$636 ( \1328 , \1326 , \1327 );
not \U$637 ( \1329 , RI994e370_16);
not \U$638 ( \1330 , \1329 );
not \U$639 ( \1331 , \840 );
or \U$640 ( \1332 , \1330 , \1331 );
nand \U$641 ( \1333 , \839 , RI994e370_16);
nand \U$642 ( \1334 , \1332 , \1333 );
nand \U$643 ( \1335 , \799 , RI98bc858_42);
nand \U$644 ( \1336 , \708 , RI994dd58_29);
nand \U$645 ( \1337 , RI995e3d8_237, RI9921910_609);
and \U$646 ( \1338 , \1335 , \1336 , \1337 );
and \U$647 ( \1339 , \722 , RI98abbc0_55);
and \U$648 ( \1340 , \727 , RI98196b8_68);
nor \U$649 ( \1341 , \1339 , \1340 );
and \U$650 ( \1342 , \735 , RI9967618_211);
and \U$651 ( \1343 , \739 , RI99669e8_224);
nor \U$652 ( \1344 , \1342 , \1343 );
and \U$653 ( \1345 , \744 , RI8946560_133);
and \U$654 ( \1346 , \748 , RI8939d38_146);
nor \U$655 ( \1347 , \1345 , \1346 );
nand \U$656 ( \1348 , \1338 , \1341 , \1344 , \1347 );
and \U$657 ( \1349 , \755 , RI8918b10_185);
and \U$658 ( \1350 , \761 , RI890fb28_198);
nor \U$659 ( \1351 , \1349 , \1350 );
and \U$660 ( \1352 , \769 , RI8930d50_159);
and \U$661 ( \1353 , \773 , RI8925338_172);
nor \U$662 ( \1354 , \1352 , \1353 );
and \U$663 ( \1355 , \779 , RI9776f08_107);
and \U$664 ( \1356 , \784 , RI9808408_94);
nor \U$665 ( \1357 , \1355 , \1356 );
and \U$666 ( \1358 , \788 , RI9808a20_81);
and \U$667 ( \1359 , \792 , RI89ec5c8_120);
nor \U$668 ( \1360 , \1358 , \1359 );
nand \U$669 ( \1361 , \1351 , \1354 , \1357 , \1360 );
nor \U$670 ( \1362 , \1348 , \1361 );
nor \U$671 ( \1363 , \1334 , \1362 );
or \U$672 ( \1364 , \1328 , \1363 );
nand \U$673 ( \1365 , \1334 , \1362 );
nand \U$674 ( \1366 , \1364 , \1365 );
not \U$675 ( \1367 , \1366 );
or \U$676 ( \1368 , \844 , \1367 );
not \U$677 ( \1369 , \842 );
nand \U$678 ( \1370 , \1369 , \835 );
nand \U$679 ( \1371 , \1368 , \1370 );
not \U$680 ( \1372 , \1371 );
or \U$681 ( \1373 , \798 , \1372 );
nand \U$682 ( \1374 , \704 , \796 );
nand \U$683 ( \1375 , \1373 , \1374 );
and \U$684 ( \1376 , RI994e460_14, \703 );
nor \U$685 ( \1377 , \1375 , \1376 );
not \U$686 ( \1378 , \1377 );
nand \U$687 ( \1379 , \1375 , \1376 );
nand \U$688 ( \1380 , \1378 , \1379 );
not \U$689 ( \1381 , \1380 );
nand \U$690 ( \1382 , \797 , \1374 );
xnor \U$691 ( \1383 , \1371 , \1382 );
not \U$692 ( \1384 , \1383 );
nand \U$693 ( \1385 , \1381 , \1384 );
nand \U$694 ( \1386 , \1380 , \1383 );
buf \U$695 ( \1387 , \1366 );
nand \U$696 ( \1388 , \843 , \1370 );
nor \U$697 ( \1389 , \1387 , \1388 );
not \U$698 ( \1390 , \1389 );
nand \U$699 ( \1391 , \1387 , \1388 );
nand \U$700 ( \1392 , \1390 , \1391 );
buf \U$701 ( \1393 , \1392 );
not \U$702 ( \1394 , \1393 );
xor \U$703 ( \1395 , \1394 , \1383 );
and \U$704 ( \1396 , \1385 , \1386 , \1395 );
not \U$705 ( \1397 , \1396 );
not \U$706 ( \1398 , \1380 );
buf \U$707 ( \1399 , \1398 );
not \U$708 ( \1400 , \1399 );
not \U$709 ( \1401 , \764 );
nor \U$710 ( \1402 , RI9921a00_607, RI9921988_608);
nor \U$711 ( \1403 , RI9921a78_606, RI9921910_609);
nor \U$712 ( \1404 , RI9921cd0_601, RI9921b68_604);
nor \U$713 ( \1405 , RI9921c58_602, RI9921af0_605);
nand \U$714 ( \1406 , \1402 , \1403 , \1404 , \1405 );
not \U$715 ( \1407 , \724 );
nand \U$716 ( \1408 , RI9921898_610, RI9921820_611);
not \U$717 ( \1409 , RI9921be0_603);
nand \U$718 ( \1410 , \1407 , \1408 , \1409 );
nor \U$719 ( \1411 , \1406 , \1410 );
not \U$720 ( \1412 , \1411 );
or \U$721 ( \1413 , \1401 , \1412 );
not \U$722 ( \1414 , \1410 );
not \U$723 ( \1415 , \1414 );
not \U$724 ( \1416 , \1406 );
not \U$725 ( \1417 , \1416 );
or \U$726 ( \1418 , \1415 , \1417 );
nand \U$727 ( \1419 , \1418 , RI9921820_611);
nand \U$728 ( \1420 , \1413 , \1419 );
not \U$729 ( \1421 , \1420 );
not \U$730 ( \1422 , RI9921c58_602);
nor \U$731 ( \1423 , RI9921af0_605, RI9921a78_606, RI9921910_609);
nand \U$732 ( \1424 , \1422 , \1423 );
not \U$733 ( \1425 , \1424 );
nor \U$734 ( \1426 , RI9921be0_603, RI9921cd0_601);
nor \U$735 ( \1427 , RI9921b68_604, RI9921a00_607, RI9921988_608);
nand \U$736 ( \1428 , \1426 , \1427 );
not \U$737 ( \1429 , \1428 );
nand \U$738 ( \1430 , RI9921898_610, RI9921820_611, RI99217a8_612, RI9921730_613);
nand \U$739 ( \1431 , \1425 , \1429 , \1430 );
and \U$740 ( \1432 , \1431 , RI9921730_613);
not \U$741 ( \1433 , \1431 );
not \U$742 ( \1434 , RI9921730_613);
and \U$743 ( \1435 , \1433 , \1434 );
nor \U$744 ( \1436 , \1432 , \1435 );
nand \U$745 ( \1437 , \1421 , \1436 );
not \U$746 ( \1438 , \1437 );
buf \U$747 ( \1439 , \1411 );
nand \U$748 ( \1440 , RI9921820_611, \1439 );
nand \U$749 ( \1441 , \1440 , \758 );
buf \U$750 ( \1442 , \1441 );
not \U$751 ( \1443 , RI99217a8_612);
not \U$752 ( \1444 , \1443 );
and \U$753 ( \1445 , \1405 , \1404 , \1403 );
nand \U$754 ( \1446 , RI9921898_610, RI9921820_611, RI99217a8_612);
not \U$755 ( \1447 , RI9921730_613);
nor \U$756 ( \1448 , \1447 , RI9921be0_603);
and \U$757 ( \1449 , \1446 , \1448 , \1402 );
nand \U$758 ( \1450 , \1445 , \1449 );
not \U$759 ( \1451 , \1450 );
not \U$760 ( \1452 , \1451 );
or \U$761 ( \1453 , \1444 , \1452 );
nand \U$762 ( \1454 , \1450 , RI99217a8_612);
nand \U$763 ( \1455 , \1453 , \1454 );
not \U$764 ( \1456 , \1455 );
not \U$765 ( \1457 , \1456 );
nor \U$766 ( \1458 , \1442 , \1457 );
not \U$767 ( \1459 , RI9921910_609);
and \U$768 ( \1460 , \1438 , \1458 , \1459 );
buf \U$769 ( \1461 , \1460 );
nand \U$770 ( \1462 , \1461 , RI994d650_248);
not \U$771 ( \1463 , \1420 );
not \U$772 ( \1464 , \1436 );
nand \U$773 ( \1465 , \1463 , \1464 );
not \U$774 ( \1466 , \1465 );
and \U$775 ( \1467 , \1466 , \1458 );
buf \U$776 ( \1468 , \1467 );
buf \U$777 ( \1469 , \1468 );
not \U$778 ( \1470 , \1469 );
not \U$779 ( \1471 , \1470 );
and \U$780 ( \1472 , \1471 , RI9931b58_268);
not \U$781 ( \1473 , RI9923878_548);
not \U$782 ( \1474 , \735 );
buf \U$783 ( \1475 , \1429 );
nand \U$784 ( \1476 , \1475 , \1425 );
not \U$785 ( \1477 , \1476 );
not \U$786 ( \1478 , \1477 );
or \U$787 ( \1479 , \1474 , \1478 );
nand \U$788 ( \1480 , \739 , \1476 );
nand \U$789 ( \1481 , \1479 , \1480 );
not \U$790 ( \1482 , \1481 );
or \U$791 ( \1483 , \1473 , \1482 );
not \U$792 ( \1484 , \1477 );
not \U$793 ( \1485 , \739 );
or \U$794 ( \1486 , \1484 , \1485 );
nand \U$795 ( \1487 , \1486 , \1459 );
nand \U$796 ( \1488 , \1487 , RI9922f18_568);
nand \U$797 ( \1489 , \1483 , \1488 );
nor \U$798 ( \1490 , \1472 , \1489 );
and \U$799 ( \1491 , \1439 , RI9921820_611);
nor \U$800 ( \1492 , \1491 , RI9921898_610);
not \U$801 ( \1493 , \1456 );
nand \U$802 ( \1494 , \1492 , \1493 );
nand \U$803 ( \1495 , \1464 , \1420 );
nor \U$804 ( \1496 , \1494 , \1495 );
not \U$805 ( \1497 , \1496 );
not \U$806 ( \1498 , \1497 );
buf \U$807 ( \1499 , \1498 );
nand \U$808 ( \1500 , \1499 , RI992a268_388);
nand \U$809 ( \1501 , \1462 , \1490 , \1500 );
nand \U$810 ( \1502 , \1492 , \1493 );
not \U$811 ( \1503 , \1502 );
nand \U$812 ( \1504 , \1503 , \1438 );
not \U$813 ( \1505 , \1504 );
not \U$814 ( \1506 , \1505 );
not \U$815 ( \1507 , \1506 );
not \U$816 ( \1508 , \1507 );
not \U$817 ( \1509 , \1508 );
not \U$818 ( \1510 , RI992f8a8_288);
not \U$819 ( \1511 , \1510 );
and \U$820 ( \1512 , \1509 , \1511 );
not \U$821 ( \1513 , \1465 );
and \U$822 ( \1514 , \1456 , \1441 );
nand \U$823 ( \1515 , \1513 , \1514 );
not \U$824 ( \1516 , \1515 );
not \U$825 ( \1517 , \1516 );
not \U$826 ( \1518 , \1517 );
buf \U$827 ( \1519 , \1518 );
and \U$828 ( \1520 , \1519 , RI9928198_428);
nor \U$829 ( \1521 , \1512 , \1520 );
not \U$830 ( \1522 , \1495 );
and \U$831 ( \1523 , \1522 , \1458 );
not \U$832 ( \1524 , \1523 );
not \U$833 ( \1525 , \1524 );
not \U$834 ( \1526 , \1525 );
not \U$835 ( \1527 , \1526 );
not \U$836 ( \1528 , RI992c6f8_348);
not \U$837 ( \1529 , \1528 );
and \U$838 ( \1530 , \1527 , \1529 );
not \U$839 ( \1531 , \1436 );
nand \U$840 ( \1532 , \1421 , \1531 );
nor \U$841 ( \1533 , \1502 , \1532 );
not \U$842 ( \1534 , \1533 );
not \U$843 ( \1535 , \1534 );
and \U$844 ( \1536 , \1535 , RI992ef48_308);
nor \U$845 ( \1537 , \1530 , \1536 );
nand \U$846 ( \1538 , \1521 , \1537 );
nor \U$847 ( \1539 , \1501 , \1538 );
and \U$848 ( \1540 , \1455 , \1441 );
not \U$849 ( \1541 , \1540 );
not \U$850 ( \1542 , \1541 );
nand \U$851 ( \1543 , \1542 , \1438 );
buf \U$852 ( \1544 , \1543 );
buf \U$853 ( \1545 , \1544 );
not \U$854 ( \1546 , RI9926de8_448);
or \U$855 ( \1547 , \1545 , \1546 );
not \U$856 ( \1548 , \1532 );
and \U$857 ( \1549 , \1540 , \1548 );
buf \U$858 ( \1550 , \1549 );
not \U$859 ( \1551 , \1550 );
not \U$860 ( \1552 , RI9926488_468);
or \U$861 ( \1553 , \1551 , \1552 );
and \U$862 ( \1554 , \1420 , \1436 );
not \U$863 ( \1555 , \1554 );
nor \U$864 ( \1556 , \1555 , \1494 );
buf \U$865 ( \1557 , \1556 );
and \U$866 ( \1558 , \1557 , RI992abc8_368);
not \U$867 ( \1559 , \1541 );
and \U$868 ( \1560 , \1420 , \1436 );
nand \U$869 ( \1561 , \1559 , \1560 );
not \U$870 ( \1562 , \1561 );
not \U$871 ( \1563 , \1562 );
not \U$872 ( \1564 , \1563 );
not \U$873 ( \1565 , \1564 );
not \U$874 ( \1566 , RI99241d8_528);
nor \U$875 ( \1567 , \1565 , \1566 );
nor \U$876 ( \1568 , \1558 , \1567 );
nand \U$877 ( \1569 , \1547 , \1553 , \1568 );
nand \U$878 ( \1570 , \1514 , \1560 );
not \U$879 ( \1571 , \1570 );
not \U$880 ( \1572 , \1571 );
not \U$881 ( \1573 , RI9925b28_488);
nor \U$882 ( \1574 , \1572 , \1573 );
not \U$883 ( \1575 , RI9928af8_408);
nand \U$884 ( \1576 , \1514 , \1438 );
not \U$885 ( \1577 , \1576 );
not \U$886 ( \1578 , \1577 );
nor \U$887 ( \1579 , \1575 , \1578 );
nor \U$888 ( \1580 , \1574 , \1579 );
not \U$889 ( \1581 , \1464 );
buf \U$890 ( \1582 , \1420 );
not \U$891 ( \1583 , \1493 );
buf \U$892 ( \1584 , \1492 );
and \U$893 ( \1585 , \1581 , \1582 , \1583 , \1584 );
buf \U$894 ( \1586 , \1585 );
not \U$895 ( \1587 , \1586 );
not \U$896 ( \1588 , \1587 );
not \U$897 ( \1589 , RI992d058_328);
not \U$898 ( \1590 , \1589 );
and \U$899 ( \1591 , \1588 , \1590 );
nand \U$900 ( \1592 , \1514 , \1522 );
not \U$901 ( \1593 , \1592 );
and \U$902 ( \1594 , \1593 , RI9924b38_508);
nor \U$903 ( \1595 , \1591 , \1594 );
nand \U$904 ( \1596 , \1580 , \1595 );
nor \U$905 ( \1597 , \1569 , \1596 );
nand \U$906 ( \1598 , \1539 , \1597 );
not \U$907 ( \1599 , \1598 );
and \U$908 ( \1600 , \1400 , \1599 );
not \U$909 ( \1601 , \1599 );
and \U$910 ( \1602 , \1399 , \1601 );
nor \U$911 ( \1603 , \1600 , \1602 );
or \U$912 ( \1604 , \1397 , \1603 );
not \U$913 ( \1605 , \1395 );
not \U$914 ( \1606 , \1605 );
or \U$915 ( \1607 , \1606 , \1399 );
nand \U$916 ( \1608 , \1604 , \1607 );
buf \U$918 ( \1609 , \1377 );
not \U$919 ( \1610 , \1609 );
nand \U$920 ( \1611 , \1380 , \1610 );
nand \U$921 ( \1612 , 1'b1 , \1611 );
buf \U$922 ( \1613 , \1612 );
buf \U$923 ( \1614 , \1610 );
not \U$924 ( \1615 , RI994d5d8_249);
not \U$925 ( \1616 , \1461 );
nor \U$926 ( \1617 , \1615 , \1616 );
not \U$927 ( \1618 , RI992a1f0_389);
nor \U$928 ( \1619 , \1497 , \1618 );
nor \U$929 ( \1620 , \1617 , \1619 );
not \U$930 ( \1621 , \1506 );
not \U$931 ( \1622 , RI992f830_289);
not \U$932 ( \1623 , \1622 );
and \U$933 ( \1624 , \1621 , \1623 );
buf \U$934 ( \1625 , \1517 );
not \U$935 ( \1626 , \1625 );
and \U$936 ( \1627 , \1626 , RI9928120_429);
nor \U$937 ( \1628 , \1624 , \1627 );
not \U$938 ( \1629 , \1535 );
not \U$939 ( \1630 , \1629 );
not \U$940 ( \1631 , RI992eed0_309);
not \U$941 ( \1632 , \1631 );
and \U$942 ( \1633 , \1630 , \1632 );
buf \U$943 ( \1634 , \1525 );
not \U$944 ( \1635 , \1634 );
not \U$945 ( \1636 , \1635 );
and \U$946 ( \1637 , \1636 , RI992b4b0_349);
nor \U$947 ( \1638 , \1633 , \1637 );
and \U$948 ( \1639 , \1469 , RI9931ae0_269);
not \U$949 ( \1640 , RI9922bd0_569);
not \U$950 ( \1641 , \1487 );
or \U$951 ( \1642 , \1640 , \1641 );
not \U$952 ( \1643 , \1481 );
not \U$953 ( \1644 , RI9923800_549);
or \U$954 ( \1645 , \1643 , \1644 );
nand \U$955 ( \1646 , \1642 , \1645 );
nor \U$956 ( \1647 , \1639 , \1646 );
nand \U$957 ( \1648 , \1620 , \1628 , \1638 , \1647 );
not \U$958 ( \1649 , \1545 );
not \U$959 ( \1650 , RI9926d70_449);
not \U$960 ( \1651 , \1650 );
and \U$961 ( \1652 , \1649 , \1651 );
buf \U$962 ( \1653 , \1551 );
not \U$963 ( \1654 , RI9926410_469);
nor \U$964 ( \1655 , \1653 , \1654 );
nor \U$965 ( \1656 , \1652 , \1655 );
not \U$966 ( \1657 , \1578 );
and \U$967 ( \1658 , \1657 , RI9928a80_409);
not \U$968 ( \1659 , \1572 );
and \U$969 ( \1660 , \1659 , RI9925ab0_489);
nor \U$970 ( \1661 , \1658 , \1660 );
not \U$971 ( \1662 , \1587 );
not \U$972 ( \1663 , RI992cfe0_329);
not \U$973 ( \1664 , \1663 );
and \U$974 ( \1665 , \1662 , \1664 );
and \U$975 ( \1666 , \1593 , RI9924ac0_509);
nor \U$976 ( \1667 , \1665 , \1666 );
not \U$977 ( \1668 , \1557 );
not \U$978 ( \1669 , \1668 );
not \U$979 ( \1670 , RI992ab50_369);
not \U$980 ( \1671 , \1670 );
and \U$981 ( \1672 , \1669 , \1671 );
not \U$982 ( \1673 , RI9924160_529);
nor \U$983 ( \1674 , \1565 , \1673 );
nor \U$984 ( \1675 , \1672 , \1674 );
nand \U$985 ( \1676 , \1656 , \1661 , \1667 , \1675 );
or \U$986 ( \1677 , \1648 , \1676 );
not \U$987 ( \1678 , \1677 );
and \U$988 ( \1679 , \1614 , \1678 );
not \U$989 ( \1680 , \1614 );
not \U$990 ( \1681 , \1678 );
and \U$991 ( \1682 , \1680 , \1681 );
nor \U$992 ( \1683 , \1679 , \1682 );
nand \U$993 ( \1684 , \1613 , \1683 );
xor \U$994 ( \1685 , \1608 , \1684 );
not \U$995 ( \1686 , \1587 );
not \U$996 ( \1687 , RI992cf68_330);
not \U$997 ( \1688 , \1687 );
and \U$998 ( \1689 , \1686 , \1688 );
and \U$999 ( \1690 , \1593 , RI9924a48_510);
nor \U$1000 ( \1691 , \1689 , \1690 );
nand \U$1001 ( \1692 , \1461 , RI994d560_250);
and \U$1002 ( \1693 , \1469 , RI9931a68_270);
not \U$1003 ( \1694 , RI9922b58_570);
not \U$1004 ( \1695 , \1487 );
or \U$1005 ( \1696 , \1694 , \1695 );
nand \U$1006 ( \1697 , \1481 , RI9923788_550);
nand \U$1007 ( \1698 , \1696 , \1697 );
nor \U$1008 ( \1699 , \1693 , \1698 );
and \U$1009 ( \1700 , \1691 , \1692 , \1699 );
not \U$1010 ( \1701 , RI992aad8_370);
not \U$1011 ( \1702 , \1701 );
nand \U$1012 ( \1703 , \1702 , \1557 );
nand \U$1013 ( \1704 , \1564 , RI99240e8_530);
nand \U$1014 ( \1705 , \1535 , RI992ee58_310);
nand \U$1015 ( \1706 , \1703 , \1704 , \1705 );
not \U$1016 ( \1707 , RI9928a08_410);
not \U$1017 ( \1708 , \1657 );
or \U$1018 ( \1709 , \1707 , \1708 );
not \U$1019 ( \1710 , \1572 );
nand \U$1020 ( \1711 , \1710 , RI9925a38_490);
nand \U$1021 ( \1712 , \1709 , \1711 );
nor \U$1022 ( \1713 , \1706 , \1712 );
not \U$1023 ( \1714 , RI9926cf8_450);
not \U$1024 ( \1715 , \1545 );
not \U$1025 ( \1716 , \1715 );
or \U$1026 ( \1717 , \1714 , \1716 );
nand \U$1027 ( \1718 , \1550 , RI9926398_470);
nand \U$1028 ( \1719 , \1717 , \1718 );
not \U$1029 ( \1720 , RI99280a8_430);
not \U$1030 ( \1721 , \1519 );
or \U$1031 ( \1722 , \1720 , \1721 );
nand \U$1032 ( \1723 , \1634 , RI992b438_350);
nand \U$1033 ( \1724 , \1722 , \1723 );
nor \U$1034 ( \1725 , \1719 , \1724 );
and \U$1035 ( \1726 , \1507 , RI992f7b8_290);
and \U$1036 ( \1727 , \1499 , RI992a178_390);
nor \U$1037 ( \1728 , \1726 , \1727 );
nand \U$1038 ( \1729 , \1700 , \1713 , \1725 , \1728 );
buf \U$1039 ( \1730 , \1729 );
not \U$1040 ( \1731 , \1730 );
and \U$1041 ( \1732 , \1614 , \1731 );
and \U$1042 ( \1733 , \1680 , \1730 );
nor \U$1043 ( \1734 , \1732 , \1733 );
and \U$1044 ( \1735 , \1613 , \1734 );
not \U$1045 ( \1736 , \1327 );
nand \U$1046 ( \1737 , \1736 , \1325 );
not \U$1047 ( \1738 , \1737 );
buf \U$1048 ( \1739 , \1295 );
not \U$1049 ( \1740 , \1739 );
or \U$1050 ( \1741 , \1738 , \1740 );
or \U$1051 ( \1742 , \1737 , \1739 );
nand \U$1052 ( \1743 , \1741 , \1742 );
buf \U$1053 ( \1744 , \1743 );
buf \U$1054 ( \1745 , \1328 );
not \U$1055 ( \1746 , \1363 );
nand \U$1056 ( \1747 , \1746 , \1365 );
and \U$1057 ( \1748 , \1745 , \1747 );
not \U$1058 ( \1749 , \1745 );
not \U$1059 ( \1750 , \1747 );
and \U$1060 ( \1751 , \1749 , \1750 );
nor \U$1061 ( \1752 , \1748 , \1751 );
not \U$1062 ( \1753 , \1752 );
and \U$1063 ( \1754 , \1744 , \1753 );
not \U$1064 ( \1755 , \1744 );
and \U$1065 ( \1756 , \1755 , \1752 );
nor \U$1066 ( \1757 , \1754 , \1756 );
not \U$1067 ( \1758 , \1757 );
not \U$1068 ( \1759 , \1758 );
not \U$1069 ( \1760 , \1759 );
not \U$1070 ( \1761 , \1393 );
nand \U$1071 ( \1762 , \1761 , \1753 );
nand \U$1072 ( \1763 , \1393 , \1752 );
and \U$1073 ( \1764 , \1762 , \1763 , \1757 );
not \U$1074 ( \1765 , \1764 );
not \U$1075 ( \1766 , \1765 );
not \U$1076 ( \1767 , \1766 );
not \U$1077 ( \1768 , \1767 );
or \U$1078 ( \1769 , \1760 , \1768 );
buf \U$1079 ( \1770 , \1393 );
nand \U$1080 ( \1771 , \1769 , \1770 );
xor \U$1081 ( \1772 , \1735 , \1771 );
and \U$1082 ( \1773 , \1400 , \1678 );
and \U$1083 ( \1774 , \1399 , \1681 );
nor \U$1084 ( \1775 , \1773 , \1774 );
or \U$1085 ( \1776 , \1397 , \1775 );
or \U$1086 ( \1777 , \1603 , \1606 );
nand \U$1087 ( \1778 , \1776 , \1777 );
and \U$1088 ( \1779 , \1772 , \1778 );
and \U$1089 ( \1780 , \1735 , \1771 );
or \U$1090 ( \1781 , \1779 , \1780 );
xor \U$1091 ( \1782 , \1685 , \1781 );
and \U$1092 ( \1783 , \1770 , \1599 );
not \U$1093 ( \1784 , \1770 );
and \U$1094 ( \1785 , \1784 , \1601 );
nor \U$1095 ( \1786 , \1783 , \1785 );
or \U$1096 ( \1787 , \1767 , \1786 );
or \U$1097 ( \1788 , \1759 , \1784 );
nand \U$1098 ( \1789 , \1787 , \1788 );
not \U$1099 ( \1790 , \1789 );
and \U$1100 ( \1791 , \1657 , RI9928990_411);
and \U$1101 ( \1792 , \1659 , RI99259c0_491);
nor \U$1102 ( \1793 , \1791 , \1792 );
and \U$1103 ( \1794 , \1557 , RI992aa60_371);
and \U$1104 ( \1795 , \1564 , RI9924070_531);
nor \U$1105 ( \1796 , \1794 , \1795 );
nand \U$1106 ( \1797 , \1535 , RI992ede0_311);
nand \U$1107 ( \1798 , \1793 , \1796 , \1797 );
and \U$1108 ( \1799 , \1626 , RI9928030_431);
and \U$1109 ( \1800 , \1636 , RI992b3c0_351);
nor \U$1110 ( \1801 , \1799 , \1800 );
and \U$1111 ( \1802 , \1715 , RI9926c80_451);
and \U$1112 ( \1803 , \1550 , RI9926320_471);
nor \U$1113 ( \1804 , \1802 , \1803 );
and \U$1114 ( \1805 , \1507 , RI992f740_291);
and \U$1115 ( \1806 , \1498 , RI992a100_391);
nor \U$1116 ( \1807 , \1805 , \1806 );
nand \U$1117 ( \1808 , \1801 , \1804 , \1807 );
nor \U$1118 ( \1809 , \1798 , \1808 );
and \U$1119 ( \1810 , \1469 , RI99319f0_271);
not \U$1120 ( \1811 , RI9922ae0_571);
not \U$1121 ( \1812 , \1487 );
or \U$1122 ( \1813 , \1811 , \1812 );
nand \U$1123 ( \1814 , \1481 , RI9923710_551);
nand \U$1124 ( \1815 , \1813 , \1814 );
nor \U$1125 ( \1816 , \1810 , \1815 );
nand \U$1126 ( \1817 , \1593 , RI99249d0_511);
nand \U$1127 ( \1818 , \1586 , RI992cef0_331);
nand \U$1128 ( \1819 , \1816 , \1817 , \1818 );
not \U$1129 ( \1820 , RI994d4e8_251);
nor \U$1130 ( \1821 , \1820 , \1616 );
nor \U$1131 ( \1822 , \1819 , \1821 );
nand \U$1132 ( \1823 , \1809 , \1822 );
not \U$1133 ( \1824 , \1823 );
and \U$1134 ( \1825 , \1614 , \1824 );
and \U$1135 ( \1826 , \1680 , \1823 );
nor \U$1136 ( \1827 , \1825 , \1826 );
and \U$1137 ( \1828 , \1613 , \1827 );
xor \U$1138 ( \1829 , \1790 , \1828 );
or \U$1139 ( \1830 , \1399 , \1730 );
or \U$1140 ( \1831 , \1400 , \1731 );
nand \U$1141 ( \1832 , \1830 , \1831 );
not \U$1142 ( \1833 , \1832 );
or \U$1143 ( \1834 , \1397 , \1833 );
or \U$1144 ( \1835 , \1775 , \1606 );
nand \U$1145 ( \1836 , \1834 , \1835 );
and \U$1146 ( \1837 , \1829 , \1836 );
and \U$1147 ( \1838 , \1790 , \1828 );
or \U$1148 ( \1839 , \1837 , \1838 );
xor \U$1149 ( \1840 , \1789 , \1839 );
xor \U$1150 ( \1841 , \1735 , \1771 );
xor \U$1151 ( \1842 , \1841 , \1778 );
and \U$1152 ( \1843 , \1840 , \1842 );
and \U$1153 ( \1844 , \1789 , \1839 );
or \U$1154 ( \1845 , \1843 , \1844 );
xor \U$1155 ( \1846 , \1782 , \1845 );
nand \U$1156 ( \1847 , \1279 , \1015 );
not \U$1157 ( \1848 , \1847 );
not \U$1158 ( \1849 , \1272 );
not \U$1159 ( \1850 , \1218 );
or \U$1160 ( \1851 , \1849 , \1850 );
not \U$1161 ( \1852 , \1280 );
nand \U$1162 ( \1853 , \1851 , \1852 );
not \U$1163 ( \1854 , \1853 );
or \U$1164 ( \1855 , \1848 , \1854 );
or \U$1165 ( \1856 , \1847 , \1853 );
nand \U$1166 ( \1857 , \1855 , \1856 );
not \U$1167 ( \1858 , \1857 );
buf \U$1168 ( \1859 , \1218 );
not \U$1169 ( \1860 , \1273 );
nand \U$1170 ( \1861 , \1860 , \1852 );
not \U$1171 ( \1862 , \1861 );
and \U$1172 ( \1863 , \1859 , \1862 );
not \U$1173 ( \1864 , \1859 );
and \U$1174 ( \1865 , \1864 , \1861 );
nor \U$1175 ( \1866 , \1863 , \1865 );
not \U$1176 ( \1867 , \1866 );
nand \U$1177 ( \1868 , \1858 , \1867 );
nand \U$1178 ( \1869 , \1857 , \1866 );
xor \U$1179 ( \1870 , \1019 , \1064 );
xor \U$1180 ( \1871 , \1870 , \1215 );
not \U$1181 ( \1872 , \1871 );
and \U$1182 ( \1873 , \1872 , \1866 );
not \U$1183 ( \1874 , \1872 );
and \U$1184 ( \1875 , \1874 , \1867 );
nor \U$1185 ( \1876 , \1873 , \1875 );
and \U$1186 ( \1877 , \1868 , \1869 , \1876 );
buf \U$1187 ( \1878 , \1877 );
not \U$1188 ( \1879 , \1878 );
and \U$1189 ( \1880 , \1519 , RI9927fb8_432);
and \U$1190 ( \1881 , \1634 , RI992b348_352);
nor \U$1191 ( \1882 , \1880 , \1881 );
and \U$1192 ( \1883 , \1715 , RI9926c08_452);
not \U$1193 ( \1884 , RI99262a8_472);
nor \U$1194 ( \1885 , \1551 , \1884 );
nor \U$1195 ( \1886 , \1883 , \1885 );
and \U$1196 ( \1887 , \1507 , RI992f6c8_292);
and \U$1197 ( \1888 , \1498 , RI9929278_392);
nor \U$1198 ( \1889 , \1887 , \1888 );
nand \U$1199 ( \1890 , \1882 , \1886 , \1889 );
and \U$1200 ( \1891 , \1657 , RI9928918_412);
and \U$1201 ( \1892 , \1659 , RI9925948_492);
nor \U$1202 ( \1893 , \1891 , \1892 );
and \U$1203 ( \1894 , \1557 , RI992a9e8_372);
and \U$1204 ( \1895 , \1564 , RI9923ff8_532);
nor \U$1205 ( \1896 , \1894 , \1895 );
nand \U$1206 ( \1897 , \1535 , RI992ed68_312);
nand \U$1207 ( \1898 , \1893 , \1896 , \1897 );
nor \U$1208 ( \1899 , \1890 , \1898 );
and \U$1209 ( \1900 , \1469 , RI9931978_272);
not \U$1210 ( \1901 , RI9922a68_572);
not \U$1211 ( \1902 , \1487 );
or \U$1212 ( \1903 , \1901 , \1902 );
nand \U$1213 ( \1904 , \1481 , RI9923698_552);
nand \U$1214 ( \1905 , \1903 , \1904 );
nor \U$1215 ( \1906 , \1900 , \1905 );
nand \U$1216 ( \1907 , \1593 , RI9924958_512);
nand \U$1217 ( \1908 , \1586 , RI992ce78_332);
nand \U$1218 ( \1909 , \1906 , \1907 , \1908 );
and \U$1219 ( \1910 , \1461 , RI994d470_252);
nor \U$1220 ( \1911 , \1909 , \1910 );
nand \U$1221 ( \1912 , \1899 , \1911 );
not \U$1222 ( \1913 , \1912 );
buf \U$1223 ( \1914 , \1857 );
not \U$1224 ( \1915 , \1914 );
and \U$1225 ( \1916 , \1913 , \1915 );
not \U$1226 ( \1917 , \1913 );
and \U$1227 ( \1918 , \1917 , \1914 );
nor \U$1228 ( \1919 , \1916 , \1918 );
not \U$1229 ( \1920 , \1919 );
or \U$1230 ( \1921 , \1879 , \1920 );
not \U$1231 ( \1922 , \1857 );
and \U$1232 ( \1923 , \1824 , \1922 );
not \U$1233 ( \1924 , \1824 );
not \U$1234 ( \1925 , \1922 );
and \U$1235 ( \1926 , \1924 , \1925 );
nor \U$1236 ( \1927 , \1923 , \1926 );
buf \U$1237 ( \1928 , \1876 );
not \U$1238 ( \1929 , \1928 );
nand \U$1239 ( \1930 , \1927 , \1929 );
nand \U$1240 ( \1931 , \1921 , \1930 );
nand \U$1241 ( \1932 , \1214 , \1116 );
buf \U$1242 ( \1933 , \1210 );
xnor \U$1243 ( \1934 , \1932 , \1933 );
and \U$1244 ( \1935 , \1871 , \1934 );
not \U$1245 ( \1936 , \1871 );
not \U$1246 ( \1937 , \1934 );
and \U$1247 ( \1938 , \1936 , \1937 );
nor \U$1248 ( \1939 , \1935 , \1938 );
and \U$1249 ( \1940 , \1209 , \1168 );
buf \U$1250 ( \1941 , \1205 );
xor \U$1251 ( \1942 , \1940 , \1941 );
and \U$1252 ( \1943 , \1934 , \1942 );
not \U$1253 ( \1944 , \1934 );
not \U$1254 ( \1945 , \1942 );
and \U$1255 ( \1946 , \1944 , \1945 );
or \U$1256 ( \1947 , \1943 , \1946 );
nand \U$1257 ( \1948 , \1939 , \1947 );
not \U$1258 ( \1949 , \1948 );
not \U$1259 ( \1950 , \1949 );
not \U$1260 ( \1951 , \1872 );
not \U$1261 ( \1952 , \1951 );
not \U$1262 ( \1953 , \1824 );
or \U$1263 ( \1954 , \1952 , \1953 );
nand \U$1264 ( \1955 , \1823 , \1872 );
nand \U$1265 ( \1956 , \1954 , \1955 );
not \U$1266 ( \1957 , \1956 );
or \U$1267 ( \1958 , \1950 , \1957 );
and \U$1268 ( \1959 , \1951 , \1730 );
not \U$1269 ( \1960 , \1951 );
and \U$1270 ( \1961 , \1960 , \1731 );
nor \U$1271 ( \1962 , \1959 , \1961 );
buf \U$1272 ( \1963 , \1947 );
not \U$1273 ( \1964 , \1963 );
nand \U$1274 ( \1965 , \1962 , \1964 );
nand \U$1275 ( \1966 , \1958 , \1965 );
not \U$1276 ( \1967 , \1945 );
not \U$1277 ( \1968 , RI994dec0_26);
not \U$1278 ( \1969 , \1203 );
not \U$1279 ( \1970 , \1969 );
or \U$1280 ( \1971 , \1968 , \1970 );
nand \U$1281 ( \1972 , \1971 , \1941 );
buf \U$1282 ( \1973 , \1972 );
not \U$1283 ( \1974 , \1973 );
and \U$1284 ( \1975 , \1967 , \1974 );
not \U$1285 ( \1976 , \1975 );
and \U$1286 ( \1977 , \1967 , \1677 );
not \U$1287 ( \1978 , \1967 );
not \U$1288 ( \1979 , \1677 );
and \U$1289 ( \1980 , \1978 , \1979 );
nor \U$1290 ( \1981 , \1977 , \1980 );
not \U$1291 ( \1982 , \1981 );
or \U$1292 ( \1983 , \1976 , \1982 );
not \U$1293 ( \1984 , \1967 );
not \U$1294 ( \1985 , \1599 );
or \U$1295 ( \1986 , \1984 , \1985 );
nand \U$1296 ( \1987 , \1598 , \1945 );
nand \U$1297 ( \1988 , \1986 , \1987 );
nand \U$1298 ( \1989 , \1988 , \1973 );
nand \U$1299 ( \1990 , \1983 , \1989 );
and \U$1300 ( \1991 , \1966 , \1990 );
xor \U$1301 ( \1992 , \1931 , \1991 );
not \U$1302 ( \1993 , \1945 );
not \U$1303 ( \1994 , \1974 );
and \U$1304 ( \1995 , \1993 , \1994 );
and \U$1305 ( \1996 , \1988 , \1975 );
nor \U$1306 ( \1997 , \1995 , \1996 );
not \U$1307 ( \1998 , \1997 );
not \U$1308 ( \1999 , \1949 );
not \U$1309 ( \2000 , \1962 );
or \U$1310 ( \2001 , \1999 , \2000 );
and \U$1311 ( \2002 , \1951 , \1677 );
not \U$1312 ( \2003 , \1951 );
and \U$1313 ( \2004 , \2003 , \1979 );
nor \U$1314 ( \2005 , \2002 , \2004 );
nand \U$1315 ( \2006 , \2005 , \1964 );
nand \U$1316 ( \2007 , \2001 , \2006 );
not \U$1317 ( \2008 , \2007 );
or \U$1318 ( \2009 , \1998 , \2008 );
or \U$1319 ( \2010 , \2007 , \1997 );
nand \U$1320 ( \2011 , \2009 , \2010 );
xor \U$1321 ( \2012 , \1992 , \2011 );
not \U$1322 ( \2013 , \966 );
not \U$1323 ( \2014 , \1015 );
not \U$1324 ( \2015 , \1853 );
or \U$1325 ( \2016 , \2014 , \2015 );
nand \U$1326 ( \2017 , \2016 , \1279 );
not \U$1327 ( \2018 , \2017 );
or \U$1328 ( \2019 , \2013 , \2018 );
not \U$1329 ( \2020 , \1284 );
nand \U$1330 ( \2021 , \2019 , \2020 );
nand \U$1331 ( \2022 , \1288 , \937 );
and \U$1332 ( \2023 , \2021 , \2022 );
not \U$1333 ( \2024 , \2021 );
not \U$1334 ( \2025 , \2022 );
and \U$1335 ( \2026 , \2024 , \2025 );
or \U$1336 ( \2027 , \2023 , \2026 );
buf \U$1337 ( \2028 , \2027 );
not \U$1338 ( \2029 , \2028 );
not \U$1339 ( \2030 , \2029 );
nand \U$1340 ( \2031 , \1461 , RI9935fc8_254);
and \U$1341 ( \2032 , \1469 , RI9931888_274);
not \U$1342 ( \2033 , RI9922978_574);
not \U$1343 ( \2034 , \1487 );
or \U$1344 ( \2035 , \2033 , \2034 );
not \U$1345 ( \2036 , RI99235a8_554);
or \U$1346 ( \2037 , \1643 , \2036 );
nand \U$1347 ( \2038 , \2035 , \2037 );
nor \U$1348 ( \2039 , \2032 , \2038 );
nand \U$1349 ( \2040 , \1498 , RI9929188_394);
nand \U$1350 ( \2041 , \2031 , \2039 , \2040 );
not \U$1351 ( \2042 , \1506 );
not \U$1352 ( \2043 , RI992f5d8_294);
not \U$1353 ( \2044 , \2043 );
and \U$1354 ( \2045 , \2042 , \2044 );
and \U$1355 ( \2046 , \1626 , RI9927ec8_434);
nor \U$1356 ( \2047 , \2045 , \2046 );
not \U$1357 ( \2048 , \1629 );
not \U$1358 ( \2049 , RI992d6e8_314);
not \U$1359 ( \2050 , \2049 );
and \U$1360 ( \2051 , \2048 , \2050 );
and \U$1361 ( \2052 , \1634 , RI992b258_354);
nor \U$1362 ( \2053 , \2051 , \2052 );
nand \U$1363 ( \2054 , \2047 , \2053 );
nor \U$1364 ( \2055 , \2041 , \2054 );
and \U$1365 ( \2056 , \1715 , RI9926b18_454);
not \U$1366 ( \2057 , RI99261b8_474);
nor \U$1367 ( \2058 , \1551 , \2057 );
nor \U$1368 ( \2059 , \2056 , \2058 );
not \U$1369 ( \2060 , \1668 );
not \U$1370 ( \2061 , RI992a8f8_374);
not \U$1371 ( \2062 , \2061 );
and \U$1372 ( \2063 , \2060 , \2062 );
not \U$1373 ( \2064 , RI9923f08_534);
nor \U$1374 ( \2065 , \1565 , \2064 );
nor \U$1375 ( \2066 , \2063 , \2065 );
nand \U$1376 ( \2067 , \2059 , \2066 );
and \U$1377 ( \2068 , \1657 , RI9928828_414);
and \U$1378 ( \2069 , \1710 , RI9925858_494);
nor \U$1379 ( \2070 , \2068 , \2069 );
and \U$1380 ( \2071 , \1586 , RI992cd88_334);
and \U$1381 ( \2072 , \1593 , RI9924868_514);
nor \U$1382 ( \2073 , \2071 , \2072 );
nand \U$1383 ( \2074 , \2070 , \2073 );
nor \U$1384 ( \2075 , \2067 , \2074 );
nand \U$1385 ( \2076 , \2055 , \2075 );
not \U$1386 ( \2077 , \2076 );
or \U$1387 ( \2078 , \2030 , \2077 );
buf \U$1388 ( \2079 , \2028 );
not \U$1389 ( \2080 , \2076 );
nand \U$1390 ( \2081 , \2079 , \2080 );
nand \U$1391 ( \2082 , \2078 , \2081 );
not \U$1392 ( \2083 , \2082 );
nand \U$1393 ( \2084 , \2020 , \966 );
not \U$1394 ( \2085 , \2084 );
not \U$1395 ( \2086 , \2017 );
or \U$1396 ( \2087 , \2085 , \2086 );
or \U$1397 ( \2088 , \2017 , \2084 );
nand \U$1398 ( \2089 , \2087 , \2088 );
and \U$1399 ( \2090 , \2028 , \2089 );
not \U$1400 ( \2091 , \2028 );
not \U$1401 ( \2092 , \2089 );
and \U$1402 ( \2093 , \2091 , \2092 );
or \U$1403 ( \2094 , \2090 , \2093 );
not \U$1404 ( \2095 , \1925 );
not \U$1405 ( \2096 , \2092 );
or \U$1406 ( \2097 , \2095 , \2096 );
nand \U$1407 ( \2098 , \2089 , \1915 );
nand \U$1408 ( \2099 , \2097 , \2098 );
nor \U$1409 ( \2100 , \2094 , \2099 );
not \U$1410 ( \2101 , \2100 );
or \U$1411 ( \2102 , \2083 , \2101 );
nand \U$1412 ( \2103 , \1461 , RI994d3f8_253);
and \U$1413 ( \2104 , \1471 , RI9931900_273);
not \U$1414 ( \2105 , RI99229f0_573);
not \U$1415 ( \2106 , \1487 );
or \U$1416 ( \2107 , \2105 , \2106 );
not \U$1417 ( \2108 , RI9923620_553);
or \U$1418 ( \2109 , \1643 , \2108 );
nand \U$1419 ( \2110 , \2107 , \2109 );
nor \U$1420 ( \2111 , \2104 , \2110 );
nand \U$1421 ( \2112 , \1499 , RI9929200_393);
nand \U$1422 ( \2113 , \2103 , \2111 , \2112 );
not \U$1423 ( \2114 , \1508 );
not \U$1424 ( \2115 , RI992f650_293);
not \U$1425 ( \2116 , \2115 );
and \U$1426 ( \2117 , \2114 , \2116 );
and \U$1427 ( \2118 , \1626 , RI9927f40_433);
nor \U$1428 ( \2119 , \2117 , \2118 );
not \U$1429 ( \2120 , \1629 );
not \U$1430 ( \2121 , RI992ecf0_313);
not \U$1431 ( \2122 , \2121 );
and \U$1432 ( \2123 , \2120 , \2122 );
and \U$1433 ( \2124 , \1634 , RI992b2d0_353);
nor \U$1434 ( \2125 , \2123 , \2124 );
nand \U$1435 ( \2126 , \2119 , \2125 );
nor \U$1436 ( \2127 , \2113 , \2126 );
and \U$1437 ( \2128 , \1715 , RI9926b90_453);
not \U$1438 ( \2129 , RI9926230_473);
nor \U$1439 ( \2130 , \1551 , \2129 );
nor \U$1440 ( \2131 , \2128 , \2130 );
not \U$1441 ( \2132 , \1668 );
not \U$1442 ( \2133 , RI992a970_373);
not \U$1443 ( \2134 , \2133 );
and \U$1444 ( \2135 , \2132 , \2134 );
not \U$1445 ( \2136 , RI9923f80_533);
nor \U$1446 ( \2137 , \1565 , \2136 );
nor \U$1447 ( \2138 , \2135 , \2137 );
nand \U$1448 ( \2139 , \2131 , \2138 );
and \U$1449 ( \2140 , \1657 , RI99288a0_413);
and \U$1450 ( \2141 , \1659 , RI99258d0_493);
nor \U$1451 ( \2142 , \2140 , \2141 );
and \U$1452 ( \2143 , \1586 , RI992ce00_333);
and \U$1453 ( \2144 , \1593 , RI99248e0_513);
nor \U$1454 ( \2145 , \2143 , \2144 );
nand \U$1455 ( \2146 , \2142 , \2145 );
nor \U$1456 ( \2147 , \2139 , \2146 );
nand \U$1457 ( \2148 , \2127 , \2147 );
not \U$1458 ( \2149 , \2148 );
buf \U$1459 ( \2150 , \2149 );
not \U$1460 ( \2151 , \2150 );
not \U$1461 ( \2152 , \2151 );
not \U$1462 ( \2153 , \2029 );
or \U$1463 ( \2154 , \2152 , \2153 );
nand \U$1464 ( \2155 , \2028 , \2150 );
nand \U$1465 ( \2156 , \2154 , \2155 );
buf \U$1466 ( \2157 , \2099 );
nand \U$1467 ( \2158 , \2156 , \2157 );
nand \U$1468 ( \2159 , \2102 , \2158 );
not \U$1469 ( \2160 , \1564 );
not \U$1470 ( \2161 , RI9923e18_536);
nor \U$1471 ( \2162 , \2160 , \2161 );
not \U$1472 ( \2163 , RI992a808_376);
nor \U$1473 ( \2164 , \1668 , \2163 );
nor \U$1474 ( \2165 , \2162 , \2164 );
and \U$1475 ( \2166 , \1657 , RI9928738_416);
and \U$1476 ( \2167 , \1710 , RI9925768_496);
nor \U$1477 ( \2168 , \2166 , \2167 );
nand \U$1478 ( \2169 , \1535 , RI992d5f8_316);
nand \U$1479 ( \2170 , \2165 , \2168 , \2169 );
and \U$1480 ( \2171 , \1715 , RI9926a28_456);
not \U$1481 ( \2172 , RI99260c8_476);
nor \U$1482 ( \2173 , \2172 , \1551 );
nor \U$1483 ( \2174 , \2171 , \2173 );
and \U$1484 ( \2175 , \1626 , RI9927dd8_436);
and \U$1485 ( \2176 , \1634 , RI992b168_356);
nor \U$1486 ( \2177 , \2175 , \2176 );
not \U$1487 ( \2178 , \1508 );
not \U$1488 ( \2179 , RI992f4e8_296);
not \U$1489 ( \2180 , \2179 );
and \U$1490 ( \2181 , \2178 , \2180 );
and \U$1491 ( \2182 , \1498 , RI9929098_396);
nor \U$1492 ( \2183 , \2181 , \2182 );
nand \U$1493 ( \2184 , \2174 , \2177 , \2183 );
nor \U$1494 ( \2185 , \2170 , \2184 );
and \U$1495 ( \2186 , \1586 , RI992cc98_336);
and \U$1496 ( \2187 , \1593 , RI9924778_516);
nor \U$1497 ( \2188 , \2186 , \2187 );
and \U$1498 ( \2189 , \1469 , RI9931798_276);
not \U$1499 ( \2190 , RI9922888_576);
not \U$1500 ( \2191 , \1487 );
or \U$1501 ( \2192 , \2190 , \2191 );
nand \U$1502 ( \2193 , \1481 , RI99234b8_556);
nand \U$1503 ( \2194 , \2192 , \2193 );
nor \U$1504 ( \2195 , \2189 , \2194 );
nand \U$1505 ( \2196 , \2188 , \2195 );
and \U$1506 ( \2197 , \1461 , RI9935ed8_256);
nor \U$1507 ( \2198 , \2196 , \2197 );
nand \U$1508 ( \2199 , \2185 , \2198 );
and \U$1509 ( \2200 , \2199 , \1744 );
not \U$1510 ( \2201 , \2199 );
not \U$1511 ( \2202 , \1744 );
and \U$1512 ( \2203 , \2201 , \2202 );
nor \U$1513 ( \2204 , \2200 , \2203 );
not \U$1514 ( \2205 , \2204 );
not \U$1515 ( \2206 , \2028 );
not \U$1516 ( \2207 , \1287 );
nand \U$1517 ( \2208 , \2207 , \1292 );
not \U$1518 ( \2209 , \2208 );
not \U$1519 ( \2210 , \937 );
not \U$1520 ( \2211 , \2021 );
or \U$1521 ( \2212 , \2210 , \2211 );
nand \U$1522 ( \2213 , \2212 , \1288 );
not \U$1523 ( \2214 , \2213 );
or \U$1524 ( \2215 , \2209 , \2214 );
or \U$1525 ( \2216 , \2213 , \2208 );
nand \U$1526 ( \2217 , \2215 , \2216 );
nand \U$1527 ( \2218 , \2206 , \2217 );
not \U$1528 ( \2219 , \2218 );
or \U$1529 ( \2220 , \1744 , \2217 );
nand \U$1530 ( \2221 , \2028 , \1744 );
nand \U$1531 ( \2222 , \2220 , \2221 );
nor \U$1532 ( \2223 , \2219 , \2222 );
not \U$1533 ( \2224 , \2223 );
or \U$1534 ( \2225 , \2205 , \2224 );
not \U$1535 ( \2226 , \2079 );
not \U$1536 ( \2227 , \2217 );
not \U$1537 ( \2228 , \2227 );
or \U$1538 ( \2229 , \2226 , \2228 );
nand \U$1539 ( \2230 , \2229 , \2218 );
not \U$1540 ( \2231 , RI9926140_475);
nor \U$1541 ( \2232 , \2231 , \1551 );
not \U$1542 ( \2233 , \1544 );
and \U$1543 ( \2234 , RI9926aa0_455, \2233 );
nor \U$1544 ( \2235 , \2232 , \2234 );
not \U$1545 ( \2236 , \1635 );
not \U$1546 ( \2237 , RI992b1e0_355);
not \U$1547 ( \2238 , \2237 );
and \U$1548 ( \2239 , \2236 , \2238 );
and \U$1549 ( \2240 , \1626 , RI9927e50_435);
nor \U$1550 ( \2241 , \2239 , \2240 );
not \U$1551 ( \2242 , RI9929110_395);
nor \U$1552 ( \2243 , \2242 , \1497 );
not \U$1553 ( \2244 , RI992f560_295);
nor \U$1554 ( \2245 , \1506 , \2244 );
nor \U$1555 ( \2246 , \2243 , \2245 );
nand \U$1556 ( \2247 , \2235 , \2241 , \2246 );
not \U$1557 ( \2248 , RI99257e0_495);
nor \U$1558 ( \2249 , \1572 , \2248 );
not \U$1559 ( \2250 , RI99287b0_415);
nor \U$1560 ( \2251 , \1578 , \2250 );
nor \U$1561 ( \2252 , \2249 , \2251 );
not \U$1562 ( \2253 , RI9923e90_535);
nor \U$1563 ( \2254 , \1563 , \2253 );
not \U$1564 ( \2255 , RI992a880_375);
nor \U$1565 ( \2256 , \1668 , \2255 );
nor \U$1566 ( \2257 , \2254 , \2256 );
nand \U$1567 ( \2258 , \1535 , RI992d670_315);
nand \U$1568 ( \2259 , \2252 , \2257 , \2258 );
nor \U$1569 ( \2260 , \2247 , \2259 );
nand \U$1570 ( \2261 , \1593 , RI99247f0_515);
nand \U$1571 ( \2262 , \1586 , RI992cd10_335);
nand \U$1572 ( \2263 , \1469 , RI9931810_275);
and \U$1573 ( \2264 , \1481 , RI9923530_555);
and \U$1574 ( \2265 , \1487 , RI9922900_575);
nor \U$1575 ( \2266 , \2264 , \2265 );
nand \U$1576 ( \2267 , \2261 , \2262 , \2263 , \2266 );
and \U$1577 ( \2268 , \1461 , RI9935f50_255);
nor \U$1578 ( \2269 , \2267 , \2268 );
nand \U$1579 ( \2270 , \2260 , \2269 );
buf \U$1580 ( \2271 , \2270 );
or \U$1581 ( \2272 , \2202 , \2271 );
not \U$1582 ( \2273 , \2271 );
or \U$1583 ( \2274 , \1744 , \2273 );
nand \U$1584 ( \2275 , \2272 , \2274 );
nand \U$1585 ( \2276 , \2230 , \2275 );
nand \U$1586 ( \2277 , \2225 , \2276 );
xor \U$1587 ( \2278 , \2159 , \2277 );
not \U$1588 ( \2279 , RI9933d18_258);
nor \U$1589 ( \2280 , \2279 , \1616 );
not \U$1590 ( \2281 , RI9928fa8_398);
nor \U$1591 ( \2282 , \1497 , \2281 );
nor \U$1592 ( \2283 , \2280 , \2282 );
not \U$1593 ( \2284 , \1625 );
not \U$1594 ( \2285 , RI9927ce8_438);
not \U$1595 ( \2286 , \2285 );
and \U$1596 ( \2287 , \2284 , \2286 );
not \U$1597 ( \2288 , \1506 );
and \U$1598 ( \2289 , \2288 , RI992f3f8_298);
nor \U$1599 ( \2290 , \2287 , \2289 );
not \U$1600 ( \2291 , \1629 );
not \U$1601 ( \2292 , RI992d508_318);
not \U$1602 ( \2293 , \2292 );
and \U$1603 ( \2294 , \2291 , \2293 );
not \U$1604 ( \2295 , \1526 );
and \U$1605 ( \2296 , \2295 , RI992b078_358);
nor \U$1606 ( \2297 , \2294 , \2296 );
and \U$1607 ( \2298 , \1471 , RI99316a8_278);
not \U$1608 ( \2299 , RI9922798_578);
not \U$1609 ( \2300 , \1487 );
or \U$1610 ( \2301 , \2299 , \2300 );
not \U$1611 ( \2302 , RI99233c8_558);
or \U$1612 ( \2303 , \1643 , \2302 );
nand \U$1613 ( \2304 , \2301 , \2303 );
nor \U$1614 ( \2305 , \2298 , \2304 );
nand \U$1615 ( \2306 , \2283 , \2290 , \2297 , \2305 );
not \U$1616 ( \2307 , \1587 );
not \U$1617 ( \2308 , RI992cba8_338);
not \U$1618 ( \2309 , \2308 );
and \U$1619 ( \2310 , \2307 , \2309 );
and \U$1620 ( \2311 , \1593 , RI9924688_518);
nor \U$1621 ( \2312 , \2310 , \2311 );
and \U$1622 ( \2313 , \1657 , RI9928648_418);
and \U$1623 ( \2314 , \1710 , RI9925678_498);
nor \U$1624 ( \2315 , \2313 , \2314 );
not \U$1625 ( \2316 , \1545 );
not \U$1626 ( \2317 , RI9926938_458);
not \U$1627 ( \2318 , \2317 );
and \U$1628 ( \2319 , \2316 , \2318 );
not \U$1629 ( \2320 , RI9925fd8_478);
nor \U$1630 ( \2321 , \1653 , \2320 );
nor \U$1631 ( \2322 , \2319 , \2321 );
not \U$1632 ( \2323 , \1668 );
not \U$1633 ( \2324 , RI992a718_378);
not \U$1634 ( \2325 , \2324 );
and \U$1635 ( \2326 , \2323 , \2325 );
not \U$1636 ( \2327 , RI9923d28_538);
nor \U$1637 ( \2328 , \1565 , \2327 );
nor \U$1638 ( \2329 , \2326 , \2328 );
nand \U$1639 ( \2330 , \2312 , \2315 , \2322 , \2329 );
nor \U$1640 ( \2331 , \2306 , \2330 );
not \U$1641 ( \2332 , \2331 );
not \U$1642 ( \2333 , \2332 );
not \U$1643 ( \2334 , \1393 );
not \U$1644 ( \2335 , \2334 );
or \U$1645 ( \2336 , \2333 , \2335 );
not \U$1646 ( \2337 , \1394 );
not \U$1647 ( \2338 , \2332 );
nand \U$1648 ( \2339 , \2337 , \2338 );
nand \U$1649 ( \2340 , \2336 , \2339 );
not \U$1650 ( \2341 , \2340 );
not \U$1651 ( \2342 , \1766 );
or \U$1652 ( \2343 , \2341 , \2342 );
not \U$1653 ( \2344 , \2334 );
not \U$1654 ( \2345 , \1545 );
not \U$1655 ( \2346 , RI99269b0_457);
not \U$1656 ( \2347 , \2346 );
and \U$1657 ( \2348 , \2345 , \2347 );
not \U$1658 ( \2349 , RI9926050_477);
nor \U$1659 ( \2350 , \1653 , \2349 );
nor \U$1660 ( \2351 , \2348 , \2350 );
and \U$1661 ( \2352 , \1657 , RI99286c0_417);
and \U$1662 ( \2353 , \1710 , RI99256f0_497);
nor \U$1663 ( \2354 , \2352 , \2353 );
not \U$1664 ( \2355 , \1587 );
not \U$1665 ( \2356 , RI992cc20_337);
not \U$1666 ( \2357 , \2356 );
and \U$1667 ( \2358 , \2355 , \2357 );
and \U$1668 ( \2359 , \1593 , RI9924700_517);
nor \U$1669 ( \2360 , \2358 , \2359 );
not \U$1670 ( \2361 , \1668 );
not \U$1671 ( \2362 , RI992a790_377);
not \U$1672 ( \2363 , \2362 );
and \U$1673 ( \2364 , \2361 , \2363 );
not \U$1674 ( \2365 , RI9923da0_537);
nor \U$1675 ( \2366 , \1565 , \2365 );
nor \U$1676 ( \2367 , \2364 , \2366 );
nand \U$1677 ( \2368 , \2351 , \2354 , \2360 , \2367 );
not \U$1678 ( \2369 , RI9933d90_257);
nor \U$1679 ( \2370 , \2369 , \1616 );
not \U$1680 ( \2371 , RI9929020_397);
nor \U$1681 ( \2372 , \1497 , \2371 );
nor \U$1682 ( \2373 , \2370 , \2372 );
not \U$1683 ( \2374 , \1519 );
not \U$1684 ( \2375 , \2374 );
not \U$1685 ( \2376 , RI9927d60_437);
not \U$1686 ( \2377 , \2376 );
and \U$1687 ( \2378 , \2375 , \2377 );
and \U$1688 ( \2379 , \1507 , RI992f470_297);
nor \U$1689 ( \2380 , \2378 , \2379 );
not \U$1690 ( \2381 , \1629 );
not \U$1691 ( \2382 , RI992d580_317);
not \U$1692 ( \2383 , \2382 );
and \U$1693 ( \2384 , \2381 , \2383 );
and \U$1694 ( \2385 , \1636 , RI992b0f0_357);
nor \U$1695 ( \2386 , \2384 , \2385 );
and \U$1696 ( \2387 , \1469 , RI9931720_277);
not \U$1697 ( \2388 , RI9922810_577);
not \U$1698 ( \2389 , \1487 );
or \U$1699 ( \2390 , \2388 , \2389 );
not \U$1700 ( \2391 , RI9923440_557);
or \U$1701 ( \2392 , \1643 , \2391 );
nand \U$1702 ( \2393 , \2390 , \2392 );
nor \U$1703 ( \2394 , \2387 , \2393 );
nand \U$1704 ( \2395 , \2373 , \2380 , \2386 , \2394 );
or \U$1705 ( \2396 , \2368 , \2395 );
not \U$1706 ( \2397 , \2396 );
not \U$1707 ( \2398 , \2397 );
not \U$1708 ( \2399 , \2398 );
or \U$1709 ( \2400 , \2344 , \2399 );
nand \U$1710 ( \2401 , \1770 , \2397 );
nand \U$1711 ( \2402 , \2400 , \2401 );
nand \U$1712 ( \2403 , \2402 , \1758 );
nand \U$1713 ( \2404 , \2343 , \2403 );
xor \U$1714 ( \2405 , \2278 , \2404 );
xor \U$1715 ( \2406 , \2012 , \2405 );
not \U$1716 ( \2407 , \2271 );
not \U$1717 ( \2408 , \2079 );
not \U$1718 ( \2409 , \2408 );
or \U$1719 ( \2410 , \2407 , \2409 );
nand \U$1720 ( \2411 , \2079 , \2273 );
nand \U$1721 ( \2412 , \2410 , \2411 );
not \U$1722 ( \2413 , \2412 );
buf \U$1723 ( \2414 , \2100 );
not \U$1724 ( \2415 , \2414 );
or \U$1725 ( \2416 , \2413 , \2415 );
nand \U$1726 ( \2417 , \2082 , \2157 );
nand \U$1727 ( \2418 , \2416 , \2417 );
nand \U$1728 ( \2419 , \1461 , RI9933ca0_259);
and \U$1729 ( \2420 , \1469 , RI9931630_279);
not \U$1730 ( \2421 , RI9922720_579);
not \U$1731 ( \2422 , \1487 );
or \U$1732 ( \2423 , \2421 , \2422 );
not \U$1733 ( \2424 , RI9923350_559);
or \U$1734 ( \2425 , \1643 , \2424 );
nand \U$1735 ( \2426 , \2423 , \2425 );
nor \U$1736 ( \2427 , \2420 , \2426 );
nand \U$1737 ( \2428 , \1498 , RI9928f30_399);
nand \U$1738 ( \2429 , \2419 , \2427 , \2428 );
not \U$1739 ( \2430 , \1506 );
not \U$1740 ( \2431 , RI992f380_299);
not \U$1741 ( \2432 , \2431 );
and \U$1742 ( \2433 , \2430 , \2432 );
and \U$1743 ( \2434 , \1519 , RI9927c70_439);
nor \U$1744 ( \2435 , \2433 , \2434 );
and \U$1745 ( \2436 , \1535 , RI992d490_319);
and \U$1746 ( \2437 , \1634 , RI992b000_359);
nor \U$1747 ( \2438 , \2436 , \2437 );
nand \U$1748 ( \2439 , \2435 , \2438 );
nor \U$1749 ( \2440 , \2429 , \2439 );
and \U$1750 ( \2441 , \2233 , RI99268c0_459);
and \U$1751 ( \2442 , \1550 , RI9925f60_479);
nor \U$1752 ( \2443 , \2441 , \2442 );
and \U$1753 ( \2444 , \1557 , RI992a6a0_379);
not \U$1754 ( \2445 , \1563 );
and \U$1755 ( \2446 , \2445 , RI9923cb0_539);
nor \U$1756 ( \2447 , \2444 , \2446 );
nand \U$1757 ( \2448 , \2443 , \2447 );
and \U$1758 ( \2449 , \1657 , RI99285d0_419);
and \U$1759 ( \2450 , \1710 , RI9925600_499);
nor \U$1760 ( \2451 , \2449 , \2450 );
and \U$1761 ( \2452 , \1586 , RI992cb30_339);
and \U$1762 ( \2453 , \1593 , RI9924610_519);
nor \U$1763 ( \2454 , \2452 , \2453 );
nand \U$1764 ( \2455 , \2451 , \2454 );
nor \U$1765 ( \2456 , \2448 , \2455 );
nand \U$1766 ( \2457 , \2440 , \2456 );
not \U$1767 ( \2458 , \2457 );
not \U$1768 ( \2459 , \1394 );
or \U$1769 ( \2460 , \2458 , \2459 );
not \U$1770 ( \2461 , \2457 );
nand \U$1771 ( \2462 , \1393 , \2461 );
nand \U$1772 ( \2463 , \2460 , \2462 );
not \U$1773 ( \2464 , \2463 );
buf \U$1774 ( \2465 , \1764 );
not \U$1775 ( \2466 , \2465 );
or \U$1776 ( \2467 , \2464 , \2466 );
nand \U$1777 ( \2468 , \2340 , \1758 );
nand \U$1778 ( \2469 , \2467 , \2468 );
xor \U$1779 ( \2470 , \2418 , \2469 );
not \U$1780 ( \2471 , \2204 );
buf \U$1781 ( \2472 , \2230 );
not \U$1782 ( \2473 , \2472 );
or \U$1783 ( \2474 , \2471 , \2473 );
and \U$1784 ( \2475 , \1744 , \2397 );
and \U$1785 ( \2476 , \2202 , \2398 );
nor \U$1786 ( \2477 , \2475 , \2476 );
not \U$1787 ( \2478 , \2477 );
buf \U$1788 ( \2479 , \2223 );
nand \U$1789 ( \2480 , \2478 , \2479 );
nand \U$1790 ( \2481 , \2474 , \2480 );
and \U$1791 ( \2482 , \2470 , \2481 );
and \U$1792 ( \2483 , \2418 , \2469 );
or \U$1793 ( \2484 , \2482 , \2483 );
xor \U$1794 ( \2485 , \2406 , \2484 );
not \U$1795 ( \2486 , \2485 );
not \U$1796 ( \2487 , \1587 );
not \U$1797 ( \2488 , RI992c9c8_342);
not \U$1798 ( \2489 , \2488 );
and \U$1799 ( \2490 , \2487 , \2489 );
and \U$1800 ( \2491 , \1593 , RI99244a8_522);
nor \U$1801 ( \2492 , \2490 , \2491 );
nand \U$1802 ( \2493 , \1461 , RI9933b38_262);
and \U$1803 ( \2494 , \1469 , RI99314c8_282);
not \U$1804 ( \2495 , RI99225b8_582);
not \U$1805 ( \2496 , \1487 );
or \U$1806 ( \2497 , \2495 , \2496 );
nand \U$1807 ( \2498 , \1481 , RI99231e8_562);
nand \U$1808 ( \2499 , \2497 , \2498 );
nor \U$1809 ( \2500 , \2494 , \2499 );
and \U$1810 ( \2501 , \2492 , \2493 , \2500 );
and \U$1811 ( \2502 , \2445 , RI9923b48_542);
and \U$1812 ( \2503 , \1557 , RI992a538_382);
and \U$1813 ( \2504 , \1535 , RI992d328_322);
nor \U$1814 ( \2505 , \2502 , \2503 , \2504 );
not \U$1815 ( \2506 , RI9925df8_482);
nor \U$1816 ( \2507 , \1551 , \2506 );
not \U$1817 ( \2508 , RI9926758_462);
nor \U$1818 ( \2509 , \1544 , \2508 );
nor \U$1819 ( \2510 , \2507 , \2509 );
not \U$1820 ( \2511 , \1635 );
not \U$1821 ( \2512 , RI992ae98_362);
not \U$1822 ( \2513 , \2512 );
and \U$1823 ( \2514 , \2511 , \2513 );
and \U$1824 ( \2515 , \1519 , RI9927b08_442);
nor \U$1825 ( \2516 , \2514 , \2515 );
not \U$1826 ( \2517 , RI9928dc8_402);
nor \U$1827 ( \2518 , \2517 , \1497 );
not \U$1828 ( \2519 , RI992f218_302);
nor \U$1829 ( \2520 , \1506 , \2519 );
nor \U$1830 ( \2521 , \2518 , \2520 );
and \U$1831 ( \2522 , \2510 , \2516 , \2521 );
and \U$1832 ( \2523 , \1657 , RI9928468_422);
and \U$1833 ( \2524 , \1710 , RI9924e08_502);
nor \U$1834 ( \2525 , \2523 , \2524 );
nand \U$1835 ( \2526 , \2501 , \2505 , \2522 , \2525 );
not \U$1836 ( \2527 , \2526 );
buf \U$1837 ( \2528 , \1380 );
not \U$1838 ( \2529 , \2528 );
not \U$1839 ( \2530 , \2529 );
or \U$1840 ( \2531 , \2527 , \2530 );
not \U$1841 ( \2532 , \2526 );
nand \U$1842 ( \2533 , \2528 , \2532 );
nand \U$1843 ( \2534 , \2531 , \2533 );
not \U$1844 ( \2535 , \2534 );
and \U$1845 ( \2536 , \1385 , \1386 , \1395 );
not \U$1846 ( \2537 , \2536 );
or \U$1847 ( \2538 , \2535 , \2537 );
not \U$1848 ( \2539 , \1398 );
not \U$1849 ( \2540 , RI9933bb0_261);
nor \U$1850 ( \2541 , \2540 , \1616 );
not \U$1851 ( \2542 , RI9928e40_401);
nor \U$1852 ( \2543 , \2542 , \1497 );
nor \U$1853 ( \2544 , \2541 , \2543 );
not \U$1854 ( \2545 , \1625 );
not \U$1855 ( \2546 , RI9927b80_441);
not \U$1856 ( \2547 , \2546 );
and \U$1857 ( \2548 , \2545 , \2547 );
and \U$1858 ( \2549 , \2288 , RI992f290_301);
nor \U$1859 ( \2550 , \2548 , \2549 );
not \U$1860 ( \2551 , \1629 );
not \U$1861 ( \2552 , RI992d3a0_321);
not \U$1862 ( \2553 , \2552 );
and \U$1863 ( \2554 , \2551 , \2553 );
and \U$1864 ( \2555 , \1636 , RI992af10_361);
nor \U$1865 ( \2556 , \2554 , \2555 );
and \U$1866 ( \2557 , \1469 , RI9931540_281);
and \U$1867 ( \2558 , RI9923260_561, \1481 );
and \U$1868 ( \2559 , \1487 , RI9922630_581);
nor \U$1869 ( \2560 , \2557 , \2558 , \2559 );
nand \U$1870 ( \2561 , \2544 , \2550 , \2556 , \2560 );
not \U$1871 ( \2562 , \1545 );
not \U$1872 ( \2563 , RI99267d0_461);
not \U$1873 ( \2564 , \2563 );
and \U$1874 ( \2565 , \2562 , \2564 );
not \U$1875 ( \2566 , RI9925e70_481);
nor \U$1876 ( \2567 , \2566 , \1551 );
nor \U$1877 ( \2568 , \2565 , \2567 );
and \U$1878 ( \2569 , \1657 , RI99284e0_421);
and \U$1879 ( \2570 , \1659 , RI9925510_501);
nor \U$1880 ( \2571 , \2569 , \2570 );
not \U$1881 ( \2572 , \1587 );
not \U$1882 ( \2573 , RI992ca40_341);
not \U$1883 ( \2574 , \2573 );
and \U$1884 ( \2575 , \2572 , \2574 );
and \U$1885 ( \2576 , \1593 , RI9924520_521);
nor \U$1886 ( \2577 , \2575 , \2576 );
not \U$1887 ( \2578 , RI9923bc0_541);
nor \U$1888 ( \2579 , \2578 , \1565 );
not \U$1889 ( \2580 , RI992a5b0_381);
nor \U$1890 ( \2581 , \2580 , \1668 );
nor \U$1891 ( \2582 , \2579 , \2581 );
nand \U$1892 ( \2583 , \2568 , \2571 , \2577 , \2582 );
or \U$1893 ( \2584 , \2561 , \2583 );
not \U$1894 ( \2585 , \2584 );
or \U$1895 ( \2586 , \2539 , \2585 );
not \U$1896 ( \2587 , \2584 );
nand \U$1897 ( \2588 , \2528 , \2587 );
nand \U$1898 ( \2589 , \2586 , \2588 );
nand \U$1899 ( \2590 , \2589 , \1605 );
nand \U$1900 ( \2591 , \2538 , \2590 );
and \U$1901 ( \2592 , \1715 , RI99266e0_463);
and \U$1902 ( \2593 , \1550 , RI9925d80_483);
nor \U$1903 ( \2594 , \2592 , \2593 );
not \U$1904 ( \2595 , \1526 );
not \U$1905 ( \2596 , RI992ae20_363);
not \U$1906 ( \2597 , \2596 );
and \U$1907 ( \2598 , \2595 , \2597 );
and \U$1908 ( \2599 , \1519 , RI9927040_443);
nor \U$1909 ( \2600 , \2598 , \2599 );
not \U$1910 ( \2601 , \1498 );
not \U$1911 ( \2602 , RI9928d50_403);
nor \U$1912 ( \2603 , \2601 , \2602 );
not \U$1913 ( \2604 , RI992f1a0_303);
nor \U$1914 ( \2605 , \1508 , \2604 );
nor \U$1915 ( \2606 , \2603 , \2605 );
and \U$1916 ( \2607 , \2594 , \2600 , \2606 );
and \U$1917 ( \2608 , \1586 , RI992c950_343);
and \U$1918 ( \2609 , \1593 , RI9924430_523);
nor \U$1919 ( \2610 , \2608 , \2609 );
nand \U$1920 ( \2611 , \1461 , RI9933ac0_263);
and \U$1921 ( \2612 , \1469 , RI9931450_283);
not \U$1922 ( \2613 , RI9922540_583);
not \U$1923 ( \2614 , \1487 );
or \U$1924 ( \2615 , \2613 , \2614 );
not \U$1925 ( \2616 , RI9923170_563);
or \U$1926 ( \2617 , \1643 , \2616 );
nand \U$1927 ( \2618 , \2615 , \2617 );
nor \U$1928 ( \2619 , \2612 , \2618 );
and \U$1929 ( \2620 , \2610 , \2611 , \2619 );
nand \U$1930 ( \2621 , \1564 , RI9923ad0_543);
not \U$1931 ( \2622 , \1668 );
nand \U$1932 ( \2623 , \2622 , RI992a4c0_383);
nand \U$1933 ( \2624 , \1535 , RI992d2b0_323);
nand \U$1934 ( \2625 , \2621 , \2623 , \2624 );
not \U$1935 ( \2626 , RI99283f0_423);
not \U$1936 ( \2627 , \1577 );
or \U$1937 ( \2628 , \2626 , \2627 );
nand \U$1938 ( \2629 , \1710 , RI9924d90_503);
nand \U$1939 ( \2630 , \2628 , \2629 );
nor \U$1940 ( \2631 , \2625 , \2630 );
nand \U$1941 ( \2632 , \2607 , \2620 , \2631 );
not \U$1942 ( \2633 , \2632 );
not \U$1943 ( \2634 , \2633 );
not \U$1944 ( \2635 , \2634 );
and \U$1945 ( \2636 , \1610 , \2635 );
not \U$1946 ( \2637 , \1614 );
and \U$1947 ( \2638 , \2637 , \2634 );
nor \U$1948 ( \2639 , \2636 , \2638 );
and \U$1949 ( \2640 , \1612 , \2639 );
or \U$1950 ( \2641 , \2591 , \2640 );
not \U$1951 ( \2642 , \1964 );
xor \U$1952 ( \2643 , \1951 , \1912 );
not \U$1953 ( \2644 , \2643 );
or \U$1954 ( \2645 , \2642 , \2644 );
not \U$1955 ( \2646 , \1951 );
not \U$1956 ( \2647 , \2149 );
or \U$1957 ( \2648 , \2646 , \2647 );
nand \U$1958 ( \2649 , \2148 , \1872 );
nand \U$1959 ( \2650 , \2648 , \2649 );
nand \U$1960 ( \2651 , \2650 , \1949 );
nand \U$1961 ( \2652 , \2645 , \2651 );
not \U$1962 ( \2653 , \1975 );
and \U$1963 ( \2654 , \1967 , \1823 );
not \U$1964 ( \2655 , \1967 );
and \U$1965 ( \2656 , \2655 , \1824 );
nor \U$1966 ( \2657 , \2654 , \2656 );
not \U$1967 ( \2658 , \2657 );
or \U$1968 ( \2659 , \2653 , \2658 );
and \U$1969 ( \2660 , \1729 , \1945 );
not \U$1970 ( \2661 , \1729 );
and \U$1971 ( \2662 , \2661 , \1967 );
or \U$1972 ( \2663 , \2660 , \2662 );
not \U$1973 ( \2664 , \2663 );
or \U$1974 ( \2665 , \2664 , \1974 );
nand \U$1975 ( \2666 , \2659 , \2665 );
xor \U$1976 ( \2667 , \2652 , \2666 );
not \U$1977 ( \2668 , \2270 );
not \U$1978 ( \2669 , \1915 );
or \U$1979 ( \2670 , \2668 , \2669 );
not \U$1980 ( \2671 , \2270 );
nand \U$1981 ( \2672 , \1914 , \2671 );
nand \U$1982 ( \2673 , \2670 , \2672 );
not \U$1983 ( \2674 , \2673 );
not \U$1984 ( \2675 , \1878 );
or \U$1985 ( \2676 , \2674 , \2675 );
and \U$1986 ( \2677 , \2076 , \1914 );
not \U$1987 ( \2678 , \2076 );
and \U$1988 ( \2679 , \2678 , \1915 );
nor \U$1989 ( \2680 , \2677 , \2679 );
nand \U$1990 ( \2681 , \2680 , \1929 );
nand \U$1991 ( \2682 , \2676 , \2681 );
not \U$1992 ( \2683 , \2682 );
not \U$1993 ( \2684 , \1975 );
xor \U$1994 ( \2685 , \1967 , \1912 );
not \U$1995 ( \2686 , \2685 );
or \U$1996 ( \2687 , \2684 , \2686 );
nand \U$1997 ( \2688 , \2657 , \1973 );
nand \U$1998 ( \2689 , \2687 , \2688 );
not \U$1999 ( \2690 , \1949 );
not \U$2000 ( \2691 , \1951 );
not \U$2001 ( \2692 , \2080 );
or \U$2002 ( \2693 , \2691 , \2692 );
nand \U$2003 ( \2694 , \2076 , \1872 );
nand \U$2004 ( \2695 , \2693 , \2694 );
not \U$2005 ( \2696 , \2695 );
or \U$2006 ( \2697 , \2690 , \2696 );
nand \U$2007 ( \2698 , \2650 , \1964 );
nand \U$2008 ( \2699 , \2697 , \2698 );
nand \U$2009 ( \2700 , \2689 , \2699 );
nand \U$2010 ( \2701 , \2683 , \2700 );
and \U$2011 ( \2702 , \2667 , \2701 );
nor \U$2012 ( \2703 , \2683 , \2700 );
nor \U$2013 ( \2704 , \2702 , \2703 );
not \U$2014 ( \2705 , \2704 );
nand \U$2015 ( \2706 , \2641 , \2705 );
nand \U$2016 ( \2707 , \2591 , \2640 );
and \U$2017 ( \2708 , \2706 , \2707 );
not \U$2018 ( \2709 , \2708 );
not \U$2019 ( \2710 , \2709 );
not \U$2020 ( \2711 , \1878 );
not \U$2021 ( \2712 , \2680 );
or \U$2022 ( \2713 , \2711 , \2712 );
not \U$2023 ( \2714 , \2148 );
not \U$2024 ( \2715 , \1915 );
or \U$2025 ( \2716 , \2714 , \2715 );
nand \U$2026 ( \2717 , \1914 , \2149 );
nand \U$2027 ( \2718 , \2716 , \2717 );
nand \U$2028 ( \2719 , \2718 , \1929 );
nand \U$2029 ( \2720 , \2713 , \2719 );
and \U$2030 ( \2721 , \2652 , \2666 );
xor \U$2031 ( \2722 , \2720 , \2721 );
not \U$2032 ( \2723 , \1964 );
not \U$2033 ( \2724 , \1956 );
or \U$2034 ( \2725 , \2723 , \2724 );
nand \U$2035 ( \2726 , \2643 , \1949 );
nand \U$2036 ( \2727 , \2725 , \2726 );
not \U$2037 ( \2728 , \1973 );
not \U$2038 ( \2729 , \1981 );
or \U$2039 ( \2730 , \2728 , \2729 );
nand \U$2040 ( \2731 , \2663 , \1975 );
nand \U$2041 ( \2732 , \2730 , \2731 );
xor \U$2042 ( \2733 , \2727 , \2732 );
and \U$2043 ( \2734 , \2722 , \2733 );
and \U$2044 ( \2735 , \2720 , \2721 );
or \U$2045 ( \2736 , \2734 , \2735 );
and \U$2046 ( \2737 , \2532 , \1610 );
not \U$2047 ( \2738 , \2532 );
and \U$2048 ( \2739 , \2738 , \2637 );
nor \U$2049 ( \2740 , \2737 , \2739 );
and \U$2050 ( \2741 , \1612 , \2740 );
xor \U$2051 ( \2742 , \2736 , \2741 );
not \U$2052 ( \2743 , \2589 );
not \U$2053 ( \2744 , \1396 );
or \U$2054 ( \2745 , \2743 , \2744 );
not \U$2055 ( \2746 , \1395 );
nand \U$2056 ( \2747 , \1461 , RI9933c28_260);
and \U$2057 ( \2748 , \1471 , RI99315b8_280);
not \U$2058 ( \2749 , RI99226a8_580);
not \U$2059 ( \2750 , \1487 );
or \U$2060 ( \2751 , \2749 , \2750 );
nand \U$2061 ( \2752 , \1481 , RI99232d8_560);
nand \U$2062 ( \2753 , \2751 , \2752 );
nor \U$2063 ( \2754 , \2748 , \2753 );
nand \U$2064 ( \2755 , \1499 , RI9928eb8_400);
nand \U$2065 ( \2756 , \2747 , \2754 , \2755 );
not \U$2066 ( \2757 , \1508 );
not \U$2067 ( \2758 , RI992f308_300);
not \U$2068 ( \2759 , \2758 );
and \U$2069 ( \2760 , \2757 , \2759 );
and \U$2070 ( \2761 , \1626 , RI9927bf8_440);
nor \U$2071 ( \2762 , \2760 , \2761 );
not \U$2072 ( \2763 , \1524 );
not \U$2073 ( \2764 , RI992af88_360);
not \U$2074 ( \2765 , \2764 );
and \U$2075 ( \2766 , \2763 , \2765 );
and \U$2076 ( \2767 , \1535 , RI992d418_320);
nor \U$2077 ( \2768 , \2766 , \2767 );
nand \U$2078 ( \2769 , \2762 , \2768 );
nor \U$2079 ( \2770 , \2756 , \2769 );
not \U$2080 ( \2771 , RI9925588_500);
or \U$2081 ( \2772 , \1572 , \2771 );
not \U$2082 ( \2773 , RI9928558_420);
or \U$2083 ( \2774 , \1578 , \2773 );
not \U$2084 ( \2775 , \1587 );
not \U$2085 ( \2776 , RI992cab8_340);
not \U$2086 ( \2777 , \2776 );
and \U$2087 ( \2778 , \2775 , \2777 );
and \U$2088 ( \2779 , \1593 , RI9924598_520);
nor \U$2089 ( \2780 , \2778 , \2779 );
nand \U$2090 ( \2781 , \2772 , \2774 , \2780 );
not \U$2091 ( \2782 , \1551 );
not \U$2092 ( \2783 , RI9925ee8_480);
not \U$2093 ( \2784 , \2783 );
and \U$2094 ( \2785 , \2782 , \2784 );
not \U$2095 ( \2786 , RI9926848_460);
nor \U$2096 ( \2787 , \1545 , \2786 );
nor \U$2097 ( \2788 , \2785 , \2787 );
and \U$2098 ( \2789 , \2622 , RI992a628_380);
not \U$2099 ( \2790 , RI9923c38_540);
nor \U$2100 ( \2791 , \2160 , \2790 );
nor \U$2101 ( \2792 , \2789 , \2791 );
nand \U$2102 ( \2793 , \2788 , \2792 );
nor \U$2103 ( \2794 , \2781 , \2793 );
nand \U$2104 ( \2795 , \2770 , \2794 );
not \U$2105 ( \2796 , \2795 );
not \U$2106 ( \2797 , \2796 );
not \U$2107 ( \2798 , \2797 );
not \U$2108 ( \2799 , \2529 );
or \U$2109 ( \2800 , \2798 , \2799 );
not \U$2110 ( \2801 , \1381 );
nand \U$2111 ( \2802 , \2801 , \2796 );
nand \U$2112 ( \2803 , \2800 , \2802 );
nand \U$2113 ( \2804 , \2746 , \2803 );
nand \U$2114 ( \2805 , \2745 , \2804 );
xor \U$2115 ( \2806 , \2742 , \2805 );
not \U$2116 ( \2807 , \2806 );
or \U$2117 ( \2808 , \2710 , \2807 );
or \U$2118 ( \2809 , \2709 , \2806 );
not \U$2119 ( \2810 , \2414 );
not \U$2120 ( \2811 , \2398 );
not \U$2121 ( \2812 , \2029 );
or \U$2122 ( \2813 , \2811 , \2812 );
not \U$2123 ( \2814 , \2029 );
nand \U$2124 ( \2815 , \2814 , \2397 );
nand \U$2125 ( \2816 , \2813 , \2815 );
not \U$2126 ( \2817 , \2816 );
or \U$2127 ( \2818 , \2810 , \2817 );
not \U$2128 ( \2819 , \2029 );
not \U$2129 ( \2820 , \2199 );
or \U$2130 ( \2821 , \2819 , \2820 );
not \U$2131 ( \2822 , \2199 );
nand \U$2132 ( \2823 , \2079 , \2822 );
nand \U$2133 ( \2824 , \2821 , \2823 );
nand \U$2134 ( \2825 , \2824 , \2157 );
nand \U$2135 ( \2826 , \2818 , \2825 );
not \U$2136 ( \2827 , \2826 );
and \U$2137 ( \2828 , \2332 , \1744 );
not \U$2138 ( \2829 , \2332 );
and \U$2139 ( \2830 , \2829 , \2202 );
nor \U$2140 ( \2831 , \2828 , \2830 );
not \U$2141 ( \2832 , \2831 );
not \U$2142 ( \2833 , \2472 );
or \U$2143 ( \2834 , \2832 , \2833 );
or \U$2144 ( \2835 , \2202 , \2457 );
or \U$2145 ( \2836 , \1744 , \2461 );
nand \U$2146 ( \2837 , \2835 , \2836 );
nand \U$2147 ( \2838 , \2479 , \2837 );
nand \U$2148 ( \2839 , \2834 , \2838 );
not \U$2149 ( \2840 , \2839 );
nand \U$2150 ( \2841 , \2827 , \2840 );
not \U$2151 ( \2842 , \2584 );
not \U$2152 ( \2843 , \1394 );
or \U$2153 ( \2844 , \2842 , \2843 );
nand \U$2154 ( \2845 , \1393 , \2587 );
nand \U$2155 ( \2846 , \2844 , \2845 );
not \U$2156 ( \2847 , \2846 );
not \U$2157 ( \2848 , \1764 );
or \U$2158 ( \2849 , \2847 , \2848 );
not \U$2159 ( \2850 , \2797 );
not \U$2160 ( \2851 , \1394 );
or \U$2161 ( \2852 , \2850 , \2851 );
nand \U$2162 ( \2853 , \1393 , \2796 );
nand \U$2163 ( \2854 , \2852 , \2853 );
nand \U$2164 ( \2855 , \2854 , \1758 );
nand \U$2165 ( \2856 , \2849 , \2855 );
and \U$2166 ( \2857 , \2841 , \2856 );
and \U$2167 ( \2858 , \2839 , \2826 );
nor \U$2168 ( \2859 , \2857 , \2858 );
not \U$2169 ( \2860 , \2859 );
not \U$2170 ( \2861 , \2860 );
not \U$2171 ( \2862 , \2854 );
not \U$2172 ( \2863 , \1764 );
or \U$2173 ( \2864 , \2862 , \2863 );
nand \U$2174 ( \2865 , \2463 , \1758 );
nand \U$2175 ( \2866 , \2864 , \2865 );
not \U$2176 ( \2867 , \2866 );
not \U$2177 ( \2868 , \2414 );
not \U$2178 ( \2869 , \2824 );
or \U$2179 ( \2870 , \2868 , \2869 );
nand \U$2180 ( \2871 , \2412 , \2157 );
nand \U$2181 ( \2872 , \2870 , \2871 );
not \U$2182 ( \2873 , \2872 );
not \U$2183 ( \2874 , \2873 );
or \U$2184 ( \2875 , \2867 , \2874 );
or \U$2185 ( \2876 , \2873 , \2866 );
nand \U$2186 ( \2877 , \2875 , \2876 );
not \U$2187 ( \2878 , \2472 );
not \U$2188 ( \2879 , \2878 );
not \U$2189 ( \2880 , \2477 );
and \U$2190 ( \2881 , \2879 , \2880 );
and \U$2191 ( \2882 , \2479 , \2831 );
nor \U$2192 ( \2883 , \2881 , \2882 );
and \U$2193 ( \2884 , \2877 , \2883 );
not \U$2194 ( \2885 , \2877 );
not \U$2195 ( \2886 , \2883 );
and \U$2196 ( \2887 , \2885 , \2886 );
nor \U$2197 ( \2888 , \2884 , \2887 );
not \U$2198 ( \2889 , \2888 );
not \U$2199 ( \2890 , \2889 );
or \U$2200 ( \2891 , \2861 , \2890 );
not \U$2201 ( \2892 , \2859 );
not \U$2202 ( \2893 , \2888 );
or \U$2203 ( \2894 , \2892 , \2893 );
xor \U$2204 ( \2895 , \2720 , \2721 );
xor \U$2205 ( \2896 , \2895 , \2733 );
nand \U$2206 ( \2897 , \2894 , \2896 );
nand \U$2207 ( \2898 , \2891 , \2897 );
nand \U$2208 ( \2899 , \2809 , \2898 );
nand \U$2209 ( \2900 , \2808 , \2899 );
not \U$2210 ( \2901 , \2900 );
or \U$2211 ( \2902 , \2486 , \2901 );
or \U$2212 ( \2903 , \2900 , \2485 );
xor \U$2213 ( \2904 , \2736 , \2741 );
and \U$2214 ( \2905 , \2904 , \2805 );
and \U$2215 ( \2906 , \2736 , \2741 );
or \U$2216 ( \2907 , \2905 , \2906 );
not \U$2217 ( \2908 , \2718 );
not \U$2218 ( \2909 , \1878 );
or \U$2219 ( \2910 , \2908 , \2909 );
nand \U$2220 ( \2911 , \1919 , \1929 );
nand \U$2221 ( \2912 , \2910 , \2911 );
and \U$2222 ( \2913 , \2727 , \2732 );
xor \U$2223 ( \2914 , \2912 , \2913 );
xor \U$2224 ( \2915 , \1966 , \1990 );
and \U$2225 ( \2916 , \2914 , \2915 );
and \U$2226 ( \2917 , \2912 , \2913 );
or \U$2227 ( \2918 , \2916 , \2917 );
not \U$2228 ( \2919 , \1610 );
and \U$2229 ( \2920 , \2584 , \2919 );
not \U$2230 ( \2921 , \2584 );
and \U$2231 ( \2922 , \2921 , \1610 );
nor \U$2232 ( \2923 , \2920 , \2922 );
and \U$2233 ( \2924 , \1612 , \2923 );
xor \U$2234 ( \2925 , \2918 , \2924 );
not \U$2235 ( \2926 , \2803 );
not \U$2236 ( \2927 , \1396 );
or \U$2237 ( \2928 , \2926 , \2927 );
not \U$2238 ( \2929 , \1395 );
not \U$2239 ( \2930 , \2457 );
not \U$2240 ( \2931 , \2801 );
not \U$2241 ( \2932 , \2931 );
or \U$2242 ( \2933 , \2930 , \2932 );
nand \U$2243 ( \2934 , \2801 , \2461 );
nand \U$2244 ( \2935 , \2933 , \2934 );
nand \U$2245 ( \2936 , \2929 , \2935 );
nand \U$2246 ( \2937 , \2928 , \2936 );
xor \U$2247 ( \2938 , \2925 , \2937 );
xor \U$2248 ( \2939 , \2907 , \2938 );
xor \U$2249 ( \2940 , \2912 , \2913 );
xor \U$2250 ( \2941 , \2940 , \2915 );
not \U$2251 ( \2942 , \2886 );
not \U$2252 ( \2943 , \2872 );
or \U$2253 ( \2944 , \2942 , \2943 );
not \U$2254 ( \2945 , \2873 );
not \U$2255 ( \2946 , \2883 );
or \U$2256 ( \2947 , \2945 , \2946 );
nand \U$2257 ( \2948 , \2947 , \2866 );
nand \U$2258 ( \2949 , \2944 , \2948 );
xor \U$2259 ( \2950 , \2941 , \2949 );
xor \U$2260 ( \2951 , \2418 , \2469 );
xor \U$2261 ( \2952 , \2951 , \2481 );
and \U$2262 ( \2953 , \2950 , \2952 );
and \U$2263 ( \2954 , \2941 , \2949 );
or \U$2264 ( \2955 , \2953 , \2954 );
xor \U$2265 ( \2956 , \2939 , \2955 );
nand \U$2266 ( \2957 , \2903 , \2956 );
nand \U$2267 ( \2958 , \2902 , \2957 );
not \U$2268 ( \2959 , \2958 );
or \U$2269 ( \2960 , \2277 , \2159 );
and \U$2270 ( \2961 , \2960 , \2404 );
and \U$2271 ( \2962 , \2277 , \2159 );
nor \U$2272 ( \2963 , \2961 , \2962 );
not \U$2273 ( \2964 , \2963 );
not \U$2274 ( \2965 , \1997 );
nand \U$2275 ( \2966 , \2965 , \2007 );
not \U$2276 ( \2967 , \1964 );
and \U$2277 ( \2968 , \1872 , \1599 );
not \U$2278 ( \2969 , \1872 );
and \U$2279 ( \2970 , \2969 , \1598 );
nor \U$2280 ( \2971 , \2968 , \2970 );
not \U$2281 ( \2972 , \2971 );
or \U$2282 ( \2973 , \2967 , \2972 );
not \U$2283 ( \2974 , \2005 );
or \U$2284 ( \2975 , \2974 , \1948 );
nand \U$2285 ( \2976 , \2973 , \2975 );
xor \U$2286 ( \2977 , \2966 , \2976 );
not \U$2287 ( \2978 , \2977 );
not \U$2288 ( \2979 , \2156 );
not \U$2289 ( \2980 , \2414 );
or \U$2290 ( \2981 , \2979 , \2980 );
not \U$2291 ( \2982 , \1913 );
not \U$2292 ( \2983 , \2982 );
not \U$2293 ( \2984 , \2029 );
or \U$2294 ( \2985 , \2983 , \2984 );
nand \U$2295 ( \2986 , \2079 , \1913 );
nand \U$2296 ( \2987 , \2985 , \2986 );
nand \U$2297 ( \2988 , \2987 , \2157 );
nand \U$2298 ( \2989 , \2981 , \2988 );
not \U$2299 ( \2990 , \2989 );
and \U$2300 ( \2991 , \2978 , \2990 );
and \U$2301 ( \2992 , \2977 , \2989 );
nor \U$2302 ( \2993 , \2991 , \2992 );
not \U$2303 ( \2994 , \2993 );
xor \U$2304 ( \2995 , \2964 , \2994 );
not \U$2305 ( \2996 , \1945 );
not \U$2306 ( \2997 , \1927 );
not \U$2307 ( \2998 , \1878 );
or \U$2308 ( \2999 , \2997 , \2998 );
and \U$2309 ( \3000 , \1731 , \1922 );
not \U$2310 ( \3001 , \1731 );
and \U$2311 ( \3002 , \3001 , \1925 );
nor \U$2312 ( \3003 , \3000 , \3002 );
nand \U$2313 ( \3004 , \3003 , \1929 );
nand \U$2314 ( \3005 , \2999 , \3004 );
not \U$2315 ( \3006 , \3005 );
or \U$2316 ( \3007 , \2996 , \3006 );
not \U$2317 ( \3008 , \3005 );
nand \U$2318 ( \3009 , \3008 , \1967 );
nand \U$2319 ( \3010 , \3007 , \3009 );
not \U$2320 ( \3011 , \2402 );
not \U$2321 ( \3012 , \2465 );
or \U$2322 ( \3013 , \3011 , \3012 );
not \U$2323 ( \3014 , \2334 );
and \U$2324 ( \3015 , \2199 , \3014 );
not \U$2325 ( \3016 , \2199 );
and \U$2326 ( \3017 , \3016 , \1784 );
nor \U$2327 ( \3018 , \3015 , \3017 );
nand \U$2328 ( \3019 , \3018 , \1758 );
nand \U$2329 ( \3020 , \3013 , \3019 );
xor \U$2330 ( \3021 , \3010 , \3020 );
not \U$2331 ( \3022 , \2275 );
not \U$2332 ( \3023 , \2479 );
or \U$2333 ( \3024 , \3022 , \3023 );
buf \U$2334 ( \3025 , \2076 );
and \U$2335 ( \3026 , \3025 , \1744 );
not \U$2336 ( \3027 , \3025 );
and \U$2337 ( \3028 , \3027 , \2202 );
nor \U$2338 ( \3029 , \3026 , \3028 );
nand \U$2339 ( \3030 , \2472 , \3029 );
nand \U$2340 ( \3031 , \3024 , \3030 );
xor \U$2341 ( \3032 , \3021 , \3031 );
buf \U$2342 ( \3033 , \3032 );
xnor \U$2343 ( \3034 , \2995 , \3033 );
not \U$2344 ( \3035 , \3034 );
xor \U$2345 ( \3036 , \2918 , \2924 );
and \U$2346 ( \3037 , \3036 , \2937 );
and \U$2347 ( \3038 , \2918 , \2924 );
or \U$2348 ( \3039 , \3037 , \3038 );
xor \U$2349 ( \3040 , \1931 , \1991 );
and \U$2350 ( \3041 , \3040 , \2011 );
and \U$2351 ( \3042 , \1931 , \1991 );
or \U$2352 ( \3043 , \3041 , \3042 );
and \U$2353 ( \3044 , \2797 , \2637 );
not \U$2354 ( \3045 , \2797 );
and \U$2355 ( \3046 , \3045 , \1610 );
nor \U$2356 ( \3047 , \3044 , \3046 );
and \U$2357 ( \3048 , \1612 , \3047 );
xor \U$2358 ( \3049 , \3043 , \3048 );
not \U$2359 ( \3050 , \2935 );
not \U$2360 ( \3051 , \1396 );
or \U$2361 ( \3052 , \3050 , \3051 );
not \U$2362 ( \3053 , \1395 );
not \U$2363 ( \3054 , \2332 );
not \U$2364 ( \3055 , \2529 );
or \U$2365 ( \3056 , \3054 , \3055 );
not \U$2366 ( \3057 , \2931 );
nand \U$2367 ( \3058 , \3057 , \2338 );
nand \U$2368 ( \3059 , \3056 , \3058 );
nand \U$2369 ( \3060 , \3053 , \3059 );
nand \U$2370 ( \3061 , \3052 , \3060 );
xor \U$2371 ( \3062 , \3049 , \3061 );
xor \U$2372 ( \3063 , \3039 , \3062 );
xor \U$2373 ( \3064 , \2012 , \2405 );
and \U$2374 ( \3065 , \3064 , \2484 );
and \U$2375 ( \3066 , \2012 , \2405 );
or \U$2376 ( \3067 , \3065 , \3066 );
xor \U$2377 ( \3068 , \3063 , \3067 );
not \U$2378 ( \3069 , \3068 );
or \U$2379 ( \3070 , \3035 , \3069 );
or \U$2380 ( \3071 , \3034 , \3068 );
nand \U$2381 ( \3072 , \3070 , \3071 );
xor \U$2382 ( \3073 , \2907 , \2938 );
and \U$2383 ( \3074 , \3073 , \2955 );
and \U$2384 ( \3075 , \2907 , \2938 );
or \U$2385 ( \3076 , \3074 , \3075 );
not \U$2386 ( \3077 , \3076 );
and \U$2387 ( \3078 , \3072 , \3077 );
not \U$2388 ( \3079 , \3072 );
and \U$2389 ( \3080 , \3079 , \3076 );
nor \U$2390 ( \3081 , \3078 , \3080 );
nand \U$2391 ( \3082 , \2959 , \3081 );
xor \U$2392 ( \3083 , \2941 , \2949 );
xor \U$2393 ( \3084 , \3083 , \2952 );
not \U$2394 ( \3085 , \3084 );
not \U$2395 ( \3086 , \2634 );
not \U$2396 ( \3087 , \2529 );
or \U$2397 ( \3088 , \3086 , \3087 );
nand \U$2398 ( \3089 , \2801 , \2635 );
nand \U$2399 ( \3090 , \3088 , \3089 );
not \U$2400 ( \3091 , \3090 );
not \U$2401 ( \3092 , \2536 );
or \U$2402 ( \3093 , \3091 , \3092 );
nand \U$2403 ( \3094 , \2534 , \1605 );
nand \U$2404 ( \3095 , \3093 , \3094 );
not \U$2405 ( \3096 , \3095 );
not \U$2406 ( \3097 , \2374 );
not \U$2407 ( \3098 , RI9926fc8_444);
not \U$2408 ( \3099 , \3098 );
and \U$2409 ( \3100 , \3097 , \3099 );
and \U$2410 ( \3101 , \1636 , RI992ada8_364);
nor \U$2411 ( \3102 , \3100 , \3101 );
not \U$2412 ( \3103 , \1551 );
not \U$2413 ( \3104 , RI9925d08_484);
not \U$2414 ( \3105 , \3104 );
and \U$2415 ( \3106 , \3103 , \3105 );
not \U$2416 ( \3107 , RI9926668_464);
nor \U$2417 ( \3108 , \3107 , \1545 );
nor \U$2418 ( \3109 , \3106 , \3108 );
and \U$2419 ( \3110 , \2288 , RI992f128_304);
and \U$2420 ( \3111 , \1498 , RI9928cd8_404);
nor \U$2421 ( \3112 , \3110 , \3111 );
nand \U$2422 ( \3113 , \3102 , \3109 , \3112 );
not \U$2423 ( \3114 , \1668 );
not \U$2424 ( \3115 , RI992a448_384);
not \U$2425 ( \3116 , \3115 );
and \U$2426 ( \3117 , \3114 , \3116 );
not \U$2427 ( \3118 , RI9923a58_544);
nor \U$2428 ( \3119 , \2160 , \3118 );
nor \U$2429 ( \3120 , \3117 , \3119 );
and \U$2430 ( \3121 , \1657 , RI9928378_424);
and \U$2431 ( \3122 , \1710 , RI9924d18_504);
nor \U$2432 ( \3123 , \3121 , \3122 );
nand \U$2433 ( \3124 , \1535 , RI992d238_324);
nand \U$2434 ( \3125 , \3120 , \3123 , \3124 );
nor \U$2435 ( \3126 , \3113 , \3125 );
not \U$2436 ( \3127 , \1587 );
not \U$2437 ( \3128 , RI992c8d8_344);
not \U$2438 ( \3129 , \3128 );
and \U$2439 ( \3130 , \3127 , \3129 );
and \U$2440 ( \3131 , \1593 , RI99243b8_524);
nor \U$2441 ( \3132 , \3130 , \3131 );
and \U$2442 ( \3133 , \1469 , RI99313d8_284);
not \U$2443 ( \3134 , RI99224c8_584);
not \U$2444 ( \3135 , \1487 );
or \U$2445 ( \3136 , \3134 , \3135 );
nand \U$2446 ( \3137 , \1481 , RI99230f8_564);
nand \U$2447 ( \3138 , \3136 , \3137 );
nor \U$2448 ( \3139 , \3133 , \3138 );
nand \U$2449 ( \3140 , \3132 , \3139 );
and \U$2450 ( \3141 , \1461 , RI9933a48_264);
nor \U$2451 ( \3142 , \3140 , \3141 );
nand \U$2452 ( \3143 , \3126 , \3142 );
not \U$2453 ( \3144 , \3143 );
not \U$2454 ( \3145 , \3144 );
buf \U$2455 ( \3146 , \3145 );
and \U$2456 ( \3147 , \3146 , \2919 );
not \U$2457 ( \3148 , \3146 );
and \U$2458 ( \3149 , \3148 , \1610 );
nor \U$2459 ( \3150 , \3147 , \3149 );
and \U$2460 ( \3151 , \1612 , \3150 );
not \U$2461 ( \3152 , \3151 );
or \U$2462 ( \3153 , \3096 , \3152 );
or \U$2463 ( \3154 , \3095 , \3151 );
not \U$2464 ( \3155 , \2199 );
not \U$2465 ( \3156 , \1915 );
or \U$2466 ( \3157 , \3155 , \3156 );
nand \U$2467 ( \3158 , \1914 , \2822 );
nand \U$2468 ( \3159 , \3157 , \3158 );
not \U$2469 ( \3160 , \3159 );
not \U$2470 ( \3161 , \1878 );
or \U$2471 ( \3162 , \3160 , \3161 );
nand \U$2472 ( \3163 , \2673 , \1929 );
nand \U$2473 ( \3164 , \3162 , \3163 );
not \U$2474 ( \3165 , \1949 );
xor \U$2475 ( \3166 , \1951 , \2270 );
not \U$2476 ( \3167 , \3166 );
or \U$2477 ( \3168 , \3165 , \3167 );
nand \U$2478 ( \3169 , \2695 , \1964 );
nand \U$2479 ( \3170 , \3168 , \3169 );
not \U$2480 ( \3171 , \1973 );
not \U$2481 ( \3172 , \2685 );
or \U$2482 ( \3173 , \3171 , \3172 );
and \U$2483 ( \3174 , \2148 , \1945 );
not \U$2484 ( \3175 , \2148 );
and \U$2485 ( \3176 , \3175 , \1967 );
or \U$2486 ( \3177 , \3174 , \3176 );
nand \U$2487 ( \3178 , \3177 , \1975 );
nand \U$2488 ( \3179 , \3173 , \3178 );
and \U$2489 ( \3180 , \3170 , \3179 );
xor \U$2490 ( \3181 , \3164 , \3180 );
xor \U$2491 ( \3182 , \2699 , \2689 );
and \U$2492 ( \3183 , \3181 , \3182 );
and \U$2493 ( \3184 , \3164 , \3180 );
or \U$2494 ( \3185 , \3183 , \3184 );
nand \U$2495 ( \3186 , \3154 , \3185 );
nand \U$2496 ( \3187 , \3153 , \3186 );
not \U$2497 ( \3188 , \3187 );
not \U$2498 ( \3189 , \2640 );
not \U$2499 ( \3190 , \2704 );
and \U$2500 ( \3191 , \3189 , \3190 );
and \U$2501 ( \3192 , \2640 , \2704 );
nor \U$2502 ( \3193 , \3191 , \3192 );
not \U$2503 ( \3194 , \2591 );
and \U$2504 ( \3195 , \3193 , \3194 );
not \U$2505 ( \3196 , \3193 );
and \U$2506 ( \3197 , \3196 , \2591 );
nor \U$2507 ( \3198 , \3195 , \3197 );
not \U$2508 ( \3199 , \3198 );
or \U$2509 ( \3200 , \3188 , \3199 );
or \U$2510 ( \3201 , \3187 , \3198 );
xor \U$2511 ( \3202 , \2700 , \2682 );
xnor \U$2512 ( \3203 , \3202 , \2667 );
not \U$2513 ( \3204 , \2526 );
not \U$2514 ( \3205 , \1394 );
or \U$2515 ( \3206 , \3204 , \3205 );
nand \U$2516 ( \3207 , \1393 , \2532 );
nand \U$2517 ( \3208 , \3206 , \3207 );
not \U$2518 ( \3209 , \3208 );
not \U$2519 ( \3210 , \1764 );
or \U$2520 ( \3211 , \3209 , \3210 );
nand \U$2521 ( \3212 , \2846 , \1758 );
nand \U$2522 ( \3213 , \3211 , \3212 );
not \U$2523 ( \3214 , \2414 );
not \U$2524 ( \3215 , \2332 );
not \U$2525 ( \3216 , \2408 );
or \U$2526 ( \3217 , \3215 , \3216 );
nand \U$2527 ( \3218 , \2079 , \2338 );
nand \U$2528 ( \3219 , \3217 , \3218 );
not \U$2529 ( \3220 , \3219 );
or \U$2530 ( \3221 , \3214 , \3220 );
nand \U$2531 ( \3222 , \2816 , \2157 );
nand \U$2532 ( \3223 , \3221 , \3222 );
xor \U$2533 ( \3224 , \3213 , \3223 );
not \U$2534 ( \3225 , \2837 );
not \U$2535 ( \3226 , \2472 );
or \U$2536 ( \3227 , \3225 , \3226 );
and \U$2537 ( \3228 , \2797 , \1744 );
not \U$2538 ( \3229 , \2797 );
and \U$2539 ( \3230 , \3229 , \2202 );
nor \U$2540 ( \3231 , \3228 , \3230 );
nand \U$2541 ( \3232 , \2479 , \3231 );
nand \U$2542 ( \3233 , \3227 , \3232 );
and \U$2543 ( \3234 , \3224 , \3233 );
and \U$2544 ( \3235 , \3213 , \3223 );
or \U$2545 ( \3236 , \3234 , \3235 );
xor \U$2546 ( \3237 , \3203 , \3236 );
xor \U$2547 ( \3238 , \2826 , \2856 );
and \U$2548 ( \3239 , \3238 , \2839 );
not \U$2549 ( \3240 , \3238 );
and \U$2550 ( \3241 , \3240 , \2840 );
nor \U$2551 ( \3242 , \3239 , \3241 );
and \U$2552 ( \3243 , \3237 , \3242 );
and \U$2553 ( \3244 , \3203 , \3236 );
or \U$2554 ( \3245 , \3243 , \3244 );
nand \U$2555 ( \3246 , \3201 , \3245 );
nand \U$2556 ( \3247 , \3200 , \3246 );
not \U$2557 ( \3248 , \3247 );
or \U$2558 ( \3249 , \3085 , \3248 );
or \U$2559 ( \3250 , \3084 , \3247 );
xor \U$2560 ( \3251 , \2708 , \2806 );
xnor \U$2561 ( \3252 , \3251 , \2898 );
nand \U$2562 ( \3253 , \3250 , \3252 );
nand \U$2563 ( \3254 , \3249 , \3253 );
not \U$2564 ( \3255 , \3254 );
xor \U$2565 ( \3256 , \2485 , \2900 );
xnor \U$2566 ( \3257 , \3256 , \2956 );
nand \U$2567 ( \3258 , \3255 , \3257 );
and \U$2568 ( \3259 , \3082 , \3258 );
not \U$2569 ( \3260 , \3003 );
not \U$2570 ( \3261 , \1878 );
or \U$2571 ( \3262 , \3260 , \3261 );
and \U$2572 ( \3263 , \1925 , \1677 );
not \U$2573 ( \3264 , \1925 );
and \U$2574 ( \3265 , \3264 , \1678 );
nor \U$2575 ( \3266 , \3263 , \3265 );
nand \U$2576 ( \3267 , \3266 , \1929 );
nand \U$2577 ( \3268 , \3262 , \3267 );
not \U$2578 ( \3269 , \3268 );
not \U$2579 ( \3270 , \2971 );
or \U$2580 ( \3271 , \3270 , \1948 );
or \U$2581 ( \3272 , \1963 , \1872 );
nand \U$2582 ( \3273 , \3271 , \3272 );
xor \U$2583 ( \3274 , \3269 , \3273 );
and \U$2584 ( \3275 , \3274 , \3009 );
and \U$2585 ( \3276 , \3269 , \3273 );
or \U$2586 ( \3277 , \3275 , \3276 );
not \U$2587 ( \3278 , \3018 );
not \U$2588 ( \3279 , \1766 );
or \U$2589 ( \3280 , \3278 , \3279 );
and \U$2590 ( \3281 , \2334 , \2271 );
not \U$2591 ( \3282 , \2334 );
and \U$2592 ( \3283 , \3282 , \2273 );
or \U$2593 ( \3284 , \3281 , \3283 );
nand \U$2594 ( \3285 , \3284 , \1758 );
nand \U$2595 ( \3286 , \3280 , \3285 );
not \U$2596 ( \3287 , \2987 );
not \U$2597 ( \3288 , \2414 );
or \U$2598 ( \3289 , \3287 , \3288 );
not \U$2599 ( \3290 , \1823 );
not \U$2600 ( \3291 , \2408 );
or \U$2601 ( \3292 , \3290 , \3291 );
nand \U$2602 ( \3293 , \2079 , \1824 );
nand \U$2603 ( \3294 , \3292 , \3293 );
nand \U$2604 ( \3295 , \3294 , \2157 );
nand \U$2605 ( \3296 , \3289 , \3295 );
xor \U$2606 ( \3297 , \3286 , \3296 );
not \U$2607 ( \3298 , \3029 );
not \U$2608 ( \3299 , \2479 );
or \U$2609 ( \3300 , \3298 , \3299 );
and \U$2610 ( \3301 , \2151 , \1744 );
not \U$2611 ( \3302 , \2151 );
and \U$2612 ( \3303 , \3302 , \2202 );
nor \U$2613 ( \3304 , \3301 , \3303 );
nand \U$2614 ( \3305 , \2472 , \3304 );
nand \U$2615 ( \3306 , \3300 , \3305 );
and \U$2616 ( \3307 , \3297 , \3306 );
and \U$2617 ( \3308 , \3286 , \3296 );
or \U$2618 ( \3309 , \3307 , \3308 );
xor \U$2619 ( \3310 , \3277 , \3309 );
not \U$2620 ( \3311 , \3284 );
not \U$2621 ( \3312 , \2465 );
or \U$2622 ( \3313 , \3311 , \3312 );
not \U$2623 ( \3314 , \1757 );
not \U$2624 ( \3315 , \3025 );
not \U$2625 ( \3316 , \1784 );
or \U$2626 ( \3317 , \3315 , \3316 );
not \U$2627 ( \3318 , \3025 );
nand \U$2628 ( \3319 , \3014 , \3318 );
nand \U$2629 ( \3320 , \3317 , \3319 );
nand \U$2630 ( \3321 , \3314 , \3320 );
nand \U$2631 ( \3322 , \3313 , \3321 );
not \U$2632 ( \3323 , \3294 );
not \U$2633 ( \3324 , \2414 );
or \U$2634 ( \3325 , \3323 , \3324 );
and \U$2635 ( \3326 , \1730 , \2079 );
not \U$2636 ( \3327 , \1730 );
and \U$2637 ( \3328 , \3327 , \2408 );
nor \U$2638 ( \3329 , \3326 , \3328 );
nand \U$2639 ( \3330 , \3329 , \2157 );
nand \U$2640 ( \3331 , \3325 , \3330 );
xor \U$2641 ( \3332 , \3322 , \3331 );
not \U$2642 ( \3333 , \3304 );
not \U$2643 ( \3334 , \2479 );
not \U$2644 ( \3335 , \3334 );
not \U$2645 ( \3336 , \3335 );
or \U$2646 ( \3337 , \3333 , \3336 );
and \U$2647 ( \3338 , \2982 , \1744 );
not \U$2648 ( \3339 , \2982 );
and \U$2649 ( \3340 , \3339 , \2202 );
nor \U$2650 ( \3341 , \3338 , \3340 );
nand \U$2651 ( \3342 , \2472 , \3341 );
nand \U$2652 ( \3343 , \3337 , \3342 );
xor \U$2653 ( \3344 , \3332 , \3343 );
xor \U$2654 ( \3345 , \3310 , \3344 );
not \U$2655 ( \3346 , \3032 );
nand \U$2656 ( \3347 , \2963 , \2993 );
not \U$2657 ( \3348 , \3347 );
or \U$2658 ( \3349 , \3346 , \3348 );
nand \U$2659 ( \3350 , \2964 , \2994 );
nand \U$2660 ( \3351 , \3349 , \3350 );
xor \U$2661 ( \3352 , \3043 , \3048 );
and \U$2662 ( \3353 , \3352 , \3061 );
and \U$2663 ( \3354 , \3043 , \3048 );
or \U$2664 ( \3355 , \3353 , \3354 );
xor \U$2665 ( \3356 , \3351 , \3355 );
nor \U$2666 ( \3357 , \2989 , \2976 );
or \U$2667 ( \3358 , \3357 , \2966 );
nand \U$2668 ( \3359 , \2989 , \2976 );
nand \U$2669 ( \3360 , \3358 , \3359 );
not \U$2670 ( \3361 , \1613 );
not \U$2671 ( \3362 , \2461 );
not \U$2672 ( \3363 , \1614 );
or \U$2673 ( \3364 , \3362 , \3363 );
nand \U$2674 ( \3365 , \1680 , \2457 );
nand \U$2675 ( \3366 , \3364 , \3365 );
nor \U$2676 ( \3367 , \3361 , \3366 );
xor \U$2677 ( \3368 , \3360 , \3367 );
not \U$2678 ( \3369 , \3059 );
not \U$2679 ( \3370 , \1396 );
or \U$2680 ( \3371 , \3369 , \3370 );
not \U$2681 ( \3372 , \2931 );
not \U$2682 ( \3373 , \2398 );
or \U$2683 ( \3374 , \3372 , \3373 );
not \U$2684 ( \3375 , \1398 );
nand \U$2685 ( \3376 , \3375 , \2397 );
nand \U$2686 ( \3377 , \3374 , \3376 );
nand \U$2687 ( \3378 , \3377 , \1605 );
nand \U$2688 ( \3379 , \3371 , \3378 );
xor \U$2689 ( \3380 , \3368 , \3379 );
and \U$2690 ( \3381 , \3356 , \3380 );
and \U$2691 ( \3382 , \3351 , \3355 );
or \U$2692 ( \3383 , \3381 , \3382 );
xor \U$2693 ( \3384 , \3345 , \3383 );
xor \U$2694 ( \3385 , \3360 , \3367 );
and \U$2695 ( \3386 , \3385 , \3379 );
and \U$2696 ( \3387 , \3360 , \3367 );
or \U$2697 ( \3388 , \3386 , \3387 );
not \U$2698 ( \3389 , \1963 );
not \U$2699 ( \3390 , \1948 );
or \U$2700 ( \3391 , \3389 , \3390 );
nand \U$2701 ( \3392 , \3391 , \1951 );
xor \U$2702 ( \3393 , \3392 , \3268 );
not \U$2703 ( \3394 , \1878 );
not \U$2704 ( \3395 , \3266 );
or \U$2705 ( \3396 , \3394 , \3395 );
and \U$2706 ( \3397 , \1599 , \1914 );
not \U$2707 ( \3398 , \1599 );
and \U$2708 ( \3399 , \3398 , \1915 );
nor \U$2709 ( \3400 , \3397 , \3399 );
or \U$2710 ( \3401 , \3400 , \1928 );
nand \U$2711 ( \3402 , \3396 , \3401 );
xor \U$2712 ( \3403 , \3393 , \3402 );
not \U$2713 ( \3404 , \3377 );
not \U$2714 ( \3405 , \1396 );
or \U$2715 ( \3406 , \3404 , \3405 );
and \U$2716 ( \3407 , \2822 , \1398 );
not \U$2717 ( \3408 , \2822 );
and \U$2718 ( \3409 , \3408 , \2528 );
nor \U$2719 ( \3410 , \3407 , \3409 );
nand \U$2720 ( \3411 , \3410 , \1605 );
nand \U$2721 ( \3412 , \3406 , \3411 );
xor \U$2722 ( \3413 , \3403 , \3412 );
and \U$2723 ( \3414 , \1614 , \2338 );
and \U$2724 ( \3415 , \2637 , \2332 );
nor \U$2725 ( \3416 , \3414 , \3415 );
and \U$2726 ( \3417 , \1613 , \3416 );
xor \U$2727 ( \3418 , \3413 , \3417 );
xor \U$2728 ( \3419 , \3388 , \3418 );
xor \U$2729 ( \3420 , \3269 , \3273 );
xor \U$2730 ( \3421 , \3420 , \3009 );
xor \U$2731 ( \3422 , \3010 , \3020 );
and \U$2732 ( \3423 , \3422 , \3031 );
and \U$2733 ( \3424 , \3010 , \3020 );
or \U$2734 ( \3425 , \3423 , \3424 );
xor \U$2735 ( \3426 , \3421 , \3425 );
xor \U$2736 ( \3427 , \3286 , \3296 );
xor \U$2737 ( \3428 , \3427 , \3306 );
and \U$2738 ( \3429 , \3426 , \3428 );
and \U$2739 ( \3430 , \3421 , \3425 );
or \U$2740 ( \3431 , \3429 , \3430 );
xor \U$2741 ( \3432 , \3419 , \3431 );
xor \U$2742 ( \3433 , \3384 , \3432 );
xor \U$2743 ( \3434 , \3421 , \3425 );
xor \U$2744 ( \3435 , \3434 , \3428 );
xor \U$2745 ( \3436 , \3039 , \3062 );
and \U$2746 ( \3437 , \3436 , \3067 );
and \U$2747 ( \3438 , \3039 , \3062 );
or \U$2748 ( \3439 , \3437 , \3438 );
xor \U$2749 ( \3440 , \3435 , \3439 );
xor \U$2750 ( \3441 , \3351 , \3355 );
xor \U$2751 ( \3442 , \3441 , \3380 );
and \U$2752 ( \3443 , \3440 , \3442 );
and \U$2753 ( \3444 , \3435 , \3439 );
or \U$2754 ( \3445 , \3443 , \3444 );
nor \U$2755 ( \3446 , \3433 , \3445 );
xor \U$2756 ( \3447 , \3435 , \3439 );
xor \U$2757 ( \3448 , \3447 , \3442 );
not \U$2758 ( \3449 , \3034 );
not \U$2759 ( \3450 , \3077 );
or \U$2760 ( \3451 , \3449 , \3450 );
nand \U$2761 ( \3452 , \3451 , \3068 );
not \U$2762 ( \3453 , \3034 );
nand \U$2763 ( \3454 , \3453 , \3076 );
nand \U$2764 ( \3455 , \3452 , \3454 );
nor \U$2765 ( \3456 , \3448 , \3455 );
nor \U$2766 ( \3457 , \3446 , \3456 );
and \U$2767 ( \3458 , \3259 , \3457 );
not \U$2768 ( \3459 , \3458 );
nand \U$2769 ( \3460 , \1461 , RI99339d0_265);
and \U$2770 ( \3461 , \1471 , RI9931360_285);
not \U$2771 ( \3462 , RI9922450_585);
not \U$2772 ( \3463 , \1487 );
or \U$2773 ( \3464 , \3462 , \3463 );
not \U$2774 ( \3465 , RI9923080_565);
or \U$2775 ( \3466 , \1643 , \3465 );
nand \U$2776 ( \3467 , \3464 , \3466 );
nor \U$2777 ( \3468 , \3461 , \3467 );
nand \U$2778 ( \3469 , \1499 , RI9928c60_405);
nand \U$2779 ( \3470 , \3460 , \3468 , \3469 );
not \U$2780 ( \3471 , \1506 );
not \U$2781 ( \3472 , RI992f0b0_305);
not \U$2782 ( \3473 , \3472 );
and \U$2783 ( \3474 , \3471 , \3473 );
and \U$2784 ( \3475 , \1626 , RI9926f50_445);
nor \U$2785 ( \3476 , \3474 , \3475 );
not \U$2786 ( \3477 , \1629 );
not \U$2787 ( \3478 , RI992d1c0_325);
not \U$2788 ( \3479 , \3478 );
and \U$2789 ( \3480 , \3477 , \3479 );
and \U$2790 ( \3481 , \2295 , RI992ad30_365);
nor \U$2791 ( \3482 , \3480 , \3481 );
nand \U$2792 ( \3483 , \3476 , \3482 );
nor \U$2793 ( \3484 , \3470 , \3483 );
not \U$2794 ( \3485 , RI99265f0_465);
or \U$2795 ( \3486 , \1545 , \3485 );
not \U$2796 ( \3487 , RI9925c90_485);
or \U$2797 ( \3488 , \1653 , \3487 );
and \U$2798 ( \3489 , \2622 , RI992a3d0_385);
not \U$2799 ( \3490 , RI99239e0_545);
nor \U$2800 ( \3491 , \2160 , \3490 );
nor \U$2801 ( \3492 , \3489 , \3491 );
nand \U$2802 ( \3493 , \3486 , \3488 , \3492 );
and \U$2803 ( \3494 , \1657 , RI9928300_425);
and \U$2804 ( \3495 , \1659 , RI9924ca0_505);
nor \U$2805 ( \3496 , \3494 , \3495 );
not \U$2806 ( \3497 , \1587 );
not \U$2807 ( \3498 , RI992c860_345);
not \U$2808 ( \3499 , \3498 );
and \U$2809 ( \3500 , \3497 , \3499 );
and \U$2810 ( \3501 , \1593 , RI9924340_525);
nor \U$2811 ( \3502 , \3500 , \3501 );
nand \U$2812 ( \3503 , \3496 , \3502 );
nor \U$2813 ( \3504 , \3493 , \3503 );
nand \U$2814 ( \3505 , \3484 , \3504 );
buf \U$2815 ( \3506 , \3505 );
and \U$2816 ( \3507 , \3506 , \1744 );
not \U$2817 ( \3508 , \3506 );
and \U$2818 ( \3509 , \3508 , \2202 );
nor \U$2819 ( \3510 , \3507 , \3509 );
not \U$2820 ( \3511 , \3510 );
not \U$2821 ( \3512 , \2479 );
or \U$2822 ( \3513 , \3511 , \3512 );
or \U$2823 ( \3514 , \2202 , \3146 );
not \U$2824 ( \3515 , \3146 );
or \U$2825 ( \3516 , \1744 , \3515 );
nand \U$2826 ( \3517 , \3514 , \3516 );
nand \U$2827 ( \3518 , \2472 , \3517 );
nand \U$2828 ( \3519 , \3513 , \3518 );
and \U$2829 ( \3520 , \2584 , \1915 );
not \U$2830 ( \3521 , \2584 );
and \U$2831 ( \3522 , \3521 , \1925 );
nor \U$2832 ( \3523 , \3520 , \3522 );
not \U$2833 ( \3524 , \3523 );
not \U$2834 ( \3525 , \3524 );
not \U$2835 ( \3526 , \1878 );
or \U$2836 ( \3527 , \3525 , \3526 );
not \U$2837 ( \3528 , \2797 );
not \U$2838 ( \3529 , \1915 );
or \U$2839 ( \3530 , \3528 , \3529 );
nand \U$2840 ( \3531 , \1925 , \2796 );
nand \U$2841 ( \3532 , \3530 , \3531 );
nand \U$2842 ( \3533 , \3532 , \1929 );
nand \U$2843 ( \3534 , \3527 , \3533 );
not \U$2844 ( \3535 , \1949 );
and \U$2845 ( \3536 , \1951 , \2457 );
not \U$2846 ( \3537 , \1951 );
and \U$2847 ( \3538 , \3537 , \2461 );
nor \U$2848 ( \3539 , \3536 , \3538 );
not \U$2849 ( \3540 , \3539 );
or \U$2850 ( \3541 , \3535 , \3540 );
and \U$2851 ( \3542 , \1951 , \2332 );
not \U$2852 ( \3543 , \1951 );
and \U$2853 ( \3544 , \3543 , \2338 );
nor \U$2854 ( \3545 , \3542 , \3544 );
nand \U$2855 ( \3546 , \1964 , \3545 );
nand \U$2856 ( \3547 , \3541 , \3546 );
xor \U$2857 ( \3548 , \3534 , \3547 );
or \U$2858 ( \3549 , \1752 , \1744 );
not \U$2859 ( \3550 , RI9926500_467);
nor \U$2860 ( \3551 , \1544 , \3550 );
not \U$2861 ( \3552 , \3551 );
not \U$2862 ( \3553 , \1653 );
nand \U$2863 ( \3554 , \3553 , RI9925ba0_487);
and \U$2864 ( \3555 , \1626 , RI9926e60_447);
and \U$2865 ( \3556 , \1634 , RI992ac40_367);
nor \U$2866 ( \3557 , \3555 , \3556 );
nand \U$2867 ( \3558 , \3552 , \3554 , \3557 );
not \U$2868 ( \3559 , RI9928b70_407);
not \U$2869 ( \3560 , \1499 );
or \U$2870 ( \3561 , \3559 , \3560 );
nand \U$2871 ( \3562 , RI992efc0_307, \1507 );
nand \U$2872 ( \3563 , \3561 , \3562 );
nor \U$2873 ( \3564 , \3558 , \3563 );
nand \U$2874 ( \3565 , \1593 , RI9924250_527);
nand \U$2875 ( \3566 , \1586 , RI992c770_347);
nand \U$2876 ( \3567 , \1469 , RI992f920_287);
and \U$2877 ( \3568 , \1481 , RI9922f90_567);
and \U$2878 ( \3569 , \1487 , RI9922360_587);
nor \U$2879 ( \3570 , \3568 , \3569 );
nand \U$2880 ( \3571 , \3565 , \3566 , \3567 , \3570 );
and \U$2881 ( \3572 , \1461 , RI99338e0_267);
nor \U$2882 ( \3573 , \3571 , \3572 );
nand \U$2883 ( \3574 , \2622 , RI992a2e0_387);
nand \U$2884 ( \3575 , \1564 , RI99238f0_547);
nand \U$2885 ( \3576 , \1535 , RI992d0d0_327);
nand \U$2886 ( \3577 , \3574 , \3575 , \3576 );
not \U$2887 ( \3578 , RI9928210_427);
not \U$2888 ( \3579 , \1657 );
or \U$2889 ( \3580 , \3578 , \3579 );
nand \U$2890 ( \3581 , \1710 , RI9924bb0_507);
nand \U$2891 ( \3582 , \3580 , \3581 );
nor \U$2892 ( \3583 , \3577 , \3582 );
nand \U$2893 ( \3584 , \3564 , \3573 , \3583 );
buf \U$2894 ( \3585 , \3584 );
nand \U$2895 ( \3586 , \3549 , \3585 );
nand \U$2896 ( \3587 , \1752 , \1744 );
and \U$2897 ( \3588 , \1393 , \3586 , \3587 );
not \U$2898 ( \3589 , \1975 );
and \U$2899 ( \3590 , \1967 , \2396 );
not \U$2900 ( \3591 , \1967 );
and \U$2901 ( \3592 , \3591 , \2397 );
nor \U$2902 ( \3593 , \3590 , \3592 );
not \U$2903 ( \3594 , \3593 );
or \U$2904 ( \3595 , \3589 , \3594 );
and \U$2905 ( \3596 , \1967 , \2199 );
not \U$2906 ( \3597 , \1967 );
and \U$2907 ( \3598 , \3597 , \2822 );
nor \U$2908 ( \3599 , \3596 , \3598 );
nand \U$2909 ( \3600 , \3599 , \1973 );
nand \U$2910 ( \3601 , \3595 , \3600 );
xnor \U$2911 ( \3602 , \3588 , \3601 );
xnor \U$2912 ( \3603 , \3548 , \3602 );
or \U$2913 ( \3604 , \3519 , \3603 );
and \U$2914 ( \3605 , \2526 , \1914 );
not \U$2915 ( \3606 , \2526 );
and \U$2916 ( \3607 , \3606 , \1922 );
nor \U$2917 ( \3608 , \3605 , \3607 );
not \U$2918 ( \3609 , \3608 );
or \U$2919 ( \3610 , \3394 , \3609 );
or \U$2920 ( \3611 , \3523 , \1928 );
nand \U$2921 ( \3612 , \3610 , \3611 );
not \U$2922 ( \3613 , \1975 );
and \U$2923 ( \3614 , \1967 , \2457 );
not \U$2924 ( \3615 , \1967 );
and \U$2925 ( \3616 , \3615 , \2461 );
nor \U$2926 ( \3617 , \3614 , \3616 );
not \U$2927 ( \3618 , \3617 );
or \U$2928 ( \3619 , \3613 , \3618 );
and \U$2929 ( \3620 , \1967 , \2332 );
not \U$2930 ( \3621 , \1967 );
and \U$2931 ( \3622 , \3621 , \2338 );
nor \U$2932 ( \3623 , \3620 , \3622 );
nand \U$2933 ( \3624 , \3623 , \1973 );
nand \U$2934 ( \3625 , \3619 , \3624 );
not \U$2935 ( \3626 , \1964 );
and \U$2936 ( \3627 , \2795 , \1951 );
not \U$2937 ( \3628 , \2795 );
and \U$2938 ( \3629 , \3628 , \1872 );
nor \U$2939 ( \3630 , \3627 , \3629 );
not \U$2940 ( \3631 , \3630 );
or \U$2941 ( \3632 , \3626 , \3631 );
and \U$2942 ( \3633 , \1951 , \2584 );
not \U$2943 ( \3634 , \1951 );
and \U$2944 ( \3635 , \3634 , \2587 );
nor \U$2945 ( \3636 , \3633 , \3635 );
nand \U$2946 ( \3637 , \3636 , \1949 );
nand \U$2947 ( \3638 , \3632 , \3637 );
and \U$2948 ( \3639 , \3625 , \3638 );
xor \U$2949 ( \3640 , \3612 , \3639 );
not \U$2950 ( \3641 , \3146 );
not \U$2951 ( \3642 , \2408 );
or \U$2952 ( \3643 , \3641 , \3642 );
nand \U$2953 ( \3644 , \2079 , \3515 );
nand \U$2954 ( \3645 , \3643 , \3644 );
not \U$2955 ( \3646 , \3645 );
not \U$2956 ( \3647 , \2414 );
or \U$2957 ( \3648 , \3646 , \3647 );
not \U$2958 ( \3649 , \2634 );
not \U$2959 ( \3650 , \2408 );
or \U$2960 ( \3651 , \3649 , \3650 );
nand \U$2961 ( \3652 , \2814 , \2633 );
nand \U$2962 ( \3653 , \3651 , \3652 );
nand \U$2963 ( \3654 , \3653 , \2157 );
nand \U$2964 ( \3655 , \3648 , \3654 );
and \U$2965 ( \3656 , \3640 , \3655 );
and \U$2966 ( \3657 , \3612 , \3639 );
or \U$2967 ( \3658 , \3656 , \3657 );
nand \U$2968 ( \3659 , \3604 , \3658 );
nand \U$2969 ( \3660 , \3519 , \3603 );
and \U$2970 ( \3661 , \3659 , \3660 );
not \U$2971 ( \3662 , \3661 );
not \U$2972 ( \3663 , \3534 );
nand \U$2973 ( \3664 , \3602 , \3663 );
and \U$2974 ( \3665 , \3664 , \3547 );
nor \U$2975 ( \3666 , \3602 , \3663 );
nor \U$2976 ( \3667 , \3665 , \3666 );
not \U$2977 ( \3668 , \3585 );
not \U$2978 ( \3669 , \2337 );
not \U$2979 ( \3670 , \3669 );
or \U$2980 ( \3671 , \3668 , \3670 );
not \U$2981 ( \3672 , \3585 );
nand \U$2982 ( \3673 , \1770 , \3672 );
nand \U$2983 ( \3674 , \3671 , \3673 );
not \U$2984 ( \3675 , \3674 );
not \U$2985 ( \3676 , \1766 );
or \U$2986 ( \3677 , \3675 , \3676 );
nand \U$2987 ( \3678 , \1461 , RI9933958_266);
and \U$2988 ( \3679 , \1469 , RI99312e8_286);
not \U$2989 ( \3680 , RI99223d8_586);
not \U$2990 ( \3681 , \1487 );
or \U$2991 ( \3682 , \3680 , \3681 );
not \U$2992 ( \3683 , RI9923008_566);
or \U$2993 ( \3684 , \1643 , \3683 );
nand \U$2994 ( \3685 , \3682 , \3684 );
nor \U$2995 ( \3686 , \3679 , \3685 );
nand \U$2996 ( \3687 , \1499 , RI9928be8_406);
nand \U$2997 ( \3688 , \3678 , \3686 , \3687 );
and \U$2998 ( \3689 , \1519 , RI9926ed8_446);
not \U$2999 ( \3690 , RI992f038_306);
nor \U$3000 ( \3691 , \1506 , \3690 );
nor \U$3001 ( \3692 , \3689 , \3691 );
and \U$3002 ( \3693 , \1535 , RI992d148_326);
and \U$3003 ( \3694 , \1636 , RI992acb8_366);
nor \U$3004 ( \3695 , \3693 , \3694 );
nand \U$3005 ( \3696 , \3692 , \3695 );
nor \U$3006 ( \3697 , \3688 , \3696 );
and \U$3007 ( \3698 , \1715 , RI9926578_466);
and \U$3008 ( \3699 , \1550 , RI9925c18_486);
nor \U$3009 ( \3700 , \3698 , \3699 );
and \U$3010 ( \3701 , \2622 , RI992a358_386);
and \U$3011 ( \3702 , \1564 , RI9923968_546);
nor \U$3012 ( \3703 , \3701 , \3702 );
nand \U$3013 ( \3704 , \3700 , \3703 );
and \U$3014 ( \3705 , \1657 , RI9928288_426);
and \U$3015 ( \3706 , \1710 , RI9924c28_506);
nor \U$3016 ( \3707 , \3705 , \3706 );
and \U$3017 ( \3708 , \1586 , RI992c7e8_346);
and \U$3018 ( \3709 , \1593 , RI99242c8_526);
nor \U$3019 ( \3710 , \3708 , \3709 );
nand \U$3020 ( \3711 , \3707 , \3710 );
nor \U$3021 ( \3712 , \3704 , \3711 );
nand \U$3022 ( \3713 , \3697 , \3712 );
not \U$3023 ( \3714 , \3713 );
not \U$3024 ( \3715 , \3714 );
not \U$3025 ( \3716 , \3715 );
not \U$3026 ( \3717 , \2334 );
or \U$3027 ( \3718 , \3716 , \3717 );
nand \U$3028 ( \3719 , \2337 , \3714 );
nand \U$3029 ( \3720 , \3718 , \3719 );
nand \U$3030 ( \3721 , \3720 , \1758 );
nand \U$3031 ( \3722 , \3677 , \3721 );
not \U$3032 ( \3723 , \3653 );
not \U$3033 ( \3724 , \2414 );
or \U$3034 ( \3725 , \3723 , \3724 );
not \U$3035 ( \3726 , \2526 );
not \U$3036 ( \3727 , \2408 );
or \U$3037 ( \3728 , \3726 , \3727 );
not \U$3038 ( \3729 , \2029 );
nand \U$3039 ( \3730 , \3729 , \2532 );
nand \U$3040 ( \3731 , \3728 , \3730 );
nand \U$3041 ( \3732 , \3731 , \2157 );
nand \U$3042 ( \3733 , \3725 , \3732 );
or \U$3043 ( \3734 , \3722 , \3733 );
not \U$3044 ( \3735 , \1973 );
not \U$3045 ( \3736 , \3593 );
or \U$3046 ( \3737 , \3735 , \3736 );
nand \U$3047 ( \3738 , \3623 , \1975 );
nand \U$3048 ( \3739 , \3737 , \3738 );
not \U$3049 ( \3740 , \1964 );
not \U$3050 ( \3741 , \3539 );
or \U$3051 ( \3742 , \3740 , \3741 );
nand \U$3052 ( \3743 , \3630 , \1949 );
nand \U$3053 ( \3744 , \3742 , \3743 );
xor \U$3054 ( \3745 , \3739 , \3744 );
and \U$3055 ( \3746 , \1758 , \3585 );
and \U$3056 ( \3747 , \3745 , \3746 );
and \U$3057 ( \3748 , \3739 , \3744 );
or \U$3058 ( \3749 , \3747 , \3748 );
nand \U$3059 ( \3750 , \3734 , \3749 );
nand \U$3060 ( \3751 , \3733 , \3722 );
and \U$3061 ( \3752 , \3750 , \3751 );
xor \U$3062 ( \3753 , \3667 , \3752 );
nand \U$3063 ( \3754 , \3588 , \3601 );
nand \U$3064 ( \3755 , \1605 , \3585 );
xor \U$3065 ( \3756 , \3754 , \3755 );
not \U$3066 ( \3757 , \3731 );
not \U$3067 ( \3758 , \2414 );
nor \U$3068 ( \3759 , \3757 , \3758 );
not \U$3069 ( \3760 , \2584 );
not \U$3070 ( \3761 , \2408 );
or \U$3071 ( \3762 , \3760 , \3761 );
nand \U$3072 ( \3763 , \2079 , \2587 );
nand \U$3073 ( \3764 , \3762 , \3763 );
not \U$3074 ( \3765 , \3764 );
not \U$3075 ( \3766 , \2157 );
nor \U$3076 ( \3767 , \3765 , \3766 );
nor \U$3077 ( \3768 , \3759 , \3767 );
xor \U$3078 ( \3769 , \3756 , \3768 );
xor \U$3079 ( \3770 , \3753 , \3769 );
not \U$3080 ( \3771 , \3770 );
or \U$3081 ( \3772 , \3662 , \3771 );
not \U$3082 ( \3773 , \3517 );
not \U$3083 ( \3774 , \2479 );
or \U$3084 ( \3775 , \3773 , \3774 );
and \U$3085 ( \3776 , \2634 , \1744 );
not \U$3086 ( \3777 , \2634 );
and \U$3087 ( \3778 , \3777 , \2202 );
nor \U$3088 ( \3779 , \3776 , \3778 );
nand \U$3089 ( \3780 , \2472 , \3779 );
nand \U$3090 ( \3781 , \3775 , \3780 );
not \U$3091 ( \3782 , \1973 );
and \U$3092 ( \3783 , \1967 , \2270 );
not \U$3093 ( \3784 , \1967 );
and \U$3094 ( \3785 , \3784 , \2671 );
nor \U$3095 ( \3786 , \3783 , \3785 );
not \U$3096 ( \3787 , \3786 );
or \U$3097 ( \3788 , \3782 , \3787 );
nand \U$3098 ( \3789 , \3599 , \1975 );
nand \U$3099 ( \3790 , \3788 , \3789 );
not \U$3100 ( \3791 , \1964 );
xor \U$3101 ( \3792 , \1951 , \2396 );
not \U$3102 ( \3793 , \3792 );
or \U$3103 ( \3794 , \3791 , \3793 );
nand \U$3104 ( \3795 , \3545 , \1949 );
nand \U$3105 ( \3796 , \3794 , \3795 );
xor \U$3106 ( \3797 , \3790 , \3796 );
not \U$3107 ( \3798 , \3532 );
not \U$3108 ( \3799 , \1878 );
or \U$3109 ( \3800 , \3798 , \3799 );
not \U$3110 ( \3801 , \2457 );
not \U$3111 ( \3802 , \1915 );
or \U$3112 ( \3803 , \3801 , \3802 );
nand \U$3113 ( \3804 , \1914 , \2461 );
nand \U$3114 ( \3805 , \3803 , \3804 );
nand \U$3115 ( \3806 , \3805 , \1929 );
nand \U$3116 ( \3807 , \3800 , \3806 );
xor \U$3117 ( \3808 , \3797 , \3807 );
xor \U$3118 ( \3809 , \3781 , \3808 );
not \U$3119 ( \3810 , \3720 );
not \U$3120 ( \3811 , \1766 );
or \U$3121 ( \3812 , \3810 , \3811 );
not \U$3122 ( \3813 , \3506 );
not \U$3123 ( \3814 , \2334 );
or \U$3124 ( \3815 , \3813 , \3814 );
not \U$3125 ( \3816 , \3506 );
nand \U$3126 ( \3817 , \3014 , \3816 );
nand \U$3127 ( \3818 , \3815 , \3817 );
nand \U$3128 ( \3819 , \3818 , \1758 );
nand \U$3129 ( \3820 , \3812 , \3819 );
xor \U$3130 ( \3821 , \3809 , \3820 );
nand \U$3131 ( \3822 , \3772 , \3821 );
not \U$3132 ( \3823 , \3661 );
not \U$3133 ( \3824 , \3770 );
nand \U$3134 ( \3825 , \3823 , \3824 );
nand \U$3135 ( \3826 , \3822 , \3825 );
not \U$3136 ( \3827 , \3826 );
not \U$3137 ( \3828 , \3779 );
not \U$3138 ( \3829 , \2479 );
or \U$3139 ( \3830 , \3828 , \3829 );
and \U$3140 ( \3831 , \2526 , \1744 );
not \U$3141 ( \3832 , \2526 );
and \U$3142 ( \3833 , \3832 , \2202 );
nor \U$3143 ( \3834 , \3831 , \3833 );
nand \U$3144 ( \3835 , \2472 , \3834 );
nand \U$3145 ( \3836 , \3830 , \3835 );
and \U$3146 ( \3837 , \3585 , \3375 );
not \U$3147 ( \3838 , \3585 );
and \U$3148 ( \3839 , \3838 , \1381 );
nor \U$3149 ( \3840 , \3837 , \3839 );
not \U$3150 ( \3841 , \3840 );
not \U$3151 ( \3842 , \2536 );
or \U$3152 ( \3843 , \3841 , \3842 );
and \U$3153 ( \3844 , \3715 , \2528 );
not \U$3154 ( \3845 , \3715 );
and \U$3155 ( \3846 , \3845 , \1381 );
nor \U$3156 ( \3847 , \3844 , \3846 );
nand \U$3157 ( \3848 , \3847 , \1605 );
nand \U$3158 ( \3849 , \3843 , \3848 );
xor \U$3159 ( \3850 , \3836 , \3849 );
xor \U$3160 ( \3851 , \3754 , \3755 );
and \U$3161 ( \3852 , \3851 , \3768 );
and \U$3162 ( \3853 , \3754 , \3755 );
or \U$3163 ( \3854 , \3852 , \3853 );
xor \U$3164 ( \3855 , \3850 , \3854 );
xor \U$3165 ( \3856 , \3667 , \3752 );
and \U$3166 ( \3857 , \3856 , \3769 );
and \U$3167 ( \3858 , \3667 , \3752 );
or \U$3168 ( \3859 , \3857 , \3858 );
xor \U$3169 ( \3860 , \3855 , \3859 );
not \U$3170 ( \3861 , \3805 );
or \U$3171 ( \3862 , \3394 , \3861 );
and \U$3172 ( \3863 , \2332 , \1915 );
not \U$3173 ( \3864 , \2332 );
and \U$3174 ( \3865 , \3864 , \1914 );
nor \U$3175 ( \3866 , \3863 , \3865 );
or \U$3176 ( \3867 , \3866 , \1928 );
nand \U$3177 ( \3868 , \3862 , \3867 );
not \U$3178 ( \3869 , \1964 );
and \U$3179 ( \3870 , \1872 , \2822 );
not \U$3180 ( \3871 , \1872 );
and \U$3181 ( \3872 , \3871 , \2199 );
nor \U$3182 ( \3873 , \3870 , \3872 );
not \U$3183 ( \3874 , \3873 );
or \U$3184 ( \3875 , \3869 , \3874 );
nand \U$3185 ( \3876 , \3792 , \1949 );
nand \U$3186 ( \3877 , \3875 , \3876 );
and \U$3187 ( \3878 , \3786 , \1975 );
not \U$3188 ( \3879 , \1967 );
not \U$3189 ( \3880 , \2080 );
or \U$3190 ( \3881 , \3879 , \3880 );
nand \U$3191 ( \3882 , \2076 , \1945 );
nand \U$3192 ( \3883 , \3881 , \3882 );
and \U$3193 ( \3884 , \3883 , \1973 );
nor \U$3194 ( \3885 , \3878 , \3884 );
xor \U$3195 ( \3886 , \3877 , \3885 );
xor \U$3196 ( \3887 , \3868 , \3886 );
nand \U$3197 ( \3888 , \1384 , \2334 );
and \U$3198 ( \3889 , \3888 , \3585 );
and \U$3199 ( \3890 , \1383 , \2337 );
nor \U$3200 ( \3891 , \3889 , \3890 );
nand \U$3201 ( \3892 , \3375 , \3891 );
xnor \U$3202 ( \3893 , \3887 , \3892 );
or \U$3203 ( \3894 , \3781 , \3820 );
nand \U$3204 ( \3895 , \3894 , \3808 );
nand \U$3205 ( \3896 , \3781 , \3820 );
and \U$3206 ( \3897 , \3895 , \3896 );
xor \U$3207 ( \3898 , \3893 , \3897 );
xor \U$3208 ( \3899 , \3790 , \3796 );
and \U$3209 ( \3900 , \3899 , \3807 );
and \U$3210 ( \3901 , \3790 , \3796 );
or \U$3211 ( \3902 , \3900 , \3901 );
not \U$3212 ( \3903 , \3764 );
not \U$3213 ( \3904 , \2414 );
or \U$3214 ( \3905 , \3903 , \3904 );
not \U$3215 ( \3906 , \2797 );
not \U$3216 ( \3907 , \2029 );
or \U$3217 ( \3908 , \3906 , \3907 );
nand \U$3218 ( \3909 , \2079 , \2796 );
nand \U$3219 ( \3910 , \3908 , \3909 );
nand \U$3220 ( \3911 , \3910 , \2157 );
nand \U$3221 ( \3912 , \3905 , \3911 );
xor \U$3222 ( \3913 , \3902 , \3912 );
not \U$3223 ( \3914 , \3818 );
not \U$3224 ( \3915 , \1766 );
or \U$3225 ( \3916 , \3914 , \3915 );
and \U$3226 ( \3917 , \3146 , \1770 );
not \U$3227 ( \3918 , \3146 );
and \U$3228 ( \3919 , \3918 , \1784 );
nor \U$3229 ( \3920 , \3917 , \3919 );
nand \U$3230 ( \3921 , \3920 , \1758 );
nand \U$3231 ( \3922 , \3916 , \3921 );
not \U$3232 ( \3923 , \3922 );
xor \U$3233 ( \3924 , \3913 , \3923 );
xor \U$3234 ( \3925 , \3898 , \3924 );
xor \U$3235 ( \3926 , \3860 , \3925 );
nand \U$3236 ( \3927 , \3827 , \3926 );
not \U$3237 ( \3928 , \3927 );
xor \U$3238 ( \3929 , \3821 , \3661 );
xor \U$3239 ( \3930 , \3929 , \3824 );
xor \U$3240 ( \3931 , \3733 , \3749 );
xor \U$3241 ( \3932 , \3931 , \3722 );
not \U$3242 ( \3933 , \3932 );
not \U$3243 ( \3934 , \3933 );
and \U$3244 ( \3935 , \3715 , \1744 );
not \U$3245 ( \3936 , \3715 );
and \U$3246 ( \3937 , \3936 , \2202 );
nor \U$3247 ( \3938 , \3935 , \3937 );
not \U$3248 ( \3939 , \3938 );
not \U$3249 ( \3940 , \3335 );
or \U$3250 ( \3941 , \3939 , \3940 );
nand \U$3251 ( \3942 , \2472 , \3510 );
nand \U$3252 ( \3943 , \3941 , \3942 );
not \U$3253 ( \3944 , \2634 );
not \U$3254 ( \3945 , \1915 );
or \U$3255 ( \3946 , \3944 , \3945 );
nand \U$3256 ( \3947 , \1925 , \2633 );
nand \U$3257 ( \3948 , \3946 , \3947 );
not \U$3258 ( \3949 , \3948 );
not \U$3259 ( \3950 , \1878 );
or \U$3260 ( \3951 , \3949 , \3950 );
nand \U$3261 ( \3952 , \3608 , \1929 );
nand \U$3262 ( \3953 , \3951 , \3952 );
xor \U$3263 ( \3954 , \3625 , \3638 );
xor \U$3264 ( \3955 , \3953 , \3954 );
buf \U$3265 ( \3956 , \2217 );
not \U$3266 ( \3957 , \3956 );
not \U$3267 ( \3958 , \3957 );
not \U$3268 ( \3959 , \2408 );
or \U$3269 ( \3960 , \3958 , \3959 );
nand \U$3270 ( \3961 , \3960 , \3585 );
and \U$3271 ( \3962 , \2814 , \3956 );
nor \U$3272 ( \3963 , \3962 , \2202 );
and \U$3273 ( \3964 , \3961 , \3963 );
and \U$3274 ( \3965 , \3955 , \3964 );
and \U$3275 ( \3966 , \3953 , \3954 );
or \U$3276 ( \3967 , \3965 , \3966 );
xor \U$3277 ( \3968 , \3943 , \3967 );
xor \U$3278 ( \3969 , \3739 , \3744 );
xor \U$3279 ( \3970 , \3969 , \3746 );
and \U$3280 ( \3971 , \3968 , \3970 );
and \U$3281 ( \3972 , \3943 , \3967 );
or \U$3282 ( \3973 , \3971 , \3972 );
not \U$3283 ( \3974 , \3973 );
not \U$3284 ( \3975 , \3974 );
or \U$3285 ( \3976 , \3934 , \3975 );
not \U$3286 ( \3977 , \3603 );
xor \U$3287 ( \3978 , \3658 , \3977 );
xnor \U$3288 ( \3979 , \3978 , \3519 );
nand \U$3289 ( \3980 , \3976 , \3979 );
nand \U$3290 ( \3981 , \3973 , \3932 );
and \U$3291 ( \3982 , \3980 , \3981 );
nor \U$3292 ( \3983 , \3930 , \3982 );
not \U$3293 ( \3984 , \3983 );
or \U$3294 ( \3985 , \3928 , \3984 );
not \U$3295 ( \3986 , \3926 );
nand \U$3296 ( \3987 , \3986 , \3826 );
nand \U$3297 ( \3988 , \3985 , \3987 );
xor \U$3298 ( \3989 , \3893 , \3897 );
and \U$3299 ( \3990 , \3989 , \3924 );
and \U$3300 ( \3991 , \3893 , \3897 );
or \U$3301 ( \3992 , \3990 , \3991 );
not \U$3302 ( \3993 , \3992 );
not \U$3303 ( \3994 , \3836 );
not \U$3304 ( \3995 , \3994 );
not \U$3305 ( \3996 , \3849 );
not \U$3306 ( \3997 , \3996 );
or \U$3307 ( \3998 , \3995 , \3997 );
not \U$3308 ( \3999 , \3854 );
nand \U$3309 ( \4000 , \3998 , \3999 );
nand \U$3310 ( \4001 , \3849 , \3836 );
nand \U$3311 ( \4002 , \4000 , \4001 );
not \U$3312 ( \4003 , \4002 );
and \U$3313 ( \4004 , \3993 , \4003 );
and \U$3314 ( \4005 , \3992 , \4002 );
nor \U$3315 ( \4006 , \4004 , \4005 );
not \U$3316 ( \4007 , \1975 );
not \U$3317 ( \4008 , \3883 );
or \U$3318 ( \4009 , \4007 , \4008 );
nand \U$3319 ( \4010 , \3177 , \1973 );
nand \U$3320 ( \4011 , \4009 , \4010 );
not \U$3321 ( \4012 , \1949 );
not \U$3322 ( \4013 , \3873 );
or \U$3323 ( \4014 , \4012 , \4013 );
nand \U$3324 ( \4015 , \3166 , \1964 );
nand \U$3325 ( \4016 , \4014 , \4015 );
xor \U$3326 ( \4017 , \4011 , \4016 );
or \U$3327 ( \4018 , \3394 , \3866 );
and \U$3328 ( \4019 , \2396 , \1925 );
not \U$3329 ( \4020 , \2396 );
and \U$3330 ( \4021 , \4020 , \1915 );
nor \U$3331 ( \4022 , \4019 , \4021 );
not \U$3332 ( \4023 , \4022 );
or \U$3333 ( \4024 , \4023 , \1928 );
nand \U$3334 ( \4025 , \4018 , \4024 );
xor \U$3335 ( \4026 , \4017 , \4025 );
not \U$3336 ( \4027 , \3920 );
not \U$3337 ( \4028 , \1766 );
or \U$3338 ( \4029 , \4027 , \4028 );
not \U$3339 ( \4030 , \2634 );
not \U$3340 ( \4031 , \1784 );
or \U$3341 ( \4032 , \4030 , \4031 );
nand \U$3342 ( \4033 , \3014 , \2633 );
nand \U$3343 ( \4034 , \4032 , \4033 );
nand \U$3344 ( \4035 , \4034 , \1758 );
nand \U$3345 ( \4036 , \4029 , \4035 );
xor \U$3346 ( \4037 , \4026 , \4036 );
not \U$3347 ( \4038 , \3834 );
not \U$3348 ( \4039 , \2479 );
or \U$3349 ( \4040 , \4038 , \4039 );
and \U$3350 ( \4041 , \2584 , \1744 );
not \U$3351 ( \4042 , \2584 );
and \U$3352 ( \4043 , \4042 , \2202 );
nor \U$3353 ( \4044 , \4041 , \4043 );
nand \U$3354 ( \4045 , \2472 , \4044 );
nand \U$3355 ( \4046 , \4040 , \4045 );
xor \U$3356 ( \4047 , \4037 , \4046 );
not \U$3357 ( \4048 , \3877 );
nor \U$3358 ( \4049 , \4048 , \3885 );
not \U$3359 ( \4050 , \3910 );
not \U$3360 ( \4051 , \2414 );
or \U$3361 ( \4052 , \4050 , \4051 );
not \U$3362 ( \4053 , \2457 );
not \U$3363 ( \4054 , \2408 );
or \U$3364 ( \4055 , \4053 , \4054 );
nand \U$3365 ( \4056 , \2079 , \2461 );
nand \U$3366 ( \4057 , \4055 , \4056 );
nand \U$3367 ( \4058 , \4057 , \2157 );
nand \U$3368 ( \4059 , \4052 , \4058 );
xor \U$3369 ( \4060 , \4049 , \4059 );
nor \U$3370 ( \4061 , \3361 , \3672 );
xor \U$3371 ( \4062 , \4060 , \4061 );
xor \U$3372 ( \4063 , \4047 , \4062 );
not \U$3373 ( \4064 , \3847 );
not \U$3374 ( \4065 , \2536 );
or \U$3375 ( \4066 , \4064 , \4065 );
and \U$3376 ( \4067 , \3506 , \2801 );
not \U$3377 ( \4068 , \3506 );
and \U$3378 ( \4069 , \4068 , \1398 );
nor \U$3379 ( \4070 , \4067 , \4069 );
nand \U$3380 ( \4071 , \4070 , \1605 );
nand \U$3381 ( \4072 , \4066 , \4071 );
not \U$3382 ( \4073 , \3868 );
not \U$3383 ( \4074 , \4073 );
not \U$3384 ( \4075 , \3892 );
or \U$3385 ( \4076 , \4074 , \4075 );
not \U$3386 ( \4077 , \3886 );
nand \U$3387 ( \4078 , \4076 , \4077 );
not \U$3388 ( \4079 , \3892 );
nand \U$3389 ( \4080 , \4079 , \3868 );
nand \U$3390 ( \4081 , \4078 , \4080 );
xor \U$3391 ( \4082 , \4072 , \4081 );
not \U$3392 ( \4083 , \3912 );
not \U$3393 ( \4084 , \3922 );
or \U$3394 ( \4085 , \4083 , \4084 );
or \U$3395 ( \4086 , \3922 , \3912 );
nand \U$3396 ( \4087 , \4086 , \3902 );
nand \U$3397 ( \4088 , \4085 , \4087 );
xor \U$3398 ( \4089 , \4082 , \4088 );
xor \U$3399 ( \4090 , \4063 , \4089 );
xor \U$3400 ( \4091 , \4006 , \4090 );
xor \U$3401 ( \4092 , \3855 , \3859 );
and \U$3402 ( \4093 , \4092 , \3925 );
and \U$3403 ( \4094 , \3855 , \3859 );
or \U$3404 ( \4095 , \4093 , \4094 );
nand \U$3405 ( \4096 , \4091 , \4095 );
nand \U$3406 ( \4097 , \3988 , \4096 );
not \U$3407 ( \4098 , \4097 );
or \U$3408 ( \4099 , \4091 , \4095 );
not \U$3409 ( \4100 , \4099 );
or \U$3410 ( \4101 , \4098 , \4100 );
not \U$3411 ( \4102 , \4002 );
nand \U$3412 ( \4103 , \4102 , \3992 );
not \U$3413 ( \4104 , \4103 );
not \U$3414 ( \4105 , \4090 );
or \U$3415 ( \4106 , \4104 , \4105 );
not \U$3416 ( \4107 , \3992 );
nand \U$3417 ( \4108 , \4107 , \4002 );
nand \U$3418 ( \4109 , \4106 , \4108 );
not \U$3419 ( \4110 , \4109 );
not \U$3420 ( \4111 , \1878 );
not \U$3421 ( \4112 , \4022 );
or \U$3422 ( \4113 , \4111 , \4112 );
nand \U$3423 ( \4114 , \3159 , \1929 );
nand \U$3424 ( \4115 , \4113 , \4114 );
not \U$3425 ( \4116 , \3170 );
not \U$3426 ( \4117 , \3179 );
not \U$3427 ( \4118 , \4117 );
or \U$3428 ( \4119 , \4116 , \4118 );
or \U$3429 ( \4120 , \4117 , \3170 );
nand \U$3430 ( \4121 , \4119 , \4120 );
xor \U$3431 ( \4122 , \4115 , \4121 );
xor \U$3433 ( \4123 , \4122 , 1'b0 );
xor \U$3434 ( \4124 , \4011 , \4016 );
and \U$3435 ( \4125 , \4124 , \4025 );
and \U$3436 ( \4126 , \4011 , \4016 );
or \U$3437 ( \4127 , \4125 , \4126 );
not \U$3438 ( \4128 , \2414 );
not \U$3439 ( \4129 , \4057 );
or \U$3440 ( \4130 , \4128 , \4129 );
nand \U$3441 ( \4131 , \3219 , \2157 );
nand \U$3442 ( \4132 , \4130 , \4131 );
xor \U$3443 ( \4133 , \4127 , \4132 );
not \U$3444 ( \4134 , \4034 );
not \U$3445 ( \4135 , \1766 );
or \U$3446 ( \4136 , \4134 , \4135 );
nand \U$3447 ( \4137 , \3208 , \1758 );
nand \U$3448 ( \4138 , \4136 , \4137 );
xor \U$3449 ( \4139 , \4133 , \4138 );
xor \U$3450 ( \4140 , \4123 , \4139 );
xor \U$3451 ( \4141 , \4049 , \4059 );
and \U$3452 ( \4142 , \4141 , \4061 );
and \U$3453 ( \4143 , \4049 , \4059 );
or \U$3454 ( \4144 , \4142 , \4143 );
xor \U$3455 ( \4145 , \4140 , \4144 );
xor \U$3456 ( \4146 , \4047 , \4062 );
and \U$3457 ( \4147 , \4146 , \4089 );
and \U$3458 ( \4148 , \4047 , \4062 );
or \U$3459 ( \4149 , \4147 , \4148 );
xor \U$3460 ( \4150 , \4145 , \4149 );
xor \U$3461 ( \4151 , \4026 , \4036 );
and \U$3462 ( \4152 , \4151 , \4046 );
and \U$3463 ( \4153 , \4026 , \4036 );
or \U$3464 ( \4154 , \4152 , \4153 );
xor \U$3465 ( \4155 , \4072 , \4081 );
and \U$3466 ( \4156 , \4155 , \4088 );
and \U$3467 ( \4157 , \4072 , \4081 );
or \U$3468 ( \4158 , \4156 , \4157 );
xor \U$3469 ( \4159 , \4154 , \4158 );
not \U$3470 ( \4160 , \4044 );
not \U$3471 ( \4161 , \2479 );
or \U$3472 ( \4162 , \4160 , \4161 );
nand \U$3473 ( \4163 , \2472 , \3231 );
nand \U$3474 ( \4164 , \4162 , \4163 );
and \U$3475 ( \4165 , \1614 , \3714 );
and \U$3476 ( \4166 , \2637 , \3715 );
nor \U$3477 ( \4167 , \4165 , \4166 );
nand \U$3478 ( \4168 , \1612 , \4167 );
xor \U$3479 ( \4169 , \4164 , \4168 );
not \U$3480 ( \4170 , \4070 );
not \U$3481 ( \4171 , \1396 );
or \U$3482 ( \4172 , \4170 , \4171 );
not \U$3483 ( \4173 , \3146 );
not \U$3484 ( \4174 , \2529 );
or \U$3485 ( \4175 , \4173 , \4174 );
nand \U$3486 ( \4176 , \2528 , \3515 );
nand \U$3487 ( \4177 , \4175 , \4176 );
nand \U$3488 ( \4178 , \4177 , \1605 );
nand \U$3489 ( \4179 , \4172 , \4178 );
xnor \U$3490 ( \4180 , \4169 , \4179 );
xnor \U$3491 ( \4181 , \4159 , \4180 );
not \U$3492 ( \4182 , \4181 );
xnor \U$3493 ( \4183 , \4150 , \4182 );
nand \U$3494 ( \4184 , \4110 , \4183 );
nand \U$3495 ( \4185 , \4101 , \4184 );
xor \U$3496 ( \4186 , \3612 , \3639 );
xor \U$3497 ( \4187 , \4186 , \3655 );
or \U$3498 ( \4188 , \2202 , \3585 );
or \U$3499 ( \4189 , \1744 , \3672 );
nand \U$3500 ( \4190 , \4188 , \4189 );
not \U$3501 ( \4191 , \4190 );
not \U$3502 ( \4192 , \2479 );
or \U$3503 ( \4193 , \4191 , \4192 );
nand \U$3504 ( \4194 , \2472 , \3938 );
nand \U$3505 ( \4195 , \4193 , \4194 );
not \U$3506 ( \4196 , \3506 );
not \U$3507 ( \4197 , \2029 );
or \U$3508 ( \4198 , \4196 , \4197 );
nand \U$3509 ( \4199 , \2079 , \3816 );
nand \U$3510 ( \4200 , \4198 , \4199 );
not \U$3511 ( \4201 , \4200 );
not \U$3512 ( \4202 , \2414 );
or \U$3513 ( \4203 , \4201 , \4202 );
nand \U$3514 ( \4204 , \3645 , \2157 );
nand \U$3515 ( \4205 , \4203 , \4204 );
xor \U$3516 ( \4206 , \4195 , \4205 );
not \U$3517 ( \4207 , \1973 );
not \U$3518 ( \4208 , \3617 );
or \U$3519 ( \4209 , \4207 , \4208 );
and \U$3520 ( \4210 , \2795 , \1945 );
not \U$3521 ( \4211 , \2795 );
and \U$3522 ( \4212 , \4211 , \1967 );
or \U$3523 ( \4213 , \4210 , \4212 );
nand \U$3524 ( \4214 , \4213 , \1975 );
nand \U$3525 ( \4215 , \4209 , \4214 );
not \U$3526 ( \4216 , \4215 );
not \U$3527 ( \4217 , \1915 );
not \U$3528 ( \4218 , \3145 );
or \U$3529 ( \4219 , \4217 , \4218 );
nand \U$3530 ( \4220 , \3144 , \1925 );
nand \U$3531 ( \4221 , \4219 , \4220 );
not \U$3532 ( \4222 , \4221 );
not \U$3533 ( \4223 , \1877 );
or \U$3534 ( \4224 , \4222 , \4223 );
nand \U$3535 ( \4225 , \3948 , \1929 );
nand \U$3536 ( \4226 , \4224 , \4225 );
not \U$3537 ( \4227 , \4226 );
or \U$3538 ( \4228 , \4216 , \4227 );
or \U$3539 ( \4229 , \4226 , \4215 );
not \U$3540 ( \4230 , \3636 );
not \U$3541 ( \4231 , \4230 );
not \U$3542 ( \4232 , \1963 );
and \U$3543 ( \4233 , \4231 , \4232 );
not \U$3544 ( \4234 , \1951 );
not \U$3545 ( \4235 , \2532 );
or \U$3546 ( \4236 , \4234 , \4235 );
nand \U$3547 ( \4237 , \2526 , \1872 );
nand \U$3548 ( \4238 , \4236 , \4237 );
and \U$3549 ( \4239 , \4238 , \1949 );
nor \U$3550 ( \4240 , \4233 , \4239 );
not \U$3551 ( \4241 , \4240 );
nand \U$3552 ( \4242 , \4229 , \4241 );
nand \U$3553 ( \4243 , \4228 , \4242 );
and \U$3554 ( \4244 , \4206 , \4243 );
and \U$3555 ( \4245 , \4195 , \4205 );
or \U$3556 ( \4246 , \4244 , \4245 );
xor \U$3557 ( \4247 , \4187 , \4246 );
xor \U$3558 ( \4248 , \3943 , \3967 );
xor \U$3559 ( \4249 , \4248 , \3970 );
and \U$3560 ( \4250 , \4247 , \4249 );
and \U$3561 ( \4251 , \4187 , \4246 );
or \U$3562 ( \4252 , \4250 , \4251 );
and \U$3563 ( \4253 , \3973 , \3933 );
not \U$3564 ( \4254 , \3973 );
and \U$3565 ( \4255 , \4254 , \3932 );
nor \U$3566 ( \4256 , \4253 , \4255 );
xnor \U$3567 ( \4257 , \4256 , \3979 );
xor \U$3568 ( \4258 , \4252 , \4257 );
xor \U$3569 ( \4259 , \3953 , \3954 );
xor \U$3570 ( \4260 , \4259 , \3964 );
nand \U$3571 ( \4261 , \2472 , \3585 );
not \U$3572 ( \4262 , \4261 );
not \U$3573 ( \4263 , \3715 );
not \U$3574 ( \4264 , \2408 );
or \U$3575 ( \4265 , \4263 , \4264 );
nand \U$3576 ( \4266 , \2814 , \3714 );
nand \U$3577 ( \4267 , \4265 , \4266 );
not \U$3578 ( \4268 , \4267 );
not \U$3579 ( \4269 , \2414 );
or \U$3580 ( \4270 , \4268 , \4269 );
nand \U$3581 ( \4271 , \4200 , \2157 );
nand \U$3582 ( \4272 , \4270 , \4271 );
not \U$3583 ( \4273 , \4272 );
not \U$3584 ( \4274 , \4273 );
or \U$3585 ( \4275 , \4262 , \4274 );
nand \U$3586 ( \4276 , \2092 , \1915 );
and \U$3587 ( \4277 , \4276 , \3585 );
and \U$3588 ( \4278 , \1925 , \2089 );
nor \U$3589 ( \4279 , \4277 , \4278 );
and \U$3590 ( \4280 , \2028 , \4279 );
not \U$3591 ( \4281 , \1964 );
not \U$3592 ( \4282 , \4238 );
or \U$3593 ( \4283 , \4281 , \4282 );
not \U$3594 ( \4284 , \1951 );
not \U$3595 ( \4285 , \2633 );
or \U$3596 ( \4286 , \4284 , \4285 );
nand \U$3597 ( \4287 , \2632 , \1872 );
nand \U$3598 ( \4288 , \4286 , \4287 );
nand \U$3599 ( \4289 , \4288 , \1949 );
nand \U$3600 ( \4290 , \4283 , \4289 );
nand \U$3601 ( \4291 , \4280 , \4290 );
not \U$3602 ( \4292 , \4291 );
nand \U$3603 ( \4293 , \4275 , \4292 );
not \U$3604 ( \4294 , \4261 );
nand \U$3605 ( \4295 , \4294 , \4272 );
nand \U$3606 ( \4296 , \4293 , \4295 );
xor \U$3607 ( \4297 , \4260 , \4296 );
xor \U$3608 ( \4298 , \4195 , \4205 );
xor \U$3609 ( \4299 , \4298 , \4243 );
and \U$3610 ( \4300 , \4297 , \4299 );
and \U$3611 ( \4301 , \4260 , \4296 );
or \U$3612 ( \4302 , \4300 , \4301 );
xor \U$3613 ( \4303 , \4187 , \4246 );
xor \U$3614 ( \4304 , \4303 , \4249 );
xor \U$3615 ( \4305 , \4302 , \4304 );
xor \U$3616 ( \4306 , \4215 , \4240 );
xor \U$3617 ( \4307 , \4306 , \4226 );
xor \U$3618 ( \4308 , \4280 , \4290 );
not \U$3619 ( \4309 , \1915 );
not \U$3620 ( \4310 , \3506 );
or \U$3621 ( \4311 , \4309 , \4310 );
not \U$3622 ( \4312 , \3505 );
nand \U$3623 ( \4313 , \4312 , \1925 );
nand \U$3624 ( \4314 , \4311 , \4313 );
not \U$3625 ( \4315 , \4314 );
not \U$3626 ( \4316 , \1878 );
or \U$3627 ( \4317 , \4315 , \4316 );
nand \U$3628 ( \4318 , \4221 , \1929 );
nand \U$3629 ( \4319 , \4317 , \4318 );
not \U$3630 ( \4320 , \4319 );
not \U$3631 ( \4321 , \1975 );
and \U$3632 ( \4322 , \1967 , \2584 );
not \U$3633 ( \4323 , \1967 );
and \U$3634 ( \4324 , \4323 , \2587 );
nor \U$3635 ( \4325 , \4322 , \4324 );
not \U$3636 ( \4326 , \4325 );
or \U$3637 ( \4327 , \4321 , \4326 );
nand \U$3638 ( \4328 , \4213 , \1973 );
nand \U$3639 ( \4329 , \4327 , \4328 );
not \U$3640 ( \4330 , \4329 );
nand \U$3641 ( \4331 , \4320 , \4330 );
and \U$3642 ( \4332 , \4308 , \4331 );
nor \U$3643 ( \4333 , \4320 , \4330 );
nor \U$3644 ( \4334 , \4332 , \4333 );
or \U$3645 ( \4335 , \4307 , \4334 );
xor \U$3646 ( \4336 , \4291 , \4261 );
xnor \U$3647 ( \4337 , \4336 , \4272 );
and \U$3648 ( \4338 , \4334 , \4307 );
or \U$3649 ( \4339 , \4337 , \4338 );
nand \U$3650 ( \4340 , \4335 , \4339 );
xor \U$3651 ( \4341 , \4260 , \4296 );
xor \U$3652 ( \4342 , \4341 , \4299 );
xor \U$3653 ( \4343 , \4340 , \4342 );
not \U$3654 ( \4344 , \1964 );
not \U$3655 ( \4345 , \4288 );
or \U$3656 ( \4346 , \4344 , \4345 );
xor \U$3657 ( \4347 , \1951 , \3143 );
nand \U$3658 ( \4348 , \4347 , \1949 );
nand \U$3659 ( \4349 , \4346 , \4348 );
and \U$3660 ( \4350 , \2099 , \3585 );
xor \U$3661 ( \4351 , \4349 , \4350 );
not \U$3662 ( \4352 , \1929 );
not \U$3663 ( \4353 , \4314 );
or \U$3664 ( \4354 , \4352 , \4353 );
not \U$3665 ( \4355 , \1925 );
not \U$3666 ( \4356 , \3714 );
or \U$3667 ( \4357 , \4355 , \4356 );
nand \U$3668 ( \4358 , \3713 , \1922 );
nand \U$3669 ( \4359 , \4357 , \4358 );
nand \U$3670 ( \4360 , \4359 , \1877 );
nand \U$3671 ( \4361 , \4354 , \4360 );
and \U$3672 ( \4362 , \4351 , \4361 );
and \U$3673 ( \4363 , \4349 , \4350 );
or \U$3674 ( \4364 , \4362 , \4363 );
and \U$3675 ( \4365 , \3585 , \2814 );
not \U$3676 ( \4366 , \3585 );
and \U$3677 ( \4367 , \4366 , \2408 );
nor \U$3678 ( \4368 , \4365 , \4367 );
not \U$3679 ( \4369 , \4368 );
not \U$3680 ( \4370 , \2414 );
or \U$3681 ( \4371 , \4369 , \4370 );
nand \U$3682 ( \4372 , \4267 , \2157 );
nand \U$3683 ( \4373 , \4371 , \4372 );
xor \U$3684 ( \4374 , \4364 , \4373 );
not \U$3685 ( \4375 , \4308 );
not \U$3686 ( \4376 , \4330 );
not \U$3687 ( \4377 , \4319 );
and \U$3688 ( \4378 , \4376 , \4377 );
and \U$3689 ( \4379 , \4319 , \4330 );
nor \U$3690 ( \4380 , \4378 , \4379 );
not \U$3691 ( \4381 , \4380 );
or \U$3692 ( \4382 , \4375 , \4381 );
or \U$3693 ( \4383 , \4308 , \4380 );
nand \U$3694 ( \4384 , \4382 , \4383 );
xor \U$3695 ( \4385 , \4374 , \4384 );
not \U$3696 ( \4386 , \1973 );
not \U$3697 ( \4387 , \4325 );
or \U$3698 ( \4388 , \4386 , \4387 );
and \U$3699 ( \4389 , \1967 , \2532 );
not \U$3700 ( \4390 , \1967 );
and \U$3701 ( \4391 , \4390 , \2526 );
nor \U$3702 ( \4392 , \4389 , \4391 );
not \U$3703 ( \4393 , \4392 );
nand \U$3704 ( \4394 , \4393 , \1975 );
nand \U$3705 ( \4395 , \4388 , \4394 );
or \U$3706 ( \4396 , \1866 , \1951 );
nand \U$3707 ( \4397 , \4396 , \3585 );
nand \U$3708 ( \4398 , \1866 , \1951 );
and \U$3709 ( \4399 , \4397 , \1914 , \4398 );
not \U$3710 ( \4400 , \1964 );
not \U$3711 ( \4401 , \4347 );
or \U$3712 ( \4402 , \4400 , \4401 );
and \U$3713 ( \4403 , \1951 , \4312 );
not \U$3714 ( \4404 , \1951 );
and \U$3715 ( \4405 , \4404 , \3505 );
or \U$3716 ( \4406 , \4403 , \4405 );
nand \U$3717 ( \4407 , \4406 , \1949 );
nand \U$3718 ( \4408 , \4402 , \4407 );
and \U$3719 ( \4409 , \4399 , \4408 );
xor \U$3720 ( \4410 , \4395 , \4409 );
xor \U$3721 ( \4411 , \4349 , \4350 );
xor \U$3722 ( \4412 , \4411 , \4361 );
and \U$3723 ( \4413 , \4410 , \4412 );
and \U$3724 ( \4414 , \4395 , \4409 );
or \U$3725 ( \4415 , \4413 , \4414 );
nor \U$3726 ( \4416 , \4385 , \4415 );
xor \U$3727 ( \4417 , \4399 , \4408 );
not \U$3728 ( \4418 , \4417 );
not \U$3729 ( \4419 , \1929 );
not \U$3730 ( \4420 , \4359 );
or \U$3731 ( \4421 , \4419 , \4420 );
not \U$3732 ( \4422 , \1922 );
not \U$3733 ( \4423 , \3585 );
or \U$3734 ( \4424 , \4422 , \4423 );
nand \U$3735 ( \4425 , \3672 , \1914 );
nand \U$3736 ( \4426 , \4424 , \4425 );
nand \U$3737 ( \4427 , \4426 , \1877 );
nand \U$3738 ( \4428 , \4421 , \4427 );
not \U$3739 ( \4429 , \4428 );
and \U$3740 ( \4430 , \2632 , \1945 );
not \U$3741 ( \4431 , \2632 );
and \U$3742 ( \4432 , \4431 , \1967 );
or \U$3743 ( \4433 , \4430 , \4432 );
and \U$3744 ( \4434 , \4433 , \1975 );
nor \U$3745 ( \4435 , \4392 , \1974 );
nor \U$3746 ( \4436 , \4434 , \4435 );
not \U$3747 ( \4437 , \4436 );
and \U$3748 ( \4438 , \4429 , \4437 );
and \U$3749 ( \4439 , \4428 , \4436 );
nor \U$3750 ( \4440 , \4438 , \4439 );
not \U$3751 ( \4441 , \4440 );
and \U$3752 ( \4442 , \4418 , \4441 );
and \U$3753 ( \4443 , \4440 , \4417 );
nor \U$3754 ( \4444 , \4442 , \4443 );
not \U$3755 ( \4445 , \1975 );
and \U$3756 ( \4446 , \3143 , \1945 );
not \U$3757 ( \4447 , \3143 );
and \U$3758 ( \4448 , \4447 , \1967 );
or \U$3759 ( \4449 , \4446 , \4448 );
not \U$3760 ( \4450 , \4449 );
or \U$3761 ( \4451 , \4445 , \4450 );
nand \U$3762 ( \4452 , \4433 , \1973 );
nand \U$3763 ( \4453 , \4451 , \4452 );
not \U$3764 ( \4454 , \1876 );
nand \U$3765 ( \4455 , \4454 , \3585 );
not \U$3766 ( \4456 , \4455 );
or \U$3767 ( \4457 , \4453 , \4456 );
not \U$3768 ( \4458 , \1949 );
and \U$3769 ( \4459 , \3713 , \1872 );
not \U$3770 ( \4460 , \3713 );
and \U$3771 ( \4461 , \4460 , \1951 );
or \U$3772 ( \4462 , \4459 , \4461 );
not \U$3773 ( \4463 , \4462 );
or \U$3774 ( \4464 , \4458 , \4463 );
nand \U$3775 ( \4465 , \4406 , \1964 );
nand \U$3776 ( \4466 , \4464 , \4465 );
nand \U$3777 ( \4467 , \4457 , \4466 );
nand \U$3778 ( \4468 , \4453 , \4456 );
and \U$3779 ( \4469 , \4467 , \4468 );
nand \U$3780 ( \4470 , \4444 , \4469 );
nand \U$3781 ( \4471 , \1937 , \1945 );
nand \U$3782 ( \4472 , \3585 , \4471 );
and \U$3783 ( \4473 , \1934 , \1967 );
nor \U$3784 ( \4474 , \4473 , \1872 );
and \U$3785 ( \4475 , \4472 , \4474 );
not \U$3786 ( \4476 , \1973 );
not \U$3787 ( \4477 , \4449 );
or \U$3788 ( \4478 , \4476 , \4477 );
and \U$3789 ( \4479 , \3505 , \1945 );
not \U$3790 ( \4480 , \3505 );
and \U$3791 ( \4481 , \4480 , \1967 );
or \U$3792 ( \4482 , \4479 , \4481 );
nand \U$3793 ( \4483 , \4482 , \1975 );
nand \U$3794 ( \4484 , \4478 , \4483 );
and \U$3795 ( \4485 , \4475 , \4484 );
xor \U$3796 ( \4486 , \4455 , \4453 );
xnor \U$3797 ( \4487 , \4486 , \4466 );
xor \U$3798 ( \4488 , \4485 , \4487 );
and \U$3799 ( \4489 , \1951 , \3672 );
not \U$3800 ( \4490 , \1951 );
and \U$3801 ( \4491 , \4490 , \3585 );
nor \U$3802 ( \4492 , \4489 , \4491 );
or \U$3803 ( \4493 , \4492 , \1948 );
not \U$3804 ( \4494 , \4462 );
or \U$3805 ( \4495 , \4494 , \1963 );
nand \U$3806 ( \4496 , \4493 , \4495 );
not \U$3807 ( \4497 , \4496 );
xor \U$3808 ( \4498 , \4475 , \4484 );
not \U$3809 ( \4499 , \4498 );
or \U$3810 ( \4500 , \4497 , \4499 );
or \U$3811 ( \4501 , \4498 , \4496 );
not \U$3812 ( \4502 , \1975 );
xor \U$3813 ( \4503 , \1967 , \3713 );
not \U$3814 ( \4504 , \4503 );
or \U$3815 ( \4505 , \4502 , \4504 );
nand \U$3816 ( \4506 , \4482 , \1973 );
nand \U$3817 ( \4507 , \4505 , \4506 );
nor \U$3818 ( \4508 , \3672 , \1963 );
nor \U$3819 ( \4509 , \4507 , \4508 );
not \U$3820 ( \4510 , \1973 );
not \U$3821 ( \4511 , \4503 );
or \U$3822 ( \4512 , \4510 , \4511 );
nand \U$3823 ( \4513 , \3672 , \1975 );
nand \U$3824 ( \4514 , \4512 , \4513 );
nand \U$3825 ( \4515 , \3585 , \1973 );
and \U$3826 ( \4516 , \4515 , \1967 );
nand \U$3827 ( \4517 , \4514 , \4516 );
or \U$3828 ( \4518 , \4509 , \4517 );
nand \U$3829 ( \4519 , \4507 , \4508 );
nand \U$3830 ( \4520 , \4518 , \4519 );
nand \U$3831 ( \4521 , \4501 , \4520 );
nand \U$3832 ( \4522 , \4500 , \4521 );
and \U$3833 ( \4523 , \4488 , \4522 );
and \U$3834 ( \4524 , \4485 , \4487 );
or \U$3835 ( \4525 , \4523 , \4524 );
and \U$3836 ( \4526 , \4470 , \4525 );
nor \U$3837 ( \4527 , \4444 , \4469 );
nor \U$3838 ( \4528 , \4526 , \4527 );
xor \U$3839 ( \4529 , \4395 , \4409 );
xor \U$3840 ( \4530 , \4529 , \4412 );
not \U$3841 ( \4531 , \4428 );
nand \U$3842 ( \4532 , \4531 , \4436 );
not \U$3843 ( \4533 , \4532 );
not \U$3844 ( \4534 , \4417 );
or \U$3845 ( \4535 , \4533 , \4534 );
not \U$3846 ( \4536 , \4436 );
nand \U$3847 ( \4537 , \4536 , \4428 );
nand \U$3848 ( \4538 , \4535 , \4537 );
nor \U$3849 ( \4539 , \4530 , \4538 );
or \U$3850 ( \4540 , \4528 , \4539 );
nand \U$3851 ( \4541 , \4538 , \4530 );
nand \U$3852 ( \4542 , \4540 , \4541 );
not \U$3853 ( \4543 , \4542 );
or \U$3854 ( \4544 , \4416 , \4543 );
nand \U$3855 ( \4545 , \4385 , \4415 );
nand \U$3856 ( \4546 , \4544 , \4545 );
xor \U$3857 ( \4547 , \4364 , \4373 );
and \U$3858 ( \4548 , \4547 , \4384 );
and \U$3859 ( \4549 , \4364 , \4373 );
or \U$3860 ( \4550 , \4548 , \4549 );
not \U$3861 ( \4551 , \4550 );
not \U$3862 ( \4552 , \4337 );
xor \U$3863 ( \4553 , \4334 , \4307 );
not \U$3864 ( \4554 , \4553 );
and \U$3865 ( \4555 , \4552 , \4554 );
and \U$3866 ( \4556 , \4337 , \4553 );
nor \U$3867 ( \4557 , \4555 , \4556 );
nand \U$3868 ( \4558 , \4551 , \4557 );
nand \U$3869 ( \4559 , \4546 , \4558 );
not \U$3870 ( \4560 , \4557 );
nand \U$3871 ( \4561 , \4560 , \4550 );
nand \U$3872 ( \4562 , \4559 , \4561 );
and \U$3873 ( \4563 , \4343 , \4562 );
and \U$3874 ( \4564 , \4340 , \4342 );
or \U$3875 ( \4565 , \4563 , \4564 );
and \U$3876 ( \4566 , \4305 , \4565 );
and \U$3877 ( \4567 , \4302 , \4304 );
or \U$3878 ( \4568 , \4566 , \4567 );
and \U$3879 ( \4569 , \4258 , \4568 );
and \U$3880 ( \4570 , \4252 , \4257 );
or \U$3881 ( \4571 , \4569 , \4570 );
not \U$3882 ( \4572 , \4096 );
nand \U$3883 ( \4573 , \3930 , \3982 );
nand \U$3884 ( \4574 , \3927 , \4573 );
nor \U$3885 ( \4575 , \4572 , \4574 );
nand \U$3886 ( \4576 , \4571 , \4184 , \4575 );
not \U$3887 ( \4577 , \4183 );
nand \U$3888 ( \4578 , \4577 , \4109 );
nand \U$3889 ( \4579 , \4185 , \4576 , \4578 );
xor \U$3890 ( \4580 , \3203 , \3236 );
xor \U$3891 ( \4581 , \4580 , \3242 );
not \U$3892 ( \4582 , \4164 );
not \U$3893 ( \4583 , \4582 );
not \U$3894 ( \4584 , \4168 );
or \U$3895 ( \4585 , \4583 , \4584 );
nand \U$3896 ( \4586 , \4585 , \4179 );
not \U$3897 ( \4587 , \4168 );
nand \U$3898 ( \4588 , \4587 , \4164 );
nand \U$3899 ( \4589 , \4586 , \4588 );
not \U$3900 ( \4590 , \4589 );
and \U$3902 ( \4591 , \4115 , \4121 );
or \U$3903 ( \4592 , 1'b0 , \4591 );
and \U$3904 ( \4593 , \3506 , \2637 );
not \U$3905 ( \4594 , \3506 );
and \U$3906 ( \4595 , \4594 , \1614 );
nor \U$3907 ( \4596 , \4593 , \4595 );
and \U$3908 ( \4597 , \1612 , \4596 );
xor \U$3909 ( \4598 , \4592 , \4597 );
not \U$3910 ( \4599 , \4177 );
not \U$3911 ( \4600 , \2536 );
or \U$3912 ( \4601 , \4599 , \4600 );
nand \U$3913 ( \4602 , \3090 , \1605 );
nand \U$3914 ( \4603 , \4601 , \4602 );
xor \U$3915 ( \4604 , \4598 , \4603 );
not \U$3916 ( \4605 , \4604 );
or \U$3917 ( \4606 , \4590 , \4605 );
or \U$3918 ( \4607 , \4604 , \4589 );
xor \U$3919 ( \4608 , \4123 , \4139 );
and \U$3920 ( \4609 , \4608 , \4144 );
and \U$3921 ( \4610 , \4123 , \4139 );
or \U$3922 ( \4611 , \4609 , \4610 );
nand \U$3923 ( \4612 , \4607 , \4611 );
nand \U$3924 ( \4613 , \4606 , \4612 );
xor \U$3925 ( \4614 , \4581 , \4613 );
not \U$3926 ( \4615 , \4603 );
not \U$3927 ( \4616 , \4597 );
or \U$3928 ( \4617 , \4615 , \4616 );
or \U$3929 ( \4618 , \4597 , \4603 );
nand \U$3930 ( \4619 , \4618 , \4592 );
nand \U$3931 ( \4620 , \4617 , \4619 );
not \U$3932 ( \4621 , \4620 );
xor \U$3933 ( \4622 , \3185 , \3151 );
xnor \U$3934 ( \4623 , \4622 , \3095 );
not \U$3935 ( \4624 , \4623 );
or \U$3936 ( \4625 , \4621 , \4624 );
or \U$3937 ( \4626 , \4623 , \4620 );
nand \U$3938 ( \4627 , \4625 , \4626 );
xor \U$3939 ( \4628 , \3164 , \3180 );
xor \U$3940 ( \4629 , \4628 , \3182 );
xor \U$3941 ( \4630 , \4127 , \4132 );
and \U$3942 ( \4631 , \4630 , \4138 );
and \U$3943 ( \4632 , \4127 , \4132 );
or \U$3944 ( \4633 , \4631 , \4632 );
xor \U$3945 ( \4634 , \4629 , \4633 );
xor \U$3946 ( \4635 , \3213 , \3223 );
xor \U$3947 ( \4636 , \4635 , \3233 );
and \U$3948 ( \4637 , \4634 , \4636 );
and \U$3949 ( \4638 , \4629 , \4633 );
or \U$3950 ( \4639 , \4637 , \4638 );
and \U$3951 ( \4640 , \4627 , \4639 );
not \U$3952 ( \4641 , \4627 );
not \U$3953 ( \4642 , \4639 );
and \U$3954 ( \4643 , \4641 , \4642 );
nor \U$3955 ( \4644 , \4640 , \4643 );
xor \U$3956 ( \4645 , \4614 , \4644 );
not \U$3957 ( \4646 , \4645 );
xor \U$3958 ( \4647 , \4629 , \4633 );
xor \U$3959 ( \4648 , \4647 , \4636 );
not \U$3960 ( \4649 , \4154 );
not \U$3961 ( \4650 , \4180 );
or \U$3962 ( \4651 , \4649 , \4650 );
or \U$3963 ( \4652 , \4180 , \4154 );
nand \U$3964 ( \4653 , \4652 , \4158 );
nand \U$3965 ( \4654 , \4651 , \4653 );
xor \U$3966 ( \4655 , \4648 , \4654 );
xor \U$3967 ( \4656 , \4589 , \4604 );
xor \U$3968 ( \4657 , \4656 , \4611 );
and \U$3969 ( \4658 , \4655 , \4657 );
and \U$3970 ( \4659 , \4648 , \4654 );
or \U$3971 ( \4660 , \4658 , \4659 );
not \U$3972 ( \4661 , \4660 );
nand \U$3973 ( \4662 , \4646 , \4661 );
xor \U$3974 ( \4663 , \4648 , \4654 );
xor \U$3975 ( \4664 , \4663 , \4657 );
not \U$3976 ( \4665 , \4182 );
not \U$3977 ( \4666 , \4145 );
or \U$3978 ( \4667 , \4665 , \4666 );
not \U$3979 ( \4668 , \4145 );
not \U$3980 ( \4669 , \4668 );
not \U$3981 ( \4670 , \4181 );
or \U$3982 ( \4671 , \4669 , \4670 );
nand \U$3983 ( \4672 , \4671 , \4149 );
nand \U$3984 ( \4673 , \4667 , \4672 );
or \U$3985 ( \4674 , \4664 , \4673 );
nand \U$3986 ( \4675 , \4662 , \4674 );
xor \U$3987 ( \4676 , \2896 , \2860 );
xor \U$3988 ( \4677 , \4676 , \2888 );
not \U$3989 ( \4678 , \4623 );
not \U$3990 ( \4679 , \4620 );
not \U$3991 ( \4680 , \4679 );
or \U$3992 ( \4681 , \4678 , \4680 );
nand \U$3993 ( \4682 , \4681 , \4639 );
not \U$3994 ( \4683 , \4623 );
nand \U$3995 ( \4684 , \4683 , \4620 );
and \U$3996 ( \4685 , \4682 , \4684 );
xor \U$3997 ( \4686 , \4677 , \4685 );
xor \U$3998 ( \4687 , \3187 , \3198 );
xnor \U$3999 ( \4688 , \4687 , \3245 );
xor \U$4000 ( \4689 , \4686 , \4688 );
not \U$4001 ( \4690 , \4581 );
not \U$4002 ( \4691 , \4644 );
nand \U$4003 ( \4692 , \4690 , \4691 );
and \U$4004 ( \4693 , \4692 , \4613 );
not \U$4005 ( \4694 , \4581 );
nor \U$4006 ( \4695 , \4694 , \4691 );
nor \U$4007 ( \4696 , \4693 , \4695 );
nand \U$4008 ( \4697 , \4689 , \4696 );
xor \U$4009 ( \4698 , \3084 , \3247 );
xnor \U$4010 ( \4699 , \4698 , \3252 );
xor \U$4011 ( \4700 , \4677 , \4685 );
and \U$4012 ( \4701 , \4700 , \4688 );
and \U$4013 ( \4702 , \4677 , \4685 );
or \U$4014 ( \4703 , \4701 , \4702 );
nand \U$4015 ( \4704 , \4699 , \4703 );
nand \U$4016 ( \4705 , \4697 , \4704 );
nor \U$4017 ( \4706 , \4675 , \4705 );
and \U$4018 ( \4707 , \4579 , \4706 );
not \U$4019 ( \4708 , \4707 );
or \U$4020 ( \4709 , \3459 , \4708 );
not \U$4021 ( \4710 , \3254 );
nor \U$4022 ( \4711 , \4710 , \3257 );
and \U$4023 ( \4712 , \3082 , \4711 );
nand \U$4024 ( \4713 , \3433 , \3445 );
not \U$4025 ( \4714 , \4713 );
nor \U$4026 ( \4715 , \4712 , \4714 );
not \U$4027 ( \4716 , \4705 );
nand \U$4028 ( \4717 , \4664 , \4673 );
nand \U$4029 ( \4718 , \4645 , \4660 );
nand \U$4030 ( \4719 , \4717 , \4718 );
and \U$4031 ( \4720 , \4719 , \4662 );
nand \U$4032 ( \4721 , \4716 , \4720 );
nor \U$4033 ( \4722 , \4689 , \4696 );
not \U$4034 ( \4723 , \4722 );
not \U$4035 ( \4724 , \4704 );
or \U$4036 ( \4725 , \4723 , \4724 );
or \U$4037 ( \4726 , \4699 , \4703 );
nand \U$4038 ( \4727 , \4725 , \4726 );
not \U$4039 ( \4728 , \3081 );
nand \U$4040 ( \4729 , \4728 , \2958 );
nand \U$4041 ( \4730 , \3448 , \3455 );
nand \U$4042 ( \4731 , \4729 , \4730 );
nor \U$4043 ( \4732 , \4727 , \4731 );
nand \U$4044 ( \4733 , \4715 , \4721 , \4732 );
nor \U$4045 ( \4734 , \3259 , \4731 );
nand \U$4046 ( \4735 , \4715 , \4734 );
and \U$4047 ( \4736 , \4713 , \3456 );
nor \U$4048 ( \4737 , \4736 , \3446 );
nand \U$4049 ( \4738 , \4733 , \4735 , \4737 );
nand \U$4050 ( \4739 , \4709 , \4738 );
not \U$4051 ( \4740 , \3320 );
not \U$4052 ( \4741 , \2465 );
or \U$4053 ( \4742 , \4740 , \4741 );
and \U$4054 ( \4743 , \2150 , \1393 );
not \U$4055 ( \4744 , \2150 );
and \U$4056 ( \4745 , \4744 , \2334 );
nor \U$4057 ( \4746 , \4743 , \4745 );
not \U$4058 ( \4747 , \4746 );
nand \U$4059 ( \4748 , \4747 , \1758 );
nand \U$4060 ( \4749 , \4742 , \4748 );
not \U$4061 ( \4750 , \3400 );
nand \U$4062 ( \4751 , \4750 , \1878 );
nand \U$4063 ( \4752 , \1914 , \1929 );
and \U$4064 ( \4753 , \4751 , \4752 );
xor \U$4065 ( \4754 , \4749 , \4753 );
not \U$4066 ( \4755 , \3329 );
not \U$4067 ( \4756 , \2414 );
or \U$4068 ( \4757 , \4755 , \4756 );
not \U$4069 ( \4758 , \1681 );
not \U$4070 ( \4759 , \2408 );
or \U$4071 ( \4760 , \4758 , \4759 );
nand \U$4072 ( \4761 , \2079 , \1678 );
nand \U$4073 ( \4762 , \4760 , \4761 );
nand \U$4074 ( \4763 , \4762 , \2157 );
nand \U$4075 ( \4764 , \4757 , \4763 );
xor \U$4076 ( \4765 , \4754 , \4764 );
not \U$4077 ( \4766 , \3410 );
not \U$4078 ( \4767 , \1397 );
not \U$4079 ( \4768 , \4767 );
or \U$4080 ( \4769 , \4766 , \4768 );
and \U$4081 ( \4770 , \2273 , \3375 );
not \U$4082 ( \4771 , \2273 );
and \U$4083 ( \4772 , \4771 , \2931 );
nor \U$4084 ( \4773 , \4770 , \4772 );
not \U$4085 ( \4774 , \4773 );
nand \U$4086 ( \4775 , \4774 , \1605 );
nand \U$4087 ( \4776 , \4769 , \4775 );
xor \U$4088 ( \4777 , \4765 , \4776 );
xor \U$4089 ( \4778 , \3322 , \3331 );
and \U$4090 ( \4779 , \4778 , \3343 );
and \U$4091 ( \4780 , \3322 , \3331 );
or \U$4092 ( \4781 , \4779 , \4780 );
xor \U$4093 ( \4782 , \4777 , \4781 );
xor \U$4094 ( \4783 , \3388 , \3418 );
and \U$4095 ( \4784 , \4783 , \3431 );
and \U$4096 ( \4785 , \3388 , \3418 );
or \U$4097 ( \4786 , \4784 , \4785 );
xor \U$4098 ( \4787 , \4782 , \4786 );
and \U$4099 ( \4788 , \2398 , \2919 );
not \U$4100 ( \4789 , \2398 );
and \U$4101 ( \4790 , \4789 , \1610 );
nor \U$4102 ( \4791 , \4788 , \4790 );
nand \U$4103 ( \4792 , \1613 , \4791 );
xor \U$4104 ( \4793 , \3392 , \3268 );
and \U$4105 ( \4794 , \4793 , \3402 );
and \U$4106 ( \4795 , \3392 , \3268 );
or \U$4107 ( \4796 , \4794 , \4795 );
not \U$4108 ( \4797 , \3341 );
not \U$4109 ( \4798 , \2479 );
or \U$4110 ( \4799 , \4797 , \4798 );
and \U$4111 ( \4800 , \1744 , \1824 );
and \U$4112 ( \4801 , \2202 , \1823 );
nor \U$4113 ( \4802 , \4800 , \4801 );
not \U$4114 ( \4803 , \4802 );
nand \U$4115 ( \4804 , \4803 , \2472 );
nand \U$4116 ( \4805 , \4799 , \4804 );
xor \U$4117 ( \4806 , \4796 , \4805 );
xnor \U$4118 ( \4807 , \4792 , \4806 );
xor \U$4119 ( \4808 , \3403 , \3412 );
and \U$4120 ( \4809 , \4808 , \3417 );
and \U$4121 ( \4810 , \3403 , \3412 );
or \U$4122 ( \4811 , \4809 , \4810 );
xor \U$4123 ( \4812 , \4807 , \4811 );
xor \U$4124 ( \4813 , \3277 , \3309 );
and \U$4125 ( \4814 , \4813 , \3344 );
and \U$4126 ( \4815 , \3277 , \3309 );
or \U$4127 ( \4816 , \4814 , \4815 );
xor \U$4128 ( \4817 , \4812 , \4816 );
and \U$4129 ( \4818 , \4787 , \4817 );
and \U$4130 ( \4819 , \4782 , \4786 );
or \U$4131 ( \4820 , \4818 , \4819 );
xor \U$4132 ( \4821 , \4765 , \4776 );
and \U$4133 ( \4822 , \4821 , \4781 );
and \U$4134 ( \4823 , \4765 , \4776 );
or \U$4135 ( \4824 , \4822 , \4823 );
and \U$4136 ( \4825 , \2199 , \2637 );
not \U$4137 ( \4826 , \2199 );
and \U$4138 ( \4827 , \4826 , \1614 );
nor \U$4139 ( \4828 , \4825 , \4827 );
and \U$4140 ( \4829 , \1613 , \4828 );
not \U$4141 ( \4830 , \3334 );
not \U$4142 ( \4831 , \4802 );
and \U$4143 ( \4832 , \4830 , \4831 );
and \U$4144 ( \4833 , \1731 , \2202 );
not \U$4145 ( \4834 , \1731 );
and \U$4146 ( \4835 , \4834 , \1744 );
nor \U$4147 ( \4836 , \4833 , \4835 );
and \U$4148 ( \4837 , \2472 , \4836 );
nor \U$4149 ( \4838 , \4832 , \4837 );
not \U$4150 ( \4839 , \4762 );
not \U$4151 ( \4840 , \2414 );
or \U$4152 ( \4841 , \4839 , \4840 );
not \U$4153 ( \4842 , \1598 );
not \U$4154 ( \4843 , \2408 );
or \U$4155 ( \4844 , \4842 , \4843 );
nand \U$4156 ( \4845 , \2079 , \1599 );
nand \U$4157 ( \4846 , \4844 , \4845 );
nand \U$4158 ( \4847 , \4846 , \2157 );
nand \U$4159 ( \4848 , \4841 , \4847 );
not \U$4160 ( \4849 , \4848 );
and \U$4161 ( \4850 , \4838 , \4849 );
not \U$4162 ( \4851 , \4838 );
and \U$4163 ( \4852 , \4851 , \4848 );
nor \U$4164 ( \4853 , \4850 , \4852 );
xor \U$4165 ( \4854 , \4829 , \4853 );
not \U$4166 ( \4855 , \4854 );
not \U$4167 ( \4856 , \4855 );
not \U$4168 ( \4857 , \4805 );
not \U$4169 ( \4858 , \4857 );
not \U$4170 ( \4859 , \4792 );
or \U$4171 ( \4860 , \4858 , \4859 );
nand \U$4172 ( \4861 , \4860 , \4796 );
not \U$4173 ( \4862 , \4792 );
nand \U$4174 ( \4863 , \4862 , \4805 );
and \U$4175 ( \4864 , \4861 , \4863 );
not \U$4176 ( \4865 , \4864 );
not \U$4177 ( \4866 , \4865 );
or \U$4178 ( \4867 , \4856 , \4866 );
nand \U$4179 ( \4868 , \4864 , \4854 );
nand \U$4180 ( \4869 , \4867 , \4868 );
and \U$4181 ( \4870 , \3394 , \1928 );
nor \U$4182 ( \4871 , \4870 , \1915 );
xor \U$4183 ( \4872 , \4753 , \4871 );
not \U$4184 ( \4873 , \1765 );
not \U$4185 ( \4874 , \4746 );
and \U$4186 ( \4875 , \4873 , \4874 );
xor \U$4187 ( \4876 , \1913 , \1393 );
nor \U$4188 ( \4877 , \4876 , \1759 );
nor \U$4189 ( \4878 , \4875 , \4877 );
xor \U$4190 ( \4879 , \4872 , \4878 );
or \U$4191 ( \4880 , \4749 , \4753 );
nand \U$4192 ( \4881 , \4880 , \4764 );
nand \U$4193 ( \4882 , \4749 , \4753 );
and \U$4194 ( \4883 , \4881 , \4882 );
xor \U$4195 ( \4884 , \4879 , \4883 );
nor \U$4196 ( \4885 , \1397 , \4773 );
not \U$4197 ( \4886 , \1605 );
and \U$4198 ( \4887 , \3318 , \3375 );
not \U$4199 ( \4888 , \3318 );
and \U$4200 ( \4889 , \4888 , \2931 );
nor \U$4201 ( \4890 , \4887 , \4889 );
nor \U$4202 ( \4891 , \4886 , \4890 );
nor \U$4203 ( \4892 , \4885 , \4891 );
xor \U$4204 ( \4893 , \4884 , \4892 );
not \U$4205 ( \4894 , \4893 );
and \U$4206 ( \4895 , \4869 , \4894 );
not \U$4207 ( \4896 , \4869 );
and \U$4208 ( \4897 , \4896 , \4893 );
nor \U$4209 ( \4898 , \4895 , \4897 );
xor \U$4210 ( \4899 , \4824 , \4898 );
xor \U$4211 ( \4900 , \4807 , \4811 );
and \U$4212 ( \4901 , \4900 , \4816 );
and \U$4213 ( \4902 , \4807 , \4811 );
or \U$4214 ( \4903 , \4901 , \4902 );
xor \U$4215 ( \4904 , \4899 , \4903 );
nor \U$4216 ( \4905 , \4820 , \4904 );
buf \U$4217 ( \4906 , \4905 );
not \U$4218 ( \4907 , \4906 );
xor \U$4219 ( \4908 , \4782 , \4786 );
xor \U$4220 ( \4909 , \4908 , \4817 );
xor \U$4221 ( \4910 , \3345 , \3383 );
and \U$4222 ( \4911 , \4910 , \3432 );
and \U$4223 ( \4912 , \3345 , \3383 );
or \U$4224 ( \4913 , \4911 , \4912 );
or \U$4225 ( \4914 , \4909 , \4913 );
xor \U$4226 ( \4915 , \4824 , \4898 );
and \U$4227 ( \4916 , \4915 , \4903 );
and \U$4228 ( \4917 , \4824 , \4898 );
or \U$4229 ( \4918 , \4916 , \4917 );
not \U$4230 ( \4919 , \4918 );
or \U$4231 ( \4920 , \1765 , \4876 );
and \U$4232 ( \4921 , \1824 , \1770 );
not \U$4233 ( \4922 , \1824 );
and \U$4234 ( \4923 , \4922 , \2334 );
nor \U$4235 ( \4924 , \4921 , \4923 );
or \U$4236 ( \4925 , \4924 , \1759 );
nand \U$4237 ( \4926 , \4920 , \4925 );
xor \U$4238 ( \4927 , \4753 , \4871 );
and \U$4239 ( \4928 , \4927 , \4878 );
and \U$4240 ( \4929 , \4753 , \4871 );
or \U$4241 ( \4930 , \4928 , \4929 );
xor \U$4242 ( \4931 , \4926 , \4930 );
not \U$4243 ( \4932 , \4890 );
and \U$4244 ( \4933 , \4767 , \4932 );
and \U$4245 ( \4934 , \2151 , \1400 );
not \U$4246 ( \4935 , \2151 );
and \U$4247 ( \4936 , \4935 , \1399 );
nor \U$4248 ( \4937 , \4934 , \4936 );
and \U$4249 ( \4938 , \4937 , \1605 );
nor \U$4250 ( \4939 , \4933 , \4938 );
xor \U$4251 ( \4940 , \4931 , \4939 );
nand \U$4252 ( \4941 , \4864 , \4855 );
nand \U$4253 ( \4942 , \4894 , \4941 );
nand \U$4254 ( \4943 , \4865 , \4854 );
and \U$4255 ( \4944 , \4942 , \4943 );
xor \U$4256 ( \4945 , \4940 , \4944 );
not \U$4257 ( \4946 , \4829 );
nand \U$4258 ( \4947 , \4946 , \4838 );
and \U$4259 ( \4948 , \4947 , \4848 );
nor \U$4260 ( \4949 , \4946 , \4838 );
nor \U$4261 ( \4950 , \4948 , \4949 );
and \U$4262 ( \4951 , \2414 , \4846 );
and \U$4263 ( \4952 , \2079 , \2157 );
nor \U$4264 ( \4953 , \4951 , \4952 );
not \U$4265 ( \4954 , \2878 );
and \U$4266 ( \4955 , \1744 , \1678 );
and \U$4267 ( \4956 , \2202 , \1681 );
nor \U$4268 ( \4957 , \4955 , \4956 );
not \U$4269 ( \4958 , \4957 );
and \U$4270 ( \4959 , \4954 , \4958 );
and \U$4271 ( \4960 , \2479 , \4836 );
nor \U$4272 ( \4961 , \4959 , \4960 );
xor \U$4273 ( \4962 , \4953 , \4961 );
and \U$4274 ( \4963 , \1614 , \2273 );
and \U$4275 ( \4964 , \1680 , \2271 );
nor \U$4276 ( \4965 , \4963 , \4964 );
nand \U$4277 ( \4966 , \1613 , \4965 );
xor \U$4278 ( \4967 , \4962 , \4966 );
xor \U$4279 ( \4968 , \4950 , \4967 );
xor \U$4280 ( \4969 , \4879 , \4883 );
and \U$4281 ( \4970 , \4969 , \4892 );
and \U$4282 ( \4971 , \4879 , \4883 );
or \U$4283 ( \4972 , \4970 , \4971 );
xor \U$4284 ( \4973 , \4968 , \4972 );
xor \U$4285 ( \4974 , \4945 , \4973 );
nand \U$4286 ( \4975 , \4919 , \4974 );
xor \U$4287 ( \4976 , \4940 , \4944 );
and \U$4288 ( \4977 , \4976 , \4973 );
and \U$4289 ( \4978 , \4940 , \4944 );
or \U$4290 ( \4979 , \4977 , \4978 );
not \U$4291 ( \4980 , \4926 );
and \U$4292 ( \4981 , \1614 , \3318 );
and \U$4293 ( \4982 , \2637 , \3025 );
nor \U$4294 ( \4983 , \4981 , \4982 );
nand \U$4295 ( \4984 , \1613 , \4983 );
xor \U$4296 ( \4985 , \4980 , \4984 );
and \U$4297 ( \4986 , \4767 , \4937 );
and \U$4298 ( \4987 , \2982 , \1399 );
not \U$4299 ( \4988 , \2982 );
and \U$4300 ( \4989 , \4988 , \1400 );
nor \U$4301 ( \4990 , \4987 , \4989 );
not \U$4302 ( \4991 , \4990 );
and \U$4303 ( \4992 , \4991 , \1605 );
nor \U$4304 ( \4993 , \4986 , \4992 );
xor \U$4305 ( \4994 , \4985 , \4993 );
xor \U$4306 ( \4995 , \4950 , \4967 );
and \U$4307 ( \4996 , \4995 , \4972 );
and \U$4308 ( \4997 , \4950 , \4967 );
or \U$4309 ( \4998 , \4996 , \4997 );
xor \U$4310 ( \4999 , \4994 , \4998 );
not \U$4311 ( \5000 , \4924 );
not \U$4312 ( \5001 , \5000 );
not \U$4313 ( \5002 , \1766 );
or \U$4314 ( \5003 , \5001 , \5002 );
and \U$4315 ( \5004 , \1730 , \1770 );
not \U$4316 ( \5005 , \1730 );
and \U$4317 ( \5006 , \5005 , \3669 );
nor \U$4318 ( \5007 , \5004 , \5006 );
nand \U$4319 ( \5008 , \5007 , \1758 );
nand \U$4320 ( \5009 , \5003 , \5008 );
nand \U$4321 ( \5010 , \3758 , \3766 );
and \U$4322 ( \5011 , \5010 , \2079 );
xor \U$4323 ( \5012 , \5009 , \5011 );
not \U$4324 ( \5013 , \2472 );
or \U$4325 ( \5014 , \2202 , \1601 );
or \U$4326 ( \5015 , \1744 , \1599 );
nand \U$4327 ( \5016 , \5014 , \5015 );
not \U$4328 ( \5017 , \5016 );
or \U$4329 ( \5018 , \5013 , \5017 );
not \U$4330 ( \5019 , \4957 );
nand \U$4331 ( \5020 , \5019 , \2479 );
nand \U$4332 ( \5021 , \5018 , \5020 );
xor \U$4333 ( \5022 , \5012 , \5021 );
xor \U$4334 ( \5023 , \4953 , \4961 );
and \U$4335 ( \5024 , \5023 , \4966 );
and \U$4336 ( \5025 , \4953 , \4961 );
or \U$4337 ( \5026 , \5024 , \5025 );
xor \U$4338 ( \5027 , \5022 , \5026 );
xor \U$4339 ( \5028 , \4926 , \4930 );
and \U$4340 ( \5029 , \5028 , \4939 );
and \U$4341 ( \5030 , \4926 , \4930 );
or \U$4342 ( \5031 , \5029 , \5030 );
xor \U$4343 ( \5032 , \5027 , \5031 );
xor \U$4344 ( \5033 , \4999 , \5032 );
nand \U$4345 ( \5034 , \4979 , \5033 );
nand \U$4346 ( \5035 , \4907 , \4914 , \4975 , \5034 );
not \U$4347 ( \5036 , \5035 );
nand \U$4348 ( \5037 , \4739 , \5036 );
xor \U$4349 ( \5038 , \1789 , \1839 );
xor \U$4350 ( \5039 , \5038 , \1842 );
not \U$4351 ( \5040 , \5007 );
or \U$4352 ( \5041 , \1767 , \5040 );
and \U$4353 ( \5042 , \3014 , \1678 );
and \U$4354 ( \5043 , \2334 , \1681 );
nor \U$4355 ( \5044 , \5042 , \5043 );
or \U$4356 ( \5045 , \5044 , \1759 );
nand \U$4357 ( \5046 , \5041 , \5045 );
or \U$4358 ( \5047 , \1767 , \5044 );
or \U$4359 ( \5048 , \1786 , \1759 );
nand \U$4360 ( \5049 , \5047 , \5048 );
xor \U$4361 ( \5050 , \5046 , \5049 );
not \U$4362 ( \5051 , \2878 );
not \U$4363 ( \5052 , \3334 );
or \U$4364 ( \5053 , \5051 , \5052 );
not \U$4365 ( \5054 , \2202 );
nand \U$4366 ( \5055 , \5053 , \5054 );
and \U$4367 ( \5056 , \5050 , \5055 );
and \U$4368 ( \5057 , \5046 , \5049 );
or \U$4369 ( \5058 , \5056 , \5057 );
xor \U$4370 ( \5059 , \1790 , \1828 );
xor \U$4371 ( \5060 , \5059 , \1836 );
xor \U$4372 ( \5061 , \5058 , \5060 );
and \U$4373 ( \5062 , \1614 , \1913 );
and \U$4374 ( \5063 , \1680 , \2982 );
nor \U$4375 ( \5064 , \5062 , \5063 );
and \U$4376 ( \5065 , \1613 , \5064 );
and \U$4377 ( \5066 , \1824 , \1399 );
not \U$4378 ( \5067 , \1824 );
and \U$4379 ( \5068 , \5067 , \1400 );
nor \U$4380 ( \5069 , \5066 , \5068 );
not \U$4381 ( \5070 , \5069 );
not \U$4382 ( \5071 , \4767 );
or \U$4383 ( \5072 , \5070 , \5071 );
nand \U$4384 ( \5073 , \1832 , \1605 );
nand \U$4385 ( \5074 , \5072 , \5073 );
xor \U$4386 ( \5075 , \5065 , \5074 );
not \U$4387 ( \5076 , \5016 );
not \U$4388 ( \5077 , \2479 );
or \U$4389 ( \5078 , \5076 , \5077 );
nand \U$4390 ( \5079 , \2472 , \5054 );
nand \U$4391 ( \5080 , \5078 , \5079 );
not \U$4392 ( \5081 , \5080 );
and \U$4393 ( \5082 , \1614 , \2150 );
and \U$4394 ( \5083 , \2637 , \2151 );
nor \U$4395 ( \5084 , \5082 , \5083 );
nand \U$4396 ( \5085 , \1613 , \5084 );
not \U$4397 ( \5086 , \5085 );
not \U$4398 ( \5087 , \5086 );
or \U$4399 ( \5088 , \5081 , \5087 );
not \U$4400 ( \5089 , \5080 );
not \U$4401 ( \5090 , \5089 );
not \U$4402 ( \5091 , \5085 );
or \U$4403 ( \5092 , \5090 , \5091 );
not \U$4404 ( \5093 , \5046 );
nand \U$4405 ( \5094 , \5092 , \5093 );
nand \U$4406 ( \5095 , \5088 , \5094 );
and \U$4407 ( \5096 , \5075 , \5095 );
and \U$4408 ( \5097 , \5065 , \5074 );
or \U$4409 ( \5098 , \5096 , \5097 );
and \U$4410 ( \5099 , \5061 , \5098 );
and \U$4411 ( \5100 , \5058 , \5060 );
or \U$4412 ( \5101 , \5099 , \5100 );
nor \U$4413 ( \5102 , \5039 , \5101 );
not \U$4414 ( \5103 , \5102 );
xor \U$4415 ( \5104 , \4994 , \4998 );
and \U$4416 ( \5105 , \5104 , \5032 );
and \U$4417 ( \5106 , \4994 , \4998 );
or \U$4418 ( \5107 , \5105 , \5106 );
xor \U$4419 ( \5108 , \5046 , \5080 );
xor \U$4420 ( \5109 , \5108 , \5086 );
xor \U$4421 ( \5110 , \4980 , \4984 );
and \U$4422 ( \5111 , \5110 , \4993 );
and \U$4423 ( \5112 , \4980 , \4984 );
or \U$4424 ( \5113 , \5111 , \5112 );
nor \U$4425 ( \5114 , \5021 , \5009 );
or \U$4426 ( \5115 , \5114 , \5011 );
nand \U$4427 ( \5116 , \5021 , \5009 );
nand \U$4428 ( \5117 , \5115 , \5116 );
not \U$4429 ( \5118 , \5117 );
not \U$4430 ( \5119 , \1397 );
not \U$4431 ( \5120 , \4990 );
and \U$4432 ( \5121 , \5119 , \5120 );
and \U$4433 ( \5122 , \5069 , \1605 );
nor \U$4434 ( \5123 , \5121 , \5122 );
not \U$4435 ( \5124 , \5123 );
or \U$4436 ( \5125 , \5118 , \5124 );
or \U$4437 ( \5126 , \5117 , \5123 );
nand \U$4438 ( \5127 , \5125 , \5126 );
xor \U$4439 ( \5128 , \5113 , \5127 );
xor \U$4440 ( \5129 , \5109 , \5128 );
xor \U$4441 ( \5130 , \5022 , \5026 );
and \U$4442 ( \5131 , \5130 , \5031 );
and \U$4443 ( \5132 , \5022 , \5026 );
or \U$4444 ( \5133 , \5131 , \5132 );
xor \U$4445 ( \5134 , \5129 , \5133 );
nand \U$4446 ( \5135 , \5107 , \5134 );
xor \U$4447 ( \5136 , \5046 , \5049 );
xor \U$4448 ( \5137 , \5136 , \5055 );
xor \U$4449 ( \5138 , \5065 , \5074 );
xor \U$4450 ( \5139 , \5138 , \5095 );
xor \U$4451 ( \5140 , \5137 , \5139 );
not \U$4452 ( \5141 , \5123 );
not \U$4453 ( \5142 , \5113 );
or \U$4454 ( \5143 , \5141 , \5142 );
nand \U$4455 ( \5144 , \5143 , \5117 );
or \U$4456 ( \5145 , \5113 , \5123 );
nand \U$4457 ( \5146 , \5144 , \5145 );
xnor \U$4458 ( \5147 , \5140 , \5146 );
xor \U$4459 ( \5148 , \5109 , \5128 );
and \U$4460 ( \5149 , \5148 , \5133 );
and \U$4461 ( \5150 , \5109 , \5128 );
or \U$4462 ( \5151 , \5149 , \5150 );
nand \U$4463 ( \5152 , \5147 , \5151 );
nand \U$4464 ( \5153 , \5135 , \5152 );
not \U$4465 ( \5154 , \5137 );
not \U$4466 ( \5155 , \5139 );
or \U$4467 ( \5156 , \5154 , \5155 );
or \U$4468 ( \5157 , \5139 , \5137 );
nand \U$4469 ( \5158 , \5157 , \5146 );
nand \U$4470 ( \5159 , \5156 , \5158 );
xor \U$4471 ( \5160 , \5058 , \5060 );
xor \U$4472 ( \5161 , \5160 , \5098 );
nor \U$4473 ( \5162 , \5159 , \5161 );
nor \U$4474 ( \5163 , \5153 , \5162 );
nand \U$4475 ( \5164 , \5103 , \5163 );
buf \U$4476 ( \5165 , \5164 );
or \U$4477 ( \5166 , \5037 , \5165 );
not \U$4478 ( \5167 , \4975 );
nand \U$4479 ( \5168 , \4909 , \4913 );
or \U$4480 ( \5169 , \5168 , \4905 );
nand \U$4481 ( \5170 , \4904 , \4820 );
nand \U$4482 ( \5171 , \5169 , \5170 );
not \U$4483 ( \5172 , \5171 );
or \U$4484 ( \5173 , \5167 , \5172 );
not \U$4485 ( \5174 , \4974 );
nand \U$4486 ( \5175 , \5174 , \4918 );
nand \U$4487 ( \5176 , \5173 , \5175 );
and \U$4488 ( \5177 , \5176 , \5034 );
nor \U$4489 ( \5178 , \4979 , \5033 );
nor \U$4490 ( \5179 , \5177 , \5178 );
not \U$4491 ( \5180 , \5179 );
not \U$4492 ( \5181 , \5164 );
and \U$4493 ( \5182 , \5180 , \5181 );
or \U$4494 ( \5183 , \5107 , \5134 );
not \U$4495 ( \5184 , \5152 );
or \U$4496 ( \5185 , \5183 , \5184 );
or \U$4497 ( \5186 , \5147 , \5151 );
nand \U$4498 ( \5187 , \5185 , \5186 );
not \U$4499 ( \5188 , \5162 );
and \U$4500 ( \5189 , \5187 , \5188 );
and \U$4501 ( \5190 , \5159 , \5161 );
nor \U$4502 ( \5191 , \5189 , \5190 );
or \U$4503 ( \5192 , \5191 , \5102 );
nand \U$4504 ( \5193 , \5039 , \5101 );
nand \U$4505 ( \5194 , \5192 , \5193 );
nor \U$4506 ( \5195 , \5182 , \5194 );
nand \U$4507 ( \5196 , \5166 , \5195 );
and \U$4508 ( \5197 , \1846 , \5196 );
and \U$4509 ( \5198 , \1782 , \1845 );
or \U$4510 ( \5199 , \5197 , \5198 );
xor \U$4511 ( \5200 , \1608 , \1684 );
and \U$4512 ( \5201 , \5200 , \1781 );
and \U$4513 ( \5202 , \1608 , \1684 );
or \U$4514 ( \5203 , \5201 , \5202 );
not \U$4515 ( \5204 , \5203 );
not \U$4516 ( \5205 , \1684 );
and \U$4517 ( \5206 , \1614 , \1599 );
and \U$4518 ( \5207 , \1680 , \1601 );
nor \U$4519 ( \5208 , \5206 , \5207 , \3361 );
not \U$4520 ( \5209 , \5208 );
and \U$4521 ( \5210 , \1397 , \1606 );
nor \U$4522 ( \5211 , \5210 , \1399 );
not \U$4523 ( \5212 , \5211 );
or \U$4524 ( \5213 , \5209 , \5212 );
or \U$4525 ( \5214 , \5211 , \5208 );
nand \U$4526 ( \5215 , \5213 , \5214 );
not \U$4527 ( \5216 , \5215 );
or \U$4528 ( \5217 , \5205 , \5216 );
or \U$4529 ( \5218 , \5215 , \1684 );
nand \U$4530 ( \5219 , \5217 , \5218 );
not \U$4531 ( \5220 , \5219 );
and \U$4532 ( \5221 , \5204 , \5220 );
and \U$4533 ( \5222 , \5203 , \5219 );
nor \U$4534 ( \5223 , \5221 , \5222 );
xnor \U$4535 ( \5224 , \5199 , \5223 );
not \U$4536 ( \5225 , RI995e978_225);
nand \U$4537 ( \5226 , \1531 , \1420 );
not \U$4538 ( \5227 , \5226 );
nand \U$4539 ( \5228 , \1540 , \5227 );
not \U$4540 ( \5229 , \5228 );
not \U$4541 ( \5230 , \5229 );
or \U$4542 ( \5231 , \5225 , \5230 );
nand \U$4543 ( \5232 , \5231 , \1312 );
not \U$4544 ( \5233 , RI89ec550_121);
nor \U$4545 ( \5234 , \5233 , \1497 );
nor \U$4546 ( \5235 , \5232 , \5234 );
and \U$4547 ( \5236 , \1461 , RI994dce0_30);
and \U$4548 ( \5237 , \1505 , RI98abb48_56);
nor \U$4549 ( \5238 , \5236 , \5237 );
nand \U$4550 ( \5239 , \5235 , \5238 );
nand \U$4551 ( \5240 , \1710 , RI8918a98_186);
nand \U$4552 ( \5241 , \1550 , RI89252c0_173);
nand \U$4553 ( \5242 , \1468 , RI98bc7e0_43);
not \U$4554 ( \5243 , \1543 );
nand \U$4555 ( \5244 , \5243 , RI8930cd8_160);
nand \U$4556 ( \5245 , \5240 , \5241 , \5242 , \5244 );
nor \U$4557 ( \5246 , \5239 , \5245 );
nand \U$4558 ( \5247 , \1525 , RI9808390_95);
nand \U$4559 ( \5248 , \1518 , RI8939cc0_147);
not \U$4560 ( \5249 , \1592 );
nand \U$4561 ( \5250 , \5249 , RI890fab0_199);
nand \U$4562 ( \5251 , \1586 , RI98089a8_82);
nand \U$4563 ( \5252 , \5247 , \5248 , \5250 , \5251 );
nand \U$4564 ( \5253 , \2445 , RI99675a0_212);
nand \U$4565 ( \5254 , \1535 , RI9819640_69);
nand \U$4566 ( \5255 , \1557 , RI9776e90_108);
nand \U$4567 ( \5256 , \1577 , RI89464e8_134);
nand \U$4568 ( \5257 , \5253 , \5254 , \5255 , \5256 );
nor \U$4569 ( \5258 , \5252 , \5257 );
nand \U$4570 ( \5259 , \5246 , \5258 );
not \U$4571 ( \5260 , \5259 );
not \U$4572 ( \5261 , RI994e2f8_17);
not \U$4573 ( \5262 , RI994dfb0_24);
not \U$4574 ( \5263 , RI99216b8_614);
nand \U$4575 ( \5264 , \5263 , RI994df38_25);
nor \U$4576 ( \5265 , \5262 , \5264 );
nand \U$4577 ( \5266 , \5265 , RI994e028_23);
nor \U$4578 ( \5267 , \5266 , \1267 );
and \U$4579 ( \5268 , \5267 , RI994e118_21);
nand \U$4580 ( \5269 , \5268 , RI994e190_20);
nor \U$4581 ( \5270 , \5269 , \934 );
nand \U$4582 ( \5271 , \5270 , RI994e280_18);
not \U$4583 ( \5272 , \5271 );
or \U$4584 ( \5273 , \5261 , \5272 );
or \U$4585 ( \5274 , \5271 , RI994e2f8_17);
nand \U$4586 ( \5275 , \5273 , \5274 );
or \U$4587 ( \5276 , \5260 , \5275 );
not \U$4588 ( \5277 , RI8930dc8_158);
nor \U$4589 ( \5278 , \1544 , \5277 );
not \U$4590 ( \5279 , RI9967078_223);
not \U$4591 ( \5280 , \5229 );
or \U$4592 ( \5281 , \5279 , \5280 );
nand \U$4593 ( \5282 , \5281 , \802 );
nor \U$4594 ( \5283 , \5278 , \5282 );
and \U$4595 ( \5284 , \1498 , RI89ec640_119);
and \U$4596 ( \5285 , \1461 , RI994ddd0_28);
nor \U$4597 ( \5286 , \5284 , \5285 );
nand \U$4598 ( \5287 , \5283 , \5286 );
and \U$4599 ( \5288 , \1469 , RI98bc8d0_41);
and \U$4600 ( \5289 , \1586 , RI9808a98_80);
nor \U$4601 ( \5290 , \5288 , \5289 );
not \U$4602 ( \5291 , RI8918b88_184);
nor \U$4603 ( \5292 , \1572 , \5291 );
not \U$4604 ( \5293 , RI89465d8_132);
nor \U$4605 ( \5294 , \1578 , \5293 );
nor \U$4606 ( \5295 , \5292 , \5294 );
nand \U$4607 ( \5296 , \5290 , \5295 );
nor \U$4608 ( \5297 , \5287 , \5296 );
not \U$4609 ( \5298 , \1668 );
not \U$4610 ( \5299 , \829 );
and \U$4611 ( \5300 , \5298 , \5299 );
not \U$4612 ( \5301 , RI9967690_210);
nor \U$4613 ( \5302 , \1565 , \5301 );
nor \U$4614 ( \5303 , \5300 , \5302 );
not \U$4615 ( \5304 , RI8939db0_145);
nor \U$4616 ( \5305 , \1625 , \5304 );
not \U$4617 ( \5306 , RI89253b0_171);
nor \U$4618 ( \5307 , \5306 , \1551 );
nor \U$4619 ( \5308 , \5305 , \5307 );
nand \U$4620 ( \5309 , \5303 , \5308 );
not \U$4621 ( \5310 , \1629 );
not \U$4622 ( \5311 , RI9819730_67);
not \U$4623 ( \5312 , \5311 );
and \U$4624 ( \5313 , \5310 , \5312 );
and \U$4625 ( \5314 , \1593 , RI890fba0_197);
nor \U$4626 ( \5315 , \5313 , \5314 );
not \U$4627 ( \5316 , \1524 );
not \U$4628 ( \5317 , RI9808480_93);
not \U$4629 ( \5318 , \5317 );
and \U$4630 ( \5319 , \5316 , \5318 );
and \U$4631 ( \5320 , \1507 , RI98abc38_54);
nor \U$4632 ( \5321 , \5319 , \5320 );
nand \U$4633 ( \5322 , \5315 , \5321 );
nor \U$4634 ( \5323 , \5309 , \5322 );
nand \U$4635 ( \5324 , \5297 , \5323 );
buf \U$4636 ( \5325 , \5324 );
not \U$4637 ( \5326 , \5271 );
nand \U$4638 ( \5327 , \5326 , RI994e2f8_17);
not \U$4639 ( \5328 , \5327 );
nand \U$4640 ( \5329 , \5328 , RI994e370_16);
and \U$4641 ( \5330 , \5329 , RI994e3e8_15);
nor \U$4642 ( \5331 , \5329 , RI994e3e8_15);
nor \U$4643 ( \5332 , \5330 , \5331 );
nand \U$4644 ( \5333 , \5325 , \5332 );
not \U$4645 ( \5334 , RI994e370_16);
not \U$4646 ( \5335 , \5327 );
or \U$4647 ( \5336 , \5334 , \5335 );
or \U$4648 ( \5337 , \5327 , RI994e370_16);
nand \U$4649 ( \5338 , \5336 , \5337 );
not \U$4650 ( \5339 , \5338 );
not \U$4651 ( \5340 , RI99669e8_224);
not \U$4652 ( \5341 , \5229 );
or \U$4653 ( \5342 , \5340 , \5341 );
nand \U$4654 ( \5343 , \5342 , \1337 );
not \U$4655 ( \5344 , RI8930d50_159);
nor \U$4656 ( \5345 , \5344 , \1544 );
nor \U$4657 ( \5346 , \5343 , \5345 );
not \U$4658 ( \5347 , \1497 );
not \U$4659 ( \5348 , RI89ec5c8_120);
not \U$4660 ( \5349 , \5348 );
and \U$4661 ( \5350 , \5347 , \5349 );
and \U$4662 ( \5351 , \1461 , RI994dd58_29);
nor \U$4663 ( \5352 , \5350 , \5351 );
nand \U$4664 ( \5353 , \5346 , \5352 );
nand \U$4665 ( \5354 , \1657 , RI8946560_133);
nand \U$4666 ( \5355 , \1710 , RI8918b10_185);
nand \U$4667 ( \5356 , \1468 , RI98bc858_42);
nand \U$4668 ( \5357 , \1586 , RI9808a20_81);
nand \U$4669 ( \5358 , \5354 , \5355 , \5356 , \5357 );
nor \U$4670 ( \5359 , \5353 , \5358 );
nand \U$4671 ( \5360 , \1507 , RI98abbc0_55);
nand \U$4672 ( \5361 , \1593 , RI890fb28_198);
nand \U$4673 ( \5362 , \1535 , RI98196b8_68);
nand \U$4674 ( \5363 , \1525 , RI9808408_94);
nand \U$4675 ( \5364 , \5360 , \5361 , \5362 , \5363 );
nand \U$4676 ( \5365 , \1518 , RI8939d38_146);
nand \U$4677 ( \5366 , \1557 , RI9776f08_107);
nand \U$4678 ( \5367 , \1564 , RI9967618_211);
nand \U$4679 ( \5368 , \1550 , RI8925338_172);
nand \U$4680 ( \5369 , \5365 , \5366 , \5367 , \5368 );
nor \U$4681 ( \5370 , \5364 , \5369 );
nand \U$4682 ( \5371 , \5359 , \5370 );
buf \U$4683 ( \5372 , \5371 );
nand \U$4684 ( \5373 , \5339 , \5372 );
nand \U$4685 ( \5374 , \5276 , \5333 , \5373 );
not \U$4686 ( \5375 , \5374 );
nand \U$4687 ( \5376 , \1461 , RI994dc68_31);
nand \U$4688 ( \5377 , \1507 , RI98abad0_57);
and \U$4689 ( \5378 , \5229 , RI995e900_226);
not \U$4690 ( \5379 , \848 );
nor \U$4691 ( \5380 , \5378 , \5379 );
nand \U$4692 ( \5381 , \1498 , RI89ec4d8_122);
nand \U$4693 ( \5382 , \5376 , \5377 , \5380 , \5381 );
nand \U$4694 ( \5383 , \1710 , RI8918a20_187);
nand \U$4695 ( \5384 , \1550 , RI8925248_174);
nand \U$4696 ( \5385 , \1468 , RI98bc768_44);
nand \U$4697 ( \5386 , \5243 , RI8930c60_161);
nand \U$4698 ( \5387 , \5383 , \5384 , \5385 , \5386 );
nor \U$4699 ( \5388 , \5382 , \5387 );
nand \U$4700 ( \5389 , \5249 , RI890fa38_200);
nand \U$4701 ( \5390 , \1518 , RI8939c48_148);
nand \U$4702 ( \5391 , \1525 , RI9808318_96);
nand \U$4703 ( \5392 , \1586 , RI9808930_83);
nand \U$4704 ( \5393 , \5389 , \5390 , \5391 , \5392 );
nand \U$4705 ( \5394 , \2445 , RI9967528_213);
nand \U$4706 ( \5395 , \1535 , RI98195c8_70);
nand \U$4707 ( \5396 , \1557 , RI9776e18_109);
nand \U$4708 ( \5397 , \1577 , RI8946470_135);
nand \U$4709 ( \5398 , \5394 , \5395 , \5396 , \5397 );
nor \U$4710 ( \5399 , \5393 , \5398 );
nand \U$4711 ( \5400 , \5388 , \5399 );
not \U$4712 ( \5401 , \5400 );
nand \U$4713 ( \5402 , \5375 , \5401 );
not \U$4714 ( \5403 , \5270 );
not \U$4715 ( \5404 , \5403 );
not \U$4716 ( \5405 , RI994e280_18);
and \U$4717 ( \5406 , \5404 , \5405 );
and \U$4718 ( \5407 , \5403 , RI994e280_18);
nor \U$4719 ( \5408 , \5406 , \5407 );
or \U$4720 ( \5409 , \5402 , \5408 );
or \U$4721 ( \5410 , \5374 , \5408 );
nand \U$4722 ( \5411 , \5410 , \5402 );
not \U$4723 ( \5412 , RI89ec370_125);
not \U$4724 ( \5413 , \1496 );
or \U$4725 ( \5414 , \5412 , \5413 );
nand \U$4726 ( \5415 , \1467 , RI98abf80_47);
nand \U$4727 ( \5416 , \5414 , \5415 );
not \U$4728 ( \5417 , RI98ab968_60);
not \U$4729 ( \5418 , \1505 );
or \U$4730 ( \5419 , \5417 , \5418 );
nand \U$4731 ( \5420 , \5243 , RI8930af8_164);
nand \U$4732 ( \5421 , \5419 , \5420 );
nor \U$4733 ( \5422 , \5416 , \5421 );
not \U$4734 ( \5423 , RI8946308_138);
not \U$4735 ( \5424 , \1577 );
or \U$4736 ( \5425 , \5423 , \5424 );
nand \U$4737 ( \5426 , \5249 , RI890f8d0_203);
nand \U$4738 ( \5427 , \5425 , \5426 );
not \U$4739 ( \5428 , RI98087c8_86);
not \U$4740 ( \5429 , \1585 );
or \U$4741 ( \5430 , \5428 , \5429 );
nand \U$4742 ( \5431 , \1523 , RI97772c8_99);
nand \U$4743 ( \5432 , \5430 , \5431 );
nor \U$4744 ( \5433 , \5427 , \5432 );
nand \U$4745 ( \5434 , \1562 , RI99673c0_216);
not \U$4746 ( \5435 , \5228 );
nand \U$4747 ( \5436 , \5435 , RI995e798_229);
nand \U$4748 ( \5437 , \5434 , \5436 , \969 );
not \U$4749 ( \5438 , RI98bcc18_34);
not \U$4750 ( \5439 , \1460 );
or \U$4751 ( \5440 , \5438 , \5439 );
nand \U$4752 ( \5441 , \1516 , RI8939ae0_151);
nand \U$4753 ( \5442 , \5440 , \5441 );
nor \U$4754 ( \5443 , \5437 , \5442 );
not \U$4755 ( \5444 , RI89188b8_190);
not \U$4756 ( \5445 , \1571 );
or \U$4757 ( \5446 , \5444 , \5445 );
nand \U$4758 ( \5447 , \1549 , RI89250e0_177);
nand \U$4759 ( \5448 , \5446 , \5447 );
not \U$4760 ( \5449 , RI89ec988_112);
not \U$4761 ( \5450 , \1556 );
or \U$4762 ( \5451 , \5449 , \5450 );
nand \U$4763 ( \5452 , \1533 , RI9819460_73);
nand \U$4764 ( \5453 , \5451 , \5452 );
nor \U$4765 ( \5454 , \5448 , \5453 );
nand \U$4766 ( \5455 , \5422 , \5433 , \5443 , \5454 );
not \U$4767 ( \5456 , \5455 );
not \U$4768 ( \5457 , \5456 );
not \U$4769 ( \5458 , \5457 );
not \U$4770 ( \5459 , RI994e118_21);
not \U$4771 ( \5460 , \5267 );
not \U$4772 ( \5461 , \5460 );
or \U$4773 ( \5462 , \5459 , \5461 );
or \U$4774 ( \5463 , \5460 , RI994e118_21);
nand \U$4775 ( \5464 , \5462 , \5463 );
and \U$4776 ( \5465 , \5458 , \5464 );
nor \U$4777 ( \5466 , \5456 , \5464 );
not \U$4778 ( \5467 , \1543 );
not \U$4779 ( \5468 , RI8930a80_165);
not \U$4780 ( \5469 , \5468 );
and \U$4781 ( \5470 , \5467 , \5469 );
and \U$4782 ( \5471 , \1467 , RI98abf08_48);
nor \U$4783 ( \5472 , \5470 , \5471 );
and \U$4784 ( \5473 , \1516 , RI8939a68_152);
and \U$4785 ( \5474 , \1571 , RI8918840_191);
nor \U$4786 ( \5475 , \5473 , \5474 );
and \U$4787 ( \5476 , RI8925068_178, \1549 );
and \U$4788 ( \5477 , \1560 , \1540 );
and \U$4789 ( \5478 , \5477 , RI9967348_217);
nor \U$4790 ( \5479 , \5476 , \5478 );
nand \U$4791 ( \5480 , \1556 , RI89ec910_113);
nand \U$4792 ( \5481 , \1533 , RI98193e8_74);
and \U$4793 ( \5482 , \5480 , \5481 );
nand \U$4794 ( \5483 , \5472 , \5475 , \5479 , \5482 );
nand \U$4795 ( \5484 , \1460 , RI98bcba0_35);
nand \U$4796 ( \5485 , \1523 , RI9777250_100);
and \U$4797 ( \5486 , \5484 , \5485 );
not \U$4798 ( \5487 , \1585 );
not \U$4799 ( \5488 , \5487 );
not \U$4800 ( \5489 , RI9808750_87);
not \U$4801 ( \5490 , \5489 );
and \U$4802 ( \5491 , \5488 , \5490 );
not \U$4803 ( \5492 , RI995e720_230);
not \U$4804 ( \5493 , \5435 );
or \U$4805 ( \5494 , \5492 , \5493 );
nand \U$4806 ( \5495 , \5494 , \1220 );
nor \U$4807 ( \5496 , \5491 , \5495 );
nand \U$4808 ( \5497 , \1505 , RI98ab8f0_61);
nand \U$4809 ( \5498 , \1496 , RI89ec2f8_126);
and \U$4810 ( \5499 , \5497 , \5498 );
and \U$4811 ( \5500 , \1577 , RI8946290_139);
and \U$4812 ( \5501 , \5249 , RI890f858_204);
nor \U$4813 ( \5502 , \5500 , \5501 );
nand \U$4814 ( \5503 , \5486 , \5496 , \5499 , \5502 );
nor \U$4815 ( \5504 , \5483 , \5503 );
not \U$4816 ( \5505 , \5504 );
buf \U$4817 ( \5506 , \5505 );
not \U$4818 ( \5507 , \5266 );
not \U$4819 ( \5508 , RI994e0a0_22);
and \U$4820 ( \5509 , \5507 , \5508 );
and \U$4821 ( \5510 , \5266 , RI994e0a0_22);
nor \U$4822 ( \5511 , \5509 , \5510 );
nor \U$4823 ( \5512 , \5466 , \5506 , \5511 );
nor \U$4824 ( \5513 , \5465 , \5512 );
not \U$4825 ( \5514 , RI98abff8_46);
not \U$4826 ( \5515 , \1467 );
or \U$4827 ( \5516 , \5514 , \5515 );
not \U$4828 ( \5517 , \1543 );
nand \U$4829 ( \5518 , \5517 , RI8930b70_163);
nand \U$4830 ( \5519 , \5516 , \5518 );
not \U$4831 ( \5520 , RI8925158_176);
not \U$4832 ( \5521 , \1549 );
or \U$4833 ( \5522 , \5520 , \5521 );
nand \U$4834 ( \5523 , \1562 , RI9967438_215);
nand \U$4835 ( \5524 , \5522 , \5523 );
nor \U$4836 ( \5525 , \5519 , \5524 );
not \U$4837 ( \5526 , RI8939b58_150);
not \U$4838 ( \5527 , \1516 );
or \U$4839 ( \5528 , \5526 , \5527 );
nand \U$4840 ( \5529 , \1571 , RI8918930_189);
nand \U$4841 ( \5530 , \5528 , \5529 );
not \U$4842 ( \5531 , RI9776d28_111);
not \U$4843 ( \5532 , \1556 );
or \U$4844 ( \5533 , \5531 , \5532 );
nand \U$4845 ( \5534 , \1533 , RI98194d8_72);
nand \U$4846 ( \5535 , \5533 , \5534 );
nor \U$4847 ( \5536 , \5530 , \5535 );
nand \U$4848 ( \5537 , \1585 , RI9808840_85);
nand \U$4849 ( \5538 , \5435 , RI995e810_228);
nand \U$4850 ( \5539 , \5537 , \5538 , \940 );
not \U$4851 ( \5540 , RI98bcc90_33);
not \U$4852 ( \5541 , \1460 );
or \U$4853 ( \5542 , \5540 , \5541 );
nand \U$4854 ( \5543 , \1523 , RI9808228_98);
nand \U$4855 ( \5544 , \5542 , \5543 );
nor \U$4856 ( \5545 , \5539 , \5544 );
not \U$4857 ( \5546 , RI8946380_137);
not \U$4858 ( \5547 , \1577 );
or \U$4859 ( \5548 , \5546 , \5547 );
nand \U$4860 ( \5549 , \5249 , RI890f948_202);
nand \U$4861 ( \5550 , \5548 , \5549 );
not \U$4862 ( \5551 , RI89ec3e8_124);
not \U$4863 ( \5552 , \1496 );
or \U$4864 ( \5553 , \5551 , \5552 );
nand \U$4865 ( \5554 , \1505 , RI98ab9e0_59);
nand \U$4866 ( \5555 , \5553 , \5554 );
nor \U$4867 ( \5556 , \5550 , \5555 );
nand \U$4868 ( \5557 , \5525 , \5536 , \5545 , \5556 );
not \U$4869 ( \5558 , \5557 );
not \U$4870 ( \5559 , RI994e190_20);
not \U$4871 ( \5560 , \5268 );
not \U$4872 ( \5561 , \5560 );
or \U$4873 ( \5562 , \5559 , \5561 );
or \U$4874 ( \5563 , \5560 , RI994e190_20);
nand \U$4875 ( \5564 , \5562 , \5563 );
or \U$4876 ( \5565 , \5558 , \5564 );
not \U$4877 ( \5566 , RI994e208_19);
not \U$4878 ( \5567 , \5269 );
or \U$4879 ( \5568 , \5566 , \5567 );
or \U$4880 ( \5569 , \5269 , RI994e208_19);
nand \U$4881 ( \5570 , \5568 , \5569 );
not \U$4882 ( \5571 , \5570 );
not \U$4883 ( \5572 , RI995e888_227);
not \U$4884 ( \5573 , \5229 );
or \U$4885 ( \5574 , \5572 , \5573 );
nand \U$4886 ( \5575 , \5574 , \901 );
not \U$4887 ( \5576 , RI89ec460_123);
nor \U$4888 ( \5577 , \5576 , \1497 );
nor \U$4889 ( \5578 , \5575 , \5577 );
not \U$4890 ( \5579 , \1506 );
not \U$4891 ( \5580 , RI98aba58_58);
not \U$4892 ( \5581 , \5580 );
and \U$4893 ( \5582 , \5579 , \5581 );
and \U$4894 ( \5583 , \1461 , RI994dbf0_32);
nor \U$4895 ( \5584 , \5582 , \5583 );
nand \U$4896 ( \5585 , \5578 , \5584 );
nand \U$4897 ( \5586 , \1571 , RI89189a8_188);
nand \U$4898 ( \5587 , \1549 , RI89251d0_175);
nand \U$4899 ( \5588 , \1467 , RI98bc6f0_45);
nand \U$4900 ( \5589 , \5243 , RI8930be8_162);
nand \U$4901 ( \5590 , \5586 , \5587 , \5588 , \5589 );
nor \U$4902 ( \5591 , \5585 , \5590 );
not \U$4903 ( \5592 , \5487 );
nand \U$4904 ( \5593 , \5592 , RI98088b8_84);
nand \U$4905 ( \5594 , \1516 , RI8939bd0_149);
nand \U$4906 ( \5595 , \5249 , RI890f9c0_201);
nand \U$4907 ( \5596 , \1523 , RI98082a0_97);
nand \U$4908 ( \5597 , \5593 , \5594 , \5595 , \5596 );
nand \U$4909 ( \5598 , \1533 , RI9819550_71);
nand \U$4910 ( \5599 , \1577 , RI89463f8_136);
nand \U$4911 ( \5600 , \1557 , RI9776da0_110);
nand \U$4912 ( \5601 , \1562 , RI99674b0_214);
nand \U$4913 ( \5602 , \5598 , \5599 , \5600 , \5601 );
nor \U$4914 ( \5603 , \5597 , \5602 );
nand \U$4915 ( \5604 , \5591 , \5603 );
buf \U$4916 ( \5605 , \5604 );
nand \U$4917 ( \5606 , \5571 , \5605 );
nand \U$4918 ( \5607 , \5565 , \5606 );
or \U$4919 ( \5608 , \5513 , \5607 );
and \U$4920 ( \5609 , \5506 , \5511 );
nor \U$4921 ( \5610 , \5609 , \5607 , \5466 );
nand \U$4922 ( \5611 , \1516 , RI8939978_154);
not \U$4923 ( \5612 , \5435 );
not \U$4924 ( \5613 , \5612 );
and \U$4925 ( \5614 , \5613 , RI995e630_232);
not \U$4926 ( \5615 , \1079 );
nor \U$4927 ( \5616 , \5614 , \5615 );
not \U$4928 ( \5617 , \1437 );
and \U$4929 ( \5618 , \5617 , \1540 );
nand \U$4930 ( \5619 , \5618 , RI8930990_167);
not \U$4931 ( \5620 , \1540 );
nor \U$4932 ( \5621 , \5620 , \1465 );
nand \U$4933 ( \5622 , \5621 , RI8924f78_180);
nand \U$4934 ( \5623 , \5611 , \5616 , \5619 , \5622 );
not \U$4935 ( \5624 , \1455 );
not \U$4936 ( \5625 , \5624 );
nor \U$4937 ( \5626 , \1442 , \5625 );
and \U$4938 ( \5627 , \5626 , \5617 , \1459 );
nand \U$4939 ( \5628 , \5627 , RI98bcab0_37);
and \U$4940 ( \5629 , \1464 , \1582 , \5625 , \1584 );
nand \U$4941 ( \5630 , \5629 , RI89ec208_128);
and \U$4942 ( \5631 , \5626 , \1548 );
nand \U$4943 ( \5632 , \5631 , RI98abe18_50);
nand \U$4944 ( \5633 , \5477 , RI9967258_219);
nand \U$4945 ( \5634 , \5628 , \5630 , \5632 , \5633 );
nor \U$4946 ( \5635 , \5623 , \5634 );
nand \U$4947 ( \5636 , \1505 , RI98ab800_63);
not \U$4948 ( \5637 , \1457 );
and \U$4949 ( \5638 , \1584 , \1582 , \5637 , \1581 );
nand \U$4950 ( \5639 , \5638 , RI9808660_89);
nor \U$4951 ( \5640 , \1494 , \1465 );
nand \U$4952 ( \5641 , \5640 , RI98192f8_76);
and \U$4953 ( \5642 , \1582 , \1464 , \5624 , \1584 );
nand \U$4954 ( \5643 , \5642 , RI9777160_102);
nand \U$4955 ( \5644 , \5636 , \5639 , \5641 , \5643 );
nand \U$4956 ( \5645 , \1577 , RI89461a0_141);
and \U$4957 ( \5646 , \1457 , \1584 , \1582 , \1581 );
nand \U$4958 ( \5647 , \5646 , RI89ec820_115);
and \U$4959 ( \5648 , \1441 , \5624 );
nand \U$4960 ( \5649 , \5648 , \5227 );
not \U$4961 ( \5650 , \5649 );
nand \U$4962 ( \5651 , \5650 , RI890f768_206);
and \U$4963 ( \5652 , \5648 , \1554 );
nand \U$4964 ( \5653 , \5652 , RI8918750_193);
nand \U$4965 ( \5654 , \5645 , \5647 , \5651 , \5653 );
nor \U$4966 ( \5655 , \5644 , \5654 );
nand \U$4967 ( \5656 , \5635 , \5655 );
not \U$4968 ( \5657 , \5656 );
buf \U$4969 ( \5658 , \5657 );
buf \U$4970 ( \5659 , \5658 );
not \U$4971 ( \5660 , RI994dfb0_24);
not \U$4972 ( \5661 , \5264 );
or \U$4973 ( \5662 , \5660 , \5661 );
or \U$4974 ( \5663 , \5264 , RI994dfb0_24);
nand \U$4975 ( \5664 , \5662 , \5663 );
or \U$4976 ( \5665 , \5659 , \5664 );
and \U$4977 ( \5666 , \1112 , RI99216b8_614);
not \U$4978 ( \5667 , \5264 );
nor \U$4979 ( \5668 , \5666 , \5667 );
nand \U$4980 ( \5669 , \5627 , RI98bca38_38);
nand \U$4981 ( \5670 , \5642 , RI97770e8_103);
nand \U$4982 ( \5671 , \5638 , RI98085e8_90);
nand \U$4983 ( \5672 , \5631 , RI98abda0_51);
nand \U$4984 ( \5673 , \5669 , \5670 , \5671 , \5672 );
not \U$4985 ( \5674 , \5673 );
not \U$4986 ( \5675 , \5617 );
nor \U$4987 ( \5676 , \5675 , \1502 );
nand \U$4988 ( \5677 , \5676 , RI98ab788_64);
nand \U$4989 ( \5678 , \5435 , RI995e5b8_233);
nand \U$4990 ( \5679 , \5677 , \5678 , \1134 );
not \U$4991 ( \5680 , RI8924f00_181);
not \U$4992 ( \5681 , \5621 );
or \U$4993 ( \5682 , \5680 , \5681 );
and \U$4994 ( \5683 , \5648 , \5617 );
nand \U$4995 ( \5684 , \5683 , RI8946128_142);
nand \U$4996 ( \5685 , \5682 , \5684 );
nor \U$4997 ( \5686 , \5679 , \5685 );
not \U$4998 ( \5687 , RI8939900_155);
and \U$4999 ( \5688 , \5648 , \1548 );
not \U$5000 ( \5689 , \5688 );
or \U$5001 ( \5690 , \5687 , \5689 );
nand \U$5002 ( \5691 , \5650 , RI890f6f0_207);
nand \U$5003 ( \5692 , \5690 , \5691 );
not \U$5004 ( \5693 , RI99671e0_220);
not \U$5005 ( \5694 , \5477 );
or \U$5006 ( \5695 , \5693 , \5694 );
nand \U$5007 ( \5696 , \5629 , RI89ec190_129);
nand \U$5008 ( \5697 , \5695 , \5696 );
nor \U$5009 ( \5698 , \5692 , \5697 );
not \U$5010 ( \5699 , RI8930918_168);
not \U$5011 ( \5700 , \5618 );
or \U$5012 ( \5701 , \5699 , \5700 );
nand \U$5013 ( \5702 , \5646 , RI89ec7a8_116);
nand \U$5014 ( \5703 , \5701 , \5702 );
not \U$5015 ( \5704 , RI89186d8_194);
not \U$5016 ( \5705 , \5652 );
or \U$5017 ( \5706 , \5704 , \5705 );
nand \U$5018 ( \5707 , \5640 , RI9819280_77);
nand \U$5019 ( \5708 , \5706 , \5707 );
nor \U$5020 ( \5709 , \5703 , \5708 );
nand \U$5021 ( \5710 , \5674 , \5686 , \5698 , \5709 );
buf \U$5022 ( \5711 , \5710 );
not \U$5023 ( \5712 , \5711 );
or \U$5024 ( \5713 , \5668 , \5712 );
not \U$5025 ( \5714 , \5612 );
and \U$5026 ( \5715 , \5714 , RI995e6a8_231);
not \U$5027 ( \5716 , \1022 );
nor \U$5028 ( \5717 , \5715 , \5716 );
nand \U$5029 ( \5718 , \1460 , RI98bcb28_36);
nand \U$5030 ( \5719 , \1516 , RI89399f0_153);
nand \U$5031 ( \5720 , \1562 , RI99672d0_218);
nand \U$5032 ( \5721 , \5717 , \5718 , \5719 , \5720 );
nand \U$5033 ( \5722 , \1549 , RI8924ff0_179);
nand \U$5034 ( \5723 , \1556 , RI89ec898_114);
nand \U$5035 ( \5724 , \1571 , RI89187c8_192);
nand \U$5036 ( \5725 , \1533 , RI9819370_75);
nand \U$5037 ( \5726 , \5722 , \5723 , \5724 , \5725 );
nor \U$5038 ( \5727 , \5721 , \5726 );
nand \U$5039 ( \5728 , \1523 , RI97771d8_101);
nand \U$5040 ( \5729 , \1577 , RI8946218_140);
nand \U$5041 ( \5730 , \5249 , RI890f7e0_205);
nand \U$5042 ( \5731 , \1585 , RI98086d8_88);
nand \U$5043 ( \5732 , \5728 , \5729 , \5730 , \5731 );
nand \U$5044 ( \5733 , \5618 , RI8930a08_166);
nand \U$5045 ( \5734 , \1467 , RI98abe90_49);
nand \U$5046 ( \5735 , \1496 , RI89ec280_127);
nand \U$5047 ( \5736 , \1505 , RI98ab878_62);
nand \U$5048 ( \5737 , \5733 , \5734 , \5735 , \5736 );
nor \U$5049 ( \5738 , \5732 , \5737 );
nand \U$5050 ( \5739 , \5727 , \5738 );
not \U$5051 ( \5740 , \5739 );
buf \U$5052 ( \5741 , \5740 );
not \U$5053 ( \5742 , \5741 );
not \U$5054 ( \5743 , \5265 );
not \U$5055 ( \5744 , \5743 );
not \U$5056 ( \5745 , RI994e028_23);
and \U$5057 ( \5746 , \5744 , \5745 );
and \U$5058 ( \5747 , \5743 , RI994e028_23);
nor \U$5059 ( \5748 , \5746 , \5747 );
nand \U$5060 ( \5749 , \5742 , \5748 );
nand \U$5061 ( \5750 , \5665 , \5713 , \5749 );
and \U$5062 ( \5751 , \5712 , \5668 );
nand \U$5063 ( \5752 , \5435 , RI995e540_234);
nand \U$5064 ( \5753 , \5688 , RI8939888_156);
nand \U$5065 ( \5754 , \5752 , \5753 , \1172 );
not \U$5066 ( \5755 , RI89460b0_143);
not \U$5067 ( \5756 , \5683 );
or \U$5068 ( \5757 , \5755 , \5756 );
nand \U$5069 ( \5758 , \5650 , RI890f678_208);
nand \U$5070 ( \5759 , \5757 , \5758 );
nor \U$5071 ( \5760 , \5754 , \5759 );
not \U$5072 ( \5761 , RI98bc9c0_39);
not \U$5073 ( \5762 , \5627 );
or \U$5074 ( \5763 , \5761 , \5762 );
nand \U$5075 ( \5764 , \5631 , RI98abd28_52);
nand \U$5076 ( \5765 , \5763 , \5764 );
not \U$5077 ( \5766 , RI9967168_221);
not \U$5078 ( \5767 , \5477 );
or \U$5079 ( \5768 , \5766 , \5767 );
nand \U$5080 ( \5769 , \5676 , RI98ab710_65);
nand \U$5081 ( \5770 , \5768 , \5769 );
nor \U$5082 ( \5771 , \5765 , \5770 );
not \U$5083 ( \5772 , RI89308a0_169);
not \U$5084 ( \5773 , \5618 );
or \U$5085 ( \5774 , \5772 , \5773 );
nand \U$5086 ( \5775 , \5621 , RI8924e88_182);
nand \U$5087 ( \5776 , \5774 , \5775 );
not \U$5088 ( \5777 , RI8918660_195);
not \U$5089 ( \5778 , \5652 );
or \U$5090 ( \5779 , \5777 , \5778 );
nand \U$5091 ( \5780 , \5646 , RI89ec730_117);
nand \U$5092 ( \5781 , \5779 , \5780 );
nor \U$5093 ( \5782 , \5776 , \5781 );
not \U$5094 ( \5783 , RI9808570_91);
not \U$5095 ( \5784 , \5638 );
or \U$5096 ( \5785 , \5783 , \5784 );
nand \U$5097 ( \5786 , \5642 , RI9777070_104);
nand \U$5098 ( \5787 , \5785 , \5786 );
not \U$5099 ( \5788 , RI89ec118_130);
not \U$5100 ( \5789 , \5629 );
or \U$5101 ( \5790 , \5788 , \5789 );
nand \U$5102 ( \5791 , \5640 , RI9819208_78);
nand \U$5103 ( \5792 , \5790 , \5791 );
nor \U$5104 ( \5793 , \5787 , \5792 );
nand \U$5105 ( \5794 , \5760 , \5771 , \5782 , \5793 );
nand \U$5106 ( \5795 , \5794 , \1204 );
buf \U$5107 ( \5796 , \5795 );
nor \U$5108 ( \5797 , \5751 , \5796 );
or \U$5109 ( \5798 , \5750 , \5797 );
and \U$5110 ( \5799 , \5749 , \5659 , \5664 );
not \U$5111 ( \5800 , \5748 );
and \U$5112 ( \5801 , \5741 , \5800 );
nor \U$5113 ( \5802 , \5799 , \5801 );
nand \U$5114 ( \5803 , \5798 , \5802 );
nand \U$5115 ( \5804 , \5610 , \5803 );
and \U$5116 ( \5805 , \5606 , \5558 , \5564 );
not \U$5117 ( \5806 , \5605 );
and \U$5118 ( \5807 , \5806 , \5570 );
nor \U$5119 ( \5808 , \5805 , \5807 );
nand \U$5120 ( \5809 , \5608 , \5804 , \5808 );
nand \U$5121 ( \5810 , \5411 , \5809 );
and \U$5122 ( \5811 , \5333 , \5373 );
and \U$5123 ( \5812 , \5811 , \5260 , \5275 );
or \U$5124 ( \5813 , \5325 , \5332 );
not \U$5125 ( \5814 , \5372 );
nand \U$5126 ( \5815 , \5814 , \5333 , \5338 );
nand \U$5127 ( \5816 , \5813 , \5815 );
nor \U$5128 ( \5817 , \5812 , \5816 );
nand \U$5129 ( \5818 , \5409 , \5810 , \5817 );
not \U$5130 ( \5819 , \5818 );
and \U$5131 ( \5820 , \1626 , RI8946038_144);
not \U$5132 ( \5821 , RI8930828_170);
nor \U$5133 ( \5822 , \5821 , \1653 );
nor \U$5134 ( \5823 , \5820 , \5822 );
and \U$5135 ( \5824 , \2622 , RI9776ff8_105);
not \U$5136 ( \5825 , RI890f600_209);
nor \U$5137 ( \5826 , \2160 , \5825 );
nor \U$5138 ( \5827 , \5824 , \5826 );
nand \U$5139 ( \5828 , \5823 , \5827 );
and \U$5140 ( \5829 , \1657 , RI89ec0a0_131);
and \U$5141 ( \5830 , \1710 , RI8924e10_183);
nor \U$5142 ( \5831 , \5829 , \5830 );
not \U$5143 ( \5832 , \1629 );
not \U$5144 ( \5833 , RI98197a8_66);
not \U$5145 ( \5834 , \5833 );
and \U$5146 ( \5835 , \5832 , \5834 );
and \U$5147 ( \5836 , \1593 , RI89185e8_196);
nor \U$5148 ( \5837 , \5835 , \5836 );
nand \U$5149 ( \5838 , \5831 , \5837 );
nor \U$5150 ( \5839 , \5828 , \5838 );
not \U$5151 ( \5840 , RI8939810_157);
nor \U$5152 ( \5841 , \1545 , \5840 );
not \U$5153 ( \5842 , RI99670f0_222);
not \U$5154 ( \5843 , \5229 );
or \U$5155 ( \5844 , \5842 , \5843 );
nand \U$5156 ( \5845 , \5844 , \716 );
nor \U$5157 ( \5846 , \5841 , \5845 );
and \U$5158 ( \5847 , \1471 , RI98bc948_40);
and \U$5159 ( \5848 , \1586 , RI9808b10_79);
nor \U$5160 ( \5849 , \5847 , \5848 );
nand \U$5161 ( \5850 , \5846 , \5849 );
and \U$5162 ( \5851 , \1461 , RI994de48_27);
and \U$5163 ( \5852 , \1499 , RI89ec6b8_118);
nor \U$5164 ( \5853 , \5851 , \5852 );
not \U$5165 ( \5854 , \1508 );
not \U$5166 ( \5855 , RI98abcb0_53);
not \U$5167 ( \5856 , \5855 );
and \U$5168 ( \5857 , \5854 , \5856 );
and \U$5169 ( \5858 , \1525 , RI98084f8_92);
nor \U$5170 ( \5859 , \5857 , \5858 );
nand \U$5171 ( \5860 , \5853 , \5859 );
nor \U$5172 ( \5861 , \5850 , \5860 );
nand \U$5173 ( \5862 , \5839 , \5861 );
not \U$5174 ( \5863 , \5862 );
nor \U$5175 ( \5864 , \5403 , \702 );
xnor \U$5176 ( \5865 , \5864 , RI994e460_14);
not \U$5177 ( \5866 , \796 );
or \U$5178 ( \5867 , \5863 , \5865 , \5866 );
not \U$5179 ( \5868 , \1213 );
not \U$5180 ( \5869 , \5659 );
not \U$5181 ( \5870 , \5869 );
or \U$5182 ( \5871 , \5868 , \5870 );
not \U$5183 ( \5872 , \1969 );
not \U$5184 ( \5873 , \5794 );
not \U$5185 ( \5874 , \5873 );
not \U$5186 ( \5875 , \5874 );
or \U$5187 ( \5876 , \5872 , \5875 );
buf \U$5188 ( \5877 , \1167 );
nand \U$5189 ( \5878 , \5876 , \5877 );
not \U$5190 ( \5879 , \5877 );
nand \U$5191 ( \5880 , \5879 , \5874 , \1969 );
nand \U$5192 ( \5881 , \5880 , \5712 );
nand \U$5193 ( \5882 , \5878 , \5881 );
nand \U$5194 ( \5883 , \5871 , \5882 );
not \U$5195 ( \5884 , \1213 );
nand \U$5196 ( \5885 , \5884 , \5659 );
nand \U$5197 ( \5886 , \5883 , \5885 , \1064 );
nand \U$5198 ( \5887 , \5886 , \5741 );
not \U$5199 ( \5888 , \5883 );
not \U$5200 ( \5889 , \5885 );
or \U$5201 ( \5890 , \5888 , \5889 );
nand \U$5202 ( \5891 , \5890 , \1063 );
nand \U$5203 ( \5892 , \5887 , \5891 );
not \U$5204 ( \5893 , \931 );
nand \U$5205 ( \5894 , \5893 , \5605 );
not \U$5206 ( \5895 , \964 );
nand \U$5207 ( \5896 , \5895 , \5557 );
and \U$5208 ( \5897 , \5894 , \5896 );
not \U$5209 ( \5898 , \1010 );
nand \U$5210 ( \5899 , \5457 , \5898 );
and \U$5211 ( \5900 , \5897 , \5899 );
not \U$5212 ( \5901 , \1266 );
nand \U$5213 ( \5902 , \5901 , \5506 );
nand \U$5214 ( \5903 , \5892 , \5900 , \5902 );
not \U$5215 ( \5904 , \5506 );
nand \U$5216 ( \5905 , \5904 , \5900 , \1266 );
not \U$5217 ( \5906 , \5898 );
and \U$5218 ( \5907 , \5897 , \5458 , \5906 );
not \U$5219 ( \5908 , \931 );
not \U$5220 ( \5909 , \5806 );
or \U$5221 ( \5910 , \5908 , \5909 );
nand \U$5222 ( \5911 , \5894 , \5558 , \964 );
nand \U$5223 ( \5912 , \5910 , \5911 );
nor \U$5224 ( \5913 , \5907 , \5912 );
and \U$5225 ( \5914 , \5903 , \5905 , \5913 );
or \U$5226 ( \5915 , \5401 , \889 );
not \U$5227 ( \5916 , \5260 );
not \U$5228 ( \5917 , \1324 );
and \U$5229 ( \5918 , \5916 , \5917 );
nand \U$5230 ( \5919 , \5372 , \1362 );
nand \U$5231 ( \5920 , \5324 , \835 );
nand \U$5232 ( \5921 , \5919 , \5920 );
nor \U$5233 ( \5922 , \5918 , \5921 );
nand \U$5234 ( \5923 , \5915 , \5922 );
nor \U$5235 ( \5924 , \5914 , \5923 );
not \U$5236 ( \5925 , \5865 );
not \U$5237 ( \5926 , \5862 );
or \U$5238 ( \5927 , \5925 , \5926 );
nor \U$5239 ( \5928 , \5400 , \1291 );
and \U$5240 ( \5929 , \5928 , \5922 );
nor \U$5241 ( \5930 , \5372 , \1362 );
and \U$5242 ( \5931 , \5920 , \5930 );
or \U$5243 ( \5932 , \5325 , \835 );
or \U$5244 ( \5933 , \5862 , \796 );
nand \U$5245 ( \5934 , \5932 , \5933 );
nor \U$5246 ( \5935 , \5931 , \5934 );
nand \U$5247 ( \5936 , \5920 , \5919 , \5260 , \1324 );
nand \U$5248 ( \5937 , \5935 , \5936 );
nor \U$5249 ( \5938 , \5929 , \5937 );
nand \U$5250 ( \5939 , \5927 , \5938 );
or \U$5251 ( \5940 , \5924 , \5939 );
nand \U$5252 ( \5941 , \5867 , \5940 );
not \U$5253 ( \5942 , \5941 );
or \U$5254 ( \5943 , \5819 , \5942 );
not \U$5255 ( \5944 , \5865 );
nand \U$5256 ( \5945 , \5944 , \5938 , \5863 );
or \U$5257 ( \5946 , \5924 , \5945 );
nand \U$5258 ( \5947 , \5943 , \5946 );
buf \U$5259 ( \5948 , \5947 );
nor \U$5260 ( \5949 , \5224 , \5948 );
not \U$5261 ( \5950 , \5949 );
xor \U$5262 ( \5951 , \704 , \5863 );
nand \U$5263 ( \5952 , \5324 , \842 );
not \U$5264 ( \5953 , \5952 );
not \U$5265 ( \5954 , \1334 );
nand \U$5266 ( \5955 , \5954 , \5371 );
nand \U$5267 ( \5956 , \5400 , \845 );
nand \U$5268 ( \5957 , \5259 , \1296 );
nand \U$5269 ( \5958 , \5955 , \5956 , \5957 );
nor \U$5270 ( \5959 , \5953 , \5958 );
not \U$5271 ( \5960 , \5959 );
not \U$5272 ( \5961 , RI994df38_25);
not \U$5273 ( \5962 , \5710 );
or \U$5274 ( \5963 , \5961 , \5962 );
nand \U$5275 ( \5964 , \5963 , \5795 );
not \U$5276 ( \5965 , \5710 );
nand \U$5277 ( \5966 , \5965 , \1112 );
nand \U$5278 ( \5967 , \5964 , \5966 );
nand \U$5279 ( \5968 , \5656 , \1115 );
not \U$5280 ( \5969 , \1019 );
nand \U$5281 ( \5970 , \5969 , \5739 );
nand \U$5282 ( \5971 , \5967 , \5968 , \5970 );
nand \U$5283 ( \5972 , \5657 , \1114 );
not \U$5284 ( \5973 , \5972 );
nand \U$5285 ( \5974 , \5973 , \5970 );
nand \U$5286 ( \5975 , \5740 , \1019 );
nand \U$5287 ( \5976 , \5971 , \5974 , \5975 );
nand \U$5288 ( \5977 , \5505 , \1271 );
nand \U$5289 ( \5978 , \5525 , \5536 , \5545 , \5556 );
nand \U$5290 ( \5979 , \5978 , \965 );
nand \U$5291 ( \5980 , \5455 , \1014 );
and \U$5292 ( \5981 , \5977 , \5979 , \5980 );
nand \U$5293 ( \5982 , \5604 , \936 );
nand \U$5294 ( \5983 , \5976 , \5981 , \5982 );
nor \U$5295 ( \5984 , \5604 , \936 );
nor \U$5296 ( \5985 , \5557 , \965 );
nor \U$5297 ( \5986 , \5984 , \5985 );
not \U$5298 ( \5987 , \5986 );
and \U$5299 ( \5988 , \5980 , \5979 );
nand \U$5300 ( \5989 , \5456 , \1278 );
not \U$5301 ( \5990 , \1271 );
nand \U$5302 ( \5991 , \5990 , \5504 );
nand \U$5303 ( \5992 , \5989 , \5991 );
nand \U$5304 ( \5993 , \5988 , \5992 );
not \U$5305 ( \5994 , \5993 );
or \U$5306 ( \5995 , \5987 , \5994 );
nand \U$5307 ( \5996 , \5995 , \5982 );
nand \U$5308 ( \5997 , \5983 , \5996 );
not \U$5309 ( \5998 , \5997 );
or \U$5310 ( \5999 , \5960 , \5998 );
nor \U$5311 ( \6000 , \5400 , \845 );
nor \U$5312 ( \6001 , \5259 , \1296 );
or \U$5313 ( \6002 , \6000 , \6001 );
nand \U$5314 ( \6003 , \6002 , \5957 );
not \U$5315 ( \6004 , \5955 );
or \U$5316 ( \6005 , \6003 , \6004 );
not \U$5317 ( \6006 , \5371 );
nand \U$5318 ( \6007 , \6006 , \1334 );
nand \U$5319 ( \6008 , \6005 , \6007 );
and \U$5320 ( \6009 , \6008 , \5952 );
nor \U$5321 ( \6010 , \5324 , \842 );
nor \U$5322 ( \6011 , \6009 , \6010 );
nand \U$5323 ( \6012 , \5999 , \6011 );
and \U$5324 ( \6013 , \5951 , \6012 );
and \U$5325 ( \6014 , \704 , \5863 );
or \U$5326 ( \6015 , \6013 , \6014 );
not \U$5327 ( \6016 , \6015 );
not \U$5328 ( \6017 , \1376 );
nand \U$5329 ( \6018 , \6016 , \6017 );
not \U$5330 ( \6019 , \6018 );
and \U$5331 ( \6020 , \6015 , \6017 );
not \U$5332 ( \6021 , \6015 );
and \U$5333 ( \6022 , \6021 , \1376 );
nor \U$5334 ( \6023 , \6020 , \6022 );
not \U$5335 ( \6024 , \6023 );
not \U$5336 ( \6025 , \6024 );
not \U$5337 ( \6026 , \6025 );
or \U$5338 ( \6027 , \6019 , \6026 );
nand \U$5340 ( \6028 , \6027 , 1'b1 );
buf \U$5341 ( \6029 , \6028 );
buf \U$5342 ( \6030 , \6029 );
buf \U$5343 ( \6031 , \6030 );
not \U$5344 ( \6032 , \6018 );
not \U$5345 ( \6033 , \6032 );
buf \U$5346 ( \6034 , \6033 );
buf \U$5347 ( \6035 , \1582 );
not \U$5348 ( \6036 , \1476 );
not \U$5349 ( \6037 , \1581 );
nand \U$5350 ( \6038 , \6036 , \6037 );
nor \U$5351 ( \6039 , \6038 , \1583 );
nand \U$5352 ( \6040 , \6035 , \6039 );
not \U$5353 ( \6041 , \6040 );
not \U$5354 ( \6042 , \6041 );
not \U$5355 ( \6043 , \1584 );
and \U$5356 ( \6044 , \6042 , \6043 );
and \U$5357 ( \6045 , \6041 , \1584 );
nor \U$5358 ( \6046 , \6044 , \6045 );
not \U$5359 ( \6047 , \6046 );
not \U$5360 ( \6048 , \6047 );
not \U$5361 ( \6049 , \1476 );
not \U$5362 ( \6050 , \6037 );
or \U$5363 ( \6051 , \6049 , \6050 );
nand \U$5364 ( \6052 , \1445 , \1449 );
nand \U$5365 ( \6053 , \6051 , \6052 );
not \U$5366 ( \6054 , \6053 );
not \U$5367 ( \6055 , \6039 );
and \U$5368 ( \6056 , \6055 , \6035 );
not \U$5369 ( \6057 , \6055 );
not \U$5370 ( \6058 , \6035 );
and \U$5371 ( \6059 , \6057 , \6058 );
nor \U$5372 ( \6060 , \6056 , \6059 );
nor \U$5373 ( \6061 , \6054 , \6060 );
not \U$5374 ( \6062 , \1583 );
or \U$5375 ( \6063 , \1476 , \1581 );
not \U$5376 ( \6064 , \6063 );
not \U$5377 ( \6065 , \6064 );
or \U$5378 ( \6066 , \6062 , \6065 );
not \U$5379 ( \6067 , \1583 );
nand \U$5380 ( \6068 , \6067 , \6063 );
nand \U$5381 ( \6069 , \6066 , \6068 );
not \U$5382 ( \6070 , \6069 );
and \U$5383 ( \6071 , \6048 , \6061 , \6070 );
buf \U$5384 ( \6072 , \6071 );
and \U$5385 ( \6073 , \6072 , RI992b4b0_349);
not \U$5386 ( \6074 , RI9922bd0_569);
not \U$5387 ( \6075 , \6041 );
or \U$5388 ( \6076 , \6075 , \1584 );
nand \U$5389 ( \6077 , \6076 , \1459 );
not \U$5390 ( \6078 , \6077 );
or \U$5391 ( \6079 , \6074 , \6078 );
not \U$5392 ( \6080 , \1617 );
nand \U$5393 ( \6081 , \6079 , \6080 );
nor \U$5394 ( \6082 , \6073 , \6081 );
nor \U$5395 ( \6083 , \6046 , \6069 );
buf \U$5396 ( \6084 , \6083 );
nand \U$5397 ( \6085 , \6084 , \6061 );
buf \U$5398 ( \6086 , \6085 );
not \U$5399 ( \6087 , \6086 );
not \U$5400 ( \6088 , RI9924ac0_509);
not \U$5401 ( \6089 , \6088 );
and \U$5402 ( \6090 , \6087 , \6089 );
not \U$5403 ( \6091 , \6060 );
nand \U$5404 ( \6092 , \6091 , \6054 );
not \U$5405 ( \6093 , \6092 );
nand \U$5406 ( \6094 , \6084 , \6093 );
buf \U$5407 ( \6095 , \6094 );
not \U$5408 ( \6096 , RI9925ab0_489);
nor \U$5409 ( \6097 , \6095 , \6096 );
nor \U$5410 ( \6098 , \6090 , \6097 );
nand \U$5411 ( \6099 , \6082 , \6098 );
nand \U$5412 ( \6100 , \6046 , \6069 );
not \U$5413 ( \6101 , \6100 );
nand \U$5414 ( \6102 , \6060 , \6053 );
not \U$5415 ( \6103 , \6102 );
nand \U$5416 ( \6104 , \6101 , \6103 );
buf \U$5417 ( \6105 , \6104 );
or \U$5418 ( \6106 , \6105 , \1631 );
nand \U$5419 ( \6107 , \6060 , \6054 );
not \U$5420 ( \6108 , \6107 );
nand \U$5421 ( \6109 , \6101 , \6108 );
buf \U$5422 ( \6110 , \6109 );
or \U$5423 ( \6111 , \6110 , \1622 );
nand \U$5424 ( \6112 , \6101 , \6093 );
buf \U$5425 ( \6113 , \6112 );
not \U$5426 ( \6114 , \6113 );
not \U$5427 ( \6115 , \1670 );
and \U$5428 ( \6116 , \6114 , \6115 );
nand \U$5429 ( \6117 , \6047 , \6069 );
not \U$5430 ( \6118 , \6117 );
nand \U$5431 ( \6119 , \6118 , \6093 );
buf \U$5432 ( \6120 , \6119 );
nor \U$5433 ( \6121 , \6120 , \1673 );
nor \U$5434 ( \6122 , \6116 , \6121 );
nand \U$5435 ( \6123 , \6106 , \6111 , \6122 );
nor \U$5436 ( \6124 , \6099 , \6123 );
and \U$5437 ( \6125 , \6103 , \6083 );
not \U$5438 ( \6126 , \6125 );
not \U$5439 ( \6127 , \6126 );
not \U$5440 ( \6128 , RI9928120_429);
not \U$5441 ( \6129 , \6128 );
and \U$5442 ( \6130 , \6127 , \6129 );
nand \U$5443 ( \6131 , \6084 , \6108 );
buf \U$5444 ( \6132 , \6131 );
not \U$5445 ( \6133 , RI9928a80_409);
nor \U$5446 ( \6134 , \6132 , \6133 );
nor \U$5447 ( \6135 , \6130 , \6134 );
not \U$5448 ( \6136 , \6117 );
nand \U$5449 ( \6137 , \6136 , \6061 );
buf \U$5450 ( \6138 , \6137 );
not \U$5451 ( \6139 , \6138 );
not \U$5452 ( \6140 , \1644 );
and \U$5453 ( \6141 , \6139 , \6140 );
not \U$5454 ( \6142 , \6117 );
nand \U$5455 ( \6143 , \6142 , \6103 );
not \U$5456 ( \6144 , \6143 );
not \U$5457 ( \6145 , \6144 );
nor \U$5458 ( \6146 , \6145 , \1654 );
nor \U$5459 ( \6147 , \6141 , \6146 );
nand \U$5460 ( \6148 , \6135 , \6147 );
nand \U$5461 ( \6149 , \6093 , \6048 , \6070 );
buf \U$5462 ( \6150 , \6149 );
or \U$5463 ( \6151 , \6150 , \1663 );
and \U$5464 ( \6152 , \6103 , \6048 , \6070 );
buf \U$5465 ( \6153 , \6152 );
not \U$5466 ( \6154 , \6153 );
not \U$5467 ( \6155 , \6154 );
nand \U$5468 ( \6156 , \6155 , RI9931ae0_269);
nand \U$5469 ( \6157 , \6101 , \6061 );
buf \U$5470 ( \6158 , \6157 );
not \U$5471 ( \6159 , \6158 );
not \U$5472 ( \6160 , \1618 );
and \U$5473 ( \6161 , \6159 , \6160 );
nand \U$5474 ( \6162 , \6047 , \6069 );
not \U$5475 ( \6163 , \6162 );
nand \U$5476 ( \6164 , \6163 , \6108 );
not \U$5477 ( \6165 , \6164 );
not \U$5478 ( \6166 , \6165 );
nor \U$5479 ( \6167 , \6166 , \1650 );
nor \U$5480 ( \6168 , \6161 , \6167 );
nand \U$5481 ( \6169 , \6151 , \6156 , \6168 );
nor \U$5482 ( \6170 , \6148 , \6169 );
nand \U$5483 ( \6171 , \6124 , \6170 );
buf \U$5484 ( \6172 , \6171 );
buf \U$5485 ( \6173 , \6172 );
not \U$5486 ( \6174 , \6173 );
and \U$5487 ( \6175 , \6034 , \6174 );
not \U$5488 ( \6176 , \6034 );
and \U$5489 ( \6177 , \6176 , \6173 );
nor \U$5490 ( \6178 , \6175 , \6177 );
nand \U$5491 ( \6179 , \6031 , \6178 );
not \U$5492 ( \6180 , \6179 );
nand \U$5493 ( \6181 , \6072 , RI992c6f8_348);
and \U$5494 ( \6182 , \6084 , \6061 );
nand \U$5495 ( \6183 , \6182 , RI9924b38_508);
not \U$5496 ( \6184 , \6094 );
nand \U$5497 ( \6185 , \6184 , RI9925b28_488);
and \U$5498 ( \6186 , \6077 , RI9922f18_568);
not \U$5499 ( \6187 , \1462 );
nor \U$5500 ( \6188 , \6186 , \6187 );
nand \U$5501 ( \6189 , \6181 , \6183 , \6185 , \6188 );
nor \U$5502 ( \6190 , \6117 , \6092 );
buf \U$5503 ( \6191 , \6190 );
nand \U$5504 ( \6192 , \6191 , RI99241d8_528);
not \U$5505 ( \6193 , \6101 );
nor \U$5506 ( \6194 , \6193 , \6092 );
buf \U$5507 ( \6195 , \6194 );
nand \U$5508 ( \6196 , \6195 , RI992abc8_368);
and \U$5509 ( \6197 , \6101 , \6103 );
nand \U$5510 ( \6198 , \6197 , RI992ef48_308);
and \U$5511 ( \6199 , \6101 , \6108 );
nand \U$5512 ( \6200 , \6199 , RI992f8a8_288);
nand \U$5513 ( \6201 , \6192 , \6196 , \6198 , \6200 );
nor \U$5514 ( \6202 , \6189 , \6201 );
not \U$5515 ( \6203 , \6125 );
not \U$5516 ( \6204 , \6203 );
nand \U$5517 ( \6205 , \6204 , RI9928198_428);
not \U$5518 ( \6206 , \6132 );
nand \U$5519 ( \6207 , \6206 , RI9928af8_408);
not \U$5520 ( \6208 , \6061 );
nor \U$5521 ( \6209 , \6208 , \6162 );
buf \U$5522 ( \6210 , \6209 );
nand \U$5523 ( \6211 , \6210 , RI9923878_548);
nor \U$5524 ( \6212 , \6162 , \6107 );
buf \U$5525 ( \6213 , \6212 );
nand \U$5526 ( \6214 , RI9926de8_448, \6213 );
nand \U$5527 ( \6215 , \6205 , \6207 , \6211 , \6214 );
and \U$5528 ( \6216 , \6093 , \6048 , \6070 );
nand \U$5529 ( \6217 , \6216 , RI992d058_328);
nand \U$5530 ( \6218 , \6153 , RI9931b58_268);
nand \U$5531 ( \6219 , \6144 , RI9926488_468);
not \U$5532 ( \6220 , \6157 );
nand \U$5533 ( \6221 , \6220 , RI992a268_388);
nand \U$5534 ( \6222 , \6217 , \6218 , \6219 , \6221 );
nor \U$5535 ( \6223 , \6215 , \6222 );
nand \U$5536 ( \6224 , \6202 , \6223 );
not \U$5537 ( \6225 , \6224 );
and \U$5538 ( \6226 , \6034 , \6225 );
not \U$5539 ( \6227 , \6225 );
and \U$5540 ( \6228 , \6176 , \6227 );
nor \U$5541 ( \6229 , \6226 , \6228 );
nand \U$5542 ( \6230 , \6031 , \6229 );
not \U$5543 ( \6231 , \6230 );
xor \U$5544 ( \6232 , \704 , \5863 );
xor \U$5545 ( \6233 , \6232 , \6012 );
not \U$5546 ( \6234 , \6233 );
not \U$5547 ( \6235 , \6234 );
not \U$5548 ( \6236 , \5958 );
not \U$5549 ( \6237 , \6236 );
not \U$5550 ( \6238 , \5997 );
or \U$5551 ( \6239 , \6237 , \6238 );
not \U$5552 ( \6240 , \6008 );
nand \U$5553 ( \6241 , \6239 , \6240 );
not \U$5554 ( \6242 , \6010 );
nand \U$5555 ( \6243 , \6242 , \5952 );
nor \U$5556 ( \6244 , \6241 , \6243 );
not \U$5557 ( \6245 , \6244 );
nand \U$5558 ( \6246 , \6241 , \6243 );
nand \U$5559 ( \6247 , \6245 , \6246 );
not \U$5560 ( \6248 , \6247 );
or \U$5561 ( \6249 , \6235 , \6248 );
not \U$5562 ( \6250 , \6247 );
nand \U$5563 ( \6251 , \6250 , \6233 );
nand \U$5564 ( \6252 , \6249 , \6251 );
buf \U$5565 ( \6253 , \6252 );
not \U$5566 ( \6254 , \6253 );
not \U$5567 ( \6255 , \6254 );
not \U$5568 ( \6256 , \6234 );
not \U$5569 ( \6257 , \6256 );
not \U$5570 ( \6258 , \6023 );
not \U$5571 ( \6259 , \6258 );
or \U$5572 ( \6260 , \6257 , \6259 );
nand \U$5573 ( \6261 , \6023 , \6234 );
nand \U$5574 ( \6262 , \6260 , \6261 );
not \U$5575 ( \6263 , \6252 );
nand \U$5576 ( \6264 , \6262 , \6263 );
not \U$5577 ( \6265 , \6264 );
buf \U$5578 ( \6266 , \6265 );
not \U$5579 ( \6267 , \6266 );
not \U$5580 ( \6268 , \6267 );
or \U$5581 ( \6269 , \6255 , \6268 );
buf \U$5582 ( \6270 , \6258 );
not \U$5583 ( \6271 , \6270 );
not \U$5584 ( \6272 , \6271 );
not \U$5585 ( \6273 , \6272 );
nand \U$5586 ( \6274 , \6269 , \6273 );
not \U$5587 ( \6275 , \6274 );
or \U$5588 ( \6276 , \6231 , \6275 );
or \U$5589 ( \6277 , \6274 , \6230 );
nand \U$5590 ( \6278 , \6276 , \6277 );
not \U$5591 ( \6279 , \6278 );
or \U$5592 ( \6280 , \6180 , \6279 );
or \U$5593 ( \6281 , \6278 , \6179 );
nand \U$5594 ( \6282 , \6280 , \6281 );
not \U$5595 ( \6283 , \6282 );
not \U$5596 ( \6284 , \6273 );
and \U$5597 ( \6285 , \6227 , \6284 );
not \U$5598 ( \6286 , \6227 );
and \U$5599 ( \6287 , \6286 , \6273 );
nor \U$5600 ( \6288 , \6285 , \6287 );
or \U$5601 ( \6289 , \6267 , \6288 );
or \U$5602 ( \6290 , \6254 , \6284 );
nand \U$5603 ( \6291 , \6289 , \6290 );
xor \U$5604 ( \6292 , \6291 , \6179 );
not \U$5605 ( \6293 , RI9924a48_510);
nor \U$5606 ( \6294 , \6293 , \6086 );
not \U$5607 ( \6295 , RI9925a38_490);
nand \U$5608 ( \6296 , \6084 , \6093 );
not \U$5609 ( \6297 , \6296 );
not \U$5610 ( \6298 , \6297 );
nor \U$5611 ( \6299 , \6295 , \6298 );
nor \U$5612 ( \6300 , \6294 , \6299 );
and \U$5613 ( \6301 , \6072 , RI992b438_350);
nand \U$5614 ( \6302 , \6077 , RI9922b58_570);
nand \U$5615 ( \6303 , \6302 , \1692 );
nor \U$5616 ( \6304 , \6301 , \6303 );
nand \U$5617 ( \6305 , \6300 , \6304 );
nand \U$5618 ( \6306 , \6191 , RI99240e8_530);
nand \U$5619 ( \6307 , \6195 , RI992aad8_370);
nand \U$5620 ( \6308 , \6197 , RI992ee58_310);
nand \U$5621 ( \6309 , \6199 , RI992f7b8_290);
nand \U$5622 ( \6310 , \6306 , \6307 , \6308 , \6309 );
nor \U$5623 ( \6311 , \6305 , \6310 );
nand \U$5624 ( \6312 , \6204 , RI99280a8_430);
not \U$5625 ( \6313 , \6132 );
nand \U$5626 ( \6314 , \6313 , RI9928a08_410);
nand \U$5627 ( \6315 , \6210 , RI9923788_550);
not \U$5628 ( \6316 , \6162 );
nand \U$5629 ( \6317 , \6316 , \6103 );
not \U$5630 ( \6318 , \6317 );
nand \U$5631 ( \6319 , \6318 , RI9926398_470);
nand \U$5632 ( \6320 , \6312 , \6314 , \6315 , \6319 );
nand \U$5633 ( \6321 , \6216 , RI992cf68_330);
nand \U$5634 ( \6322 , \6153 , RI9931a68_270);
nand \U$5635 ( \6323 , \6220 , RI992a178_390);
nand \U$5636 ( \6324 , \6213 , RI9926cf8_450);
nand \U$5637 ( \6325 , \6321 , \6322 , \6323 , \6324 );
nor \U$5638 ( \6326 , \6320 , \6325 );
nand \U$5639 ( \6327 , \6311 , \6326 );
not \U$5640 ( \6328 , \6327 );
and \U$5641 ( \6329 , \6034 , \6328 );
not \U$5642 ( \6330 , \6328 );
and \U$5643 ( \6331 , \6176 , \6330 );
nor \U$5644 ( \6332 , \6329 , \6331 );
nand \U$5645 ( \6333 , \6031 , \6332 );
not \U$5646 ( \6334 , \6333 );
not \U$5647 ( \6335 , \6334 );
not \U$5648 ( \6336 , \6173 );
not \U$5649 ( \6337 , \6284 );
or \U$5650 ( \6338 , \6336 , \6337 );
nand \U$5651 ( \6339 , \6273 , \6174 );
nand \U$5652 ( \6340 , \6338 , \6339 );
not \U$5653 ( \6341 , \6340 );
not \U$5654 ( \6342 , \6341 );
not \U$5655 ( \6343 , \6267 );
and \U$5656 ( \6344 , \6342 , \6343 );
nor \U$5657 ( \6345 , \6288 , \6254 );
nor \U$5658 ( \6346 , \6344 , \6345 );
not \U$5659 ( \6347 , \6346 );
not \U$5660 ( \6348 , \6347 );
or \U$5661 ( \6349 , \6335 , \6348 );
or \U$5662 ( \6350 , \6347 , \6334 );
not \U$5663 ( \6351 , \5956 );
not \U$5664 ( \6352 , \5997 );
or \U$5665 ( \6353 , \6351 , \6352 );
buf \U$5666 ( \6354 , \6000 );
not \U$5667 ( \6355 , \6354 );
nand \U$5668 ( \6356 , \6353 , \6355 );
not \U$5669 ( \6357 , \6001 );
buf \U$5670 ( \6358 , \5957 );
nand \U$5671 ( \6359 , \6357 , \6358 );
nor \U$5672 ( \6360 , \6356 , \6359 );
not \U$5673 ( \6361 , \6360 );
nand \U$5674 ( \6362 , \6356 , \6359 );
nand \U$5675 ( \6363 , \6361 , \6362 );
and \U$5676 ( \6364 , \5956 , \6358 );
not \U$5677 ( \6365 , \6364 );
buf \U$5678 ( \6366 , \5997 );
not \U$5679 ( \6367 , \6366 );
or \U$5680 ( \6368 , \6365 , \6367 );
buf \U$5681 ( \6369 , \6003 );
nand \U$5682 ( \6370 , \6368 , \6369 );
not \U$5683 ( \6371 , \6004 );
nand \U$5684 ( \6372 , \6371 , \6007 );
not \U$5685 ( \6373 , \6372 );
and \U$5686 ( \6374 , \6370 , \6373 );
not \U$5687 ( \6375 , \6370 );
and \U$5688 ( \6376 , \6375 , \6372 );
nor \U$5689 ( \6377 , \6374 , \6376 );
and \U$5690 ( \6378 , \6363 , \6377 );
not \U$5691 ( \6379 , \6363 );
not \U$5692 ( \6380 , \6377 );
and \U$5693 ( \6381 , \6379 , \6380 );
nor \U$5694 ( \6382 , \6378 , \6381 );
buf \U$5695 ( \6383 , \6382 );
buf \U$5696 ( \6384 , \6383 );
not \U$5697 ( \6385 , \6384 );
not \U$5698 ( \6386 , \6385 );
not \U$5699 ( \6387 , \6382 );
not \U$5700 ( \6388 , \6250 );
not \U$5701 ( \6389 , \6377 );
or \U$5702 ( \6390 , \6388 , \6389 );
not \U$5703 ( \6391 , \6247 );
not \U$5704 ( \6392 , \6380 );
or \U$5705 ( \6393 , \6391 , \6392 );
nand \U$5706 ( \6394 , \6390 , \6393 );
nand \U$5707 ( \6395 , \6387 , \6394 );
buf \U$5708 ( \6396 , \6395 );
not \U$5709 ( \6397 , \6396 );
buf \U$5710 ( \6398 , \6397 );
not \U$5711 ( \6399 , \6398 );
not \U$5712 ( \6400 , \6399 );
or \U$5713 ( \6401 , \6386 , \6400 );
not \U$5714 ( \6402 , \6250 );
not \U$5715 ( \6403 , \6402 );
not \U$5716 ( \6404 , \6403 );
nand \U$5717 ( \6405 , \6401 , \6404 );
nand \U$5718 ( \6406 , \6350 , \6405 );
nand \U$5719 ( \6407 , \6349 , \6406 );
and \U$5720 ( \6408 , \6292 , \6407 );
and \U$5721 ( \6409 , \6291 , \6179 );
or \U$5722 ( \6410 , \6408 , \6409 );
not \U$5723 ( \6411 , \6410 );
or \U$5724 ( \6412 , \6283 , \6411 );
or \U$5725 ( \6413 , \6410 , \6282 );
nand \U$5726 ( \6414 , \6412 , \6413 );
not \U$5727 ( \6415 , \6414 );
and \U$5728 ( \6416 , \6225 , \6404 );
not \U$5729 ( \6417 , \6225 );
and \U$5730 ( \6418 , \6417 , \6403 );
nor \U$5731 ( \6419 , \6416 , \6418 );
not \U$5732 ( \6420 , \6419 );
not \U$5733 ( \6421 , \6420 );
not \U$5734 ( \6422 , \6399 );
not \U$5735 ( \6423 , \6422 );
or \U$5736 ( \6424 , \6421 , \6423 );
nand \U$5737 ( \6425 , \6384 , \6404 );
nand \U$5738 ( \6426 , \6424 , \6425 );
not \U$5739 ( \6427 , \6426 );
and \U$5740 ( \6428 , \6405 , \6333 );
not \U$5741 ( \6429 , \6405 );
and \U$5742 ( \6430 , \6429 , \6334 );
or \U$5743 ( \6431 , \6428 , \6430 );
and \U$5744 ( \6432 , \6431 , \6346 );
not \U$5745 ( \6433 , \6431 );
and \U$5746 ( \6434 , \6433 , \6347 );
nor \U$5747 ( \6435 , \6432 , \6434 );
not \U$5748 ( \6436 , \6435 );
not \U$5749 ( \6437 , \6436 );
or \U$5750 ( \6438 , \6427 , \6437 );
not \U$5751 ( \6439 , \6426 );
nand \U$5752 ( \6440 , \6435 , \6439 );
nand \U$5753 ( \6441 , \6125 , RI9928030_431);
not \U$5754 ( \6442 , \6132 );
nand \U$5755 ( \6443 , \6442 , RI9928990_411);
nand \U$5756 ( \6444 , \6210 , RI9923710_551);
nand \U$5757 ( \6445 , \6144 , RI9926320_471);
nand \U$5758 ( \6446 , \6441 , \6443 , \6444 , \6445 );
nand \U$5759 ( \6447 , \6216 , RI992cef0_331);
nand \U$5760 ( \6448 , \6153 , RI99319f0_271);
nand \U$5761 ( \6449 , \6220 , RI992a100_391);
nand \U$5762 ( \6450 , \6213 , RI9926c80_451);
nand \U$5763 ( \6451 , \6447 , \6448 , \6449 , \6450 );
nor \U$5764 ( \6452 , \6446 , \6451 );
nand \U$5765 ( \6453 , \6191 , RI9924070_531);
nand \U$5766 ( \6454 , \6195 , RI992aa60_371);
nand \U$5767 ( \6455 , \6197 , RI992ede0_311);
nand \U$5768 ( \6456 , \6199 , RI992f740_291);
nand \U$5769 ( \6457 , \6453 , \6454 , \6455 , \6456 );
nand \U$5770 ( \6458 , \6184 , RI99259c0_491);
nand \U$5771 ( \6459 , \6182 , RI99249d0_511);
nand \U$5772 ( \6460 , \6072 , RI992b3c0_351);
and \U$5773 ( \6461 , \6077 , RI9922ae0_571);
nor \U$5774 ( \6462 , \6461 , \1821 );
nand \U$5775 ( \6463 , \6458 , \6459 , \6460 , \6462 );
nor \U$5776 ( \6464 , \6457 , \6463 );
nand \U$5777 ( \6465 , \6452 , \6464 );
not \U$5778 ( \6466 , \6465 );
not \U$5779 ( \6467 , \6466 );
and \U$5780 ( \6468 , \6467 , \6176 );
not \U$5781 ( \6469 , \6467 );
and \U$5782 ( \6470 , \6469 , \6034 );
nor \U$5783 ( \6471 , \6468 , \6470 );
and \U$5784 ( \6472 , \6031 , \6471 );
xor \U$5785 ( \6473 , \6472 , \6439 );
not \U$5786 ( \6474 , \6330 );
not \U$5787 ( \6475 , \6272 );
or \U$5788 ( \6476 , \6474 , \6475 );
buf \U$5789 ( \6477 , \6270 );
not \U$5790 ( \6478 , \6477 );
nand \U$5791 ( \6479 , \6478 , \6328 );
nand \U$5792 ( \6480 , \6476 , \6479 );
not \U$5793 ( \6481 , \6480 );
not \U$5794 ( \6482 , \6266 );
or \U$5795 ( \6483 , \6481 , \6482 );
nand \U$5796 ( \6484 , \6340 , \6253 );
nand \U$5797 ( \6485 , \6483 , \6484 );
and \U$5798 ( \6486 , \6473 , \6485 );
and \U$5799 ( \6487 , \6472 , \6439 );
or \U$5800 ( \6488 , \6486 , \6487 );
nand \U$5801 ( \6489 , \6440 , \6488 );
nand \U$5802 ( \6490 , \6438 , \6489 );
xor \U$5803 ( \6491 , \6291 , \6179 );
xor \U$5804 ( \6492 , \6491 , \6407 );
or \U$5805 ( \6493 , \6490 , \6492 );
not \U$5806 ( \6494 , \6493 );
not \U$5807 ( \6495 , \6227 );
buf \U$5808 ( \6496 , \6363 );
buf \U$5809 ( \6497 , \6496 );
not \U$5810 ( \6498 , \6497 );
not \U$5811 ( \6499 , \6498 );
or \U$5812 ( \6500 , \6495 , \6499 );
nand \U$5813 ( \6501 , \6497 , \6225 );
nand \U$5814 ( \6502 , \6500 , \6501 );
not \U$5815 ( \6503 , \6502 );
not \U$5816 ( \6504 , \5956 );
nor \U$5817 ( \6505 , \6504 , \6354 );
not \U$5818 ( \6506 , \6505 );
not \U$5819 ( \6507 , \6366 );
not \U$5820 ( \6508 , \6507 );
or \U$5821 ( \6509 , \6506 , \6508 );
not \U$5822 ( \6510 , \6505 );
not \U$5823 ( \6511 , \6507 );
nand \U$5824 ( \6512 , \6510 , \6511 );
nand \U$5825 ( \6513 , \6509 , \6512 );
not \U$5826 ( \6514 , \6513 );
not \U$5827 ( \6515 , \5982 );
nor \U$5828 ( \6516 , \6515 , \5984 );
not \U$5829 ( \6517 , \6516 );
not \U$5830 ( \6518 , \6517 );
not \U$5831 ( \6519 , \5993 );
nor \U$5832 ( \6520 , \6519 , \5985 );
buf \U$5833 ( \6521 , \5976 );
nand \U$5834 ( \6522 , \5981 , \6521 );
nand \U$5835 ( \6523 , \6520 , \6522 );
not \U$5836 ( \6524 , \6523 );
or \U$5837 ( \6525 , \6518 , \6524 );
nand \U$5838 ( \6526 , \6522 , \6520 , \6516 );
nand \U$5839 ( \6527 , \6525 , \6526 );
not \U$5840 ( \6528 , \6527 );
not \U$5841 ( \6529 , \6528 );
or \U$5842 ( \6530 , \6514 , \6529 );
not \U$5843 ( \6531 , \6513 );
nand \U$5844 ( \6532 , \6527 , \6531 );
nand \U$5845 ( \6533 , \6530 , \6532 );
not \U$5846 ( \6534 , \6533 );
not \U$5847 ( \6535 , \6363 );
not \U$5848 ( \6536 , \6535 );
not \U$5849 ( \6537 , \6513 );
or \U$5850 ( \6538 , \6536 , \6537 );
nand \U$5851 ( \6539 , \6363 , \6531 );
nand \U$5852 ( \6540 , \6538 , \6539 );
nand \U$5853 ( \6541 , \6534 , \6540 );
not \U$5854 ( \6542 , \6541 );
not \U$5855 ( \6543 , \6542 );
or \U$5856 ( \6544 , \6503 , \6543 );
not \U$5857 ( \6545 , \6534 );
buf \U$5858 ( \6546 , \6545 );
not \U$5859 ( \6547 , \6496 );
not \U$5860 ( \6548 , \6547 );
nand \U$5861 ( \6549 , \6546 , \6548 );
nand \U$5862 ( \6550 , \6544 , \6549 );
nand \U$5863 ( \6551 , \6216 , RI992ce00_333);
nand \U$5864 ( \6552 , \6153 , RI9931900_273);
and \U$5865 ( \6553 , \6551 , \6552 );
nand \U$5866 ( \6554 , \6184 , RI99258d0_493);
and \U$5867 ( \6555 , \6072 , RI992b2d0_353);
not \U$5868 ( \6556 , RI99229f0_573);
not \U$5869 ( \6557 , \6077 );
or \U$5870 ( \6558 , \6556 , \6557 );
nand \U$5871 ( \6559 , \6558 , \2103 );
nor \U$5872 ( \6560 , \6555 , \6559 );
nand \U$5873 ( \6561 , \6182 , RI99248e0_513);
nand \U$5874 ( \6562 , \6553 , \6554 , \6560 , \6561 );
not \U$5875 ( \6563 , \6113 );
not \U$5876 ( \6564 , \2133 );
and \U$5877 ( \6565 , \6563 , \6564 );
nor \U$5878 ( \6566 , \6120 , \2136 );
nor \U$5879 ( \6567 , \6565 , \6566 );
not \U$5880 ( \6568 , RI9929200_393);
nor \U$5881 ( \6569 , \6568 , \6158 );
buf \U$5882 ( \6570 , \6164 );
not \U$5883 ( \6571 , RI9926b90_453);
nor \U$5884 ( \6572 , \6570 , \6571 );
nor \U$5885 ( \6573 , \6569 , \6572 );
nand \U$5886 ( \6574 , \6567 , \6573 );
nor \U$5887 ( \6575 , \6562 , \6574 );
not \U$5888 ( \6576 , \6105 );
not \U$5889 ( \6577 , \2121 );
and \U$5890 ( \6578 , \6576 , \6577 );
nor \U$5891 ( \6579 , \6110 , \2115 );
nor \U$5892 ( \6580 , \6578 , \6579 );
not \U$5893 ( \6581 , \6137 );
not \U$5894 ( \6582 , \6581 );
not \U$5895 ( \6583 , \6582 );
not \U$5896 ( \6584 , \2108 );
and \U$5897 ( \6585 , \6583 , \6584 );
nor \U$5898 ( \6586 , \6145 , \2129 );
nor \U$5899 ( \6587 , \6585 , \6586 );
nand \U$5900 ( \6588 , \6580 , \6587 );
not \U$5901 ( \6589 , RI99288a0_413);
not \U$5902 ( \6590 , \6206 );
or \U$5903 ( \6591 , \6589 , \6590 );
nand \U$5904 ( \6592 , \6204 , RI9927f40_433);
nand \U$5905 ( \6593 , \6591 , \6592 );
nor \U$5906 ( \6594 , \6588 , \6593 );
nand \U$5907 ( \6595 , \6575 , \6594 );
buf \U$5908 ( \6596 , \6595 );
not \U$5909 ( \6597 , \6034 );
and \U$5910 ( \6598 , \6596 , \6597 );
not \U$5911 ( \6599 , \6596 );
and \U$5912 ( \6600 , \6599 , \6034 );
nor \U$5913 ( \6601 , \6598 , \6600 );
and \U$5914 ( \6602 , \6031 , \6601 );
xor \U$5915 ( \6603 , \6550 , \6602 );
nand \U$5916 ( \6604 , \6184 , RI9925948_492);
nand \U$5917 ( \6605 , \6182 , RI9924958_512);
nand \U$5918 ( \6606 , \6072 , RI992b348_352);
and \U$5919 ( \6607 , \6077 , RI9922a68_572);
nor \U$5920 ( \6608 , \6607 , \1910 );
nand \U$5921 ( \6609 , \6604 , \6605 , \6606 , \6608 );
nand \U$5922 ( \6610 , \6191 , RI9923ff8_532);
nand \U$5923 ( \6611 , \6195 , RI992a9e8_372);
nand \U$5924 ( \6612 , \6197 , RI992ed68_312);
nand \U$5925 ( \6613 , \6199 , RI992f6c8_292);
nand \U$5926 ( \6614 , \6610 , \6611 , \6612 , \6613 );
nor \U$5927 ( \6615 , \6609 , \6614 );
nand \U$5928 ( \6616 , \6125 , RI9927fb8_432);
nand \U$5929 ( \6617 , \6442 , RI9928918_412);
nand \U$5930 ( \6618 , \6210 , RI9923698_552);
nand \U$5931 ( \6619 , \6144 , RI99262a8_472);
nand \U$5932 ( \6620 , \6616 , \6617 , \6618 , \6619 );
nand \U$5933 ( \6621 , \6216 , RI992ce78_332);
nand \U$5934 ( \6622 , \6153 , RI9931978_272);
nand \U$5935 ( \6623 , \6220 , RI9929278_392);
nand \U$5936 ( \6624 , \6213 , RI9926c08_452);
nand \U$5937 ( \6625 , \6621 , \6622 , \6623 , \6624 );
nor \U$5938 ( \6626 , \6620 , \6625 );
nand \U$5939 ( \6627 , \6615 , \6626 );
buf \U$5940 ( \6628 , \6627 );
not \U$5941 ( \6629 , \6628 );
not \U$5942 ( \6630 , \6272 );
or \U$5943 ( \6631 , \6629 , \6630 );
not \U$5944 ( \6632 , \6628 );
nand \U$5945 ( \6633 , \6478 , \6632 );
nand \U$5946 ( \6634 , \6631 , \6633 );
not \U$5947 ( \6635 , \6634 );
not \U$5948 ( \6636 , \6266 );
or \U$5949 ( \6637 , \6635 , \6636 );
not \U$5950 ( \6638 , \6467 );
not \U$5951 ( \6639 , \6272 );
or \U$5952 ( \6640 , \6638 , \6639 );
nand \U$5953 ( \6641 , \6478 , \6466 );
nand \U$5954 ( \6642 , \6640 , \6641 );
nand \U$5955 ( \6643 , \6642 , \6253 );
nand \U$5956 ( \6644 , \6637 , \6643 );
and \U$5957 ( \6645 , \6603 , \6644 );
and \U$5958 ( \6646 , \6550 , \6602 );
or \U$5959 ( \6647 , \6645 , \6646 );
not \U$5960 ( \6648 , \6330 );
not \U$5961 ( \6649 , \6403 );
or \U$5962 ( \6650 , \6648 , \6649 );
buf \U$5963 ( \6651 , \6391 );
not \U$5964 ( \6652 , \6651 );
nand \U$5965 ( \6653 , \6652 , \6328 );
nand \U$5966 ( \6654 , \6650 , \6653 );
not \U$5967 ( \6655 , \6654 );
not \U$5968 ( \6656 , \6422 );
or \U$5969 ( \6657 , \6655 , \6656 );
and \U$5970 ( \6658 , \6173 , \6403 );
not \U$5971 ( \6659 , \6173 );
and \U$5972 ( \6660 , \6659 , \6652 );
nor \U$5973 ( \6661 , \6658 , \6660 );
not \U$5974 ( \6662 , \6661 );
nand \U$5975 ( \6663 , \6662 , \6384 );
nand \U$5976 ( \6664 , \6657 , \6663 );
not \U$5977 ( \6665 , \6664 );
not \U$5978 ( \6666 , \5992 );
not \U$5979 ( \6667 , \6666 );
buf \U$5980 ( \6668 , \5977 );
nand \U$5981 ( \6669 , \5976 , \6668 );
not \U$5982 ( \6670 , \6669 );
or \U$5983 ( \6671 , \6667 , \6670 );
buf \U$5984 ( \6672 , \5980 );
nand \U$5985 ( \6673 , \6671 , \6672 );
not \U$5986 ( \6674 , \5985 );
nand \U$5987 ( \6675 , \5978 , \965 );
nand \U$5988 ( \6676 , \6674 , \6675 );
and \U$5989 ( \6677 , \6673 , \6676 );
not \U$5990 ( \6678 , \6673 );
not \U$5991 ( \6679 , \6676 );
and \U$5992 ( \6680 , \6678 , \6679 );
nor \U$5993 ( \6681 , \6677 , \6680 );
buf \U$5994 ( \6682 , \5991 );
nand \U$5995 ( \6683 , \6669 , \6682 );
and \U$5996 ( \6684 , \5989 , \6672 );
xor \U$5997 ( \6685 , \6683 , \6684 );
buf \U$5998 ( \6686 , \6685 );
not \U$5999 ( \6687 , \6686 );
and \U$6000 ( \6688 , \6681 , \6687 );
not \U$6001 ( \6689 , \6681 );
and \U$6002 ( \6690 , \6689 , \6686 );
nor \U$6003 ( \6691 , \6688 , \6690 );
buf \U$6004 ( \6692 , \6691 );
not \U$6005 ( \6693 , \6692 );
not \U$6006 ( \6694 , \6527 );
not \U$6007 ( \6695 , \6681 );
nand \U$6008 ( \6696 , \6694 , \6695 );
not \U$6009 ( \6697 , \6528 );
not \U$6010 ( \6698 , \6695 );
nand \U$6011 ( \6699 , \6697 , \6698 );
nand \U$6012 ( \6700 , \6696 , \6699 , \6691 );
not \U$6013 ( \6701 , \6700 );
or \U$6014 ( \6702 , \6693 , \6701 );
buf \U$6015 ( \6703 , \6527 );
nand \U$6016 ( \6704 , \6702 , \6703 );
not \U$6017 ( \6705 , \6173 );
buf \U$6018 ( \6706 , \6535 );
not \U$6019 ( \6707 , \6706 );
or \U$6020 ( \6708 , \6705 , \6707 );
nand \U$6021 ( \6709 , \6548 , \6174 );
nand \U$6022 ( \6710 , \6708 , \6709 );
not \U$6023 ( \6711 , \6710 );
not \U$6024 ( \6712 , \6542 );
or \U$6025 ( \6713 , \6711 , \6712 );
nand \U$6026 ( \6714 , \6546 , \6502 );
nand \U$6027 ( \6715 , \6713 , \6714 );
xor \U$6028 ( \6716 , \6704 , \6715 );
not \U$6029 ( \6717 , \6467 );
not \U$6030 ( \6718 , \6651 );
or \U$6031 ( \6719 , \6717 , \6718 );
nand \U$6032 ( \6720 , \6402 , \6466 );
nand \U$6033 ( \6721 , \6719 , \6720 );
not \U$6034 ( \6722 , \6721 );
not \U$6035 ( \6723 , \6397 );
or \U$6036 ( \6724 , \6722 , \6723 );
nand \U$6037 ( \6725 , \6384 , \6654 );
nand \U$6038 ( \6726 , \6724 , \6725 );
and \U$6039 ( \6727 , \6716 , \6726 );
and \U$6040 ( \6728 , \6704 , \6715 );
or \U$6041 ( \6729 , \6727 , \6728 );
xor \U$6042 ( \6730 , \6665 , \6729 );
not \U$6043 ( \6731 , \6477 );
not \U$6044 ( \6732 , \6596 );
or \U$6045 ( \6733 , \6731 , \6732 );
not \U$6046 ( \6734 , \6596 );
nand \U$6047 ( \6735 , \6271 , \6734 );
nand \U$6048 ( \6736 , \6733 , \6735 );
not \U$6049 ( \6737 , \6736 );
not \U$6050 ( \6738 , \6266 );
or \U$6051 ( \6739 , \6737 , \6738 );
nand \U$6052 ( \6740 , \6634 , \6253 );
nand \U$6053 ( \6741 , \6739 , \6740 );
not \U$6054 ( \6742 , \6741 );
not \U$6055 ( \6743 , \6105 );
not \U$6056 ( \6744 , \2049 );
and \U$6057 ( \6745 , \6743 , \6744 );
nor \U$6058 ( \6746 , \6110 , \2043 );
nor \U$6059 ( \6747 , \6745 , \6746 );
not \U$6060 ( \6748 , \6113 );
not \U$6061 ( \6749 , \2061 );
and \U$6062 ( \6750 , \6748 , \6749 );
nor \U$6063 ( \6751 , \6120 , \2064 );
nor \U$6064 ( \6752 , \6750 , \6751 );
nand \U$6065 ( \6753 , \6747 , \6752 );
and \U$6066 ( \6754 , \6072 , RI992b258_354);
not \U$6067 ( \6755 , RI9922978_574);
not \U$6068 ( \6756 , \6077 );
or \U$6069 ( \6757 , \6755 , \6756 );
nand \U$6070 ( \6758 , \6757 , \2031 );
nor \U$6071 ( \6759 , \6754 , \6758 );
not \U$6072 ( \6760 , \6086 );
not \U$6073 ( \6761 , RI9924868_514);
not \U$6074 ( \6762 , \6761 );
and \U$6075 ( \6763 , \6760 , \6762 );
not \U$6076 ( \6764 , RI9925858_494);
nor \U$6077 ( \6765 , \6764 , \6095 );
nor \U$6078 ( \6766 , \6763 , \6765 );
nand \U$6079 ( \6767 , \6759 , \6766 );
nor \U$6080 ( \6768 , \6753 , \6767 );
and \U$6081 ( \6769 , \6216 , RI992cd88_334);
not \U$6082 ( \6770 , RI9931888_274);
not \U$6083 ( \6771 , \6153 );
nor \U$6084 ( \6772 , \6770 , \6771 );
nor \U$6085 ( \6773 , \6769 , \6772 );
not \U$6086 ( \6774 , \6166 );
not \U$6087 ( \6775 , RI9926b18_454);
not \U$6088 ( \6776 , \6775 );
and \U$6089 ( \6777 , \6774 , \6776 );
not \U$6090 ( \6778 , \6158 );
and \U$6091 ( \6779 , \6778 , RI9929188_394);
nor \U$6092 ( \6780 , \6777 , \6779 );
nand \U$6093 ( \6781 , \6773 , \6780 );
not \U$6094 ( \6782 , \6126 );
not \U$6095 ( \6783 , RI9927ec8_434);
not \U$6096 ( \6784 , \6783 );
and \U$6097 ( \6785 , \6782 , \6784 );
not \U$6098 ( \6786 , \6313 );
not \U$6099 ( \6787 , RI9928828_414);
nor \U$6100 ( \6788 , \6786 , \6787 );
nor \U$6101 ( \6789 , \6785 , \6788 );
and \U$6102 ( \6790 , RI99261b8_474, \6144 );
nor \U$6103 ( \6791 , \6138 , \2036 );
nor \U$6104 ( \6792 , \6790 , \6791 );
nand \U$6105 ( \6793 , \6789 , \6792 );
nor \U$6106 ( \6794 , \6781 , \6793 );
nand \U$6107 ( \6795 , \6768 , \6794 );
not \U$6108 ( \6796 , \6033 );
and \U$6109 ( \6797 , \6795 , \6796 );
not \U$6110 ( \6798 , \6795 );
and \U$6111 ( \6799 , \6798 , \6033 );
nor \U$6112 ( \6800 , \6797 , \6799 );
nand \U$6113 ( \6801 , \6030 , \6800 );
not \U$6114 ( \6802 , \6692 );
not \U$6115 ( \6803 , \6703 );
not \U$6116 ( \6804 , \6803 );
and \U$6117 ( \6805 , \6802 , \6804 );
not \U$6118 ( \6806 , \6227 );
not \U$6119 ( \6807 , \6703 );
not \U$6120 ( \6808 , \6807 );
or \U$6121 ( \6809 , \6806 , \6808 );
nand \U$6122 ( \6810 , \6703 , \6225 );
nand \U$6123 ( \6811 , \6809 , \6810 );
not \U$6124 ( \6812 , \6811 );
nor \U$6125 ( \6813 , \6812 , \6700 );
nor \U$6126 ( \6814 , \6805 , \6813 );
nand \U$6127 ( \6815 , \6801 , \6814 );
not \U$6128 ( \6816 , \6815 );
or \U$6129 ( \6817 , \6742 , \6816 );
not \U$6130 ( \6818 , \6801 );
not \U$6131 ( \6819 , \6814 );
nand \U$6132 ( \6820 , \6818 , \6819 );
nand \U$6133 ( \6821 , \6817 , \6820 );
and \U$6134 ( \6822 , \6730 , \6821 );
and \U$6135 ( \6823 , \6665 , \6729 );
or \U$6136 ( \6824 , \6822 , \6823 );
xor \U$6137 ( \6825 , \6647 , \6824 );
and \U$6138 ( \6826 , \6034 , \6632 );
and \U$6139 ( \6827 , \6176 , \6628 );
nor \U$6140 ( \6828 , \6826 , \6827 );
nand \U$6141 ( \6829 , \6031 , \6828 );
not \U$6142 ( \6830 , \6829 );
not \U$6143 ( \6831 , \6664 );
or \U$6144 ( \6832 , \6830 , \6831 );
not \U$6145 ( \6833 , \6829 );
nand \U$6146 ( \6834 , \6833 , \6665 );
nand \U$6147 ( \6835 , \6832 , \6834 );
not \U$6148 ( \6836 , \6835 );
not \U$6149 ( \6837 , \6399 );
not \U$6150 ( \6838 , \6661 );
and \U$6151 ( \6839 , \6837 , \6838 );
nor \U$6152 ( \6840 , \6385 , \6419 );
nor \U$6153 ( \6841 , \6839 , \6840 );
not \U$6154 ( \6842 , \6546 );
not \U$6155 ( \6843 , \6842 );
not \U$6156 ( \6844 , \6541 );
or \U$6157 ( \6845 , \6843 , \6844 );
nand \U$6158 ( \6846 , \6845 , \6548 );
not \U$6159 ( \6847 , \6846 );
and \U$6160 ( \6848 , \6841 , \6847 );
not \U$6161 ( \6849 , \6841 );
and \U$6162 ( \6850 , \6849 , \6846 );
nor \U$6163 ( \6851 , \6848 , \6850 );
not \U$6164 ( \6852 , \6642 );
not \U$6165 ( \6853 , \6266 );
or \U$6166 ( \6854 , \6852 , \6853 );
nand \U$6167 ( \6855 , \6480 , \6253 );
nand \U$6168 ( \6856 , \6854 , \6855 );
not \U$6169 ( \6857 , \6856 );
and \U$6170 ( \6858 , \6851 , \6857 );
not \U$6171 ( \6859 , \6851 );
and \U$6172 ( \6860 , \6859 , \6856 );
nor \U$6173 ( \6861 , \6858 , \6860 );
not \U$6174 ( \6862 , \6861 );
or \U$6175 ( \6863 , \6836 , \6862 );
or \U$6176 ( \6864 , \6835 , \6861 );
nand \U$6177 ( \6865 , \6863 , \6864 );
xor \U$6178 ( \6866 , \6825 , \6865 );
xor \U$6179 ( \6867 , \6550 , \6602 );
xor \U$6180 ( \6868 , \6867 , \6644 );
not \U$6181 ( \6869 , \6868 );
xor \U$6182 ( \6870 , \6665 , \6729 );
xor \U$6183 ( \6871 , \6870 , \6821 );
not \U$6184 ( \6872 , \6871 );
or \U$6185 ( \6873 , \6869 , \6872 );
or \U$6186 ( \6874 , \6871 , \6868 );
xor \U$6187 ( \6875 , \6704 , \6715 );
xor \U$6188 ( \6876 , \6875 , \6726 );
not \U$6189 ( \6877 , \6876 );
not \U$6190 ( \6878 , \6877 );
xor \U$6191 ( \6879 , \6814 , \6818 );
xor \U$6192 ( \6880 , \6879 , \6741 );
not \U$6193 ( \6881 , \6880 );
or \U$6194 ( \6882 , \6878 , \6881 );
not \U$6195 ( \6883 , \6330 );
not \U$6196 ( \6884 , \6547 );
or \U$6197 ( \6885 , \6883 , \6884 );
nand \U$6198 ( \6886 , \6548 , \6328 );
nand \U$6199 ( \6887 , \6885 , \6886 );
not \U$6200 ( \6888 , \6887 );
not \U$6201 ( \6889 , \6542 );
or \U$6202 ( \6890 , \6888 , \6889 );
nand \U$6203 ( \6891 , \6710 , \6546 );
nand \U$6204 ( \6892 , \6890 , \6891 );
not \U$6205 ( \6893 , \6628 );
not \U$6206 ( \6894 , \6391 );
or \U$6207 ( \6895 , \6893 , \6894 );
not \U$6208 ( \6896 , \6651 );
nand \U$6209 ( \6897 , \6896 , \6632 );
nand \U$6210 ( \6898 , \6895 , \6897 );
not \U$6211 ( \6899 , \6898 );
not \U$6212 ( \6900 , \6396 );
not \U$6213 ( \6901 , \6900 );
or \U$6214 ( \6902 , \6899 , \6901 );
not \U$6215 ( \6903 , \6383 );
not \U$6216 ( \6904 , \6903 );
nand \U$6217 ( \6905 , \6904 , \6721 );
nand \U$6218 ( \6906 , \6902 , \6905 );
xor \U$6219 ( \6907 , \6892 , \6906 );
not \U$6220 ( \6908 , \6795 );
not \U$6221 ( \6909 , \6477 );
or \U$6222 ( \6910 , \6908 , \6909 );
buf \U$6223 ( \6911 , \6023 );
not \U$6224 ( \6912 , \6795 );
nand \U$6225 ( \6913 , \6911 , \6912 );
nand \U$6226 ( \6914 , \6910 , \6913 );
not \U$6227 ( \6915 , \6914 );
not \U$6228 ( \6916 , \6265 );
or \U$6229 ( \6917 , \6915 , \6916 );
buf \U$6230 ( \6918 , \6263 );
not \U$6231 ( \6919 , \6918 );
nand \U$6232 ( \6920 , \6736 , \6919 );
nand \U$6233 ( \6921 , \6917 , \6920 );
and \U$6234 ( \6922 , \6907 , \6921 );
and \U$6235 ( \6923 , \6892 , \6906 );
or \U$6236 ( \6924 , \6922 , \6923 );
nand \U$6237 ( \6925 , \6882 , \6924 );
or \U$6238 ( \6926 , \6880 , \6877 );
nand \U$6239 ( \6927 , \6925 , \6926 );
nand \U$6240 ( \6928 , \6874 , \6927 );
nand \U$6241 ( \6929 , \6873 , \6928 );
nor \U$6242 ( \6930 , \6866 , \6929 );
not \U$6243 ( \6931 , \6930 );
not \U$6244 ( \6932 , \6176 );
nand \U$6245 ( \6933 , \6216 , RI992cd10_335);
nand \U$6246 ( \6934 , \6153 , RI9931810_275);
nand \U$6247 ( \6935 , \6220 , RI9929110_395);
nand \U$6248 ( \6936 , \6213 , RI9926aa0_455);
nand \U$6249 ( \6937 , \6933 , \6934 , \6935 , \6936 );
nand \U$6250 ( \6938 , \6125 , RI9927e50_435);
nand \U$6251 ( \6939 , \6318 , RI9926140_475);
nand \U$6252 ( \6940 , \6210 , RI9923530_555);
not \U$6253 ( \6941 , \6132 );
nand \U$6254 ( \6942 , \6941 , RI99287b0_415);
nand \U$6255 ( \6943 , \6938 , \6939 , \6940 , \6942 );
nor \U$6256 ( \6944 , \6937 , \6943 );
nand \U$6257 ( \6945 , \6072 , RI992b1e0_355);
nand \U$6258 ( \6946 , \6182 , RI99247f0_515);
nand \U$6259 ( \6947 , \6297 , RI99257e0_495);
and \U$6260 ( \6948 , \6077 , RI9922900_575);
nor \U$6261 ( \6949 , \6948 , \2268 );
nand \U$6262 ( \6950 , \6945 , \6946 , \6947 , \6949 );
or \U$6263 ( \6951 , \6112 , \2255 );
or \U$6264 ( \6952 , \6119 , \2253 );
not \U$6265 ( \6953 , RI992d670_315);
nor \U$6266 ( \6954 , \6104 , \6953 );
nor \U$6267 ( \6955 , \6109 , \2244 );
nor \U$6268 ( \6956 , \6954 , \6955 );
nand \U$6269 ( \6957 , \6951 , \6952 , \6956 );
nor \U$6270 ( \6958 , \6950 , \6957 );
nand \U$6271 ( \6959 , \6944 , \6958 );
buf \U$6272 ( \6960 , \6959 );
not \U$6273 ( \6961 , \6960 );
and \U$6274 ( \6962 , \6932 , \6961 );
and \U$6275 ( \6963 , \6597 , \6960 );
nor \U$6276 ( \6964 , \6962 , \6963 );
nand \U$6277 ( \6965 , \6031 , \6964 );
not \U$6278 ( \6966 , \6965 );
not \U$6279 ( \6967 , \6819 );
and \U$6280 ( \6968 , \6966 , \6967 );
not \U$6281 ( \6969 , \6172 );
not \U$6282 ( \6970 , \6703 );
not \U$6283 ( \6971 , \6970 );
or \U$6284 ( \6972 , \6969 , \6971 );
not \U$6285 ( \6973 , \6528 );
not \U$6286 ( \6974 , \6172 );
nand \U$6287 ( \6975 , \6973 , \6974 );
nand \U$6288 ( \6976 , \6972 , \6975 );
not \U$6289 ( \6977 , \6976 );
and \U$6290 ( \6978 , \6699 , \6696 , \6691 );
not \U$6291 ( \6979 , \6978 );
or \U$6292 ( \6980 , \6977 , \6979 );
not \U$6293 ( \6981 , \6692 );
nand \U$6294 ( \6982 , \6811 , \6981 );
nand \U$6295 ( \6983 , \6980 , \6982 );
not \U$6296 ( \6984 , \6983 );
nand \U$6297 ( \6985 , \5975 , \5970 );
not \U$6298 ( \6986 , \6985 );
buf \U$6299 ( \6987 , \5967 );
not \U$6300 ( \6988 , \6987 );
not \U$6301 ( \6989 , \5968 );
or \U$6302 ( \6990 , \6988 , \6989 );
nand \U$6303 ( \6991 , \5658 , \1114 );
nand \U$6304 ( \6992 , \6990 , \6991 );
not \U$6305 ( \6993 , \6992 );
or \U$6306 ( \6994 , \6986 , \6993 );
or \U$6307 ( \6995 , \6992 , \6985 );
nand \U$6308 ( \6996 , \6994 , \6995 );
not \U$6309 ( \6997 , \6996 );
not \U$6310 ( \6998 , \6997 );
not \U$6311 ( \6999 , \6998 );
nand \U$6312 ( \7000 , \6682 , \6668 );
not \U$6313 ( \7001 , \7000 );
and \U$6314 ( \7002 , \6521 , \7001 );
not \U$6315 ( \7003 , \6521 );
and \U$6316 ( \7004 , \7003 , \7000 );
nor \U$6317 ( \7005 , \7002 , \7004 );
not \U$6318 ( \7006 , \7005 );
not \U$6319 ( \7007 , \7006 );
or \U$6320 ( \7008 , \6999 , \7007 );
nand \U$6321 ( \7009 , \7005 , \6997 );
nand \U$6322 ( \7010 , \7008 , \7009 );
buf \U$6323 ( \7011 , \7010 );
buf \U$6324 ( \7012 , \7011 );
not \U$6325 ( \7013 , \7010 );
nand \U$6326 ( \7014 , \6686 , \7005 );
not \U$6327 ( \7015 , \7005 );
nand \U$6328 ( \7016 , \7015 , \6687 );
and \U$6329 ( \7017 , \7013 , \7014 , \7016 );
buf \U$6330 ( \7018 , \7017 );
or \U$6331 ( \7019 , \7012 , \7018 );
buf \U$6332 ( \7020 , \6686 );
not \U$6333 ( \7021 , \7020 );
not \U$6334 ( \7022 , \7021 );
nand \U$6335 ( \7023 , \7019 , \7022 );
not \U$6336 ( \7024 , \7023 );
nand \U$6337 ( \7025 , \6984 , \7024 );
not \U$6338 ( \7026 , \7025 );
not \U$6339 ( \7027 , \6403 );
not \U$6340 ( \7028 , \6596 );
or \U$6341 ( \7029 , \7027 , \7028 );
nand \U$6342 ( \7030 , \6402 , \6734 );
nand \U$6343 ( \7031 , \7029 , \7030 );
not \U$6344 ( \7032 , \7031 );
not \U$6345 ( \7033 , \6395 );
buf \U$6346 ( \7034 , \7033 );
not \U$6347 ( \7035 , \7034 );
or \U$6348 ( \7036 , \7032 , \7035 );
nand \U$6349 ( \7037 , \6383 , \6898 );
nand \U$6350 ( \7038 , \7036 , \7037 );
not \U$6351 ( \7039 , \7038 );
or \U$6352 ( \7040 , \7026 , \7039 );
nand \U$6353 ( \7041 , \6983 , \7023 );
nand \U$6354 ( \7042 , \7040 , \7041 );
nand \U$6355 ( \7043 , \6965 , \6819 );
and \U$6356 ( \7044 , \7042 , \7043 );
nor \U$6357 ( \7045 , \6968 , \7044 );
xor \U$6358 ( \7046 , \6876 , \6924 );
xor \U$6359 ( \7047 , \7046 , \6880 );
xor \U$6360 ( \7048 , \7045 , \7047 );
not \U$6361 ( \7049 , \6265 );
not \U$6362 ( \7050 , \6477 );
not \U$6363 ( \7051 , \6960 );
or \U$6364 ( \7052 , \7050 , \7051 );
not \U$6365 ( \7053 , \6911 );
not \U$6366 ( \7054 , \7053 );
not \U$6367 ( \7055 , \6960 );
nand \U$6368 ( \7056 , \7054 , \7055 );
nand \U$6369 ( \7057 , \7052 , \7056 );
not \U$6370 ( \7058 , \7057 );
or \U$6371 ( \7059 , \7049 , \7058 );
nand \U$6372 ( \7060 , \6914 , \6919 );
nand \U$6373 ( \7061 , \7059 , \7060 );
not \U$6374 ( \7062 , \7061 );
and \U$6375 ( \7063 , \6983 , \7024 );
not \U$6376 ( \7064 , \6983 );
and \U$6377 ( \7065 , \7064 , \7023 );
or \U$6378 ( \7066 , \7063 , \7065 );
xor \U$6379 ( \7067 , \7066 , \7038 );
not \U$6380 ( \7068 , \7067 );
or \U$6381 ( \7069 , \7062 , \7068 );
or \U$6382 ( \7070 , \7067 , \7061 );
not \U$6383 ( \7071 , \6330 );
not \U$6384 ( \7072 , \6528 );
or \U$6385 ( \7073 , \7071 , \7072 );
nand \U$6386 ( \7074 , \6703 , \6328 );
nand \U$6387 ( \7075 , \7073 , \7074 );
not \U$6388 ( \7076 , \7075 );
not \U$6389 ( \7077 , \6978 );
or \U$6390 ( \7078 , \7076 , \7077 );
nand \U$6391 ( \7079 , \6976 , \6981 );
nand \U$6392 ( \7080 , \7078 , \7079 );
not \U$6393 ( \7081 , \6628 );
not \U$6394 ( \7082 , \6706 );
or \U$6395 ( \7083 , \7081 , \7082 );
buf \U$6396 ( \7084 , \6363 );
nand \U$6397 ( \7085 , \7084 , \6632 );
nand \U$6398 ( \7086 , \7083 , \7085 );
not \U$6399 ( \7087 , \7086 );
nand \U$6400 ( \7088 , \6540 , \6534 );
not \U$6401 ( \7089 , \7088 );
not \U$6402 ( \7090 , \7089 );
or \U$6403 ( \7091 , \7087 , \7090 );
not \U$6404 ( \7092 , \6467 );
not \U$6405 ( \7093 , \7084 );
not \U$6406 ( \7094 , \7093 );
or \U$6407 ( \7095 , \7092 , \7094 );
nand \U$6408 ( \7096 , \6496 , \6466 );
nand \U$6409 ( \7097 , \7095 , \7096 );
nand \U$6410 ( \7098 , \7097 , \6545 );
nand \U$6411 ( \7099 , \7091 , \7098 );
xor \U$6412 ( \7100 , \7080 , \7099 );
not \U$6413 ( \7101 , \6795 );
not \U$6414 ( \7102 , \6403 );
or \U$6415 ( \7103 , \7101 , \7102 );
nand \U$6416 ( \7104 , \6402 , \6912 );
nand \U$6417 ( \7105 , \7103 , \7104 );
not \U$6418 ( \7106 , \7105 );
not \U$6419 ( \7107 , \6397 );
or \U$6420 ( \7108 , \7106 , \7107 );
nand \U$6421 ( \7109 , \7031 , \6383 );
nand \U$6422 ( \7110 , \7108 , \7109 );
and \U$6423 ( \7111 , \7100 , \7110 );
and \U$6424 ( \7112 , \7080 , \7099 );
or \U$6425 ( \7113 , \7111 , \7112 );
nand \U$6426 ( \7114 , \7070 , \7113 );
nand \U$6427 ( \7115 , \7069 , \7114 );
xor \U$6428 ( \7116 , \6892 , \6906 );
xor \U$6429 ( \7117 , \7116 , \6921 );
not \U$6430 ( \7118 , \7117 );
not \U$6431 ( \7119 , RI9924778_516);
nor \U$6432 ( \7120 , \7119 , \6086 );
not \U$6433 ( \7121 , RI9925768_496);
nor \U$6434 ( \7122 , \7121 , \6095 );
nor \U$6435 ( \7123 , \7120 , \7122 );
and \U$6436 ( \7124 , \6072 , RI992b168_356);
not \U$6437 ( \7125 , \2197 );
nand \U$6438 ( \7126 , \6077 , RI9922888_576);
nand \U$6439 ( \7127 , \7125 , \7126 );
nor \U$6440 ( \7128 , \7124 , \7127 );
nand \U$6441 ( \7129 , \7123 , \7128 );
nand \U$6442 ( \7130 , \6191 , RI9923e18_536);
nand \U$6443 ( \7131 , \6195 , RI992a808_376);
nand \U$6444 ( \7132 , \6197 , RI992d5f8_316);
nand \U$6445 ( \7133 , \6199 , RI992f4e8_296);
nand \U$6446 ( \7134 , \7130 , \7131 , \7132 , \7133 );
nor \U$6447 ( \7135 , \7129 , \7134 );
nand \U$6448 ( \7136 , \6204 , RI9927dd8_436);
nand \U$6449 ( \7137 , \6206 , RI9928738_416);
nand \U$6450 ( \7138 , \6210 , RI99234b8_556);
nand \U$6451 ( \7139 , RI99260c8_476, \6144 );
nand \U$6452 ( \7140 , \7136 , \7137 , \7138 , \7139 );
nand \U$6453 ( \7141 , \6216 , RI992cc98_336);
nand \U$6454 ( \7142 , \6153 , RI9931798_276);
nand \U$6455 ( \7143 , \6778 , RI9929098_396);
nand \U$6456 ( \7144 , \6213 , RI9926a28_456);
nand \U$6457 ( \7145 , \7141 , \7142 , \7143 , \7144 );
nor \U$6458 ( \7146 , \7140 , \7145 );
nand \U$6459 ( \7147 , \7135 , \7146 );
not \U$6460 ( \7148 , \7147 );
buf \U$6461 ( \7149 , \7148 );
not \U$6462 ( \7150 , \7149 );
and \U$6463 ( \7151 , \7150 , \6597 );
not \U$6464 ( \7152 , \7150 );
buf \U$6465 ( \7153 , \6032 );
not \U$6466 ( \7154 , \7153 );
and \U$6467 ( \7155 , \7152 , \7154 );
nor \U$6468 ( \7156 , \7151 , \7155 );
nand \U$6469 ( \7157 , \6030 , \7156 );
not \U$6470 ( \7158 , \7157 );
not \U$6471 ( \7159 , \7097 );
not \U$6472 ( \7160 , \6542 );
or \U$6473 ( \7161 , \7159 , \7160 );
buf \U$6474 ( \7162 , \6534 );
not \U$6475 ( \7163 , \7162 );
nand \U$6476 ( \7164 , \6887 , \7163 );
nand \U$6477 ( \7165 , \7161 , \7164 );
not \U$6478 ( \7166 , \7165 );
not \U$6479 ( \7167 , \7166 );
or \U$6480 ( \7168 , \7158 , \7167 );
not \U$6481 ( \7169 , \6227 );
not \U$6482 ( \7170 , \7020 );
not \U$6483 ( \7171 , \7170 );
or \U$6484 ( \7172 , \7169 , \7171 );
nand \U$6485 ( \7173 , \7020 , \6225 );
nand \U$6486 ( \7174 , \7172 , \7173 );
not \U$6487 ( \7175 , \7174 );
buf \U$6488 ( \7176 , \7018 );
not \U$6489 ( \7177 , \7176 );
or \U$6490 ( \7178 , \7175 , \7177 );
nand \U$6491 ( \7179 , \7012 , \7022 );
nand \U$6492 ( \7180 , \7178 , \7179 );
nand \U$6493 ( \7181 , \7168 , \7180 );
not \U$6494 ( \7182 , \7157 );
nand \U$6495 ( \7183 , \7182 , \7165 );
and \U$6496 ( \7184 , \7181 , \7183 );
nand \U$6497 ( \7185 , \7118 , \7184 );
and \U$6498 ( \7186 , \7115 , \7185 );
nor \U$6499 ( \7187 , \7118 , \7184 );
nor \U$6500 ( \7188 , \7186 , \7187 );
and \U$6501 ( \7189 , \7048 , \7188 );
and \U$6502 ( \7190 , \7045 , \7047 );
or \U$6503 ( \7191 , \7189 , \7190 );
xor \U$6504 ( \7192 , \6868 , \6871 );
xnor \U$6505 ( \7193 , \7192 , \6927 );
nand \U$6506 ( \7194 , \7191 , \7193 );
nand \U$6507 ( \7195 , \6931 , \7194 );
xor \U$6508 ( \7196 , \6647 , \6824 );
and \U$6509 ( \7197 , \7196 , \6865 );
and \U$6510 ( \7198 , \6647 , \6824 );
or \U$6511 ( \7199 , \7197 , \7198 );
not \U$6512 ( \7200 , \6846 );
not \U$6513 ( \7201 , \6856 );
or \U$6514 ( \7202 , \7200 , \7201 );
or \U$6515 ( \7203 , \6856 , \6846 );
not \U$6516 ( \7204 , \6841 );
nand \U$6517 ( \7205 , \7203 , \7204 );
nand \U$6518 ( \7206 , \7202 , \7205 );
not \U$6519 ( \7207 , \7206 );
xor \U$6520 ( \7208 , \6472 , \6439 );
xor \U$6521 ( \7209 , \7208 , \6485 );
not \U$6522 ( \7210 , \7209 );
not \U$6523 ( \7211 , \7210 );
or \U$6524 ( \7212 , \7207 , \7211 );
not \U$6525 ( \7213 , \7206 );
nand \U$6526 ( \7214 , \7209 , \7213 );
nand \U$6527 ( \7215 , \7212 , \7214 );
nand \U$6528 ( \7216 , \6665 , \6829 );
not \U$6529 ( \7217 , \7216 );
not \U$6530 ( \7218 , \6861 );
not \U$6531 ( \7219 , \7218 );
or \U$6532 ( \7220 , \7217 , \7219 );
not \U$6533 ( \7221 , \6829 );
nand \U$6534 ( \7222 , \7221 , \6664 );
nand \U$6535 ( \7223 , \7220 , \7222 );
xor \U$6536 ( \7224 , \7215 , \7223 );
nor \U$6537 ( \7225 , \7199 , \7224 );
nor \U$6538 ( \7226 , \7195 , \7225 );
nand \U$6539 ( \7227 , \7210 , \7213 );
nand \U$6540 ( \7228 , \7223 , \7227 );
nand \U$6541 ( \7229 , \7209 , \7206 );
and \U$6542 ( \7230 , \7228 , \7229 );
not \U$6543 ( \7231 , \6439 );
not \U$6544 ( \7232 , \6436 );
or \U$6545 ( \7233 , \7231 , \7232 );
nand \U$6546 ( \7234 , \6435 , \6426 );
nand \U$6547 ( \7235 , \7233 , \7234 );
xnor \U$6548 ( \7236 , \7235 , \6488 );
nand \U$6549 ( \7237 , \7230 , \7236 );
and \U$6550 ( \7238 , \7226 , \7237 );
not \U$6551 ( \7239 , \7238 );
xor \U$6552 ( \7240 , \7042 , \6965 );
xor \U$6553 ( \7241 , \7240 , \6814 );
and \U$6554 ( \7242 , \7184 , \7117 );
not \U$6555 ( \7243 , \7184 );
and \U$6556 ( \7244 , \7243 , \7118 );
nor \U$6557 ( \7245 , \7242 , \7244 );
not \U$6558 ( \7246 , \7245 );
not \U$6559 ( \7247 , \7115 );
and \U$6560 ( \7248 , \7246 , \7247 );
and \U$6561 ( \7249 , \7115 , \7245 );
nor \U$6562 ( \7250 , \7248 , \7249 );
xor \U$6563 ( \7251 , \7241 , \7250 );
xor \U$6564 ( \7252 , \7061 , \7113 );
xnor \U$6565 ( \7253 , \7252 , \7067 );
not \U$6566 ( \7254 , \7253 );
buf \U$6567 ( \7255 , \7254 );
nor \U$6568 ( \7256 , \6150 , \2356 );
not \U$6569 ( \7257 , RI9931720_277);
nor \U$6570 ( \7258 , \7257 , \6154 );
nor \U$6571 ( \7259 , \7256 , \7258 );
nor \U$6572 ( \7260 , \6158 , \2371 );
nor \U$6573 ( \7261 , \6570 , \2346 );
nor \U$6574 ( \7262 , \7260 , \7261 );
nand \U$6575 ( \7263 , \7259 , \7262 );
not \U$6576 ( \7264 , \6126 );
not \U$6577 ( \7265 , \2376 );
and \U$6578 ( \7266 , \7264 , \7265 );
not \U$6579 ( \7267 , \6206 );
not \U$6580 ( \7268 , RI99286c0_417);
nor \U$6581 ( \7269 , \7267 , \7268 );
nor \U$6582 ( \7270 , \7266 , \7269 );
nor \U$6583 ( \7271 , \6138 , \2391 );
nor \U$6584 ( \7272 , \6317 , \2349 );
nor \U$6585 ( \7273 , \7271 , \7272 );
nand \U$6586 ( \7274 , \7270 , \7273 );
nor \U$6587 ( \7275 , \7263 , \7274 );
and \U$6588 ( \7276 , \6072 , RI992b0f0_357);
not \U$6589 ( \7277 , RI9922810_577);
not \U$6590 ( \7278 , \6077 );
or \U$6591 ( \7279 , \7277 , \7278 );
not \U$6592 ( \7280 , \2370 );
nand \U$6593 ( \7281 , \7279 , \7280 );
nor \U$6594 ( \7282 , \7276 , \7281 );
not \U$6595 ( \7283 , RI9924700_517);
nor \U$6596 ( \7284 , \6086 , \7283 );
not \U$6597 ( \7285 , RI99256f0_497);
nor \U$6598 ( \7286 , \6298 , \7285 );
nor \U$6599 ( \7287 , \7284 , \7286 );
nand \U$6600 ( \7288 , \7282 , \7287 );
not \U$6601 ( \7289 , \6105 );
not \U$6602 ( \7290 , \2382 );
and \U$6603 ( \7291 , \7289 , \7290 );
not \U$6604 ( \7292 , RI992f470_297);
nor \U$6605 ( \7293 , \7292 , \6110 );
nor \U$6606 ( \7294 , \7291 , \7293 );
not \U$6607 ( \7295 , \6113 );
not \U$6608 ( \7296 , \2362 );
and \U$6609 ( \7297 , \7295 , \7296 );
nor \U$6610 ( \7298 , \6120 , \2365 );
nor \U$6611 ( \7299 , \7297 , \7298 );
nand \U$6612 ( \7300 , \7294 , \7299 );
nor \U$6613 ( \7301 , \7288 , \7300 );
nand \U$6614 ( \7302 , \7275 , \7301 );
not \U$6615 ( \7303 , \7302 );
not \U$6616 ( \7304 , \7303 );
and \U$6617 ( \7305 , \7304 , \6597 );
not \U$6618 ( \7306 , \7304 );
and \U$6619 ( \7307 , \7306 , \6034 );
nor \U$6620 ( \7308 , \7305 , \7307 );
nand \U$6621 ( \7309 , \6030 , \7308 );
not \U$6622 ( \7310 , \7309 );
not \U$6623 ( \7311 , \7180 );
or \U$6624 ( \7312 , \7310 , \7311 );
not \U$6625 ( \7313 , \7150 );
not \U$6626 ( \7314 , \7053 );
or \U$6627 ( \7315 , \7313 , \7314 );
not \U$6628 ( \7316 , \6270 );
nand \U$6629 ( \7317 , \7316 , \7149 );
nand \U$6630 ( \7318 , \7315 , \7317 );
not \U$6631 ( \7319 , \7318 );
not \U$6632 ( \7320 , \6265 );
or \U$6633 ( \7321 , \7319 , \7320 );
nand \U$6634 ( \7322 , \7057 , \6919 );
nand \U$6635 ( \7323 , \7321 , \7322 );
nand \U$6636 ( \7324 , \7312 , \7323 );
not \U$6637 ( \7325 , \7180 );
not \U$6638 ( \7326 , \7309 );
nand \U$6639 ( \7327 , \7325 , \7326 );
nand \U$6640 ( \7328 , \7324 , \7327 );
xor \U$6641 ( \7329 , \7180 , \7165 );
xnor \U$6642 ( \7330 , \7329 , \7157 );
or \U$6643 ( \7331 , \7328 , \7330 );
and \U$6644 ( \7332 , \7255 , \7331 );
and \U$6645 ( \7333 , \7330 , \7328 );
nor \U$6646 ( \7334 , \7332 , \7333 );
xor \U$6647 ( \7335 , \7251 , \7334 );
xor \U$6648 ( \7336 , \1112 , \5711 );
xnor \U$6649 ( \7337 , \7336 , \5796 );
nand \U$6650 ( \7338 , \5968 , \6991 );
buf \U$6651 ( \7339 , \6987 );
not \U$6652 ( \7340 , \7339 );
and \U$6653 ( \7341 , \7338 , \7340 );
not \U$6654 ( \7342 , \7338 );
and \U$6655 ( \7343 , \7342 , \7339 );
nor \U$6656 ( \7344 , \7341 , \7343 );
xnor \U$6657 ( \7345 , \7337 , \7344 );
buf \U$6658 ( \7346 , \7345 );
not \U$6659 ( \7347 , \7346 );
not \U$6660 ( \7348 , \7344 );
not \U$6661 ( \7349 , \7348 );
not \U$6662 ( \7350 , \7349 );
not \U$6663 ( \7351 , \6997 );
or \U$6664 ( \7352 , \7350 , \7351 );
nand \U$6665 ( \7353 , \7348 , \6996 );
nand \U$6666 ( \7354 , \7352 , \7353 );
nand \U$6667 ( \7355 , \7354 , \7345 );
not \U$6668 ( \7356 , \7355 );
or \U$6669 ( \7357 , \7347 , \7356 );
buf \U$6670 ( \7358 , \6997 );
not \U$6671 ( \7359 , \7358 );
nand \U$6672 ( \7360 , \7357 , \7359 );
not \U$6673 ( \7361 , \6172 );
not \U$6674 ( \7362 , \7021 );
or \U$6675 ( \7363 , \7361 , \7362 );
nand \U$6676 ( \7364 , \7022 , \6974 );
nand \U$6677 ( \7365 , \7363 , \7364 );
not \U$6678 ( \7366 , \7365 );
not \U$6679 ( \7367 , \7176 );
or \U$6680 ( \7368 , \7366 , \7367 );
nand \U$6681 ( \7369 , \7174 , \7012 );
nand \U$6682 ( \7370 , \7368 , \7369 );
xor \U$6683 ( \7371 , \7360 , \7370 );
not \U$6684 ( \7372 , \6467 );
buf \U$6685 ( \7373 , \6528 );
not \U$6686 ( \7374 , \7373 );
or \U$6687 ( \7375 , \7372 , \7374 );
nand \U$6688 ( \7376 , \6703 , \6466 );
nand \U$6689 ( \7377 , \7375 , \7376 );
not \U$6690 ( \7378 , \7377 );
not \U$6691 ( \7379 , \6700 );
not \U$6692 ( \7380 , \7379 );
or \U$6693 ( \7381 , \7378 , \7380 );
nand \U$6694 ( \7382 , \7075 , \6981 );
nand \U$6695 ( \7383 , \7381 , \7382 );
and \U$6696 ( \7384 , \7371 , \7383 );
and \U$6697 ( \7385 , \7360 , \7370 );
or \U$6698 ( \7386 , \7384 , \7385 );
xor \U$6699 ( \7387 , \7080 , \7099 );
xor \U$6700 ( \7388 , \7387 , \7110 );
xor \U$6701 ( \7389 , \7386 , \7388 );
not \U$6702 ( \7390 , \6545 );
not \U$6703 ( \7391 , \7086 );
or \U$6704 ( \7392 , \7390 , \7391 );
not \U$6705 ( \7393 , \6596 );
not \U$6706 ( \7394 , \6547 );
or \U$6707 ( \7395 , \7393 , \7394 );
nand \U$6708 ( \7396 , \6496 , \6734 );
nand \U$6709 ( \7397 , \7395 , \7396 );
nand \U$6710 ( \7398 , \7397 , \6540 , \7162 );
nand \U$6711 ( \7399 , \7392 , \7398 );
not \U$6712 ( \7400 , \7399 );
not \U$6713 ( \7401 , \6224 );
not \U$6714 ( \7402 , \7358 );
or \U$6715 ( \7403 , \7401 , \7402 );
nand \U$6716 ( \7404 , \7359 , \6225 );
nand \U$6717 ( \7405 , \7403 , \7404 );
not \U$6718 ( \7406 , \7405 );
nor \U$6719 ( \7407 , \7406 , \7355 );
nor \U$6720 ( \7408 , \7346 , \7358 );
nor \U$6721 ( \7409 , \7407 , \7408 );
buf \U$6722 ( \7410 , \7409 );
nand \U$6723 ( \7411 , \7400 , \7410 );
not \U$6724 ( \7412 , \7411 );
not \U$6725 ( \7413 , \6960 );
not \U$6726 ( \7414 , \6651 );
or \U$6727 ( \7415 , \7413 , \7414 );
nand \U$6728 ( \7416 , \6402 , \7055 );
nand \U$6729 ( \7417 , \7415 , \7416 );
not \U$6730 ( \7418 , \7417 );
not \U$6731 ( \7419 , \6398 );
or \U$6732 ( \7420 , \7418 , \7419 );
nand \U$6733 ( \7421 , \6384 , \7105 );
nand \U$6734 ( \7422 , \7420 , \7421 );
not \U$6735 ( \7423 , \7422 );
or \U$6736 ( \7424 , \7412 , \7423 );
not \U$6737 ( \7425 , \7410 );
nand \U$6738 ( \7426 , \7425 , \7399 );
nand \U$6739 ( \7427 , \7424 , \7426 );
and \U$6740 ( \7428 , \7389 , \7427 );
and \U$6741 ( \7429 , \7386 , \7388 );
or \U$6742 ( \7430 , \7428 , \7429 );
xor \U$6743 ( \7431 , \7330 , \7328 );
not \U$6744 ( \7432 , \7431 );
nand \U$6745 ( \7433 , \7254 , \7432 );
nand \U$6746 ( \7434 , \7253 , \7431 );
nand \U$6747 ( \7435 , \7433 , \7434 );
or \U$6748 ( \7436 , \7430 , \7435 );
xor \U$6749 ( \7437 , \7386 , \7388 );
xor \U$6750 ( \7438 , \7437 , \7427 );
not \U$6751 ( \7439 , \7438 );
and \U$6752 ( \7440 , \6072 , RI992b078_358);
not \U$6753 ( \7441 , RI9922798_578);
not \U$6754 ( \7442 , \6077 );
or \U$6755 ( \7443 , \7441 , \7442 );
not \U$6756 ( \7444 , \2280 );
nand \U$6757 ( \7445 , \7443 , \7444 );
nor \U$6758 ( \7446 , \7440 , \7445 );
not \U$6759 ( \7447 , \6086 );
not \U$6760 ( \7448 , RI9924688_518);
not \U$6761 ( \7449 , \7448 );
and \U$6762 ( \7450 , \7447 , \7449 );
not \U$6763 ( \7451 , RI9925678_498);
nor \U$6764 ( \7452 , \6298 , \7451 );
nor \U$6765 ( \7453 , \7450 , \7452 );
nand \U$6766 ( \7454 , \7446 , \7453 );
nand \U$6767 ( \7455 , \6195 , RI992a718_378);
nand \U$6768 ( \7456 , \6197 , RI992d508_318);
nand \U$6769 ( \7457 , \6191 , RI9923d28_538);
nand \U$6770 ( \7458 , \6199 , RI992f3f8_298);
nand \U$6771 ( \7459 , \7455 , \7456 , \7457 , \7458 );
nor \U$6772 ( \7460 , \7454 , \7459 );
not \U$6773 ( \7461 , RI99316a8_278);
nor \U$6774 ( \7462 , \7461 , \6154 );
not \U$6775 ( \7463 , RI992cba8_338);
nor \U$6776 ( \7464 , \7463 , \6150 );
nor \U$6777 ( \7465 , \7462 , \7464 );
not \U$6778 ( \7466 , \6166 );
not \U$6779 ( \7467 , \2317 );
and \U$6780 ( \7468 , \7466 , \7467 );
nor \U$6781 ( \7469 , \6158 , \2281 );
nor \U$6782 ( \7470 , \7468 , \7469 );
nand \U$6783 ( \7471 , \7465 , \7470 );
not \U$6784 ( \7472 , \6203 );
not \U$6785 ( \7473 , \2285 );
and \U$6786 ( \7474 , \7472 , \7473 );
not \U$6787 ( \7475 , \6131 );
not \U$6788 ( \7476 , \7475 );
not \U$6789 ( \7477 , RI9928648_418);
nor \U$6790 ( \7478 , \7476 , \7477 );
nor \U$6791 ( \7479 , \7474 , \7478 );
not \U$6792 ( \7480 , \6137 );
not \U$6793 ( \7481 , \2302 );
and \U$6794 ( \7482 , \7480 , \7481 );
nor \U$6795 ( \7483 , \6317 , \2320 );
nor \U$6796 ( \7484 , \7482 , \7483 );
nand \U$6797 ( \7485 , \7479 , \7484 );
nor \U$6798 ( \7486 , \7471 , \7485 );
nand \U$6799 ( \7487 , \7460 , \7486 );
buf \U$6800 ( \7488 , \7487 );
and \U$6801 ( \7489 , \7488 , \6597 );
not \U$6802 ( \7490 , \7488 );
and \U$6803 ( \7491 , \7490 , \6034 );
nor \U$6804 ( \7492 , \7489 , \7491 );
nand \U$6805 ( \7493 , \6030 , \7492 );
not \U$6806 ( \7494 , \7493 );
not \U$6807 ( \7495 , \7494 );
not \U$6808 ( \7496 , \6265 );
not \U$6809 ( \7497 , \7304 );
not \U$6810 ( \7498 , \6477 );
or \U$6811 ( \7499 , \7497 , \7498 );
nand \U$6812 ( \7500 , \6271 , \7303 );
nand \U$6813 ( \7501 , \7499 , \7500 );
not \U$6814 ( \7502 , \7501 );
or \U$6815 ( \7503 , \7496 , \7502 );
nand \U$6816 ( \7504 , \6919 , \7318 );
nand \U$6817 ( \7505 , \7503 , \7504 );
not \U$6818 ( \7506 , \7505 );
or \U$6819 ( \7507 , \7495 , \7506 );
not \U$6820 ( \7508 , \7505 );
not \U$6821 ( \7509 , \7508 );
not \U$6822 ( \7510 , \7493 );
or \U$6823 ( \7511 , \7509 , \7510 );
not \U$6824 ( \7512 , \6330 );
not \U$6825 ( \7513 , \7170 );
or \U$6826 ( \7514 , \7512 , \7513 );
nand \U$6827 ( \7515 , \7022 , \6328 );
nand \U$6828 ( \7516 , \7514 , \7515 );
not \U$6829 ( \7517 , \7516 );
not \U$6830 ( \7518 , \7176 );
or \U$6831 ( \7519 , \7517 , \7518 );
nand \U$6832 ( \7520 , \7365 , \7012 );
nand \U$6833 ( \7521 , \7519 , \7520 );
xor \U$6834 ( \7522 , \7409 , \7521 );
not \U$6835 ( \7523 , \6628 );
not \U$6836 ( \7524 , \6807 );
or \U$6837 ( \7525 , \7523 , \7524 );
nand \U$6838 ( \7526 , \6703 , \6632 );
nand \U$6839 ( \7527 , \7525 , \7526 );
not \U$6840 ( \7528 , \7527 );
not \U$6841 ( \7529 , \7379 );
or \U$6842 ( \7530 , \7528 , \7529 );
not \U$6843 ( \7531 , \6692 );
nand \U$6844 ( \7532 , \7377 , \7531 );
nand \U$6845 ( \7533 , \7530 , \7532 );
and \U$6846 ( \7534 , \7522 , \7533 );
and \U$6847 ( \7535 , \7409 , \7521 );
or \U$6848 ( \7536 , \7534 , \7535 );
nand \U$6849 ( \7537 , \7511 , \7536 );
nand \U$6850 ( \7538 , \7507 , \7537 );
not \U$6851 ( \7539 , \7538 );
xor \U$6852 ( \7540 , \7180 , \7323 );
xor \U$6853 ( \7541 , \7540 , \7326 );
buf \U$6854 ( \7542 , \7541 );
nand \U$6855 ( \7543 , \7539 , \7542 );
not \U$6856 ( \7544 , \7543 );
or \U$6857 ( \7545 , \7439 , \7544 );
not \U$6858 ( \7546 , \7542 );
nand \U$6859 ( \7547 , \7546 , \7538 );
nand \U$6860 ( \7548 , \7545 , \7547 );
and \U$6861 ( \7549 , \7436 , \7548 );
and \U$6862 ( \7550 , \7435 , \7430 );
nor \U$6863 ( \7551 , \7549 , \7550 );
nand \U$6864 ( \7552 , \7335 , \7551 );
xor \U$6865 ( \7553 , \7241 , \7250 );
and \U$6866 ( \7554 , \7553 , \7334 );
and \U$6867 ( \7555 , \7241 , \7250 );
or \U$6868 ( \7556 , \7554 , \7555 );
xor \U$6869 ( \7557 , \7045 , \7047 );
xor \U$6870 ( \7558 , \7557 , \7188 );
nand \U$6871 ( \7559 , \7556 , \7558 );
and \U$6872 ( \7560 , \7552 , \7559 );
xor \U$6873 ( \7561 , \7430 , \7435 );
not \U$6874 ( \7562 , \7548 );
xnor \U$6875 ( \7563 , \7561 , \7562 );
xor \U$6876 ( \7564 , \7410 , \7399 );
xnor \U$6877 ( \7565 , \7564 , \7422 );
xor \U$6878 ( \7566 , \7360 , \7370 );
xor \U$6879 ( \7567 , \7566 , \7383 );
or \U$6880 ( \7568 , \7565 , \7567 );
not \U$6881 ( \7569 , \6795 );
not \U$6882 ( \7570 , \6547 );
or \U$6883 ( \7571 , \7569 , \7570 );
nand \U$6884 ( \7572 , \6497 , \6912 );
nand \U$6885 ( \7573 , \7571 , \7572 );
not \U$6886 ( \7574 , \7573 );
not \U$6887 ( \7575 , \6542 );
or \U$6888 ( \7576 , \7574 , \7575 );
nand \U$6889 ( \7577 , \7163 , \7397 );
nand \U$6890 ( \7578 , \7576 , \7577 );
not \U$6891 ( \7579 , \7578 );
not \U$6892 ( \7580 , \7150 );
not \U$6893 ( \7581 , \6651 );
or \U$6894 ( \7582 , \7580 , \7581 );
nand \U$6895 ( \7583 , \6402 , \7149 );
nand \U$6896 ( \7584 , \7582 , \7583 );
not \U$6897 ( \7585 , \7584 );
not \U$6898 ( \7586 , \7033 );
or \U$6899 ( \7587 , \7585 , \7586 );
nand \U$6900 ( \7588 , \6383 , \7417 );
nand \U$6901 ( \7589 , \7587 , \7588 );
not \U$6902 ( \7590 , \7589 );
or \U$6903 ( \7591 , \7579 , \7590 );
or \U$6904 ( \7592 , \7578 , \7589 );
not \U$6905 ( \7593 , \6171 );
buf \U$6906 ( \7594 , \6997 );
not \U$6907 ( \7595 , \7594 );
or \U$6908 ( \7596 , \7593 , \7595 );
not \U$6909 ( \7597 , \6171 );
nand \U$6910 ( \7598 , \7359 , \7597 );
nand \U$6911 ( \7599 , \7596 , \7598 );
not \U$6912 ( \7600 , \7599 );
not \U$6913 ( \7601 , \7355 );
not \U$6914 ( \7602 , \7601 );
or \U$6915 ( \7603 , \7600 , \7602 );
not \U$6916 ( \7604 , \7346 );
nand \U$6917 ( \7605 , \7405 , \7604 );
nand \U$6918 ( \7606 , \7603 , \7605 );
buf \U$6919 ( \7607 , \7337 );
not \U$6920 ( \7608 , \7607 );
nor \U$6921 ( \7609 , \7606 , \7608 );
not \U$6922 ( \7610 , \7609 );
nand \U$6923 ( \7611 , \7592 , \7610 );
nand \U$6924 ( \7612 , \7591 , \7611 );
nand \U$6925 ( \7613 , \7568 , \7612 );
nand \U$6926 ( \7614 , \7565 , \7567 );
nand \U$6927 ( \7615 , \7613 , \7614 );
not \U$6928 ( \7616 , \7488 );
not \U$6929 ( \7617 , \6270 );
or \U$6930 ( \7618 , \7616 , \7617 );
not \U$6931 ( \7619 , \7488 );
nand \U$6932 ( \7620 , \6911 , \7619 );
nand \U$6933 ( \7621 , \7618 , \7620 );
not \U$6934 ( \7622 , \7621 );
not \U$6935 ( \7623 , \6265 );
or \U$6936 ( \7624 , \7622 , \7623 );
nand \U$6937 ( \7625 , \7501 , \6919 );
nand \U$6938 ( \7626 , \7624 , \7625 );
not \U$6939 ( \7627 , \6145 );
not \U$6940 ( \7628 , RI9925f60_479);
not \U$6941 ( \7629 , \7628 );
and \U$6942 ( \7630 , \7627 , \7629 );
nor \U$6943 ( \7631 , \6582 , \2424 );
nor \U$6944 ( \7632 , \7630 , \7631 );
not \U$6945 ( \7633 , \6105 );
not \U$6946 ( \7634 , RI992d490_319);
not \U$6947 ( \7635 , \7634 );
and \U$6948 ( \7636 , \7633 , \7635 );
nor \U$6949 ( \7637 , \6110 , \2431 );
nor \U$6950 ( \7638 , \7636 , \7637 );
nand \U$6951 ( \7639 , \7632 , \7638 );
not \U$6952 ( \7640 , RI99285d0_419);
not \U$6953 ( \7641 , \6206 );
or \U$6954 ( \7642 , \7640 , \7641 );
nand \U$6955 ( \7643 , \6204 , RI9927c70_439);
nand \U$6956 ( \7644 , \7642 , \7643 );
nor \U$6957 ( \7645 , \7639 , \7644 );
and \U$6958 ( \7646 , \6072 , RI992b000_359);
not \U$6959 ( \7647 , RI9922720_579);
not \U$6960 ( \7648 , \6077 );
or \U$6961 ( \7649 , \7647 , \7648 );
nand \U$6962 ( \7650 , \7649 , \2419 );
nor \U$6963 ( \7651 , \7646 , \7650 );
not \U$6964 ( \7652 , RI9931630_279);
nor \U$6965 ( \7653 , \7652 , \6154 );
not \U$6966 ( \7654 , RI992cb30_339);
nor \U$6967 ( \7655 , \7654 , \6150 );
nor \U$6968 ( \7656 , \7653 , \7655 );
nand \U$6969 ( \7657 , \7651 , \7656 );
not \U$6970 ( \7658 , RI9925600_499);
not \U$6971 ( \7659 , \6184 );
or \U$6972 ( \7660 , \7658 , \7659 );
nand \U$6973 ( \7661 , \6182 , RI9924610_519);
nand \U$6974 ( \7662 , \7660 , \7661 );
nor \U$6975 ( \7663 , \7657 , \7662 );
not \U$6976 ( \7664 , RI992a6a0_379);
not \U$6977 ( \7665 , \6195 );
or \U$6978 ( \7666 , \7664 , \7665 );
nand \U$6979 ( \7667 , \6191 , RI9923cb0_539);
nand \U$6980 ( \7668 , \7666 , \7667 );
not \U$6981 ( \7669 , RI9928f30_399);
not \U$6982 ( \7670 , \6778 );
or \U$6983 ( \7671 , \7669 , \7670 );
nand \U$6984 ( \7672 , \6213 , RI99268c0_459);
nand \U$6985 ( \7673 , \7671 , \7672 );
nor \U$6986 ( \7674 , \7668 , \7673 );
nand \U$6987 ( \7675 , \7645 , \7663 , \7674 );
not \U$6988 ( \7676 , \7675 );
buf \U$6989 ( \7677 , \7676 );
not \U$6990 ( \7678 , \7677 );
and \U$6991 ( \7679 , \7678 , \6796 );
not \U$6992 ( \7680 , \7678 );
and \U$6993 ( \7681 , \7680 , \7154 );
nor \U$6994 ( \7682 , \7679 , \7681 );
nand \U$6995 ( \7683 , \6029 , \7682 );
not \U$6996 ( \7684 , \7683 );
or \U$6997 ( \7685 , \7626 , \7684 );
not \U$6998 ( \7686 , \6596 );
not \U$6999 ( \7687 , \6970 );
or \U$7000 ( \7688 , \7686 , \7687 );
nand \U$7001 ( \7689 , \6703 , \6734 );
nand \U$7002 ( \7690 , \7688 , \7689 );
not \U$7003 ( \7691 , \7690 );
not \U$7004 ( \7692 , \6978 );
or \U$7005 ( \7693 , \7691 , \7692 );
nand \U$7006 ( \7694 , \7527 , \6981 );
nand \U$7007 ( \7695 , \7693 , \7694 );
not \U$7008 ( \7696 , \7695 );
not \U$7009 ( \7697 , \6467 );
not \U$7010 ( \7698 , \6686 );
not \U$7011 ( \7699 , \7698 );
not \U$7012 ( \7700 , \7699 );
not \U$7013 ( \7701 , \7700 );
or \U$7014 ( \7702 , \7697 , \7701 );
nand \U$7015 ( \7703 , \7020 , \6466 );
nand \U$7016 ( \7704 , \7702 , \7703 );
not \U$7017 ( \7705 , \7704 );
not \U$7018 ( \7706 , \7018 );
or \U$7019 ( \7707 , \7705 , \7706 );
nand \U$7020 ( \7708 , \7516 , \7012 );
nand \U$7021 ( \7709 , \7707 , \7708 );
not \U$7022 ( \7710 , \7709 );
nand \U$7023 ( \7711 , \7696 , \7710 );
and \U$7024 ( \7712 , \6327 , \7594 );
not \U$7025 ( \7713 , \6327 );
not \U$7026 ( \7714 , \7594 );
and \U$7027 ( \7715 , \7713 , \7714 );
or \U$7028 ( \7716 , \7712 , \7715 );
not \U$7029 ( \7717 , \7716 );
and \U$7030 ( \7718 , \7354 , \7345 );
not \U$7031 ( \7719 , \7718 );
or \U$7032 ( \7720 , \7717 , \7719 );
nand \U$7033 ( \7721 , \7599 , \7604 );
nand \U$7034 ( \7722 , \7720 , \7721 );
not \U$7035 ( \7723 , RI994dec0_26);
not \U$7036 ( \7724 , \5873 );
or \U$7037 ( \7725 , \7723 , \7724 );
nand \U$7038 ( \7726 , \7725 , \5796 );
not \U$7039 ( \7727 , \7726 );
nand \U$7040 ( \7728 , \7727 , \7607 );
not \U$7041 ( \7729 , \7728 );
not \U$7042 ( \7730 , \7729 );
and \U$7043 ( \7731 , \6224 , \7608 );
not \U$7044 ( \7732 , \6224 );
and \U$7045 ( \7733 , \7732 , \7607 );
or \U$7046 ( \7734 , \7731 , \7733 );
not \U$7047 ( \7735 , \7734 );
or \U$7048 ( \7736 , \7730 , \7735 );
buf \U$7049 ( \7737 , \7726 );
nand \U$7050 ( \7738 , \7607 , \7737 );
nand \U$7051 ( \7739 , \7736 , \7738 );
nand \U$7052 ( \7740 , \7722 , \7739 );
not \U$7053 ( \7741 , \7740 );
and \U$7054 ( \7742 , \7711 , \7741 );
and \U$7055 ( \7743 , \7695 , \7709 );
nor \U$7056 ( \7744 , \7742 , \7743 );
not \U$7057 ( \7745 , \7744 );
nand \U$7058 ( \7746 , \7685 , \7745 );
nand \U$7059 ( \7747 , \7626 , \7684 );
nand \U$7060 ( \7748 , \7746 , \7747 );
xor \U$7061 ( \7749 , \7493 , \7505 );
not \U$7062 ( \7750 , \7536 );
xor \U$7063 ( \7751 , \7749 , \7750 );
xor \U$7064 ( \7752 , \7748 , \7751 );
xor \U$7065 ( \7753 , \7610 , \7589 );
xnor \U$7066 ( \7754 , \7753 , \7578 );
xor \U$7067 ( \7755 , \7409 , \7521 );
xor \U$7068 ( \7756 , \7755 , \7533 );
not \U$7069 ( \7757 , \7756 );
nand \U$7070 ( \7758 , \7754 , \7757 );
not \U$7071 ( \7759 , \7758 );
not \U$7072 ( \7760 , \7606 );
not \U$7073 ( \7761 , \7608 );
or \U$7074 ( \7762 , \7760 , \7761 );
nand \U$7075 ( \7763 , \7762 , \7610 );
not \U$7076 ( \7764 , \6960 );
not \U$7077 ( \7765 , \6547 );
or \U$7078 ( \7766 , \7764 , \7765 );
nand \U$7079 ( \7767 , \7084 , \7055 );
nand \U$7080 ( \7768 , \7766 , \7767 );
not \U$7081 ( \7769 , \7768 );
not \U$7082 ( \7770 , \6542 );
or \U$7083 ( \7771 , \7769 , \7770 );
nand \U$7084 ( \7772 , \7573 , \6546 );
nand \U$7085 ( \7773 , \7771 , \7772 );
xor \U$7086 ( \7774 , \7763 , \7773 );
not \U$7087 ( \7775 , \7304 );
not \U$7088 ( \7776 , \6651 );
or \U$7089 ( \7777 , \7775 , \7776 );
nand \U$7090 ( \7778 , \6652 , \7303 );
nand \U$7091 ( \7779 , \7777 , \7778 );
not \U$7092 ( \7780 , \7779 );
not \U$7093 ( \7781 , \6900 );
or \U$7094 ( \7782 , \7780 , \7781 );
nand \U$7095 ( \7783 , \6384 , \7584 );
nand \U$7096 ( \7784 , \7782 , \7783 );
and \U$7097 ( \7785 , \7774 , \7784 );
and \U$7098 ( \7786 , \7763 , \7773 );
or \U$7099 ( \7787 , \7785 , \7786 );
not \U$7100 ( \7788 , \7787 );
or \U$7101 ( \7789 , \7759 , \7788 );
not \U$7102 ( \7790 , \7757 );
not \U$7103 ( \7791 , \7754 );
nand \U$7104 ( \7792 , \7790 , \7791 );
nand \U$7105 ( \7793 , \7789 , \7792 );
and \U$7106 ( \7794 , \7752 , \7793 );
and \U$7107 ( \7795 , \7748 , \7751 );
or \U$7108 ( \7796 , \7794 , \7795 );
xor \U$7109 ( \7797 , \7615 , \7796 );
not \U$7110 ( \7798 , \7438 );
not \U$7111 ( \7799 , \7538 );
not \U$7112 ( \7800 , \7541 );
and \U$7113 ( \7801 , \7799 , \7800 );
and \U$7114 ( \7802 , \7541 , \7538 );
nor \U$7115 ( \7803 , \7801 , \7802 );
not \U$7116 ( \7804 , \7803 );
or \U$7117 ( \7805 , \7798 , \7804 );
or \U$7118 ( \7806 , \7803 , \7438 );
nand \U$7119 ( \7807 , \7805 , \7806 );
and \U$7120 ( \7808 , \7797 , \7807 );
and \U$7121 ( \7809 , \7615 , \7796 );
or \U$7122 ( \7810 , \7808 , \7809 );
nor \U$7123 ( \7811 , \7563 , \7810 );
xor \U$7124 ( \7812 , \7615 , \7796 );
xor \U$7125 ( \7813 , \7812 , \7807 );
xor \U$7126 ( \7814 , \7748 , \7751 );
xor \U$7127 ( \7815 , \7814 , \7793 );
xor \U$7128 ( \7816 , \7567 , \7612 );
xnor \U$7129 ( \7817 , \7816 , \7565 );
not \U$7130 ( \7818 , \7817 );
or \U$7131 ( \7819 , \7815 , \7818 );
not \U$7132 ( \7820 , \7678 );
not \U$7133 ( \7821 , \7053 );
or \U$7134 ( \7822 , \7820 , \7821 );
nand \U$7135 ( \7823 , \6911 , \7677 );
nand \U$7136 ( \7824 , \7822 , \7823 );
not \U$7137 ( \7825 , \7824 );
and \U$7138 ( \7826 , \6262 , \6263 );
not \U$7139 ( \7827 , \7826 );
or \U$7140 ( \7828 , \7825 , \7827 );
nand \U$7141 ( \7829 , \7621 , \6253 );
nand \U$7142 ( \7830 , \7828 , \7829 );
not \U$7143 ( \7831 , \7830 );
nand \U$7144 ( \7832 , \6210 , RI99232d8_560);
nand \U$7145 ( \7833 , \6318 , RI9925ee8_480);
and \U$7146 ( \7834 , \7475 , RI9928558_420);
and \U$7147 ( \7835 , \6204 , RI9927bf8_440);
nor \U$7148 ( \7836 , \7834 , \7835 );
nand \U$7149 ( \7837 , \7832 , \7833 , \7836 );
not \U$7150 ( \7838 , \6150 );
not \U$7151 ( \7839 , \2776 );
and \U$7152 ( \7840 , \7838 , \7839 );
not \U$7153 ( \7841 , RI99315b8_280);
not \U$7154 ( \7842 , \6153 );
nor \U$7155 ( \7843 , \7841 , \7842 );
nor \U$7156 ( \7844 , \7840 , \7843 );
not \U$7157 ( \7845 , \6164 );
not \U$7158 ( \7846 , \2786 );
and \U$7159 ( \7847 , \7845 , \7846 );
and \U$7160 ( \7848 , \6220 , RI9928eb8_400);
nor \U$7161 ( \7849 , \7847 , \7848 );
nand \U$7162 ( \7850 , \7844 , \7849 );
nor \U$7163 ( \7851 , \7837 , \7850 );
not \U$7164 ( \7852 , \6086 );
not \U$7165 ( \7853 , RI9924598_520);
not \U$7166 ( \7854 , \7853 );
and \U$7167 ( \7855 , \7852 , \7854 );
nor \U$7168 ( \7856 , \6298 , \2771 );
nor \U$7169 ( \7857 , \7855 , \7856 );
and \U$7170 ( \7858 , \6072 , RI992af88_360);
not \U$7171 ( \7859 , RI99226a8_580);
not \U$7172 ( \7860 , \6077 );
or \U$7173 ( \7861 , \7859 , \7860 );
nand \U$7174 ( \7862 , \7861 , \2747 );
nor \U$7175 ( \7863 , \7858 , \7862 );
nand \U$7176 ( \7864 , \7857 , \7863 );
and \U$7177 ( \7865 , \6197 , RI992d418_320);
and \U$7178 ( \7866 , \6199 , RI992f308_300);
nor \U$7179 ( \7867 , \7865 , \7866 );
and \U$7180 ( \7868 , \6195 , RI992a628_380);
and \U$7181 ( \7869 , \6191 , RI9923c38_540);
nor \U$7182 ( \7870 , \7868 , \7869 );
nand \U$7183 ( \7871 , \7867 , \7870 );
nor \U$7184 ( \7872 , \7864 , \7871 );
nand \U$7185 ( \7873 , \7851 , \7872 );
not \U$7186 ( \7874 , \7873 );
buf \U$7187 ( \7875 , \7874 );
and \U$7188 ( \7876 , \7875 , \6033 );
not \U$7189 ( \7877 , \7875 );
and \U$7190 ( \7878 , \7877 , \6032 );
nor \U$7191 ( \7879 , \7876 , \7878 );
nand \U$7192 ( \7880 , \6028 , \7879 );
buf \U$7193 ( \7881 , \7880 );
nand \U$7194 ( \7882 , \7831 , \7881 );
and \U$7195 ( \7883 , \6465 , \7358 );
not \U$7196 ( \7884 , \6465 );
and \U$7197 ( \7885 , \7884 , \7714 );
or \U$7198 ( \7886 , \7883 , \7885 );
not \U$7199 ( \7887 , \7886 );
not \U$7200 ( \7888 , \7718 );
or \U$7201 ( \7889 , \7887 , \7888 );
not \U$7202 ( \7890 , \7346 );
nand \U$7203 ( \7891 , \7716 , \7890 );
nand \U$7204 ( \7892 , \7889 , \7891 );
not \U$7205 ( \7893 , \7729 );
not \U$7206 ( \7894 , \7607 );
not \U$7207 ( \7895 , \7597 );
or \U$7208 ( \7896 , \7894 , \7895 );
not \U$7209 ( \7897 , \7607 );
nand \U$7210 ( \7898 , \6171 , \7897 );
nand \U$7211 ( \7899 , \7896 , \7898 );
not \U$7212 ( \7900 , \7899 );
or \U$7213 ( \7901 , \7893 , \7900 );
not \U$7214 ( \7902 , \7737 );
not \U$7215 ( \7903 , \7902 );
nand \U$7216 ( \7904 , \7734 , \7903 );
nand \U$7217 ( \7905 , \7901 , \7904 );
and \U$7218 ( \7906 , \7892 , \7905 );
not \U$7219 ( \7907 , \6628 );
not \U$7220 ( \7908 , \7700 );
or \U$7221 ( \7909 , \7907 , \7908 );
nand \U$7222 ( \7910 , \7020 , \6632 );
nand \U$7223 ( \7911 , \7909 , \7910 );
not \U$7224 ( \7912 , \7911 );
not \U$7225 ( \7913 , \7018 );
or \U$7226 ( \7914 , \7912 , \7913 );
nand \U$7227 ( \7915 , \7704 , \7012 );
nand \U$7228 ( \7916 , \7914 , \7915 );
xor \U$7229 ( \7917 , \7906 , \7916 );
not \U$7230 ( \7918 , \6795 );
not \U$7231 ( \7919 , \6528 );
or \U$7232 ( \7920 , \7918 , \7919 );
nand \U$7233 ( \7921 , \6703 , \6912 );
nand \U$7234 ( \7922 , \7920 , \7921 );
not \U$7235 ( \7923 , \7922 );
not \U$7236 ( \7924 , \6978 );
or \U$7237 ( \7925 , \7923 , \7924 );
nand \U$7238 ( \7926 , \7690 , \7531 );
nand \U$7239 ( \7927 , \7925 , \7926 );
and \U$7240 ( \7928 , \7917 , \7927 );
and \U$7241 ( \7929 , \7906 , \7916 );
or \U$7242 ( \7930 , \7928 , \7929 );
buf \U$7243 ( \7931 , \7930 );
and \U$7244 ( \7932 , \7882 , \7931 );
not \U$7245 ( \7933 , \7830 );
nor \U$7246 ( \7934 , \7933 , \7881 );
nor \U$7247 ( \7935 , \7932 , \7934 );
not \U$7248 ( \7936 , \7935 );
xor \U$7249 ( \7937 , \7683 , \7626 );
xnor \U$7250 ( \7938 , \7937 , \7744 );
not \U$7251 ( \7939 , \7938 );
or \U$7252 ( \7940 , \7936 , \7939 );
xor \U$7253 ( \7941 , \7740 , \7709 );
xnor \U$7254 ( \7942 , \7941 , \7695 );
not \U$7255 ( \7943 , \7942 );
not \U$7256 ( \7944 , \7739 );
not \U$7257 ( \7945 , \7944 );
not \U$7258 ( \7946 , \7722 );
or \U$7259 ( \7947 , \7945 , \7946 );
or \U$7260 ( \7948 , \7722 , \7944 );
nand \U$7261 ( \7949 , \7947 , \7948 );
not \U$7262 ( \7950 , \7150 );
not \U$7263 ( \7951 , \7093 );
or \U$7264 ( \7952 , \7950 , \7951 );
nand \U$7265 ( \7953 , \7084 , \7149 );
nand \U$7266 ( \7954 , \7952 , \7953 );
not \U$7267 ( \7955 , \7954 );
not \U$7268 ( \7956 , \7089 );
or \U$7269 ( \7957 , \7955 , \7956 );
nand \U$7270 ( \7958 , \7768 , \6545 );
nand \U$7271 ( \7959 , \7957 , \7958 );
xor \U$7272 ( \7960 , \7949 , \7959 );
not \U$7273 ( \7961 , \7488 );
not \U$7274 ( \7962 , \6391 );
or \U$7275 ( \7963 , \7961 , \7962 );
nand \U$7276 ( \7964 , \6652 , \7619 );
nand \U$7277 ( \7965 , \7963 , \7964 );
not \U$7278 ( \7966 , \7965 );
not \U$7279 ( \7967 , \7034 );
or \U$7280 ( \7968 , \7966 , \7967 );
nand \U$7281 ( \7969 , \6383 , \7779 );
nand \U$7282 ( \7970 , \7968 , \7969 );
and \U$7283 ( \7971 , \7960 , \7970 );
and \U$7284 ( \7972 , \7949 , \7959 );
or \U$7285 ( \7973 , \7971 , \7972 );
not \U$7286 ( \7974 , \7973 );
or \U$7287 ( \7975 , \7943 , \7974 );
or \U$7288 ( \7976 , \7942 , \7973 );
xor \U$7289 ( \7977 , \7763 , \7773 );
xor \U$7290 ( \7978 , \7977 , \7784 );
nand \U$7291 ( \7979 , \7976 , \7978 );
nand \U$7292 ( \7980 , \7975 , \7979 );
nand \U$7293 ( \7981 , \7940 , \7980 );
not \U$7294 ( \7982 , \7938 );
not \U$7295 ( \7983 , \7935 );
nand \U$7296 ( \7984 , \7982 , \7983 );
nand \U$7297 ( \7985 , \7981 , \7984 );
nand \U$7298 ( \7986 , \7819 , \7985 );
nand \U$7299 ( \7987 , \7815 , \7818 );
nand \U$7300 ( \7988 , \7986 , \7987 );
nor \U$7301 ( \7989 , \7813 , \7988 );
nor \U$7302 ( \7990 , \7811 , \7989 );
nand \U$7303 ( \7991 , \7560 , \7990 );
not \U$7304 ( \7992 , \7991 );
not \U$7305 ( \7993 , \7992 );
nor \U$7306 ( \7994 , \7239 , \7993 );
not \U$7307 ( \7995 , \7994 );
nand \U$7308 ( \7996 , \6768 , \6794 );
and \U$7309 ( \7997 , \7996 , \7594 );
not \U$7310 ( \7998 , \7996 );
not \U$7311 ( \7999 , \7594 );
and \U$7312 ( \8000 , \7998 , \7999 );
or \U$7313 ( \8001 , \7997 , \8000 );
not \U$7314 ( \8002 , \8001 );
not \U$7315 ( \8003 , \7601 );
or \U$7316 ( \8004 , \8002 , \8003 );
and \U$7317 ( \8005 , \6595 , \7594 );
not \U$7318 ( \8006 , \6595 );
and \U$7319 ( \8007 , \8006 , \7999 );
or \U$7320 ( \8008 , \8005 , \8007 );
nand \U$7321 ( \8009 , \8008 , \7604 );
nand \U$7322 ( \8010 , \8004 , \8009 );
and \U$7323 ( \8011 , \7607 , \6467 );
not \U$7324 ( \8012 , \7607 );
and \U$7325 ( \8013 , \8012 , \6466 );
nor \U$7326 ( \8014 , \8011 , \8013 );
not \U$7327 ( \8015 , \8014 );
not \U$7328 ( \8016 , \7903 );
or \U$7329 ( \8017 , \8015 , \8016 );
and \U$7330 ( \8018 , \7897 , \6627 );
not \U$7331 ( \8019 , \7897 );
not \U$7332 ( \8020 , \6627 );
and \U$7333 ( \8021 , \8019 , \8020 );
nor \U$7334 ( \8022 , \8018 , \8021 );
not \U$7335 ( \8023 , \8022 );
nand \U$7336 ( \8024 , \8023 , \7729 );
nand \U$7337 ( \8025 , \8017 , \8024 );
nand \U$7338 ( \8026 , \8010 , \8025 );
not \U$7339 ( \8027 , \6960 );
not \U$7340 ( \8028 , \7700 );
or \U$7341 ( \8029 , \8027 , \8028 );
not \U$7342 ( \8030 , \7698 );
nand \U$7343 ( \8031 , \8030 , \7055 );
nand \U$7344 ( \8032 , \8029 , \8031 );
not \U$7345 ( \8033 , \8032 );
not \U$7346 ( \8034 , \7018 );
or \U$7347 ( \8035 , \8033 , \8034 );
not \U$7348 ( \8036 , \6795 );
not \U$7349 ( \8037 , \7170 );
or \U$7350 ( \8038 , \8036 , \8037 );
nand \U$7351 ( \8039 , \8030 , \6912 );
nand \U$7352 ( \8040 , \8038 , \8039 );
nand \U$7353 ( \8041 , \8040 , \7012 );
nand \U$7354 ( \8042 , \8035 , \8041 );
xor \U$7355 ( \8043 , \8026 , \8042 );
not \U$7356 ( \8044 , \6970 );
not \U$7357 ( \8045 , \7304 );
or \U$7358 ( \8046 , \8044 , \8045 );
nand \U$7359 ( \8047 , \6703 , \7303 );
nand \U$7360 ( \8048 , \8046 , \8047 );
not \U$7361 ( \8049 , \8048 );
not \U$7362 ( \8050 , \7379 );
or \U$7363 ( \8051 , \8049 , \8050 );
not \U$7364 ( \8052 , \7150 );
not \U$7365 ( \8053 , \6803 );
or \U$7366 ( \8054 , \8052 , \8053 );
nand \U$7367 ( \8055 , \6703 , \7149 );
nand \U$7368 ( \8056 , \8054 , \8055 );
nand \U$7369 ( \8057 , \8056 , \6981 );
nand \U$7370 ( \8058 , \8051 , \8057 );
xor \U$7371 ( \8059 , \8043 , \8058 );
and \U$7372 ( \8060 , \6197 , RI992d328_322);
and \U$7373 ( \8061 , \6199 , RI992f218_302);
nor \U$7374 ( \8062 , \8060 , \8061 );
and \U$7375 ( \8063 , \6195 , RI992a538_382);
and \U$7376 ( \8064 , \6191 , RI9923b48_542);
nor \U$7377 ( \8065 , \8063 , \8064 );
nand \U$7378 ( \8066 , \8062 , \8065 );
not \U$7379 ( \8067 , RI99244a8_522);
nor \U$7380 ( \8068 , \6086 , \8067 );
not \U$7381 ( \8069 , RI9924e08_502);
nor \U$7382 ( \8070 , \8069 , \6296 );
nor \U$7383 ( \8071 , \8068 , \8070 );
and \U$7384 ( \8072 , \6072 , RI992ae98_362);
not \U$7385 ( \8073 , RI99225b8_582);
not \U$7386 ( \8074 , \6077 );
or \U$7387 ( \8075 , \8073 , \8074 );
nand \U$7388 ( \8076 , \8075 , \2493 );
nor \U$7389 ( \8077 , \8072 , \8076 );
nand \U$7390 ( \8078 , \8071 , \8077 );
nor \U$7391 ( \8079 , \8066 , \8078 );
and \U$7392 ( \8080 , \6210 , RI99231e8_562);
and \U$7393 ( \8081 , \6318 , RI9925df8_482);
nor \U$7394 ( \8082 , \8080 , \8081 );
and \U$7395 ( \8083 , \7475 , RI9928468_422);
and \U$7396 ( \8084 , \6204 , RI9927b08_442);
nor \U$7397 ( \8085 , \8083 , \8084 );
nand \U$7398 ( \8086 , \8082 , \8085 );
not \U$7399 ( \8087 , \6150 );
not \U$7400 ( \8088 , \2488 );
and \U$7401 ( \8089 , \8087 , \8088 );
not \U$7402 ( \8090 , RI99314c8_282);
nor \U$7403 ( \8091 , \8090 , \7842 );
nor \U$7404 ( \8092 , \8089 , \8091 );
not \U$7405 ( \8093 , \6164 );
not \U$7406 ( \8094 , \2508 );
and \U$7407 ( \8095 , \8093 , \8094 );
and \U$7408 ( \8096 , \6220 , RI9928dc8_402);
nor \U$7409 ( \8097 , \8095 , \8096 );
nand \U$7410 ( \8098 , \8092 , \8097 );
nor \U$7411 ( \8099 , \8086 , \8098 );
nand \U$7412 ( \8100 , \8079 , \8099 );
not \U$7413 ( \8101 , \8100 );
not \U$7414 ( \8102 , \8101 );
and \U$7415 ( \8103 , \8102 , \6250 );
not \U$7416 ( \8104 , \8102 );
not \U$7417 ( \8105 , \6391 );
and \U$7418 ( \8106 , \8104 , \8105 );
nor \U$7419 ( \8107 , \8103 , \8106 );
not \U$7420 ( \8108 , \8107 );
not \U$7421 ( \8109 , \8108 );
not \U$7422 ( \8110 , \6900 );
or \U$7423 ( \8111 , \8109 , \8110 );
not \U$7424 ( \8112 , RI9924520_521);
nor \U$7425 ( \8113 , \8112 , \6086 );
not \U$7426 ( \8114 , RI9925510_501);
nor \U$7427 ( \8115 , \8114 , \6298 );
nor \U$7428 ( \8116 , \8113 , \8115 );
and \U$7429 ( \8117 , \6072 , RI992af10_361);
not \U$7430 ( \8118 , \2541 );
nand \U$7431 ( \8119 , \6077 , RI9922630_581);
nand \U$7432 ( \8120 , \8118 , \8119 );
nor \U$7433 ( \8121 , \8117 , \8120 );
nand \U$7434 ( \8122 , \8116 , \8121 );
nand \U$7435 ( \8123 , \6191 , RI9923bc0_541);
nand \U$7436 ( \8124 , \6195 , RI992a5b0_381);
nand \U$7437 ( \8125 , \6197 , RI992d3a0_321);
nand \U$7438 ( \8126 , \6199 , RI992f290_301);
nand \U$7439 ( \8127 , \8123 , \8124 , \8125 , \8126 );
nor \U$7440 ( \8128 , \8122 , \8127 );
nand \U$7441 ( \8129 , \6204 , RI9927b80_441);
nand \U$7442 ( \8130 , \6442 , RI99284e0_421);
nand \U$7443 ( \8131 , \6210 , RI9923260_561);
nand \U$7444 ( \8132 , \6318 , RI9925e70_481);
nand \U$7445 ( \8133 , \8129 , \8130 , \8131 , \8132 );
nand \U$7446 ( \8134 , \6216 , RI992ca40_341);
nand \U$7447 ( \8135 , \6153 , RI9931540_281);
nand \U$7448 ( \8136 , \6220 , RI9928e40_401);
nand \U$7449 ( \8137 , \6213 , RI99267d0_461);
nand \U$7450 ( \8138 , \8134 , \8135 , \8136 , \8137 );
nor \U$7451 ( \8139 , \8133 , \8138 );
nand \U$7452 ( \8140 , \8128 , \8139 );
buf \U$7453 ( \8141 , \8140 );
not \U$7454 ( \8142 , \8141 );
not \U$7455 ( \8143 , \8142 );
not \U$7456 ( \8144 , \6652 );
or \U$7457 ( \8145 , \8143 , \8144 );
not \U$7458 ( \8146 , \6402 );
nand \U$7459 ( \8147 , \8146 , \8141 );
nand \U$7460 ( \8148 , \8145 , \8147 );
nand \U$7461 ( \8149 , \6383 , \8148 );
nand \U$7462 ( \8150 , \8111 , \8149 );
not \U$7463 ( \8151 , \8150 );
not \U$7464 ( \8152 , \7875 );
not \U$7465 ( \8153 , \8152 );
not \U$7466 ( \8154 , \7093 );
or \U$7467 ( \8155 , \8153 , \8154 );
nand \U$7468 ( \8156 , \6496 , \7875 );
nand \U$7469 ( \8157 , \8155 , \8156 );
not \U$7470 ( \8158 , \8157 );
not \U$7471 ( \8159 , \6542 );
or \U$7472 ( \8160 , \8158 , \8159 );
not \U$7473 ( \8161 , \7678 );
not \U$7474 ( \8162 , \6547 );
or \U$7475 ( \8163 , \8161 , \8162 );
not \U$7476 ( \8164 , \7093 );
nand \U$7477 ( \8165 , \8164 , \7677 );
nand \U$7478 ( \8166 , \8163 , \8165 );
nand \U$7479 ( \8167 , \8166 , \7163 );
nand \U$7480 ( \8168 , \8160 , \8167 );
not \U$7481 ( \8169 , \8168 );
nand \U$7482 ( \8170 , \8151 , \8169 );
xor \U$7483 ( \8171 , \8010 , \8025 );
and \U$7484 ( \8172 , \8170 , \8171 );
and \U$7485 ( \8173 , \8150 , \8168 );
nor \U$7486 ( \8174 , \8172 , \8173 );
not \U$7487 ( \8175 , \8174 );
xor \U$7488 ( \8176 , \8059 , \8175 );
not \U$7489 ( \8177 , \7729 );
not \U$7490 ( \8178 , \8014 );
or \U$7491 ( \8179 , \8177 , \8178 );
not \U$7492 ( \8180 , \7607 );
not \U$7493 ( \8181 , \6328 );
or \U$7494 ( \8182 , \8180 , \8181 );
nand \U$7495 ( \8183 , \6327 , \7608 );
nand \U$7496 ( \8184 , \8182 , \8183 );
nand \U$7497 ( \8185 , \8184 , \7737 );
nand \U$7498 ( \8186 , \8179 , \8185 );
not \U$7499 ( \8187 , \8008 );
not \U$7500 ( \8188 , \7601 );
or \U$7501 ( \8189 , \8187 , \8188 );
not \U$7502 ( \8190 , \6627 );
not \U$7503 ( \8191 , \7594 );
or \U$7504 ( \8192 , \8190 , \8191 );
nand \U$7505 ( \8193 , \7714 , \8020 );
nand \U$7506 ( \8194 , \8192 , \8193 );
nand \U$7507 ( \8195 , \8194 , \7890 );
nand \U$7508 ( \8196 , \8189 , \8195 );
xor \U$7509 ( \8197 , \8186 , \8196 );
not \U$7510 ( \8198 , \8148 );
not \U$7511 ( \8199 , \6397 );
or \U$7512 ( \8200 , \8198 , \8199 );
not \U$7513 ( \8201 , \8152 );
not \U$7514 ( \8202 , \6651 );
or \U$7515 ( \8203 , \8201 , \8202 );
nand \U$7516 ( \8204 , \8105 , \7875 );
nand \U$7517 ( \8205 , \8203 , \8204 );
nand \U$7518 ( \8206 , \6383 , \8205 );
nand \U$7519 ( \8207 , \8200 , \8206 );
xor \U$7520 ( \8208 , \8197 , \8207 );
not \U$7521 ( \8209 , \8166 );
not \U$7522 ( \8210 , \6542 );
or \U$7523 ( \8211 , \8209 , \8210 );
not \U$7524 ( \8212 , \7488 );
not \U$7525 ( \8213 , \6547 );
or \U$7526 ( \8214 , \8212 , \8213 );
nand \U$7527 ( \8215 , \6496 , \7619 );
nand \U$7528 ( \8216 , \8214 , \8215 );
nand \U$7529 ( \8217 , \8216 , \7163 );
nand \U$7530 ( \8218 , \8211 , \8217 );
xor \U$7531 ( \8219 , \8208 , \8218 );
xnor \U$7532 ( \8220 , \8176 , \8219 );
nor \U$7533 ( \8221 , \6150 , \3498 );
not \U$7534 ( \8222 , RI9931360_285);
nor \U$7535 ( \8223 , \8222 , \6771 );
nor \U$7536 ( \8224 , \8221 , \8223 );
not \U$7537 ( \8225 , RI9928c60_405);
nor \U$7538 ( \8226 , \8225 , \6158 );
nor \U$7539 ( \8227 , \6570 , \3485 );
nor \U$7540 ( \8228 , \8226 , \8227 );
nand \U$7541 ( \8229 , \8224 , \8228 );
not \U$7542 ( \8230 , \6582 );
not \U$7543 ( \8231 , \3465 );
and \U$7544 ( \8232 , \8230 , \8231 );
not \U$7545 ( \8233 , \6144 );
nor \U$7546 ( \8234 , \8233 , \3487 );
nor \U$7547 ( \8235 , \8232 , \8234 );
not \U$7548 ( \8236 , \6126 );
not \U$7549 ( \8237 , RI9926f50_445);
not \U$7550 ( \8238 , \8237 );
and \U$7551 ( \8239 , \8236 , \8238 );
not \U$7552 ( \8240 , RI9928300_425);
nor \U$7553 ( \8241 , \7476 , \8240 );
nor \U$7554 ( \8242 , \8239 , \8241 );
nand \U$7555 ( \8243 , \8235 , \8242 );
nor \U$7556 ( \8244 , \8229 , \8243 );
not \U$7557 ( \8245 , RI992a3d0_385);
nor \U$7558 ( \8246 , \8245 , \6113 );
nor \U$7559 ( \8247 , \6120 , \3490 );
nor \U$7560 ( \8248 , \8246 , \8247 );
not \U$7561 ( \8249 , \6105 );
not \U$7562 ( \8250 , \3478 );
and \U$7563 ( \8251 , \8249 , \8250 );
nor \U$7564 ( \8252 , \6110 , \3472 );
nor \U$7565 ( \8253 , \8251 , \8252 );
nand \U$7566 ( \8254 , \8248 , \8253 );
and \U$7567 ( \8255 , \6072 , RI992ad30_365);
not \U$7568 ( \8256 , RI9922450_585);
not \U$7569 ( \8257 , \6077 );
or \U$7570 ( \8258 , \8256 , \8257 );
nand \U$7571 ( \8259 , \8258 , \3460 );
nor \U$7572 ( \8260 , \8255 , \8259 );
not \U$7573 ( \8261 , \6086 );
not \U$7574 ( \8262 , RI9924340_525);
not \U$7575 ( \8263 , \8262 );
and \U$7576 ( \8264 , \8261 , \8263 );
not \U$7577 ( \8265 , RI9924ca0_505);
nor \U$7578 ( \8266 , \6094 , \8265 );
nor \U$7579 ( \8267 , \8264 , \8266 );
nand \U$7580 ( \8268 , \8260 , \8267 );
nor \U$7581 ( \8269 , \8254 , \8268 );
nand \U$7582 ( \8270 , \8244 , \8269 );
buf \U$7583 ( \8271 , \8270 );
not \U$7584 ( \8272 , \8271 );
and \U$7585 ( \8273 , \6034 , \8272 );
and \U$7586 ( \8274 , \7153 , \8271 );
nor \U$7587 ( \8275 , \8273 , \8274 );
nand \U$7588 ( \8276 , \6029 , \8275 );
not \U$7589 ( \8277 , \8276 );
not \U$7590 ( \8278 , \6095 );
not \U$7591 ( \8279 , RI9924d18_504);
not \U$7592 ( \8280 , \8279 );
and \U$7593 ( \8281 , \8278 , \8280 );
not \U$7594 ( \8282 , RI99243b8_524);
nor \U$7595 ( \8283 , \6086 , \8282 );
nor \U$7596 ( \8284 , \8281 , \8283 );
and \U$7597 ( \8285 , \6072 , RI992ada8_364);
not \U$7598 ( \8286 , \3141 );
nand \U$7599 ( \8287 , \6077 , RI99224c8_584);
nand \U$7600 ( \8288 , \8286 , \8287 );
nor \U$7601 ( \8289 , \8285 , \8288 );
nand \U$7602 ( \8290 , \8284 , \8289 );
nand \U$7603 ( \8291 , \6191 , RI9923a58_544);
nand \U$7604 ( \8292 , \6195 , RI992a448_384);
nand \U$7605 ( \8293 , \6197 , RI992d238_324);
nand \U$7606 ( \8294 , \6199 , RI992f128_304);
nand \U$7607 ( \8295 , \8291 , \8292 , \8293 , \8294 );
nor \U$7608 ( \8296 , \8290 , \8295 );
nand \U$7609 ( \8297 , \6204 , RI9926fc8_444);
nand \U$7610 ( \8298 , \6442 , RI9928378_424);
nand \U$7611 ( \8299 , \6210 , RI99230f8_564);
nand \U$7612 ( \8300 , \6318 , RI9925d08_484);
nand \U$7613 ( \8301 , \8297 , \8298 , \8299 , \8300 );
nand \U$7614 ( \8302 , \6216 , RI992c8d8_344);
nand \U$7615 ( \8303 , \6153 , RI99313d8_284);
nand \U$7616 ( \8304 , \6220 , RI9928cd8_404);
nand \U$7617 ( \8305 , \6213 , RI9926668_464);
nand \U$7618 ( \8306 , \8302 , \8303 , \8304 , \8305 );
nor \U$7619 ( \8307 , \8301 , \8306 );
nand \U$7620 ( \8308 , \8296 , \8307 );
not \U$7621 ( \8309 , \8308 );
not \U$7622 ( \8310 , \8309 );
not \U$7623 ( \8311 , \8310 );
not \U$7624 ( \8312 , \6477 );
or \U$7625 ( \8313 , \8311 , \8312 );
nand \U$7626 ( \8314 , \6911 , \8309 );
nand \U$7627 ( \8315 , \8313 , \8314 );
not \U$7628 ( \8316 , \8315 );
not \U$7629 ( \8317 , \6265 );
or \U$7630 ( \8318 , \8316 , \8317 );
and \U$7631 ( \8319 , \6072 , RI992ae20_363);
nand \U$7632 ( \8320 , \6077 , RI9922540_583);
nand \U$7633 ( \8321 , \8320 , \2611 );
nor \U$7634 ( \8322 , \8319 , \8321 );
not \U$7635 ( \8323 , \6086 );
not \U$7636 ( \8324 , RI9924430_523);
not \U$7637 ( \8325 , \8324 );
and \U$7638 ( \8326 , \8323 , \8325 );
not \U$7639 ( \8327 , RI9924d90_503);
nor \U$7640 ( \8328 , \6298 , \8327 );
nor \U$7641 ( \8329 , \8326 , \8328 );
nand \U$7642 ( \8330 , \8322 , \8329 );
not \U$7643 ( \8331 , \6105 );
not \U$7644 ( \8332 , RI992d2b0_323);
not \U$7645 ( \8333 , \8332 );
and \U$7646 ( \8334 , \8331 , \8333 );
nor \U$7647 ( \8335 , \6109 , \2604 );
nor \U$7648 ( \8336 , \8334 , \8335 );
not \U$7649 ( \8337 , RI992a4c0_383);
nor \U$7650 ( \8338 , \8337 , \6113 );
not \U$7651 ( \8339 , RI9923ad0_543);
nor \U$7652 ( \8340 , \6120 , \8339 );
nor \U$7653 ( \8341 , \8338 , \8340 );
nand \U$7654 ( \8342 , \8336 , \8341 );
nor \U$7655 ( \8343 , \8330 , \8342 );
not \U$7656 ( \8344 , \6150 );
not \U$7657 ( \8345 , RI992c950_343);
not \U$7658 ( \8346 , \8345 );
and \U$7659 ( \8347 , \8344 , \8346 );
not \U$7660 ( \8348 , RI9931450_283);
nor \U$7661 ( \8349 , \8348 , \7842 );
nor \U$7662 ( \8350 , \8347 , \8349 );
not \U$7663 ( \8351 , \6570 );
not \U$7664 ( \8352 , RI99266e0_463);
not \U$7665 ( \8353 , \8352 );
and \U$7666 ( \8354 , \8351 , \8353 );
nor \U$7667 ( \8355 , \6158 , \2602 );
nor \U$7668 ( \8356 , \8354 , \8355 );
nand \U$7669 ( \8357 , \8350 , \8356 );
not \U$7670 ( \8358 , \6203 );
not \U$7671 ( \8359 , RI9927040_443);
not \U$7672 ( \8360 , \8359 );
and \U$7673 ( \8361 , \8358 , \8360 );
not \U$7674 ( \8362 , RI99283f0_423);
nor \U$7675 ( \8363 , \6132 , \8362 );
nor \U$7676 ( \8364 , \8361 , \8363 );
not \U$7677 ( \8365 , \6138 );
not \U$7678 ( \8366 , \2616 );
and \U$7679 ( \8367 , \8365 , \8366 );
not \U$7680 ( \8368 , RI9925d80_483);
nor \U$7681 ( \8369 , \6317 , \8368 );
nor \U$7682 ( \8370 , \8367 , \8369 );
nand \U$7683 ( \8371 , \8364 , \8370 );
nor \U$7684 ( \8372 , \8357 , \8371 );
nand \U$7685 ( \8373 , \8343 , \8372 );
buf \U$7686 ( \8374 , \8373 );
not \U$7687 ( \8375 , \8374 );
not \U$7688 ( \8376 , \7053 );
or \U$7689 ( \8377 , \8375 , \8376 );
not \U$7690 ( \8378 , \8374 );
nand \U$7691 ( \8379 , \7316 , \8378 );
nand \U$7692 ( \8380 , \8377 , \8379 );
nand \U$7693 ( \8381 , \8380 , \6919 );
nand \U$7694 ( \8382 , \8318 , \8381 );
not \U$7695 ( \8383 , \8382 );
not \U$7696 ( \8384 , \8383 );
or \U$7697 ( \8385 , \8277 , \8384 );
buf \U$7698 ( \8386 , \7302 );
and \U$7699 ( \8387 , \8386 , \7700 );
not \U$7700 ( \8388 , \8386 );
and \U$7701 ( \8389 , \8388 , \7699 );
or \U$7702 ( \8390 , \8387 , \8389 );
not \U$7703 ( \8391 , \8390 );
not \U$7704 ( \8392 , \7018 );
or \U$7705 ( \8393 , \8391 , \8392 );
and \U$7706 ( \8394 , \7148 , \7699 );
not \U$7707 ( \8395 , \7148 );
and \U$7708 ( \8396 , \8395 , \7170 );
or \U$7709 ( \8397 , \8394 , \8396 );
nand \U$7710 ( \8398 , \8397 , \7012 );
nand \U$7711 ( \8399 , \8393 , \8398 );
xor \U$7713 ( \8400 , \8399 , 1'b0 );
not \U$7714 ( \8401 , \7678 );
not \U$7715 ( \8402 , \6803 );
or \U$7716 ( \8403 , \8401 , \8402 );
nand \U$7717 ( \8404 , \6703 , \7677 );
nand \U$7718 ( \8405 , \8403 , \8404 );
not \U$7719 ( \8406 , \8405 );
not \U$7720 ( \8407 , \7379 );
or \U$7721 ( \8408 , \8406 , \8407 );
not \U$7722 ( \8409 , \7488 );
not \U$7723 ( \8410 , \6970 );
or \U$7724 ( \8411 , \8409 , \8410 );
nand \U$7725 ( \8412 , \6703 , \7619 );
nand \U$7726 ( \8413 , \8411 , \8412 );
nand \U$7727 ( \8414 , \8413 , \6981 );
nand \U$7728 ( \8415 , \8408 , \8414 );
and \U$7729 ( \8416 , \8400 , \8415 );
or \U$7731 ( \8417 , \8416 , 1'b0 );
nand \U$7732 ( \8418 , \8385 , \8417 );
not \U$7733 ( \8419 , \8276 );
nand \U$7734 ( \8420 , \8419 , \8382 );
nand \U$7735 ( \8421 , \8418 , \8420 );
and \U$7736 ( \8422 , \8309 , \6034 );
not \U$7737 ( \8423 , \8309 );
and \U$7738 ( \8424 , \8423 , \6796 );
nor \U$7739 ( \8425 , \8422 , \8424 );
and \U$7740 ( \8426 , \6029 , \8425 );
not \U$7741 ( \8427 , \7018 );
not \U$7742 ( \8428 , \8397 );
or \U$7743 ( \8429 , \8427 , \8428 );
nand \U$7744 ( \8430 , \8032 , \7012 );
nand \U$7745 ( \8431 , \8429 , \8430 );
and \U$7746 ( \8432 , \6959 , \7594 );
not \U$7747 ( \8433 , \6959 );
and \U$7748 ( \8434 , \8433 , \7714 );
or \U$7749 ( \8435 , \8432 , \8434 );
not \U$7750 ( \8436 , \8435 );
not \U$7751 ( \8437 , \7718 );
or \U$7752 ( \8438 , \8436 , \8437 );
nand \U$7753 ( \8439 , \8001 , \7890 );
nand \U$7754 ( \8440 , \8438 , \8439 );
not \U$7755 ( \8441 , \8440 );
and \U$7756 ( \8442 , \6595 , \7608 );
not \U$7757 ( \8443 , \6595 );
and \U$7758 ( \8444 , \8443 , \7607 );
or \U$7759 ( \8445 , \8442 , \8444 );
and \U$7760 ( \8446 , \8445 , \7729 );
nor \U$7761 ( \8447 , \8022 , \7902 );
nor \U$7762 ( \8448 , \8446 , \8447 );
nor \U$7763 ( \8449 , \8441 , \8448 );
xor \U$7764 ( \8450 , \8431 , \8449 );
not \U$7765 ( \8451 , \8413 );
not \U$7766 ( \8452 , \6978 );
or \U$7767 ( \8453 , \8451 , \8452 );
not \U$7768 ( \8454 , \6692 );
nand \U$7769 ( \8455 , \8454 , \8048 );
nand \U$7770 ( \8456 , \8453 , \8455 );
and \U$7771 ( \8457 , \8450 , \8456 );
and \U$7772 ( \8458 , \8431 , \8449 );
or \U$7773 ( \8459 , \8457 , \8458 );
xor \U$7774 ( \8460 , \8426 , \8459 );
not \U$7775 ( \8461 , \8102 );
not \U$7776 ( \8462 , \7053 );
or \U$7777 ( \8463 , \8461 , \8462 );
not \U$7778 ( \8464 , \8102 );
nand \U$7779 ( \8465 , \7316 , \8464 );
nand \U$7780 ( \8466 , \8463 , \8465 );
not \U$7781 ( \8467 , \8466 );
or \U$7782 ( \8468 , \8467 , \6254 );
buf \U$7783 ( \8469 , \6262 );
nand \U$7784 ( \8470 , \8380 , \8469 , \6918 );
nand \U$7785 ( \8471 , \8468 , \8470 );
xor \U$7786 ( \8472 , \8460 , \8471 );
xor \U$7787 ( \8473 , \8421 , \8472 );
xor \U$7788 ( \8474 , \8431 , \8449 );
xor \U$7789 ( \8475 , \8474 , \8456 );
not \U$7790 ( \8476 , \8448 );
not \U$7791 ( \8477 , \8440 );
or \U$7792 ( \8478 , \8476 , \8477 );
or \U$7793 ( \8479 , \8440 , \8448 );
nand \U$7794 ( \8480 , \8478 , \8479 );
not \U$7795 ( \8481 , \8142 );
not \U$7796 ( \8482 , \6496 );
or \U$7797 ( \8483 , \8481 , \8482 );
not \U$7798 ( \8484 , \7084 );
nand \U$7799 ( \8485 , \8484 , \8141 );
nand \U$7800 ( \8486 , \8483 , \8485 );
not \U$7801 ( \8487 , \8486 );
not \U$7802 ( \8488 , \7089 );
or \U$7803 ( \8489 , \8487 , \8488 );
nand \U$7804 ( \8490 , \8157 , \6545 );
nand \U$7805 ( \8491 , \8489 , \8490 );
xor \U$7806 ( \8492 , \8480 , \8491 );
and \U$7807 ( \8493 , \8378 , \6402 );
not \U$7808 ( \8494 , \8378 );
and \U$7809 ( \8495 , \8494 , \6651 );
nor \U$7810 ( \8496 , \8493 , \8495 );
or \U$7811 ( \8497 , \8496 , \6396 );
or \U$7812 ( \8498 , \6903 , \8107 );
nand \U$7813 ( \8499 , \8497 , \8498 );
and \U$7814 ( \8500 , \8492 , \8499 );
and \U$7815 ( \8501 , \8480 , \8491 );
or \U$7816 ( \8502 , \8500 , \8501 );
xor \U$7817 ( \8503 , \8475 , \8502 );
not \U$7818 ( \8504 , \6253 );
not \U$7819 ( \8505 , \8315 );
or \U$7820 ( \8506 , \8504 , \8505 );
not \U$7821 ( \8507 , \7053 );
not \U$7822 ( \8508 , \8271 );
or \U$7823 ( \8509 , \8507 , \8508 );
nand \U$7824 ( \8510 , \7316 , \8272 );
nand \U$7825 ( \8511 , \8509 , \8510 );
nand \U$7826 ( \8512 , \8511 , \8469 , \6918 );
nand \U$7827 ( \8513 , \8506 , \8512 );
not \U$7828 ( \8514 , RI99312e8_286);
nor \U$7829 ( \8515 , \8514 , \6771 );
not \U$7830 ( \8516 , RI992c7e8_346);
nor \U$7831 ( \8517 , \8516 , \6150 );
nor \U$7832 ( \8518 , \8515 , \8517 );
not \U$7833 ( \8519 , \6145 );
not \U$7834 ( \8520 , RI9925c18_486);
not \U$7835 ( \8521 , \8520 );
and \U$7836 ( \8522 , \8519 , \8521 );
not \U$7837 ( \8523 , RI9926578_466);
nor \U$7838 ( \8524 , \6570 , \8523 );
nor \U$7839 ( \8525 , \8522 , \8524 );
and \U$7840 ( \8526 , \6072 , RI992acb8_366);
not \U$7841 ( \8527 , RI99223d8_586);
not \U$7842 ( \8528 , \6077 );
or \U$7843 ( \8529 , \8527 , \8528 );
nand \U$7844 ( \8530 , \8529 , \3678 );
nor \U$7845 ( \8531 , \8526 , \8530 );
nand \U$7846 ( \8532 , \8518 , \8525 , \8531 );
not \U$7847 ( \8533 , RI992a358_386);
nor \U$7848 ( \8534 , \8533 , \6113 );
not \U$7849 ( \8535 , RI9923968_546);
nor \U$7850 ( \8536 , \6120 , \8535 );
nor \U$7851 ( \8537 , \8534 , \8536 );
not \U$7852 ( \8538 , \6126 );
not \U$7853 ( \8539 , RI9926ed8_446);
not \U$7854 ( \8540 , \8539 );
and \U$7855 ( \8541 , \8538 , \8540 );
not \U$7856 ( \8542 , RI9928288_426);
nor \U$7857 ( \8543 , \7476 , \8542 );
nor \U$7858 ( \8544 , \8541 , \8543 );
nand \U$7859 ( \8545 , \8537 , \8544 );
nor \U$7860 ( \8546 , \8532 , \8545 );
not \U$7861 ( \8547 , RI9928be8_406);
nor \U$7862 ( \8548 , \8547 , \6158 );
nor \U$7863 ( \8549 , \6582 , \3683 );
nor \U$7864 ( \8550 , \8548 , \8549 );
not \U$7865 ( \8551 , RI992d148_326);
nor \U$7866 ( \8552 , \8551 , \6105 );
nor \U$7867 ( \8553 , \6110 , \3690 );
nor \U$7868 ( \8554 , \8552 , \8553 );
nand \U$7869 ( \8555 , \8550 , \8554 );
not \U$7870 ( \8556 , RI9924c28_506);
not \U$7871 ( \8557 , \6184 );
or \U$7872 ( \8558 , \8556 , \8557 );
nand \U$7873 ( \8559 , \6182 , RI99242c8_526);
nand \U$7874 ( \8560 , \8558 , \8559 );
nor \U$7875 ( \8561 , \8555 , \8560 );
nand \U$7876 ( \8562 , \8546 , \8561 );
buf \U$7877 ( \8563 , \8562 );
and \U$7878 ( \8564 , \8563 , \7153 );
not \U$7879 ( \8565 , \8563 );
and \U$7880 ( \8566 , \8565 , \6033 );
nor \U$7881 ( \8567 , \8564 , \8566 );
nand \U$7882 ( \8568 , \6029 , \8567 );
not \U$7883 ( \8569 , \8568 );
or \U$7884 ( \8570 , \8513 , \8569 );
not \U$7885 ( \8571 , \7729 );
xor \U$7886 ( \8572 , \7607 , \7996 );
not \U$7887 ( \8573 , \8572 );
or \U$7888 ( \8574 , \8571 , \8573 );
nand \U$7889 ( \8575 , \8445 , \7737 );
nand \U$7890 ( \8576 , \8574 , \8575 );
and \U$7891 ( \8577 , \7147 , \7594 );
not \U$7892 ( \8578 , \7147 );
and \U$7893 ( \8579 , \8578 , \7714 );
or \U$7894 ( \8580 , \8577 , \8579 );
not \U$7895 ( \8581 , \8580 );
not \U$7896 ( \8582 , \7601 );
or \U$7897 ( \8583 , \8581 , \8582 );
nand \U$7898 ( \8584 , \8435 , \7604 );
nand \U$7899 ( \8585 , \8583 , \8584 );
or \U$7900 ( \8586 , \8576 , \8585 );
not \U$7901 ( \8587 , \7488 );
not \U$7902 ( \8588 , \7021 );
or \U$7903 ( \8589 , \8587 , \8588 );
nand \U$7904 ( \8590 , \7020 , \7619 );
nand \U$7905 ( \8591 , \8589 , \8590 );
not \U$7906 ( \8592 , \8591 );
not \U$7907 ( \8593 , \7018 );
or \U$7908 ( \8594 , \8592 , \8593 );
nand \U$7909 ( \8595 , \8390 , \7012 );
nand \U$7910 ( \8596 , \8594 , \8595 );
nand \U$7911 ( \8597 , \8586 , \8596 );
nand \U$7912 ( \8598 , \8585 , \8576 );
nand \U$7913 ( \8599 , \8597 , \8598 );
nand \U$7914 ( \8600 , \8570 , \8599 );
nand \U$7915 ( \8601 , \8513 , \8569 );
nand \U$7916 ( \8602 , \8600 , \8601 );
and \U$7917 ( \8603 , \8503 , \8602 );
and \U$7918 ( \8604 , \8475 , \8502 );
or \U$7919 ( \8605 , \8603 , \8604 );
xor \U$7920 ( \8606 , \8473 , \8605 );
xor \U$7921 ( \8607 , \8220 , \8606 );
xor \U$7922 ( \8608 , \8171 , \8150 );
xnor \U$7923 ( \8609 , \8608 , \8169 );
xor \U$7924 ( \8610 , \8276 , \8417 );
xor \U$7925 ( \8611 , \8610 , \8383 );
xor \U$7926 ( \8612 , \8609 , \8611 );
xor \U$7927 ( \8613 , \8475 , \8502 );
xor \U$7928 ( \8614 , \8613 , \8602 );
and \U$7929 ( \8615 , \8612 , \8614 );
and \U$7930 ( \8616 , \8609 , \8611 );
or \U$7931 ( \8617 , \8615 , \8616 );
and \U$7932 ( \8618 , \8607 , \8617 );
not \U$7933 ( \8619 , \8607 );
not \U$7934 ( \8620 , \8617 );
and \U$7935 ( \8621 , \8619 , \8620 );
nor \U$7936 ( \8622 , \8618 , \8621 );
not \U$7937 ( \8623 , \8622 );
xor \U$7938 ( \8624 , \8399 , 1'b0 );
xor \U$7939 ( \8625 , \8624 , \8415 );
not \U$7940 ( \8626 , \8152 );
not \U$7941 ( \8627 , \7373 );
or \U$7942 ( \8628 , \8626 , \8627 );
nand \U$7943 ( \8629 , \6703 , \7875 );
nand \U$7944 ( \8630 , \8628 , \8629 );
not \U$7945 ( \8631 , \8630 );
not \U$7946 ( \8632 , \7379 );
or \U$7947 ( \8633 , \8631 , \8632 );
nand \U$7948 ( \8634 , \8405 , \7531 );
nand \U$7949 ( \8635 , \8633 , \8634 );
not \U$7950 ( \8636 , \8635 );
not \U$7951 ( \8637 , \8636 );
not \U$7952 ( \8638 , \6150 );
not \U$7953 ( \8639 , RI992c770_347);
not \U$7954 ( \8640 , \8639 );
and \U$7955 ( \8641 , \8638 , \8640 );
not \U$7956 ( \8642 , RI992f920_287);
nor \U$7957 ( \8643 , \6771 , \8642 );
nor \U$7958 ( \8644 , \8641 , \8643 );
not \U$7959 ( \8645 , \6166 );
not \U$7960 ( \8646 , \3550 );
and \U$7961 ( \8647 , \8645 , \8646 );
and \U$7962 ( \8648 , \6778 , RI9928b70_407);
nor \U$7963 ( \8649 , \8647 , \8648 );
not \U$7964 ( \8650 , \6203 );
not \U$7965 ( \8651 , RI9926e60_447);
not \U$7966 ( \8652 , \8651 );
and \U$7967 ( \8653 , \8650 , \8652 );
not \U$7968 ( \8654 , \7475 );
not \U$7969 ( \8655 , RI9928210_427);
nor \U$7970 ( \8656 , \8654 , \8655 );
nor \U$7971 ( \8657 , \8653 , \8656 );
not \U$7972 ( \8658 , \6582 );
not \U$7973 ( \8659 , RI9922f90_567);
not \U$7974 ( \8660 , \8659 );
and \U$7975 ( \8661 , \8658 , \8660 );
not \U$7976 ( \8662 , RI9925ba0_487);
nor \U$7977 ( \8663 , \6317 , \8662 );
nor \U$7978 ( \8664 , \8661 , \8663 );
nand \U$7979 ( \8665 , \8644 , \8649 , \8657 , \8664 );
not \U$7980 ( \8666 , RI9924250_527);
nor \U$7981 ( \8667 , \6086 , \8666 );
not \U$7982 ( \8668 , RI9924bb0_507);
nor \U$7983 ( \8669 , \6296 , \8668 );
nor \U$7984 ( \8670 , \8667 , \8669 );
not \U$7985 ( \8671 , \6105 );
not \U$7986 ( \8672 , RI992d0d0_327);
not \U$7987 ( \8673 , \8672 );
and \U$7988 ( \8674 , \8671 , \8673 );
not \U$7989 ( \8675 , RI992efc0_307);
nor \U$7990 ( \8676 , \6110 , \8675 );
nor \U$7991 ( \8677 , \8674 , \8676 );
not \U$7992 ( \8678 , \6113 );
not \U$7993 ( \8679 , RI992a2e0_387);
not \U$7994 ( \8680 , \8679 );
and \U$7995 ( \8681 , \8678 , \8680 );
not \U$7996 ( \8682 , RI99238f0_547);
nor \U$7997 ( \8683 , \6120 , \8682 );
nor \U$7998 ( \8684 , \8681 , \8683 );
and \U$7999 ( \8685 , \6072 , RI992ac40_367);
not \U$8000 ( \8686 , \3572 );
nand \U$8001 ( \8687 , \6077 , RI9922360_587);
nand \U$8002 ( \8688 , \8686 , \8687 );
nor \U$8003 ( \8689 , \8685 , \8688 );
nand \U$8004 ( \8690 , \8670 , \8677 , \8684 , \8689 );
or \U$8005 ( \8691 , \8665 , \8690 );
buf \U$8006 ( \8692 , \8691 );
nand \U$8007 ( \8693 , \6029 , \8692 );
not \U$8008 ( \8694 , \8693 );
or \U$8009 ( \8695 , \8637 , \8694 );
and \U$8010 ( \8696 , \7302 , \7358 );
not \U$8011 ( \8697 , \7302 );
and \U$8012 ( \8698 , \8697 , \7714 );
or \U$8013 ( \8699 , \8696 , \8698 );
not \U$8014 ( \8700 , \8699 );
not \U$8015 ( \8701 , \7718 );
or \U$8016 ( \8702 , \8700 , \8701 );
nand \U$8017 ( \8703 , \8580 , \7890 );
nand \U$8018 ( \8704 , \8702 , \8703 );
not \U$8019 ( \8705 , \7737 );
not \U$8020 ( \8706 , \8572 );
or \U$8021 ( \8707 , \8705 , \8706 );
not \U$8022 ( \8708 , \7607 );
not \U$8023 ( \8709 , \6959 );
not \U$8024 ( \8710 , \8709 );
or \U$8025 ( \8711 , \8708 , \8710 );
nand \U$8026 ( \8712 , \6959 , \7897 );
nand \U$8027 ( \8713 , \8711 , \8712 );
nand \U$8028 ( \8714 , \8713 , \7729 );
nand \U$8029 ( \8715 , \8707 , \8714 );
nand \U$8030 ( \8716 , \8704 , \8715 );
not \U$8031 ( \8717 , \8716 );
nand \U$8032 ( \8718 , \8695 , \8717 );
not \U$8033 ( \8719 , \8693 );
nand \U$8034 ( \8720 , \8719 , \8635 );
nand \U$8035 ( \8721 , \8718 , \8720 );
xor \U$8036 ( \8722 , \8625 , \8721 );
not \U$8037 ( \8723 , \8102 );
not \U$8038 ( \8724 , \6706 );
or \U$8039 ( \8725 , \8723 , \8724 );
nand \U$8040 ( \8726 , \6496 , \8464 );
nand \U$8041 ( \8727 , \8725 , \8726 );
not \U$8042 ( \8728 , \8727 );
not \U$8043 ( \8729 , \7089 );
or \U$8044 ( \8730 , \8728 , \8729 );
nand \U$8045 ( \8731 , \8486 , \7163 );
nand \U$8046 ( \8732 , \8730 , \8731 );
not \U$8047 ( \8733 , \8310 );
not \U$8048 ( \8734 , \6403 );
or \U$8049 ( \8735 , \8733 , \8734 );
not \U$8050 ( \8736 , \6651 );
nand \U$8051 ( \8737 , \8736 , \8309 );
nand \U$8052 ( \8738 , \8735 , \8737 );
not \U$8053 ( \8739 , \8738 );
not \U$8054 ( \8740 , \7034 );
or \U$8055 ( \8741 , \8739 , \8740 );
not \U$8056 ( \8742 , \8496 );
nand \U$8057 ( \8743 , \8742 , \6383 );
nand \U$8058 ( \8744 , \8741 , \8743 );
xor \U$8059 ( \8745 , \8732 , \8744 );
not \U$8060 ( \8746 , \8563 );
not \U$8061 ( \8747 , \7053 );
or \U$8062 ( \8748 , \8746 , \8747 );
not \U$8063 ( \8749 , \8563 );
nand \U$8064 ( \8750 , \7316 , \8749 );
nand \U$8065 ( \8751 , \8748 , \8750 );
not \U$8066 ( \8752 , \8751 );
not \U$8067 ( \8753 , \6265 );
or \U$8068 ( \8754 , \8752 , \8753 );
nand \U$8069 ( \8755 , \8511 , \6253 );
nand \U$8070 ( \8756 , \8754 , \8755 );
and \U$8071 ( \8757 , \8745 , \8756 );
and \U$8072 ( \8758 , \8732 , \8744 );
or \U$8073 ( \8759 , \8757 , \8758 );
and \U$8074 ( \8760 , \8722 , \8759 );
and \U$8075 ( \8761 , \8625 , \8721 );
or \U$8076 ( \8762 , \8760 , \8761 );
not \U$8077 ( \8763 , \8762 );
xor \U$8078 ( \8764 , \8599 , \8569 );
xnor \U$8079 ( \8765 , \8764 , \8513 );
not \U$8080 ( \8766 , \8765 );
not \U$8081 ( \8767 , \8766 );
xor \U$8082 ( \8768 , \8480 , \8491 );
xor \U$8083 ( \8769 , \8768 , \8499 );
not \U$8084 ( \8770 , \8769 );
or \U$8085 ( \8771 , \8767 , \8770 );
not \U$8086 ( \8772 , \8769 );
not \U$8087 ( \8773 , \8772 );
not \U$8088 ( \8774 , \8765 );
or \U$8089 ( \8775 , \8773 , \8774 );
not \U$8090 ( \8776 , \7675 );
not \U$8091 ( \8777 , \7698 );
or \U$8092 ( \8778 , \8776 , \8777 );
nand \U$8093 ( \8779 , \8030 , \7676 );
nand \U$8094 ( \8780 , \8778 , \8779 );
not \U$8095 ( \8781 , \8780 );
not \U$8096 ( \8782 , \7018 );
or \U$8097 ( \8783 , \8781 , \8782 );
nand \U$8098 ( \8784 , \8591 , \7012 );
nand \U$8099 ( \8785 , \8783 , \8784 );
buf \U$8100 ( \8786 , \6025 );
not \U$8101 ( \8787 , \6234 );
not \U$8102 ( \8788 , \6391 );
or \U$8103 ( \8789 , \8787 , \8788 );
nand \U$8104 ( \8790 , \8789 , \8692 );
nand \U$8105 ( \8791 , \6402 , \6256 );
and \U$8106 ( \8792 , \8786 , \8790 , \8791 );
xor \U$8107 ( \8793 , \8785 , \8792 );
not \U$8108 ( \8794 , \8141 );
not \U$8109 ( \8795 , \6807 );
or \U$8110 ( \8796 , \8794 , \8795 );
not \U$8111 ( \8797 , \6807 );
nand \U$8112 ( \8798 , \8797 , \8142 );
nand \U$8113 ( \8799 , \8796 , \8798 );
not \U$8114 ( \8800 , \8799 );
not \U$8115 ( \8801 , \7379 );
or \U$8116 ( \8802 , \8800 , \8801 );
nand \U$8117 ( \8803 , \8630 , \7531 );
nand \U$8118 ( \8804 , \8802 , \8803 );
and \U$8119 ( \8805 , \8793 , \8804 );
and \U$8120 ( \8806 , \8785 , \8792 );
or \U$8121 ( \8807 , \8805 , \8806 );
not \U$8122 ( \8808 , \8807 );
xor \U$8123 ( \8809 , \8585 , \8576 );
buf \U$8124 ( \8810 , \8596 );
xnor \U$8125 ( \8811 , \8809 , \8810 );
nand \U$8126 ( \8812 , \8808 , \8811 );
not \U$8127 ( \8813 , \8812 );
xor \U$8128 ( \8814 , \8715 , \8704 );
not \U$8129 ( \8815 , \7089 );
not \U$8130 ( \8816 , \8374 );
not \U$8131 ( \8817 , \6706 );
or \U$8132 ( \8818 , \8816 , \8817 );
nand \U$8133 ( \8819 , \6496 , \8378 );
nand \U$8134 ( \8820 , \8818 , \8819 );
not \U$8135 ( \8821 , \8820 );
or \U$8136 ( \8822 , \8815 , \8821 );
nand \U$8137 ( \8823 , \8727 , \6545 );
nand \U$8138 ( \8824 , \8822 , \8823 );
xor \U$8139 ( \8825 , \8814 , \8824 );
not \U$8140 ( \8826 , \8271 );
not \U$8141 ( \8827 , \6651 );
or \U$8142 ( \8828 , \8826 , \8827 );
nand \U$8143 ( \8829 , \6402 , \8272 );
nand \U$8144 ( \8830 , \8828 , \8829 );
not \U$8145 ( \8831 , \8830 );
not \U$8146 ( \8832 , \6900 );
or \U$8147 ( \8833 , \8831 , \8832 );
nand \U$8148 ( \8834 , \6383 , \8738 );
nand \U$8149 ( \8835 , \8833 , \8834 );
and \U$8150 ( \8836 , \8825 , \8835 );
and \U$8151 ( \8837 , \8814 , \8824 );
or \U$8152 ( \8838 , \8836 , \8837 );
not \U$8153 ( \8839 , \8838 );
or \U$8154 ( \8840 , \8813 , \8839 );
not \U$8155 ( \8841 , \8811 );
nand \U$8156 ( \8842 , \8841 , \8807 );
nand \U$8157 ( \8843 , \8840 , \8842 );
nand \U$8158 ( \8844 , \8775 , \8843 );
nand \U$8159 ( \8845 , \8771 , \8844 );
not \U$8160 ( \8846 , \8845 );
nand \U$8161 ( \8847 , \8763 , \8846 );
not \U$8162 ( \8848 , \8847 );
xor \U$8163 ( \8849 , \8609 , \8611 );
xor \U$8164 ( \8850 , \8849 , \8614 );
not \U$8165 ( \8851 , \8850 );
or \U$8166 ( \8852 , \8848 , \8851 );
nand \U$8167 ( \8853 , \8762 , \8845 );
nand \U$8168 ( \8854 , \8852 , \8853 );
not \U$8169 ( \8855 , \8854 );
nand \U$8170 ( \8856 , \8623 , \8855 );
nand \U$8171 ( \8857 , \8622 , \8854 );
not \U$8172 ( \8858 , \8850 );
not \U$8173 ( \8859 , \8762 );
not \U$8174 ( \8860 , \8846 );
and \U$8175 ( \8861 , \8859 , \8860 );
and \U$8176 ( \8862 , \8762 , \8846 );
nor \U$8177 ( \8863 , \8861 , \8862 );
not \U$8178 ( \8864 , \8863 );
or \U$8179 ( \8865 , \8858 , \8864 );
or \U$8180 ( \8866 , \8863 , \8850 );
nand \U$8181 ( \8867 , \8865 , \8866 );
xor \U$8182 ( \8868 , \8625 , \8721 );
xor \U$8183 ( \8869 , \8868 , \8759 );
xor \U$8184 ( \8870 , \8716 , \8635 );
xnor \U$8185 ( \8871 , \8870 , \8693 );
not \U$8186 ( \8872 , \8871 );
not \U$8187 ( \8873 , \8872 );
xor \U$8188 ( \8874 , \8732 , \8744 );
xor \U$8189 ( \8875 , \8874 , \8756 );
not \U$8190 ( \8876 , \8875 );
or \U$8191 ( \8877 , \8873 , \8876 );
or \U$8192 ( \8878 , \8875 , \8872 );
not \U$8193 ( \8879 , \7729 );
and \U$8194 ( \8880 , \7147 , \7608 );
not \U$8195 ( \8881 , \7147 );
and \U$8196 ( \8882 , \8881 , \7607 );
or \U$8197 ( \8883 , \8880 , \8882 );
not \U$8198 ( \8884 , \8883 );
or \U$8199 ( \8885 , \8879 , \8884 );
nand \U$8200 ( \8886 , \8713 , \7737 );
nand \U$8201 ( \8887 , \8885 , \8886 );
not \U$8202 ( \8888 , \8887 );
not \U$8203 ( \8889 , \8888 );
nand \U$8204 ( \8890 , \8692 , \6252 );
not \U$8205 ( \8891 , \8890 );
or \U$8206 ( \8892 , \8889 , \8891 );
and \U$8207 ( \8893 , \7487 , \7594 );
not \U$8208 ( \8894 , \7487 );
and \U$8209 ( \8895 , \8894 , \7714 );
or \U$8210 ( \8896 , \8893 , \8895 );
not \U$8211 ( \8897 , \8896 );
not \U$8212 ( \8898 , \7718 );
or \U$8213 ( \8899 , \8897 , \8898 );
not \U$8214 ( \8900 , \7346 );
nand \U$8215 ( \8901 , \8900 , \8699 );
nand \U$8216 ( \8902 , \8899 , \8901 );
nand \U$8217 ( \8903 , \8892 , \8902 );
not \U$8218 ( \8904 , \8890 );
nand \U$8219 ( \8905 , \8904 , \8887 );
nand \U$8220 ( \8906 , \8903 , \8905 );
not \U$8221 ( \8907 , \8152 );
not \U$8222 ( \8908 , \7698 );
or \U$8223 ( \8909 , \8907 , \8908 );
nand \U$8224 ( \8910 , \7699 , \7875 );
nand \U$8225 ( \8911 , \8909 , \8910 );
not \U$8226 ( \8912 , \8911 );
not \U$8227 ( \8913 , \7018 );
or \U$8228 ( \8914 , \8912 , \8913 );
nand \U$8229 ( \8915 , \8780 , \7012 );
nand \U$8230 ( \8916 , \8914 , \8915 );
buf \U$8231 ( \8917 , \7594 );
and \U$8232 ( \8918 , \7675 , \8917 );
not \U$8233 ( \8919 , \7675 );
not \U$8234 ( \8920 , \8917 );
and \U$8235 ( \8921 , \8919 , \8920 );
or \U$8236 ( \8922 , \8918 , \8921 );
not \U$8237 ( \8923 , \8922 );
not \U$8238 ( \8924 , \7601 );
or \U$8239 ( \8925 , \8923 , \8924 );
nand \U$8240 ( \8926 , \8896 , \7604 );
nand \U$8241 ( \8927 , \8925 , \8926 );
not \U$8242 ( \8928 , \7729 );
not \U$8243 ( \8929 , \7607 );
not \U$8244 ( \8930 , \7303 );
or \U$8245 ( \8931 , \8929 , \8930 );
nand \U$8246 ( \8932 , \8386 , \7608 );
nand \U$8247 ( \8933 , \8931 , \8932 );
not \U$8248 ( \8934 , \8933 );
or \U$8249 ( \8935 , \8928 , \8934 );
nand \U$8250 ( \8936 , \8883 , \7903 );
nand \U$8251 ( \8937 , \8935 , \8936 );
and \U$8252 ( \8938 , \8927 , \8937 );
xor \U$8253 ( \8939 , \8916 , \8938 );
not \U$8254 ( \8940 , \8102 );
not \U$8255 ( \8941 , \7373 );
or \U$8256 ( \8942 , \8940 , \8941 );
nand \U$8257 ( \8943 , \8797 , \8464 );
nand \U$8258 ( \8944 , \8942 , \8943 );
not \U$8259 ( \8945 , \8944 );
not \U$8260 ( \8946 , \7379 );
or \U$8261 ( \8947 , \8945 , \8946 );
nand \U$8262 ( \8948 , \8799 , \6981 );
nand \U$8263 ( \8949 , \8947 , \8948 );
and \U$8264 ( \8950 , \8939 , \8949 );
and \U$8265 ( \8951 , \8916 , \8938 );
or \U$8266 ( \8952 , \8950 , \8951 );
xor \U$8267 ( \8953 , \8906 , \8952 );
not \U$8268 ( \8954 , \8692 );
and \U$8269 ( \8955 , \8954 , \6272 );
not \U$8270 ( \8956 , \8954 );
and \U$8271 ( \8957 , \8956 , \6478 );
nor \U$8272 ( \8958 , \8955 , \8957 );
not \U$8273 ( \8959 , \8958 );
not \U$8274 ( \8960 , \6265 );
or \U$8275 ( \8961 , \8959 , \8960 );
nand \U$8276 ( \8962 , \8751 , \6253 );
nand \U$8277 ( \8963 , \8961 , \8962 );
and \U$8278 ( \8964 , \8953 , \8963 );
and \U$8279 ( \8965 , \8906 , \8952 );
or \U$8280 ( \8966 , \8964 , \8965 );
nand \U$8281 ( \8967 , \8878 , \8966 );
nand \U$8282 ( \8968 , \8877 , \8967 );
xor \U$8283 ( \8969 , \8869 , \8968 );
xor \U$8284 ( \8970 , \8769 , \8766 );
xor \U$8285 ( \8971 , \8970 , \8843 );
and \U$8286 ( \8972 , \8969 , \8971 );
and \U$8287 ( \8973 , \8869 , \8968 );
or \U$8288 ( \8974 , \8972 , \8973 );
nand \U$8289 ( \8975 , \8867 , \8974 );
nand \U$8290 ( \8976 , \8857 , \8975 );
nand \U$8291 ( \8977 , \8856 , \8976 );
and \U$8292 ( \8978 , \8196 , \8186 );
not \U$8293 ( \8979 , \8040 );
not \U$8294 ( \8980 , \7176 );
or \U$8295 ( \8981 , \8979 , \8980 );
not \U$8296 ( \8982 , \7021 );
not \U$8297 ( \8983 , \6596 );
or \U$8298 ( \8984 , \8982 , \8983 );
nand \U$8299 ( \8985 , \7022 , \6734 );
nand \U$8300 ( \8986 , \8984 , \8985 );
nand \U$8301 ( \8987 , \8986 , \7012 );
nand \U$8302 ( \8988 , \8981 , \8987 );
xor \U$8303 ( \8989 , \8978 , \8988 );
not \U$8304 ( \8990 , \8056 );
not \U$8305 ( \8991 , \7379 );
or \U$8306 ( \8992 , \8990 , \8991 );
not \U$8307 ( \8993 , \6960 );
not \U$8308 ( \8994 , \6970 );
or \U$8309 ( \8995 , \8993 , \8994 );
nand \U$8310 ( \8996 , \6703 , \7055 );
nand \U$8311 ( \8997 , \8995 , \8996 );
nand \U$8312 ( \8998 , \8997 , \6981 );
nand \U$8313 ( \8999 , \8992 , \8998 );
xor \U$8314 ( \9000 , \8989 , \8999 );
or \U$8315 ( \9001 , \8218 , \8207 );
nand \U$8316 ( \9002 , \9001 , \8197 );
nand \U$8317 ( \9003 , \8207 , \8218 );
and \U$8318 ( \9004 , \9002 , \9003 );
not \U$8319 ( \9005 , \9004 );
xor \U$8320 ( \9006 , \9000 , \9005 );
not \U$8321 ( \9007 , \7737 );
not \U$8322 ( \9008 , \7899 );
or \U$8323 ( \9009 , \9007 , \9008 );
nand \U$8324 ( \9010 , \8184 , \7729 );
nand \U$8325 ( \9011 , \9009 , \9010 );
not \U$8326 ( \9012 , \8194 );
not \U$8327 ( \9013 , \7601 );
or \U$8328 ( \9014 , \9012 , \9013 );
not \U$8329 ( \9015 , \7346 );
nand \U$8330 ( \9016 , \7886 , \9015 );
nand \U$8331 ( \9017 , \9014 , \9016 );
xor \U$8332 ( \9018 , \9011 , \9017 );
not \U$8333 ( \9019 , \8216 );
not \U$8334 ( \9020 , \6542 );
or \U$8335 ( \9021 , \9019 , \9020 );
not \U$8336 ( \9022 , \6547 );
not \U$8337 ( \9023 , \7304 );
or \U$8338 ( \9024 , \9022 , \9023 );
not \U$8339 ( \9025 , \6706 );
nand \U$8340 ( \9026 , \9025 , \7303 );
nand \U$8341 ( \9027 , \9024 , \9026 );
nand \U$8342 ( \9028 , \9027 , \6545 );
nand \U$8343 ( \9029 , \9021 , \9028 );
xor \U$8344 ( \9030 , \9018 , \9029 );
not \U$8345 ( \9031 , \8205 );
or \U$8346 ( \9032 , \9031 , \6396 );
and \U$8347 ( \9033 , \7677 , \6402 );
not \U$8348 ( \9034 , \7677 );
and \U$8349 ( \9035 , \9034 , \6391 );
nor \U$8350 ( \9036 , \9033 , \9035 );
or \U$8351 ( \9037 , \6903 , \9036 );
nand \U$8352 ( \9038 , \9032 , \9037 );
xor \U$8353 ( \9039 , \9030 , \9038 );
xnor \U$8354 ( \9040 , \9006 , \9039 );
xor \U$8355 ( \9041 , \8421 , \8472 );
and \U$8356 ( \9042 , \9041 , \8605 );
and \U$8357 ( \9043 , \8421 , \8472 );
or \U$8358 ( \9044 , \9042 , \9043 );
not \U$8359 ( \9045 , \9044 );
xor \U$8360 ( \9046 , \9040 , \9045 );
xor \U$8361 ( \9047 , \8426 , \8459 );
and \U$8362 ( \9048 , \9047 , \8471 );
and \U$8363 ( \9049 , \8426 , \8459 );
or \U$8364 ( \9050 , \9048 , \9049 );
not \U$8365 ( \9051 , \9050 );
and \U$8366 ( \9052 , \8378 , \6034 );
not \U$8367 ( \9053 , \8378 );
and \U$8368 ( \9054 , \9053 , \7153 );
nor \U$8369 ( \9055 , \9052 , \9054 );
and \U$8370 ( \9056 , \6029 , \9055 );
not \U$8371 ( \9057 , \8466 );
not \U$8372 ( \9058 , \6265 );
or \U$8373 ( \9059 , \9057 , \9058 );
not \U$8374 ( \9060 , \8141 );
not \U$8375 ( \9061 , \6477 );
or \U$8376 ( \9062 , \9060 , \9061 );
nand \U$8377 ( \9063 , \6911 , \8142 );
nand \U$8378 ( \9064 , \9062 , \9063 );
nand \U$8379 ( \9065 , \9064 , \6919 );
nand \U$8380 ( \9066 , \9059 , \9065 );
xor \U$8381 ( \9067 , \9056 , \9066 );
nor \U$8382 ( \9068 , \8058 , \8042 );
buf \U$8383 ( \9069 , \8026 );
or \U$8384 ( \9070 , \9068 , \9069 );
nand \U$8385 ( \9071 , \8058 , \8042 );
nand \U$8386 ( \9072 , \9070 , \9071 );
xor \U$8387 ( \9073 , \9067 , \9072 );
not \U$8388 ( \9074 , \9073 );
not \U$8389 ( \9075 , \9074 );
or \U$8390 ( \9076 , \9051 , \9075 );
not \U$8391 ( \9077 , \9050 );
nand \U$8392 ( \9078 , \9073 , \9077 );
nand \U$8393 ( \9079 , \9076 , \9078 );
not \U$8394 ( \9080 , \8059 );
not \U$8395 ( \9081 , \9080 );
not \U$8396 ( \9082 , \8175 );
or \U$8397 ( \9083 , \9081 , \9082 );
not \U$8398 ( \9084 , \8059 );
not \U$8399 ( \9085 , \8174 );
or \U$8400 ( \9086 , \9084 , \9085 );
nand \U$8401 ( \9087 , \9086 , \8219 );
nand \U$8402 ( \9088 , \9083 , \9087 );
not \U$8403 ( \9089 , \9088 );
and \U$8404 ( \9090 , \9079 , \9089 );
not \U$8405 ( \9091 , \9079 );
and \U$8406 ( \9092 , \9091 , \9088 );
nor \U$8407 ( \9093 , \9090 , \9092 );
xor \U$8408 ( \9094 , \9046 , \9093 );
or \U$8409 ( \9095 , \8606 , \8220 );
and \U$8410 ( \9096 , \9095 , \8617 );
and \U$8411 ( \9097 , \8220 , \8606 );
nor \U$8412 ( \9098 , \9096 , \9097 );
nand \U$8413 ( \9099 , \9094 , \9098 );
nand \U$8414 ( \9100 , \9017 , \9011 );
not \U$8415 ( \9101 , \8986 );
not \U$8416 ( \9102 , \7018 );
or \U$8417 ( \9103 , \9101 , \9102 );
nand \U$8418 ( \9104 , \7911 , \7012 );
nand \U$8419 ( \9105 , \9103 , \9104 );
xor \U$8420 ( \9106 , \9100 , \9105 );
not \U$8421 ( \9107 , \8997 );
not \U$8422 ( \9108 , \6978 );
or \U$8423 ( \9109 , \9107 , \9108 );
nand \U$8424 ( \9110 , \7922 , \6981 );
nand \U$8425 ( \9111 , \9109 , \9110 );
xnor \U$8426 ( \9112 , \9106 , \9111 );
xor \U$8427 ( \9113 , \9018 , \9029 );
and \U$8428 ( \9114 , \9113 , \9038 );
and \U$8429 ( \9115 , \9018 , \9029 );
or \U$8430 ( \9116 , \9114 , \9115 );
xor \U$8431 ( \9117 , \9112 , \9116 );
xor \U$8432 ( \9118 , \7905 , \7892 );
not \U$8433 ( \9119 , \9027 );
not \U$8434 ( \9120 , \7089 );
or \U$8435 ( \9121 , \9119 , \9120 );
nand \U$8436 ( \9122 , \7954 , \6545 );
nand \U$8437 ( \9123 , \9121 , \9122 );
xor \U$8438 ( \9124 , \9118 , \9123 );
not \U$8439 ( \9125 , \9036 );
not \U$8440 ( \9126 , \9125 );
not \U$8441 ( \9127 , \7034 );
or \U$8442 ( \9128 , \9126 , \9127 );
nand \U$8443 ( \9129 , \6383 , \7965 );
nand \U$8444 ( \9130 , \9128 , \9129 );
xor \U$8445 ( \9131 , \9124 , \9130 );
xnor \U$8446 ( \9132 , \9117 , \9131 );
not \U$8447 ( \9133 , \9077 );
not \U$8448 ( \9134 , \9074 );
or \U$8449 ( \9135 , \9133 , \9134 );
nand \U$8450 ( \9136 , \9135 , \9088 );
nand \U$8451 ( \9137 , \9073 , \9050 );
nand \U$8452 ( \9138 , \9136 , \9137 );
not \U$8453 ( \9139 , \9138 );
xor \U$8454 ( \9140 , \9132 , \9139 );
and \U$8455 ( \9141 , \8102 , \7153 );
not \U$8456 ( \9142 , \8102 );
and \U$8457 ( \9143 , \9142 , \6034 );
nor \U$8458 ( \9144 , \9141 , \9143 );
and \U$8459 ( \9145 , \6029 , \9144 );
not \U$8460 ( \9146 , \9064 );
not \U$8461 ( \9147 , \6265 );
or \U$8462 ( \9148 , \9146 , \9147 );
not \U$8463 ( \9149 , \8152 );
not \U$8464 ( \9150 , \6270 );
or \U$8465 ( \9151 , \9149 , \9150 );
nand \U$8466 ( \9152 , \8786 , \7875 );
nand \U$8467 ( \9153 , \9151 , \9152 );
nand \U$8468 ( \9154 , \9153 , \6919 );
nand \U$8469 ( \9155 , \9148 , \9154 );
xor \U$8470 ( \9156 , \9145 , \9155 );
xor \U$8471 ( \9157 , \8978 , \8988 );
and \U$8472 ( \9158 , \9157 , \8999 );
and \U$8473 ( \9159 , \8978 , \8988 );
or \U$8474 ( \9160 , \9158 , \9159 );
xor \U$8475 ( \9161 , \9156 , \9160 );
xor \U$8476 ( \9162 , \9056 , \9066 );
and \U$8477 ( \9163 , \9162 , \9072 );
and \U$8478 ( \9164 , \9056 , \9066 );
or \U$8479 ( \9165 , \9163 , \9164 );
and \U$8480 ( \9166 , \9161 , \9165 );
not \U$8481 ( \9167 , \9161 );
not \U$8482 ( \9168 , \9165 );
and \U$8483 ( \9169 , \9167 , \9168 );
nor \U$8484 ( \9170 , \9166 , \9169 );
not \U$8485 ( \9171 , \9000 );
nand \U$8486 ( \9172 , \9171 , \9004 );
not \U$8487 ( \9173 , \9172 );
not \U$8488 ( \9174 , \9039 );
or \U$8489 ( \9175 , \9173 , \9174 );
nand \U$8490 ( \9176 , \9005 , \9000 );
nand \U$8491 ( \9177 , \9175 , \9176 );
not \U$8492 ( \9178 , \9177 );
and \U$8493 ( \9179 , \9170 , \9178 );
not \U$8494 ( \9180 , \9170 );
and \U$8495 ( \9181 , \9180 , \9177 );
nor \U$8496 ( \9182 , \9179 , \9181 );
xor \U$8497 ( \9183 , \9140 , \9182 );
xor \U$8498 ( \9184 , \9040 , \9045 );
and \U$8499 ( \9185 , \9184 , \9093 );
and \U$8500 ( \9186 , \9040 , \9045 );
or \U$8501 ( \9187 , \9185 , \9186 );
nand \U$8502 ( \9188 , \9183 , \9187 );
nand \U$8503 ( \9189 , \9099 , \9188 );
nor \U$8504 ( \9190 , \8977 , \9189 );
not \U$8505 ( \9191 , \9190 );
nor \U$8506 ( \9192 , \9098 , \9094 );
not \U$8507 ( \9193 , \9192 );
not \U$8508 ( \9194 , \9188 );
or \U$8509 ( \9195 , \9193 , \9194 );
or \U$8510 ( \9196 , \9183 , \9187 );
nand \U$8511 ( \9197 , \9195 , \9196 );
not \U$8512 ( \9198 , \9197 );
nand \U$8513 ( \9199 , \9191 , \9198 );
xor \U$8514 ( \9200 , \7942 , \7973 );
xnor \U$8515 ( \9201 , \9200 , \7978 );
xor \U$8516 ( \9202 , \7906 , \7916 );
xor \U$8517 ( \9203 , \9202 , \7927 );
xor \U$8518 ( \9204 , \9118 , \9123 );
and \U$8519 ( \9205 , \9204 , \9130 );
and \U$8520 ( \9206 , \9118 , \9123 );
or \U$8521 ( \9207 , \9205 , \9206 );
or \U$8522 ( \9208 , \9203 , \9207 );
xor \U$8523 ( \9209 , \7949 , \7959 );
xor \U$8524 ( \9210 , \9209 , \7970 );
nand \U$8525 ( \9211 , \9208 , \9210 );
nand \U$8526 ( \9212 , \9207 , \9203 );
nand \U$8527 ( \9213 , \9211 , \9212 );
not \U$8528 ( \9214 , \9213 );
xor \U$8529 ( \9215 , \7880 , \7830 );
xnor \U$8530 ( \9216 , \9215 , \7930 );
not \U$8531 ( \9217 , \9216 );
and \U$8532 ( \9218 , \8141 , \6032 );
not \U$8533 ( \9219 , \8141 );
and \U$8534 ( \9220 , \9219 , \6033 );
nor \U$8535 ( \9221 , \9218 , \9220 );
and \U$8536 ( \9222 , \6028 , \9221 );
not \U$8537 ( \9223 , \9153 );
not \U$8538 ( \9224 , \7826 );
or \U$8539 ( \9225 , \9223 , \9224 );
nand \U$8540 ( \9226 , \7824 , \6253 );
nand \U$8541 ( \9227 , \9225 , \9226 );
xor \U$8542 ( \9228 , \9222 , \9227 );
nor \U$8543 ( \9229 , \9111 , \9105 );
or \U$8544 ( \9230 , \9229 , \9100 );
nand \U$8545 ( \9231 , \9111 , \9105 );
nand \U$8546 ( \9232 , \9230 , \9231 );
and \U$8547 ( \9233 , \9228 , \9232 );
and \U$8548 ( \9234 , \9222 , \9227 );
or \U$8549 ( \9235 , \9233 , \9234 );
not \U$8550 ( \9236 , \9235 );
not \U$8551 ( \9237 , \9236 );
and \U$8552 ( \9238 , \9217 , \9237 );
and \U$8553 ( \9239 , \9216 , \9236 );
nor \U$8554 ( \9240 , \9238 , \9239 );
not \U$8555 ( \9241 , \9240 );
or \U$8556 ( \9242 , \9214 , \9241 );
not \U$8557 ( \9243 , \9213 );
not \U$8558 ( \9244 , \9240 );
nand \U$8559 ( \9245 , \9243 , \9244 );
nand \U$8560 ( \9246 , \9242 , \9245 );
xor \U$8561 ( \9247 , \9201 , \9246 );
xor \U$8562 ( \9248 , \9145 , \9155 );
and \U$8563 ( \9249 , \9248 , \9160 );
and \U$8564 ( \9250 , \9145 , \9155 );
or \U$8565 ( \9251 , \9249 , \9250 );
not \U$8566 ( \9252 , \9251 );
xor \U$8567 ( \9253 , \9222 , \9227 );
xor \U$8568 ( \9254 , \9253 , \9232 );
not \U$8569 ( \9255 , \9254 );
or \U$8570 ( \9256 , \9252 , \9255 );
not \U$8571 ( \9257 , \9112 );
not \U$8572 ( \9258 , \9257 );
not \U$8573 ( \9259 , \9116 );
not \U$8574 ( \9260 , \9259 );
or \U$8575 ( \9261 , \9258 , \9260 );
nand \U$8576 ( \9262 , \9261 , \9131 );
nand \U$8577 ( \9263 , \9116 , \9112 );
nand \U$8578 ( \9264 , \9262 , \9263 );
not \U$8579 ( \9265 , \9254 );
not \U$8580 ( \9266 , \9251 );
nand \U$8581 ( \9267 , \9265 , \9266 );
nand \U$8582 ( \9268 , \9264 , \9267 );
nand \U$8583 ( \9269 , \9256 , \9268 );
xor \U$8584 ( \9270 , \9247 , \9269 );
buf \U$8585 ( \9271 , \9207 );
xor \U$8586 ( \9272 , \9203 , \9271 );
xnor \U$8587 ( \9273 , \9272 , \9210 );
not \U$8588 ( \9274 , \9161 );
not \U$8589 ( \9275 , \9274 );
not \U$8590 ( \9276 , \9168 );
or \U$8591 ( \9277 , \9275 , \9276 );
nand \U$8592 ( \9278 , \9277 , \9177 );
not \U$8593 ( \9279 , \9274 );
nand \U$8594 ( \9280 , \9279 , \9165 );
and \U$8595 ( \9281 , \9278 , \9280 );
xor \U$8596 ( \9282 , \9273 , \9281 );
not \U$8597 ( \9283 , \9251 );
not \U$8598 ( \9284 , \9265 );
or \U$8599 ( \9285 , \9283 , \9284 );
nand \U$8600 ( \9286 , \9254 , \9266 );
nand \U$8601 ( \9287 , \9285 , \9286 );
not \U$8602 ( \9288 , \9264 );
and \U$8603 ( \9289 , \9287 , \9288 );
not \U$8604 ( \9290 , \9287 );
and \U$8605 ( \9291 , \9290 , \9264 );
nor \U$8606 ( \9292 , \9289 , \9291 );
and \U$8607 ( \9293 , \9282 , \9292 );
and \U$8608 ( \9294 , \9273 , \9281 );
or \U$8609 ( \9295 , \9293 , \9294 );
nand \U$8610 ( \9296 , \9270 , \9295 );
xor \U$8611 ( \9297 , \7756 , \7791 );
xnor \U$8612 ( \9298 , \9297 , \7787 );
not \U$8613 ( \9299 , \9216 );
nand \U$8614 ( \9300 , \9299 , \9236 );
and \U$8615 ( \9301 , \9213 , \9300 );
nor \U$8616 ( \9302 , \9299 , \9236 );
nor \U$8617 ( \9303 , \9301 , \9302 );
xor \U$8618 ( \9304 , \9298 , \9303 );
not \U$8619 ( \9305 , \7983 );
not \U$8620 ( \9306 , \7938 );
or \U$8621 ( \9307 , \9305 , \9306 );
nand \U$8622 ( \9308 , \7982 , \7935 );
nand \U$8623 ( \9309 , \9307 , \9308 );
not \U$8624 ( \9310 , \7980 );
and \U$8625 ( \9311 , \9309 , \9310 );
not \U$8626 ( \9312 , \9309 );
and \U$8627 ( \9313 , \9312 , \7980 );
nor \U$8628 ( \9314 , \9311 , \9313 );
xor \U$8629 ( \9315 , \9304 , \9314 );
not \U$8630 ( \9316 , \9246 );
nand \U$8631 ( \9317 , \9316 , \9201 );
and \U$8632 ( \9318 , \9317 , \9269 );
nor \U$8633 ( \9319 , \9316 , \9201 );
nor \U$8634 ( \9320 , \9318 , \9319 );
nand \U$8635 ( \9321 , \9315 , \9320 );
xor \U$8636 ( \9322 , \9273 , \9281 );
xor \U$8637 ( \9323 , \9322 , \9292 );
xor \U$8638 ( \9324 , \9132 , \9139 );
and \U$8639 ( \9325 , \9324 , \9182 );
and \U$8640 ( \9326 , \9132 , \9139 );
or \U$8641 ( \9327 , \9325 , \9326 );
nand \U$8642 ( \9328 , \9323 , \9327 );
not \U$8643 ( \9329 , \7985 );
xor \U$8644 ( \9330 , \7817 , \9329 );
xnor \U$8645 ( \9331 , \9330 , \7815 );
xor \U$8646 ( \9332 , \9298 , \9303 );
and \U$8647 ( \9333 , \9332 , \9314 );
and \U$8648 ( \9334 , \9298 , \9303 );
or \U$8649 ( \9335 , \9333 , \9334 );
nand \U$8650 ( \9336 , \9331 , \9335 );
nand \U$8651 ( \9337 , \9296 , \9321 , \9328 , \9336 );
not \U$8652 ( \9338 , \9337 );
nand \U$8653 ( \9339 , \9199 , \9338 );
xor \U$8654 ( \9340 , \8785 , \8792 );
xor \U$8655 ( \9341 , \9340 , \8804 );
xor \U$8656 ( \9342 , \8814 , \8824 );
xor \U$8657 ( \9343 , \9342 , \8835 );
xor \U$8658 ( \9344 , \9341 , \9343 );
not \U$8659 ( \9345 , \8890 );
and \U$8660 ( \9346 , \8902 , \8887 );
not \U$8661 ( \9347 , \8902 );
and \U$8662 ( \9348 , \9347 , \8888 );
nor \U$8663 ( \9349 , \9346 , \9348 );
not \U$8664 ( \9350 , \9349 );
or \U$8665 ( \9351 , \9345 , \9350 );
or \U$8666 ( \9352 , \8890 , \9349 );
nand \U$8667 ( \9353 , \9351 , \9352 );
and \U$8668 ( \9354 , \8310 , \6547 );
not \U$8669 ( \9355 , \8310 );
and \U$8670 ( \9356 , \9355 , \6497 );
or \U$8671 ( \9357 , \9354 , \9356 );
not \U$8672 ( \9358 , \9357 );
not \U$8673 ( \9359 , \6542 );
or \U$8674 ( \9360 , \9358 , \9359 );
nand \U$8675 ( \9361 , \8820 , \7163 );
nand \U$8676 ( \9362 , \9360 , \9361 );
xor \U$8677 ( \9363 , \9353 , \9362 );
not \U$8678 ( \9364 , \8563 );
not \U$8679 ( \9365 , \6651 );
or \U$8680 ( \9366 , \9364 , \9365 );
nand \U$8681 ( \9367 , \6652 , \8749 );
nand \U$8682 ( \9368 , \9366 , \9367 );
not \U$8683 ( \9369 , \9368 );
not \U$8684 ( \9370 , \6398 );
or \U$8685 ( \9371 , \9369 , \9370 );
nand \U$8686 ( \9372 , \6384 , \8830 );
nand \U$8687 ( \9373 , \9371 , \9372 );
and \U$8688 ( \9374 , \9363 , \9373 );
and \U$8689 ( \9375 , \9353 , \9362 );
or \U$8690 ( \9376 , \9374 , \9375 );
and \U$8691 ( \9377 , \9344 , \9376 );
and \U$8692 ( \9378 , \9341 , \9343 );
or \U$8693 ( \9379 , \9377 , \9378 );
not \U$8694 ( \9380 , \9379 );
not \U$8695 ( \9381 , \8807 );
not \U$8696 ( \9382 , \8811 );
and \U$8697 ( \9383 , \9381 , \9382 );
and \U$8698 ( \9384 , \8807 , \8811 );
nor \U$8699 ( \9385 , \9383 , \9384 );
xor \U$8700 ( \9386 , \9385 , \8838 );
not \U$8701 ( \9387 , \9386 );
and \U$8702 ( \9388 , \9380 , \9387 );
and \U$8703 ( \9389 , \9379 , \9386 );
nor \U$8704 ( \9390 , \9388 , \9389 );
not \U$8705 ( \9391 , \9390 );
xor \U$8706 ( \9392 , \8871 , \8875 );
xor \U$8707 ( \9393 , \9392 , \8966 );
not \U$8708 ( \9394 , \9393 );
not \U$8709 ( \9395 , \9394 );
and \U$8710 ( \9396 , \9391 , \9395 );
and \U$8711 ( \9397 , \9394 , \9390 );
nor \U$8712 ( \9398 , \9396 , \9397 );
xor \U$8713 ( \9399 , \8906 , \8952 );
xor \U$8714 ( \9400 , \9399 , \8963 );
not \U$8715 ( \9401 , \8141 );
not \U$8716 ( \9402 , \7700 );
or \U$8717 ( \9403 , \9401 , \9402 );
nand \U$8718 ( \9404 , \8030 , \8142 );
nand \U$8719 ( \9405 , \9403 , \9404 );
not \U$8720 ( \9406 , \9405 );
not \U$8721 ( \9407 , \7018 );
or \U$8722 ( \9408 , \9406 , \9407 );
nand \U$8723 ( \9409 , \8911 , \7012 );
nand \U$8724 ( \9410 , \9408 , \9409 );
or \U$8725 ( \9411 , \7084 , \6392 );
and \U$8726 ( \9412 , \9411 , \8692 );
not \U$8727 ( \9413 , \6392 );
not \U$8728 ( \9414 , \7084 );
or \U$8729 ( \9415 , \9413 , \9414 );
nand \U$8730 ( \9416 , \9415 , \6402 );
nor \U$8731 ( \9417 , \9412 , \9416 );
xor \U$8732 ( \9418 , \9410 , \9417 );
not \U$8733 ( \9419 , \8374 );
not \U$8734 ( \9420 , \6803 );
or \U$8735 ( \9421 , \9419 , \9420 );
not \U$8736 ( \9422 , \7373 );
not \U$8737 ( \9423 , \8374 );
nand \U$8738 ( \9424 , \9422 , \9423 );
nand \U$8739 ( \9425 , \9421 , \9424 );
not \U$8740 ( \9426 , \9425 );
not \U$8741 ( \9427 , \7379 );
or \U$8742 ( \9428 , \9426 , \9427 );
nand \U$8743 ( \9429 , \8944 , \6981 );
nand \U$8744 ( \9430 , \9428 , \9429 );
and \U$8745 ( \9431 , \9418 , \9430 );
and \U$8746 ( \9432 , \9410 , \9417 );
or \U$8747 ( \9433 , \9431 , \9432 );
xor \U$8748 ( \9434 , \8916 , \8938 );
xor \U$8749 ( \9435 , \9434 , \8949 );
xor \U$8750 ( \9436 , \9433 , \9435 );
xor \U$8751 ( \9437 , \8937 , \8927 );
not \U$8752 ( \9438 , \8272 );
not \U$8753 ( \9439 , \6548 );
or \U$8754 ( \9440 , \9438 , \9439 );
not \U$8755 ( \9441 , \6497 );
nand \U$8756 ( \9442 , \9441 , \8271 );
nand \U$8757 ( \9443 , \9440 , \9442 );
not \U$8758 ( \9444 , \9443 );
not \U$8759 ( \9445 , \6542 );
or \U$8760 ( \9446 , \9444 , \9445 );
nand \U$8761 ( \9447 , \9357 , \6546 );
nand \U$8762 ( \9448 , \9446 , \9447 );
xor \U$8763 ( \9449 , \9437 , \9448 );
not \U$8764 ( \9450 , \8692 );
not \U$8765 ( \9451 , \6403 );
or \U$8766 ( \9452 , \9450 , \9451 );
nand \U$8767 ( \9453 , \6402 , \8954 );
nand \U$8768 ( \9454 , \9452 , \9453 );
not \U$8769 ( \9455 , \9454 );
not \U$8770 ( \9456 , \6397 );
or \U$8771 ( \9457 , \9455 , \9456 );
nand \U$8772 ( \9458 , \6384 , \9368 );
nand \U$8773 ( \9459 , \9457 , \9458 );
and \U$8774 ( \9460 , \9449 , \9459 );
and \U$8775 ( \9461 , \9437 , \9448 );
or \U$8776 ( \9462 , \9460 , \9461 );
and \U$8777 ( \9463 , \9436 , \9462 );
and \U$8778 ( \9464 , \9433 , \9435 );
or \U$8779 ( \9465 , \9463 , \9464 );
xor \U$8780 ( \9466 , \9400 , \9465 );
xor \U$8781 ( \9467 , \9341 , \9343 );
xor \U$8782 ( \9468 , \9467 , \9376 );
and \U$8783 ( \9469 , \9466 , \9468 );
and \U$8784 ( \9470 , \9400 , \9465 );
or \U$8785 ( \9471 , \9469 , \9470 );
not \U$8786 ( \9472 , \9471 );
nand \U$8787 ( \9473 , \9398 , \9472 );
not \U$8788 ( \9474 , \9473 );
xor \U$8789 ( \9475 , \9400 , \9465 );
xor \U$8790 ( \9476 , \9475 , \9468 );
xor \U$8791 ( \9477 , \9433 , \9435 );
xor \U$8792 ( \9478 , \9477 , \9462 );
not \U$8793 ( \9479 , \9478 );
not \U$8794 ( \9480 , \7729 );
and \U$8795 ( \9481 , \7607 , \7488 );
not \U$8796 ( \9482 , \7607 );
and \U$8797 ( \9483 , \9482 , \7619 );
nor \U$8798 ( \9484 , \9481 , \9483 );
not \U$8799 ( \9485 , \9484 );
or \U$8800 ( \9486 , \9480 , \9485 );
nand \U$8801 ( \9487 , \8933 , \7903 );
nand \U$8802 ( \9488 , \9486 , \9487 );
not \U$8803 ( \9489 , \8917 );
not \U$8804 ( \9490 , \8152 );
or \U$8805 ( \9491 , \9489 , \9490 );
nand \U$8806 ( \9492 , \7714 , \7875 );
nand \U$8807 ( \9493 , \9491 , \9492 );
not \U$8808 ( \9494 , \9493 );
not \U$8809 ( \9495 , \7601 );
or \U$8810 ( \9496 , \9494 , \9495 );
nand \U$8811 ( \9497 , \8922 , \7890 );
nand \U$8812 ( \9498 , \9496 , \9497 );
xor \U$8813 ( \9499 , \9488 , \9498 );
and \U$8814 ( \9500 , \6383 , \8692 );
and \U$8815 ( \9501 , \9499 , \9500 );
and \U$8816 ( \9502 , \9488 , \9498 );
or \U$8817 ( \9503 , \9501 , \9502 );
xor \U$8818 ( \9504 , \9410 , \9417 );
xor \U$8819 ( \9505 , \9504 , \9430 );
xor \U$8820 ( \9506 , \9503 , \9505 );
not \U$8821 ( \9507 , \8141 );
not \U$8822 ( \9508 , \7358 );
or \U$8823 ( \9509 , \9507 , \9508 );
nand \U$8824 ( \9510 , \7714 , \8142 );
nand \U$8825 ( \9511 , \9509 , \9510 );
not \U$8826 ( \9512 , \9511 );
not \U$8827 ( \9513 , \7601 );
or \U$8828 ( \9514 , \9512 , \9513 );
nand \U$8829 ( \9515 , \9493 , \7604 );
nand \U$8830 ( \9516 , \9514 , \9515 );
not \U$8831 ( \9517 , \7903 );
not \U$8832 ( \9518 , \9484 );
or \U$8833 ( \9519 , \9517 , \9518 );
not \U$8834 ( \9520 , \7607 );
not \U$8835 ( \9521 , \7676 );
or \U$8836 ( \9522 , \9520 , \9521 );
nand \U$8837 ( \9523 , \7675 , \7608 );
nand \U$8838 ( \9524 , \9522 , \9523 );
nand \U$8839 ( \9525 , \9524 , \7729 );
nand \U$8840 ( \9526 , \9519 , \9525 );
and \U$8841 ( \9527 , \9516 , \9526 );
not \U$8842 ( \9528 , \8102 );
not \U$8843 ( \9529 , \7698 );
or \U$8844 ( \9530 , \9528 , \9529 );
nand \U$8845 ( \9531 , \7699 , \8101 );
nand \U$8846 ( \9532 , \9530 , \9531 );
not \U$8847 ( \9533 , \9532 );
not \U$8848 ( \9534 , \7018 );
or \U$8849 ( \9535 , \9533 , \9534 );
nand \U$8850 ( \9536 , \9405 , \7012 );
nand \U$8851 ( \9537 , \9535 , \9536 );
xor \U$8852 ( \9538 , \9527 , \9537 );
not \U$8853 ( \9539 , \7379 );
and \U$8854 ( \9540 , \7373 , \8310 );
not \U$8855 ( \9541 , \7373 );
and \U$8856 ( \9542 , \9541 , \8309 );
or \U$8857 ( \9543 , \9540 , \9542 );
not \U$8858 ( \9544 , \9543 );
or \U$8859 ( \9545 , \9539 , \9544 );
not \U$8860 ( \9546 , \9425 );
or \U$8861 ( \9547 , \9546 , \6692 );
nand \U$8862 ( \9548 , \9545 , \9547 );
and \U$8863 ( \9549 , \9538 , \9548 );
and \U$8864 ( \9550 , \9527 , \9537 );
or \U$8865 ( \9551 , \9549 , \9550 );
and \U$8866 ( \9552 , \9506 , \9551 );
and \U$8867 ( \9553 , \9503 , \9505 );
or \U$8868 ( \9554 , \9552 , \9553 );
not \U$8869 ( \9555 , \9554 );
xor \U$8870 ( \9556 , \9353 , \9362 );
xor \U$8871 ( \9557 , \9556 , \9373 );
not \U$8872 ( \9558 , \9557 );
nand \U$8873 ( \9559 , \9555 , \9558 );
not \U$8874 ( \9560 , \9559 );
or \U$8875 ( \9561 , \9479 , \9560 );
nand \U$8876 ( \9562 , \9554 , \9557 );
nand \U$8877 ( \9563 , \9561 , \9562 );
or \U$8878 ( \9564 , \9476 , \9563 );
and \U$8879 ( \9565 , \9554 , \9557 );
not \U$8880 ( \9566 , \9554 );
and \U$8881 ( \9567 , \9566 , \9558 );
nor \U$8882 ( \9568 , \9565 , \9567 );
and \U$8883 ( \9569 , \9568 , \9478 );
not \U$8884 ( \9570 , \9568 );
not \U$8885 ( \9571 , \9478 );
and \U$8886 ( \9572 , \9570 , \9571 );
nor \U$8887 ( \9573 , \9569 , \9572 );
xor \U$8888 ( \9574 , \9437 , \9448 );
xor \U$8889 ( \9575 , \9574 , \9459 );
not \U$8890 ( \9576 , \8563 );
not \U$8891 ( \9577 , \6706 );
or \U$8892 ( \9578 , \9576 , \9577 );
nand \U$8893 ( \9579 , \9025 , \8749 );
nand \U$8894 ( \9580 , \9578 , \9579 );
not \U$8895 ( \9581 , \9580 );
not \U$8896 ( \9582 , \6542 );
or \U$8897 ( \9583 , \9581 , \9582 );
nand \U$8898 ( \9584 , \9443 , \6546 );
nand \U$8899 ( \9585 , \9583 , \9584 );
not \U$8900 ( \9586 , \7093 );
not \U$8901 ( \9587 , \6531 );
not \U$8902 ( \9588 , \7373 );
or \U$8903 ( \9589 , \9587 , \9588 );
nand \U$8904 ( \9590 , \9589 , \8692 );
nand \U$8905 ( \9591 , \8797 , \6513 );
nand \U$8906 ( \9592 , \9586 , \9590 , \9591 );
not \U$8907 ( \9593 , \9592 );
not \U$8908 ( \9594 , \8374 );
not \U$8909 ( \9595 , \7698 );
or \U$8910 ( \9596 , \9594 , \9595 );
nand \U$8911 ( \9597 , \7699 , \8378 );
nand \U$8912 ( \9598 , \9596 , \9597 );
not \U$8913 ( \9599 , \9598 );
not \U$8914 ( \9600 , \7018 );
or \U$8915 ( \9601 , \9599 , \9600 );
nand \U$8916 ( \9602 , \9532 , \7012 );
nand \U$8917 ( \9603 , \9601 , \9602 );
not \U$8918 ( \9604 , \9603 );
not \U$8919 ( \9605 , \9604 );
or \U$8920 ( \9606 , \9593 , \9605 );
xor \U$8921 ( \9607 , \9526 , \9516 );
nand \U$8922 ( \9608 , \9606 , \9607 );
not \U$8923 ( \9609 , \9592 );
nand \U$8924 ( \9610 , \9609 , \9603 );
nand \U$8925 ( \9611 , \9608 , \9610 );
xor \U$8926 ( \9612 , \9585 , \9611 );
xor \U$8927 ( \9613 , \9488 , \9498 );
xor \U$8928 ( \9614 , \9613 , \9500 );
and \U$8929 ( \9615 , \9612 , \9614 );
and \U$8930 ( \9616 , \9585 , \9611 );
or \U$8931 ( \9617 , \9615 , \9616 );
xor \U$8932 ( \9618 , \9575 , \9617 );
xor \U$8933 ( \9619 , \9503 , \9505 );
xor \U$8934 ( \9620 , \9619 , \9551 );
and \U$8935 ( \9621 , \9618 , \9620 );
and \U$8936 ( \9622 , \9575 , \9617 );
or \U$8937 ( \9623 , \9621 , \9622 );
nand \U$8938 ( \9624 , \9573 , \9623 );
nand \U$8939 ( \9625 , \9476 , \9563 );
nand \U$8940 ( \9626 , \9624 , \9625 );
nand \U$8941 ( \9627 , \9564 , \9626 );
nor \U$8942 ( \9628 , \9474 , \9627 );
not \U$8943 ( \9629 , \9398 );
nand \U$8944 ( \9630 , \9629 , \9471 );
xor \U$8945 ( \9631 , \8869 , \8968 );
xor \U$8946 ( \9632 , \9631 , \8971 );
not \U$8947 ( \9633 , \9386 );
not \U$8948 ( \9634 , \9633 );
not \U$8949 ( \9635 , \9394 );
or \U$8950 ( \9636 , \9634 , \9635 );
not \U$8951 ( \9637 , \9386 );
not \U$8952 ( \9638 , \9393 );
or \U$8953 ( \9639 , \9637 , \9638 );
nand \U$8954 ( \9640 , \9639 , \9379 );
nand \U$8955 ( \9641 , \9636 , \9640 );
nand \U$8956 ( \9642 , \9632 , \9641 );
nand \U$8957 ( \9643 , \9630 , \9642 );
or \U$8958 ( \9644 , \9628 , \9643 );
or \U$8959 ( \9645 , \9632 , \9641 );
nand \U$8960 ( \9646 , \9644 , \9645 );
xor \U$8961 ( \9647 , \9575 , \9617 );
xor \U$8962 ( \9648 , \9647 , \9620 );
xor \U$8963 ( \9649 , \9527 , \9537 );
xor \U$8964 ( \9650 , \9649 , \9548 );
not \U$8965 ( \9651 , \8271 );
not \U$8966 ( \9652 , \6803 );
or \U$8967 ( \9653 , \9651 , \9652 );
nand \U$8968 ( \9654 , \9422 , \8272 );
nand \U$8969 ( \9655 , \9653 , \9654 );
not \U$8970 ( \9656 , \9655 );
not \U$8971 ( \9657 , \7379 );
or \U$8972 ( \9658 , \9656 , \9657 );
nand \U$8973 ( \9659 , \9543 , \6981 );
nand \U$8974 ( \9660 , \9658 , \9659 );
not \U$8975 ( \9661 , \9660 );
not \U$8976 ( \9662 , \9661 );
and \U$8977 ( \9663 , \8954 , \6498 );
not \U$8978 ( \9664 , \8954 );
and \U$8979 ( \9665 , \9664 , \6548 );
nor \U$8980 ( \9666 , \9663 , \9665 );
not \U$8981 ( \9667 , \9666 );
not \U$8982 ( \9668 , \6542 );
or \U$8983 ( \9669 , \9667 , \9668 );
nand \U$8984 ( \9670 , \9580 , \6546 );
nand \U$8985 ( \9671 , \9669 , \9670 );
not \U$8986 ( \9672 , \9671 );
not \U$8987 ( \9673 , \9672 );
or \U$8988 ( \9674 , \9662 , \9673 );
not \U$8989 ( \9675 , \7737 );
not \U$8990 ( \9676 , \9524 );
or \U$8991 ( \9677 , \9675 , \9676 );
not \U$8992 ( \9678 , \7607 );
not \U$8993 ( \9679 , \7874 );
or \U$8994 ( \9680 , \9678 , \9679 );
nand \U$8995 ( \9681 , \7873 , \7608 );
nand \U$8996 ( \9682 , \9680 , \9681 );
nand \U$8997 ( \9683 , \9682 , \7729 );
nand \U$8998 ( \9684 , \9677 , \9683 );
not \U$8999 ( \9685 , \8102 );
not \U$9000 ( \9686 , \7358 );
or \U$9001 ( \9687 , \9685 , \9686 );
nand \U$9002 ( \9688 , \8920 , \8101 );
nand \U$9003 ( \9689 , \9687 , \9688 );
not \U$9004 ( \9690 , \9689 );
not \U$9005 ( \9691 , \7601 );
or \U$9006 ( \9692 , \9690 , \9691 );
nand \U$9007 ( \9693 , \9511 , \7604 );
nand \U$9008 ( \9694 , \9692 , \9693 );
xor \U$9009 ( \9695 , \9684 , \9694 );
nor \U$9010 ( \9696 , \7162 , \8954 );
and \U$9011 ( \9697 , \9695 , \9696 );
and \U$9012 ( \9698 , \9684 , \9694 );
or \U$9013 ( \9699 , \9697 , \9698 );
nand \U$9014 ( \9700 , \9674 , \9699 );
nand \U$9015 ( \9701 , \9671 , \9660 );
nand \U$9016 ( \9702 , \9700 , \9701 );
xor \U$9017 ( \9703 , \9650 , \9702 );
xor \U$9018 ( \9704 , \9585 , \9611 );
xor \U$9019 ( \9705 , \9704 , \9614 );
and \U$9020 ( \9706 , \9703 , \9705 );
and \U$9021 ( \9707 , \9650 , \9702 );
or \U$9022 ( \9708 , \9706 , \9707 );
nor \U$9023 ( \9709 , \9648 , \9708 );
not \U$9024 ( \9710 , \9709 );
not \U$9025 ( \9711 , \8310 );
not \U$9026 ( \9712 , \7170 );
or \U$9027 ( \9713 , \9711 , \9712 );
not \U$9028 ( \9714 , \7700 );
nand \U$9029 ( \9715 , \9714 , \8309 );
nand \U$9030 ( \9716 , \9713 , \9715 );
not \U$9031 ( \9717 , \9716 );
not \U$9032 ( \9718 , \7018 );
or \U$9033 ( \9719 , \9717 , \9718 );
nand \U$9034 ( \9720 , \9598 , \7012 );
nand \U$9035 ( \9721 , \9719 , \9720 );
not \U$9036 ( \9722 , \6695 );
not \U$9037 ( \9723 , \7698 );
or \U$9038 ( \9724 , \9722 , \9723 );
nand \U$9039 ( \9725 , \9724 , \8691 );
nand \U$9040 ( \9726 , \7020 , \6698 );
and \U$9041 ( \9727 , \6527 , \9725 , \9726 );
not \U$9042 ( \9728 , \7729 );
not \U$9043 ( \9729 , \7607 );
not \U$9044 ( \9730 , \8140 );
not \U$9045 ( \9731 , \9730 );
or \U$9046 ( \9732 , \9729 , \9731 );
nand \U$9047 ( \9733 , \7608 , \8140 );
nand \U$9048 ( \9734 , \9732 , \9733 );
not \U$9049 ( \9735 , \9734 );
or \U$9050 ( \9736 , \9728 , \9735 );
nand \U$9051 ( \9737 , \9682 , \7737 );
nand \U$9052 ( \9738 , \9736 , \9737 );
nand \U$9053 ( \9739 , \9727 , \9738 );
xor \U$9054 ( \9740 , \9721 , \9739 );
not \U$9055 ( \9741 , \8563 );
not \U$9056 ( \9742 , \7373 );
or \U$9057 ( \9743 , \9741 , \9742 );
nand \U$9058 ( \9744 , \8797 , \8749 );
nand \U$9059 ( \9745 , \9743 , \9744 );
not \U$9060 ( \9746 , \9745 );
not \U$9061 ( \9747 , \7379 );
or \U$9062 ( \9748 , \9746 , \9747 );
nand \U$9063 ( \9749 , \9655 , \6981 );
nand \U$9064 ( \9750 , \9748 , \9749 );
xor \U$9065 ( \9751 , \9740 , \9750 );
not \U$9066 ( \9752 , \9751 );
not \U$9067 ( \9753 , \9752 );
xor \U$9068 ( \9754 , \9684 , \9694 );
xor \U$9069 ( \9755 , \9754 , \9696 );
not \U$9070 ( \9756 , \9755 );
or \U$9071 ( \9757 , \9753 , \9756 );
not \U$9072 ( \9758 , \9755 );
not \U$9073 ( \9759 , \9758 );
not \U$9074 ( \9760 , \9751 );
or \U$9075 ( \9761 , \9759 , \9760 );
not \U$9076 ( \9762 , \9738 );
and \U$9077 ( \9763 , \9727 , \9762 );
not \U$9078 ( \9764 , \9727 );
and \U$9079 ( \9765 , \9764 , \9738 );
nor \U$9080 ( \9766 , \9763 , \9765 );
not \U$9081 ( \9767 , \8374 );
not \U$9082 ( \9768 , \7358 );
or \U$9083 ( \9769 , \9767 , \9768 );
nand \U$9084 ( \9770 , \7999 , \9423 );
nand \U$9085 ( \9771 , \9769 , \9770 );
not \U$9086 ( \9772 , \9771 );
not \U$9087 ( \9773 , \7601 );
or \U$9088 ( \9774 , \9772 , \9773 );
nand \U$9089 ( \9775 , \9689 , \9015 );
nand \U$9090 ( \9776 , \9774 , \9775 );
not \U$9091 ( \9777 , \9776 );
nand \U$9092 ( \9778 , \9766 , \9777 );
not \U$9093 ( \9779 , \8272 );
not \U$9094 ( \9780 , \7022 );
or \U$9095 ( \9781 , \9779 , \9780 );
not \U$9096 ( \9782 , \7020 );
nand \U$9097 ( \9783 , \9782 , \8271 );
nand \U$9098 ( \9784 , \9781 , \9783 );
not \U$9099 ( \9785 , \9784 );
not \U$9100 ( \9786 , \7018 );
or \U$9101 ( \9787 , \9785 , \9786 );
nand \U$9102 ( \9788 , \9716 , \7012 );
nand \U$9103 ( \9789 , \9787 , \9788 );
and \U$9104 ( \9790 , \9778 , \9789 );
nor \U$9105 ( \9791 , \9766 , \9777 );
nor \U$9106 ( \9792 , \9790 , \9791 );
not \U$9107 ( \9793 , \9792 );
nand \U$9108 ( \9794 , \9761 , \9793 );
nand \U$9109 ( \9795 , \9757 , \9794 );
not \U$9110 ( \9796 , \9661 );
not \U$9111 ( \9797 , \9699 );
or \U$9112 ( \9798 , \9796 , \9797 );
or \U$9113 ( \9799 , \9661 , \9699 );
nand \U$9114 ( \9800 , \9798 , \9799 );
xor \U$9115 ( \9801 , \9800 , \9672 );
not \U$9116 ( \9802 , \9801 );
not \U$9117 ( \9803 , \9721 );
nand \U$9118 ( \9804 , \9803 , \9739 );
not \U$9119 ( \9805 , \9804 );
not \U$9120 ( \9806 , \9750 );
or \U$9121 ( \9807 , \9805 , \9806 );
not \U$9122 ( \9808 , \9739 );
nand \U$9123 ( \9809 , \9808 , \9721 );
nand \U$9124 ( \9810 , \9807 , \9809 );
not \U$9125 ( \9811 , \9810 );
not \U$9126 ( \9812 , \9604 );
not \U$9127 ( \9813 , \9609 );
or \U$9128 ( \9814 , \9812 , \9813 );
nand \U$9129 ( \9815 , \9603 , \9592 );
nand \U$9130 ( \9816 , \9814 , \9815 );
not \U$9131 ( \9817 , \9607 );
and \U$9132 ( \9818 , \9816 , \9817 );
not \U$9133 ( \9819 , \9816 );
and \U$9134 ( \9820 , \9819 , \9607 );
nor \U$9135 ( \9821 , \9818 , \9820 );
not \U$9136 ( \9822 , \9821 );
or \U$9137 ( \9823 , \9811 , \9822 );
or \U$9138 ( \9824 , \9810 , \9821 );
nand \U$9139 ( \9825 , \9823 , \9824 );
not \U$9140 ( \9826 , \9825 );
or \U$9141 ( \9827 , \9802 , \9826 );
or \U$9142 ( \9828 , \9801 , \9825 );
nand \U$9143 ( \9829 , \9827 , \9828 );
xor \U$9144 ( \9830 , \9795 , \9829 );
and \U$9145 ( \9831 , \7373 , \8692 );
not \U$9146 ( \9832 , \7373 );
and \U$9147 ( \9833 , \9832 , \8954 );
or \U$9148 ( \9834 , \9831 , \9833 );
not \U$9149 ( \9835 , \9834 );
not \U$9150 ( \9836 , \7379 );
or \U$9151 ( \9837 , \9835 , \9836 );
nand \U$9152 ( \9838 , \9745 , \7531 );
nand \U$9153 ( \9839 , \9837 , \9838 );
not \U$9154 ( \9840 , \9839 );
not \U$9155 ( \9841 , \7729 );
not \U$9156 ( \9842 , \7607 );
not \U$9157 ( \9843 , \8101 );
or \U$9158 ( \9844 , \9842 , \9843 );
nand \U$9159 ( \9845 , \8100 , \7897 );
nand \U$9160 ( \9846 , \9844 , \9845 );
not \U$9161 ( \9847 , \9846 );
or \U$9162 ( \9848 , \9841 , \9847 );
nand \U$9163 ( \9849 , \9734 , \7737 );
nand \U$9164 ( \9850 , \9848 , \9849 );
not \U$9165 ( \9851 , \9850 );
not \U$9166 ( \9852 , \8691 );
or \U$9167 ( \9853 , \6691 , \9852 );
nand \U$9168 ( \9854 , \9851 , \9853 );
not \U$9169 ( \9855 , \8917 );
not \U$9170 ( \9856 , \8310 );
or \U$9171 ( \9857 , \9855 , \9856 );
nand \U$9172 ( \9858 , \7359 , \8309 );
nand \U$9173 ( \9859 , \9857 , \9858 );
not \U$9174 ( \9860 , \9859 );
not \U$9175 ( \9861 , \7601 );
or \U$9176 ( \9862 , \9860 , \9861 );
nand \U$9177 ( \9863 , \9771 , \7604 );
nand \U$9178 ( \9864 , \9862 , \9863 );
and \U$9179 ( \9865 , \9854 , \9864 );
nor \U$9180 ( \9866 , \9851 , \9853 );
nor \U$9181 ( \9867 , \9865 , \9866 );
nand \U$9182 ( \9868 , \9840 , \9867 );
not \U$9183 ( \9869 , \9868 );
not \U$9184 ( \9870 , \9789 );
not \U$9185 ( \9871 , \9766 );
and \U$9186 ( \9872 , \9777 , \9871 );
not \U$9187 ( \9873 , \9777 );
and \U$9188 ( \9874 , \9873 , \9766 );
nor \U$9189 ( \9875 , \9872 , \9874 );
not \U$9190 ( \9876 , \9875 );
or \U$9191 ( \9877 , \9870 , \9876 );
or \U$9192 ( \9878 , \9875 , \9789 );
nand \U$9193 ( \9879 , \9877 , \9878 );
not \U$9194 ( \9880 , \9879 );
or \U$9195 ( \9881 , \9869 , \9880 );
not \U$9196 ( \9882 , \9867 );
nand \U$9197 ( \9883 , \9882 , \9839 );
nand \U$9198 ( \9884 , \9881 , \9883 );
not \U$9199 ( \9885 , \9884 );
and \U$9200 ( \9886 , \9792 , \9758 );
not \U$9201 ( \9887 , \9792 );
and \U$9202 ( \9888 , \9887 , \9755 );
nor \U$9203 ( \9889 , \9886 , \9888 );
and \U$9204 ( \9890 , \9889 , \9751 );
not \U$9205 ( \9891 , \9889 );
and \U$9206 ( \9892 , \9891 , \9752 );
nor \U$9207 ( \9893 , \9890 , \9892 );
nand \U$9208 ( \9894 , \9885 , \9893 );
not \U$9209 ( \9895 , \9894 );
not \U$9210 ( \9896 , \9879 );
not \U$9211 ( \9897 , \9839 );
not \U$9212 ( \9898 , \9867 );
and \U$9213 ( \9899 , \9897 , \9898 );
and \U$9214 ( \9900 , \9839 , \9867 );
nor \U$9215 ( \9901 , \9899 , \9900 );
not \U$9216 ( \9902 , \9901 );
and \U$9217 ( \9903 , \9896 , \9902 );
and \U$9218 ( \9904 , \9879 , \9901 );
nor \U$9219 ( \9905 , \9903 , \9904 );
xor \U$9220 ( \9906 , \9850 , \9853 );
xnor \U$9221 ( \9907 , \9906 , \9864 );
not \U$9222 ( \9908 , \8563 );
not \U$9223 ( \9909 , \7700 );
or \U$9224 ( \9910 , \9908 , \9909 );
not \U$9225 ( \9911 , \8562 );
nand \U$9226 ( \9912 , \9911 , \7022 );
nand \U$9227 ( \9913 , \9910 , \9912 );
not \U$9228 ( \9914 , \9913 );
not \U$9229 ( \9915 , \7018 );
or \U$9230 ( \9916 , \9914 , \9915 );
nand \U$9231 ( \9917 , \9784 , \7012 );
nand \U$9232 ( \9918 , \9916 , \9917 );
not \U$9233 ( \9919 , \9918 );
not \U$9234 ( \9920 , \7594 );
not \U$9235 ( \9921 , \7005 );
not \U$9236 ( \9922 , \9921 );
or \U$9237 ( \9923 , \9920 , \9922 );
nand \U$9238 ( \9924 , \9923 , \8691 );
not \U$9239 ( \9925 , \9921 );
nand \U$9240 ( \9926 , \9925 , \7999 );
nand \U$9241 ( \9927 , \8030 , \9924 , \9926 );
not \U$9242 ( \9928 , \9927 );
not \U$9243 ( \9929 , \7737 );
not \U$9244 ( \9930 , \9846 );
or \U$9245 ( \9931 , \9929 , \9930 );
and \U$9246 ( \9932 , \8373 , \7608 );
not \U$9247 ( \9933 , \8373 );
and \U$9248 ( \9934 , \9933 , \7607 );
or \U$9249 ( \9935 , \9932 , \9934 );
nand \U$9250 ( \9936 , \9935 , \7729 );
nand \U$9251 ( \9937 , \9931 , \9936 );
nand \U$9252 ( \9938 , \9928 , \9937 );
nand \U$9253 ( \9939 , \9919 , \9938 );
and \U$9254 ( \9940 , \9907 , \9939 );
nor \U$9255 ( \9941 , \9919 , \9938 );
nor \U$9256 ( \9942 , \9940 , \9941 );
nand \U$9257 ( \9943 , \9905 , \9942 );
not \U$9258 ( \9944 , \9943 );
nand \U$9259 ( \9945 , \7011 , \8692 );
not \U$9260 ( \9946 , \9945 );
not \U$9261 ( \9947 , \7729 );
not \U$9262 ( \9948 , \7607 );
not \U$9263 ( \9949 , \8309 );
or \U$9264 ( \9950 , \9948 , \9949 );
nand \U$9265 ( \9951 , \8308 , \7897 );
nand \U$9266 ( \9952 , \9950 , \9951 );
not \U$9267 ( \9953 , \9952 );
or \U$9268 ( \9954 , \9947 , \9953 );
nand \U$9269 ( \9955 , \9935 , \7737 );
nand \U$9270 ( \9956 , \9954 , \9955 );
not \U$9271 ( \9957 , \9956 );
not \U$9272 ( \9958 , \9957 );
or \U$9273 ( \9959 , \9946 , \9958 );
and \U$9274 ( \9960 , \8562 , \7594 );
not \U$9275 ( \9961 , \8562 );
and \U$9276 ( \9962 , \9961 , \7359 );
or \U$9277 ( \9963 , \9960 , \9962 );
and \U$9278 ( \9964 , \7601 , \9963 );
and \U$9279 ( \9965 , \8270 , \7594 );
not \U$9280 ( \9966 , \8270 );
and \U$9281 ( \9967 , \9966 , \7999 );
or \U$9282 ( \9968 , \9965 , \9967 );
and \U$9283 ( \9969 , \9968 , \9015 );
nor \U$9284 ( \9970 , \9964 , \9969 );
not \U$9285 ( \9971 , \9970 );
nand \U$9286 ( \9972 , \9959 , \9971 );
not \U$9287 ( \9973 , \9945 );
nand \U$9288 ( \9974 , \9973 , \9956 );
nand \U$9289 ( \9975 , \9972 , \9974 );
not \U$9290 ( \9976 , \9975 );
and \U$9291 ( \9977 , \7601 , \9968 );
and \U$9292 ( \9978 , \9859 , \9015 );
nor \U$9293 ( \9979 , \9977 , \9978 );
not \U$9294 ( \9980 , \9937 );
not \U$9295 ( \9981 , \9927 );
and \U$9296 ( \9982 , \9980 , \9981 );
and \U$9297 ( \9983 , \9937 , \9927 );
nor \U$9298 ( \9984 , \9982 , \9983 );
xor \U$9299 ( \9985 , \9979 , \9984 );
not \U$9300 ( \9986 , \8692 );
not \U$9301 ( \9987 , \7700 );
or \U$9302 ( \9988 , \9986 , \9987 );
nand \U$9303 ( \9989 , \7699 , \9852 );
nand \U$9304 ( \9990 , \9988 , \9989 );
not \U$9305 ( \9991 , \9990 );
not \U$9306 ( \9992 , \7018 );
or \U$9307 ( \9993 , \9991 , \9992 );
nand \U$9308 ( \9994 , \9913 , \7012 );
nand \U$9309 ( \9995 , \9993 , \9994 );
not \U$9310 ( \9996 , \9995 );
xor \U$9311 ( \9997 , \9985 , \9996 );
nand \U$9312 ( \9998 , \9976 , \9997 );
not \U$9313 ( \9999 , \9998 );
not \U$9314 ( \10000 , \7608 );
not \U$9315 ( \10001 , \7348 );
or \U$9316 ( \10002 , \10000 , \10001 );
nand \U$9317 ( \10003 , \10002 , \8691 );
nand \U$9318 ( \10004 , \7349 , \7607 );
and \U$9319 ( \10005 , \8920 , \10003 , \10004 );
not \U$9320 ( \10006 , \7737 );
not \U$9321 ( \10007 , \9952 );
or \U$9322 ( \10008 , \10006 , \10007 );
and \U$9323 ( \10009 , \8270 , \7608 );
not \U$9324 ( \10010 , \8270 );
and \U$9325 ( \10011 , \10010 , \7607 );
or \U$9326 ( \10012 , \10009 , \10011 );
nand \U$9327 ( \10013 , \10012 , \7729 );
nand \U$9328 ( \10014 , \10008 , \10013 );
xor \U$9329 ( \10015 , \10005 , \10014 );
and \U$9330 ( \10016 , \9852 , \7358 );
not \U$9331 ( \10017 , \9852 );
and \U$9332 ( \10018 , \10017 , \7359 );
nor \U$9333 ( \10019 , \10016 , \10018 );
not \U$9334 ( \10020 , \10019 );
not \U$9335 ( \10021 , \7601 );
or \U$9336 ( \10022 , \10020 , \10021 );
nand \U$9337 ( \10023 , \9963 , \9015 );
nand \U$9338 ( \10024 , \10022 , \10023 );
nor \U$9339 ( \10025 , \10015 , \10024 );
not \U$9340 ( \10026 , \7737 );
not \U$9341 ( \10027 , \10012 );
or \U$9342 ( \10028 , \10026 , \10027 );
not \U$9343 ( \10029 , \7607 );
not \U$9344 ( \10030 , \8562 );
not \U$9345 ( \10031 , \10030 );
or \U$9346 ( \10032 , \10029 , \10031 );
nand \U$9347 ( \10033 , \8562 , \7608 );
nand \U$9348 ( \10034 , \10032 , \10033 );
nand \U$9349 ( \10035 , \10034 , \7729 );
nand \U$9350 ( \10036 , \10028 , \10035 );
not \U$9351 ( \10037 , \10036 );
nor \U$9352 ( \10038 , \8954 , \7346 );
not \U$9353 ( \10039 , \10038 );
nand \U$9354 ( \10040 , \10037 , \10039 );
not \U$9355 ( \10041 , \8692 );
not \U$9356 ( \10042 , \7728 );
and \U$9357 ( \10043 , \10041 , \10042 );
and \U$9358 ( \10044 , \10034 , \7903 );
nor \U$9359 ( \10045 , \10043 , \10044 );
nand \U$9360 ( \10046 , \8692 , \7737 );
nand \U$9361 ( \10047 , \10046 , \7607 );
nor \U$9362 ( \10048 , \10045 , \10047 );
and \U$9363 ( \10049 , \10040 , \10048 );
and \U$9364 ( \10050 , \10036 , \10038 );
nor \U$9365 ( \10051 , \10049 , \10050 );
or \U$9366 ( \10052 , \10025 , \10051 );
nand \U$9367 ( \10053 , \10015 , \10024 );
nand \U$9368 ( \10054 , \10052 , \10053 );
not \U$9369 ( \10055 , \10054 );
and \U$9370 ( \10056 , \10005 , \10014 );
not \U$9371 ( \10057 , \10056 );
xor \U$9372 ( \10058 , \9945 , \9956 );
xnor \U$9373 ( \10059 , \10058 , \9970 );
nand \U$9374 ( \10060 , \10057 , \10059 );
not \U$9375 ( \10061 , \10060 );
or \U$9376 ( \10062 , \10055 , \10061 );
not \U$9377 ( \10063 , \10059 );
nand \U$9378 ( \10064 , \10063 , \10056 );
nand \U$9379 ( \10065 , \10062 , \10064 );
not \U$9380 ( \10066 , \10065 );
or \U$9381 ( \10067 , \9999 , \10066 );
not \U$9382 ( \10068 , \9997 );
nand \U$9383 ( \10069 , \10068 , \9975 );
nand \U$9384 ( \10070 , \10067 , \10069 );
not \U$9385 ( \10071 , \10070 );
not \U$9386 ( \10072 , \9907 );
xor \U$9387 ( \10073 , \9918 , \9938 );
not \U$9388 ( \10074 , \10073 );
and \U$9389 ( \10075 , \10072 , \10074 );
and \U$9390 ( \10076 , \9907 , \10073 );
nor \U$9391 ( \10077 , \10075 , \10076 );
xor \U$9392 ( \10078 , \9979 , \9984 );
and \U$9393 ( \10079 , \10078 , \9996 );
and \U$9394 ( \10080 , \9979 , \9984 );
or \U$9395 ( \10081 , \10079 , \10080 );
nand \U$9396 ( \10082 , \10077 , \10081 );
not \U$9397 ( \10083 , \10082 );
or \U$9398 ( \10084 , \10071 , \10083 );
not \U$9399 ( \10085 , \10077 );
not \U$9400 ( \10086 , \10081 );
nand \U$9401 ( \10087 , \10085 , \10086 );
nand \U$9402 ( \10088 , \10084 , \10087 );
not \U$9403 ( \10089 , \10088 );
or \U$9404 ( \10090 , \9944 , \10089 );
not \U$9405 ( \10091 , \9905 );
not \U$9406 ( \10092 , \9942 );
nand \U$9407 ( \10093 , \10091 , \10092 );
nand \U$9408 ( \10094 , \10090 , \10093 );
not \U$9409 ( \10095 , \10094 );
or \U$9410 ( \10096 , \9895 , \10095 );
not \U$9411 ( \10097 , \9893 );
nand \U$9412 ( \10098 , \10097 , \9884 );
nand \U$9413 ( \10099 , \10096 , \10098 );
and \U$9414 ( \10100 , \9830 , \10099 );
and \U$9415 ( \10101 , \9795 , \9829 );
or \U$9416 ( \10102 , \10100 , \10101 );
xor \U$9417 ( \10103 , \9650 , \9702 );
xor \U$9418 ( \10104 , \10103 , \9705 );
not \U$9419 ( \10105 , \9810 );
nand \U$9420 ( \10106 , \10105 , \9821 );
not \U$9421 ( \10107 , \10106 );
not \U$9422 ( \10108 , \9801 );
not \U$9423 ( \10109 , \10108 );
or \U$9424 ( \10110 , \10107 , \10109 );
not \U$9425 ( \10111 , \9821 );
nand \U$9426 ( \10112 , \10111 , \9810 );
nand \U$9427 ( \10113 , \10110 , \10112 );
or \U$9428 ( \10114 , \10104 , \10113 );
nand \U$9429 ( \10115 , \9710 , \10102 , \10114 );
and \U$9430 ( \10116 , \10104 , \10113 );
nand \U$9431 ( \10117 , \9710 , \10116 );
nand \U$9432 ( \10118 , \9648 , \9708 );
nand \U$9433 ( \10119 , \10115 , \10117 , \10118 );
not \U$9434 ( \10120 , \9573 );
not \U$9435 ( \10121 , \9623 );
nand \U$9436 ( \10122 , \10120 , \10121 );
and \U$9437 ( \10123 , \9564 , \10122 );
nand \U$9438 ( \10124 , \10119 , \9645 , \10123 , \9473 );
nand \U$9439 ( \10125 , \9646 , \10124 );
not \U$9440 ( \10126 , \8867 );
not \U$9441 ( \10127 , \8974 );
nand \U$9442 ( \10128 , \10126 , \10127 );
nand \U$9443 ( \10129 , \8856 , \10128 );
nor \U$9444 ( \10130 , \10129 , \9189 );
nand \U$9445 ( \10131 , \10125 , \9338 , \10130 );
and \U$9446 ( \10132 , \9321 , \9336 );
nor \U$9447 ( \10133 , \9323 , \9327 );
nand \U$9448 ( \10134 , \9296 , \10133 );
nor \U$9449 ( \10135 , \9315 , \9320 );
nor \U$9450 ( \10136 , \9270 , \9295 );
nor \U$9451 ( \10137 , \10135 , \10136 );
nand \U$9452 ( \10138 , \10134 , \10137 );
nand \U$9453 ( \10139 , \10132 , \10138 );
nor \U$9454 ( \10140 , \9331 , \9335 );
not \U$9455 ( \10141 , \10140 );
nand \U$9456 ( \10142 , \9339 , \10131 , \10139 , \10141 );
not \U$9457 ( \10143 , \10142 );
or \U$9458 ( \10144 , \7995 , \10143 );
not \U$9459 ( \10145 , \7238 );
buf \U$9460 ( \10146 , \7559 );
not \U$9461 ( \10147 , \10146 );
and \U$9462 ( \10148 , \7563 , \7810 );
and \U$9463 ( \10149 , \7813 , \7988 );
or \U$9464 ( \10150 , \10148 , \10149 );
not \U$9465 ( \10151 , \7811 );
nand \U$9466 ( \10152 , \10150 , \10151 );
not \U$9467 ( \10153 , \7552 );
or \U$9468 ( \10154 , \10152 , \10153 );
not \U$9469 ( \10155 , \7335 );
not \U$9470 ( \10156 , \7551 );
nand \U$9471 ( \10157 , \10155 , \10156 );
nand \U$9472 ( \10158 , \10154 , \10157 );
not \U$9473 ( \10159 , \10158 );
or \U$9474 ( \10160 , \10147 , \10159 );
or \U$9475 ( \10161 , \7558 , \7556 );
nand \U$9476 ( \10162 , \10160 , \10161 );
not \U$9477 ( \10163 , \10162 );
or \U$9478 ( \10164 , \10145 , \10163 );
not \U$9479 ( \10165 , \7225 );
not \U$9480 ( \10166 , \10165 );
not \U$9481 ( \10167 , \7191 );
not \U$9482 ( \10168 , \7193 );
nand \U$9483 ( \10169 , \10167 , \10168 );
buf \U$9484 ( \10170 , \6930 );
or \U$9485 ( \10171 , \10169 , \10170 );
nand \U$9486 ( \10172 , \6866 , \6929 );
nand \U$9487 ( \10173 , \10171 , \10172 );
not \U$9488 ( \10174 , \10173 );
or \U$9489 ( \10175 , \10166 , \10174 );
nand \U$9490 ( \10176 , \7199 , \7224 );
nand \U$9491 ( \10177 , \10175 , \10176 );
and \U$9492 ( \10178 , \10177 , \7237 );
nor \U$9493 ( \10179 , \7230 , \7236 );
nor \U$9494 ( \10180 , \10178 , \10179 );
nand \U$9495 ( \10181 , \10164 , \10180 );
not \U$9496 ( \10182 , \10181 );
nand \U$9497 ( \10183 , \10144 , \10182 );
not \U$9498 ( \10184 , \10183 );
or \U$9499 ( \10185 , \6494 , \10184 );
nand \U$9500 ( \10186 , \6490 , \6492 );
nand \U$9501 ( \10187 , \10185 , \10186 );
not \U$9502 ( \10188 , \10187 );
or \U$9503 ( \10189 , \6415 , \10188 );
or \U$9504 ( \10190 , \6414 , \10187 );
nand \U$9505 ( \10191 , \10189 , \10190 );
not \U$9506 ( \10192 , \5948 );
not \U$9507 ( \10193 , \10192 );
nand \U$9508 ( \10194 , \10191 , \10193 );
nand \U$9509 ( \10195 , \5950 , \10194 );
buf \U$9510 ( \10196 , \10195 );
xor \U$9511 ( \10197 , \1782 , \1845 );
xor \U$9512 ( \10198 , \10197 , \5196 );
and \U$9513 ( \10199 , \10192 , \10198 );
not \U$9514 ( \10200 , \10192 );
nand \U$9515 ( \10201 , \10186 , \6493 );
xnor \U$9516 ( \10202 , \10183 , \10201 );
and \U$9517 ( \10203 , \10200 , \10202 );
or \U$9518 ( \10204 , \10199 , \10203 );
buf \U$9519 ( \10205 , \10204 );
buf \U$9520 ( \10206 , \5179 );
not \U$9521 ( \10207 , \10206 );
not \U$9522 ( \10208 , \5037 );
or \U$9523 ( \10209 , \10207 , \10208 );
nand \U$9524 ( \10210 , \10209 , \5163 );
nand \U$9525 ( \10211 , \10210 , \5191 );
not \U$9526 ( \10212 , \5102 );
nand \U$9527 ( \10213 , \10212 , \5193 );
xor \U$9528 ( \10214 , \10211 , \10213 );
and \U$9529 ( \10215 , \10192 , \10214 );
not \U$9530 ( \10216 , \10192 );
and \U$9531 ( \10217 , \7992 , \7226 );
not \U$9532 ( \10218 , \9646 );
and \U$9533 ( \10219 , \10218 , \10130 , \9338 );
buf \U$9534 ( \10220 , \10219 );
and \U$9535 ( \10221 , \10217 , \10220 );
nand \U$9536 ( \10222 , \9190 , \9338 );
not \U$9537 ( \10223 , \10222 );
and \U$9538 ( \10224 , \10223 , \10217 );
nor \U$9539 ( \10225 , \10221 , \10224 );
not \U$9540 ( \10226 , \7226 );
not \U$9541 ( \10227 , \10226 );
not \U$9542 ( \10228 , \10146 );
not \U$9543 ( \10229 , \10158 );
or \U$9544 ( \10230 , \10228 , \10229 );
nand \U$9545 ( \10231 , \10230 , \10161 );
and \U$9546 ( \10232 , \10227 , \10231 );
nor \U$9547 ( \10233 , \10232 , \10177 );
nand \U$9548 ( \10234 , \7992 , \10140 );
not \U$9549 ( \10235 , \10234 );
not \U$9550 ( \10236 , \10226 );
and \U$9551 ( \10237 , \10235 , \10236 );
and \U$9552 ( \10238 , \9338 , \9197 );
and \U$9553 ( \10239 , \10217 , \10238 );
nor \U$9554 ( \10240 , \10237 , \10239 );
and \U$9555 ( \10241 , \10119 , \9645 , \10123 , \9473 );
and \U$9556 ( \10242 , \7992 , \10130 , \10241 );
and \U$9557 ( \10243 , \9338 , \7226 );
and \U$9558 ( \10244 , \10242 , \10243 );
nand \U$9559 ( \10245 , \7992 , \10132 );
nand \U$9560 ( \10246 , \10138 , \7226 );
nor \U$9561 ( \10247 , \10245 , \10246 );
nor \U$9562 ( \10248 , \10244 , \10247 );
nand \U$9563 ( \10249 , \10225 , \10233 , \10240 , \10248 );
not \U$9564 ( \10250 , \10179 );
nand \U$9565 ( \10251 , \10250 , \7237 );
xor \U$9566 ( \10252 , \10249 , \10251 );
and \U$9567 ( \10253 , \10216 , \10252 );
nor \U$9568 ( \10254 , \10215 , \10253 );
buf \U$9569 ( \10255 , \10254 );
nand \U$9570 ( \10256 , \10165 , \10176 );
not \U$9571 ( \10257 , \10256 );
not \U$9572 ( \10258 , \7195 );
not \U$9573 ( \10259 , \10258 );
not \U$9574 ( \10260 , \10222 );
not \U$9575 ( \10261 , \7993 );
and \U$9576 ( \10262 , \10260 , \10261 );
buf \U$9577 ( \10263 , \9338 );
and \U$9578 ( \10264 , \10242 , \10263 );
nor \U$9579 ( \10265 , \10262 , \10264 );
not \U$9580 ( \10266 , \10234 );
nor \U$9581 ( \10267 , \10266 , \10162 );
or \U$9582 ( \10268 , \10219 , \10238 );
not \U$9583 ( \10269 , \7993 );
nand \U$9584 ( \10270 , \10268 , \10269 );
not \U$9585 ( \10271 , \10245 );
nand \U$9586 ( \10272 , \10271 , \10138 );
nand \U$9587 ( \10273 , \10265 , \10267 , \10270 , \10272 );
not \U$9588 ( \10274 , \10273 );
or \U$9589 ( \10275 , \10259 , \10274 );
not \U$9590 ( \10276 , \10173 );
nand \U$9591 ( \10277 , \10275 , \10276 );
not \U$9592 ( \10278 , \10277 );
or \U$9593 ( \10279 , \10257 , \10278 );
or \U$9594 ( \10280 , \10256 , \10277 );
nand \U$9595 ( \10281 , \10279 , \10280 );
nand \U$9596 ( \10282 , \10281 , \10193 );
not \U$9597 ( \10283 , \5948 );
not \U$9598 ( \10284 , \5153 );
not \U$9599 ( \10285 , \10284 );
not \U$9600 ( \10286 , \4712 );
buf \U$9601 ( \10287 , \4729 );
nand \U$9602 ( \10288 , \10286 , \10287 );
not \U$9603 ( \10289 , \3456 );
nand \U$9604 ( \10290 , \10288 , \10289 );
and \U$9605 ( \10291 , \10290 , \4730 );
buf \U$9606 ( \10292 , \3446 );
nor \U$9607 ( \10293 , \10291 , \10292 );
or \U$9608 ( \10294 , \10293 , \4714 );
nand \U$9609 ( \10295 , \10294 , \5036 );
not \U$9610 ( \10296 , \4707 );
not \U$9611 ( \10297 , \4727 );
nand \U$9612 ( \10298 , \10296 , \4721 , \10297 );
not \U$9613 ( \10299 , \3458 );
nor \U$9614 ( \10300 , \10299 , \5035 );
nand \U$9615 ( \10301 , \10298 , \10300 );
nand \U$9616 ( \10302 , \10295 , \10301 , \10206 );
not \U$9617 ( \10303 , \10302 );
or \U$9618 ( \10304 , \10285 , \10303 );
not \U$9619 ( \10305 , \5187 );
nand \U$9620 ( \10306 , \10304 , \10305 );
nor \U$9621 ( \10307 , \5190 , \5162 );
and \U$9622 ( \10308 , \10306 , \10307 );
not \U$9623 ( \10309 , \10306 );
not \U$9624 ( \10310 , \10307 );
and \U$9625 ( \10311 , \10309 , \10310 );
nor \U$9626 ( \10312 , \10308 , \10311 );
nand \U$9627 ( \10313 , \10283 , \10312 );
nand \U$9628 ( \10314 , \10282 , \10313 );
buf \U$9629 ( \10315 , \10314 );
not \U$9630 ( \10316 , \5135 );
not \U$9631 ( \10317 , \10302 );
or \U$9632 ( \10318 , \10316 , \10317 );
nand \U$9633 ( \10319 , \10318 , \5183 );
nand \U$9634 ( \10320 , \5186 , \5152 );
xor \U$9635 ( \10321 , \10319 , \10320 );
and \U$9636 ( \10322 , \10192 , \10321 );
not \U$9637 ( \10323 , \10192 );
not \U$9638 ( \10324 , \7194 );
not \U$9639 ( \10325 , \10273 );
or \U$9640 ( \10326 , \10324 , \10325 );
nand \U$9641 ( \10327 , \10326 , \10169 );
not \U$9642 ( \10328 , \10172 );
nor \U$9643 ( \10329 , \10328 , \10170 );
xnor \U$9644 ( \10330 , \10327 , \10329 );
and \U$9645 ( \10331 , \10323 , \10330 );
nor \U$9646 ( \10332 , \10322 , \10331 );
buf \U$9647 ( \10333 , \10332 );
not \U$9648 ( \10334 , \5948 );
nand \U$9649 ( \10335 , \7194 , \10169 );
xnor \U$9650 ( \10336 , \10273 , \10335 );
not \U$9651 ( \10337 , \10336 );
or \U$9652 ( \10338 , \10334 , \10337 );
nand \U$9653 ( \10339 , \5183 , \5135 );
not \U$9654 ( \10340 , \10339 );
not \U$9655 ( \10341 , \10302 );
or \U$9656 ( \10342 , \10340 , \10341 );
or \U$9657 ( \10343 , \10339 , \10302 );
nand \U$9658 ( \10344 , \10342 , \10343 );
nand \U$9659 ( \10345 , \10344 , \10192 );
nand \U$9660 ( \10346 , \10338 , \10345 );
buf \U$9661 ( \10347 , \10346 );
nand \U$9662 ( \10348 , \4739 , \4914 );
not \U$9663 ( \10349 , \10348 );
not \U$9664 ( \10350 , \4906 );
and \U$9665 ( \10351 , \10349 , \10350 );
nor \U$9666 ( \10352 , \10351 , \5171 );
not \U$9667 ( \10353 , \10352 );
and \U$9668 ( \10354 , \10353 , \4975 );
not \U$9669 ( \10355 , \5175 );
nor \U$9670 ( \10356 , \10354 , \10355 );
not \U$9671 ( \10357 , \5178 );
nand \U$9672 ( \10358 , \10357 , \5034 );
xnor \U$9673 ( \10359 , \10356 , \10358 );
and \U$9674 ( \10360 , \10192 , \10359 );
not \U$9675 ( \10361 , \10192 );
not \U$9676 ( \10362 , \10153 );
not \U$9677 ( \10363 , \10362 );
not \U$9678 ( \10364 , \7990 );
not \U$9679 ( \10365 , \10142 );
or \U$9680 ( \10366 , \10364 , \10365 );
buf \U$9681 ( \10367 , \10152 );
nand \U$9682 ( \10368 , \10366 , \10367 );
not \U$9683 ( \10369 , \10368 );
or \U$9684 ( \10370 , \10363 , \10369 );
buf \U$9685 ( \10371 , \10157 );
nand \U$9686 ( \10372 , \10370 , \10371 );
nand \U$9687 ( \10373 , \10161 , \10146 );
xor \U$9688 ( \10374 , \10372 , \10373 );
and \U$9689 ( \10375 , \10361 , \10374 );
nor \U$9690 ( \10376 , \10360 , \10375 );
buf \U$9691 ( \10377 , \10376 );
nand \U$9692 ( \10378 , \5175 , \4975 );
xor \U$9693 ( \10379 , \10353 , \10378 );
and \U$9694 ( \10380 , \10192 , \10379 );
not \U$9695 ( \10381 , \10192 );
nand \U$9696 ( \10382 , \10371 , \10362 );
xor \U$9697 ( \10383 , \10368 , \10382 );
and \U$9698 ( \10384 , \10381 , \10383 );
nor \U$9699 ( \10385 , \10380 , \10384 );
buf \U$9700 ( \10386 , \10385 );
nand \U$9701 ( \10387 , \10348 , \5168 );
nand \U$9702 ( \10388 , \5170 , \4907 );
xor \U$9703 ( \10389 , \10387 , \10388 );
and \U$9704 ( \10390 , \10192 , \10389 );
not \U$9705 ( \10391 , \10192 );
not \U$9706 ( \10392 , \7989 );
not \U$9707 ( \10393 , \10392 );
buf \U$9708 ( \10394 , \10142 );
not \U$9709 ( \10395 , \10394 );
or \U$9710 ( \10396 , \10393 , \10395 );
not \U$9711 ( \10397 , \10149 );
nand \U$9712 ( \10398 , \10396 , \10397 );
not \U$9713 ( \10399 , \10148 );
nand \U$9714 ( \10400 , \10399 , \10151 );
xor \U$9715 ( \10401 , \10398 , \10400 );
and \U$9716 ( \10402 , \10391 , \10401 );
nor \U$9717 ( \10403 , \10390 , \10402 );
buf \U$9718 ( \10404 , \10403 );
not \U$9719 ( \10405 , \5948 );
not \U$9720 ( \10406 , \7989 );
nand \U$9721 ( \10407 , \10406 , \10397 );
not \U$9722 ( \10408 , \10407 );
not \U$9723 ( \10409 , \10394 );
or \U$9724 ( \10410 , \10408 , \10409 );
or \U$9725 ( \10411 , \10407 , \10394 );
nand \U$9726 ( \10412 , \10410 , \10411 );
not \U$9727 ( \10413 , \10412 );
or \U$9728 ( \10414 , \10405 , \10413 );
nand \U$9729 ( \10415 , \5168 , \4914 );
xnor \U$9730 ( \10416 , \4739 , \10415 );
nand \U$9731 ( \10417 , \10416 , \10192 );
nand \U$9732 ( \10418 , \10414 , \10417 );
buf \U$9733 ( \10419 , \10418 );
not \U$9734 ( \10420 , \10289 );
not \U$9735 ( \10421 , \3259 );
not \U$9736 ( \10422 , \10298 );
or \U$9737 ( \10423 , \10421 , \10422 );
not \U$9738 ( \10424 , \10288 );
nand \U$9739 ( \10425 , \10423 , \10424 );
not \U$9740 ( \10426 , \10425 );
or \U$9741 ( \10427 , \10420 , \10426 );
nand \U$9742 ( \10428 , \10427 , \4730 );
nor \U$9743 ( \10429 , \4714 , \10292 );
xnor \U$9744 ( \10430 , \10428 , \10429 );
and \U$9745 ( \10431 , \10192 , \10430 );
not \U$9746 ( \10432 , \10192 );
not \U$9747 ( \10433 , \9321 );
buf \U$9748 ( \10434 , \9296 );
and \U$9749 ( \10435 , \10434 , \9328 );
not \U$9750 ( \10436 , \10435 );
not \U$9751 ( \10437 , \10129 );
nand \U$9752 ( \10438 , \10437 , \10125 );
buf \U$9753 ( \10439 , \9189 );
or \U$9754 ( \10440 , \10438 , \10439 );
not \U$9755 ( \10441 , \9199 );
nand \U$9756 ( \10442 , \10440 , \10441 );
not \U$9757 ( \10443 , \10442 );
or \U$9758 ( \10444 , \10436 , \10443 );
not \U$9759 ( \10445 , \10134 );
nor \U$9760 ( \10446 , \10445 , \10136 );
nand \U$9761 ( \10447 , \10444 , \10446 );
not \U$9762 ( \10448 , \10447 );
or \U$9763 ( \10449 , \10433 , \10448 );
not \U$9764 ( \10450 , \10135 );
nand \U$9765 ( \10451 , \10449 , \10450 );
nand \U$9766 ( \10452 , \10141 , \9336 );
xor \U$9767 ( \10453 , \10451 , \10452 );
and \U$9768 ( \10454 , \10432 , \10453 );
nor \U$9769 ( \10455 , \10431 , \10454 );
buf \U$9770 ( \10456 , \10455 );
nand \U$9771 ( \10457 , \4730 , \10289 );
xor \U$9772 ( \10458 , \10425 , \10457 );
and \U$9773 ( \10459 , \10192 , \10458 );
not \U$9774 ( \10460 , \10192 );
nand \U$9775 ( \10461 , \10450 , \9321 );
xor \U$9776 ( \10462 , \10461 , \10447 );
and \U$9777 ( \10463 , \10460 , \10462 );
nor \U$9778 ( \10464 , \10459 , \10463 );
buf \U$9779 ( \10465 , \10464 );
not \U$9780 ( \10466 , \3258 );
not \U$9781 ( \10467 , \10298 );
or \U$9782 ( \10468 , \10466 , \10467 );
not \U$9783 ( \10469 , \4711 );
nand \U$9784 ( \10470 , \10468 , \10469 );
nand \U$9785 ( \10471 , \3082 , \10287 );
xor \U$9786 ( \10472 , \10470 , \10471 );
and \U$9787 ( \10473 , \10192 , \10472 );
not \U$9788 ( \10474 , \10192 );
not \U$9789 ( \10475 , \9328 );
not \U$9790 ( \10476 , \10442 );
or \U$9791 ( \10477 , \10475 , \10476 );
buf \U$9792 ( \10478 , \10133 );
not \U$9793 ( \10479 , \10478 );
nand \U$9794 ( \10480 , \10477 , \10479 );
not \U$9795 ( \10481 , \10434 );
nor \U$9796 ( \10482 , \10481 , \10136 );
and \U$9797 ( \10483 , \10480 , \10482 );
not \U$9798 ( \10484 , \10480 );
not \U$9799 ( \10485 , \10482 );
and \U$9800 ( \10486 , \10484 , \10485 );
or \U$9801 ( \10487 , \10483 , \10486 );
and \U$9802 ( \10488 , \10474 , \10487 );
nor \U$9803 ( \10489 , \10473 , \10488 );
buf \U$9804 ( \10490 , \10489 );
nand \U$9805 ( \10491 , \10469 , \3258 );
xnor \U$9806 ( \10492 , \10298 , \10491 );
and \U$9807 ( \10493 , \10192 , \10492 );
not \U$9808 ( \10494 , \10192 );
not \U$9809 ( \10495 , \9328 );
nor \U$9810 ( \10496 , \10495 , \10478 );
xor \U$9811 ( \10497 , \10496 , \10442 );
and \U$9812 ( \10498 , \10494 , \10497 );
or \U$9813 ( \10499 , \10493 , \10498 );
buf \U$9814 ( \10500 , \10499 );
not \U$9815 ( \10501 , \4697 );
not \U$9816 ( \10502 , \4662 );
buf \U$9817 ( \10503 , \4579 );
and \U$9818 ( \10504 , \10503 , \4674 );
not \U$9819 ( \10505 , \10504 );
or \U$9820 ( \10506 , \10502 , \10505 );
not \U$9821 ( \10507 , \4720 );
nand \U$9822 ( \10508 , \10506 , \10507 );
not \U$9823 ( \10509 , \10508 );
or \U$9824 ( \10510 , \10501 , \10509 );
not \U$9825 ( \10511 , \4722 );
nand \U$9826 ( \10512 , \10510 , \10511 );
nand \U$9827 ( \10513 , \4726 , \4704 );
xor \U$9828 ( \10514 , \10512 , \10513 );
and \U$9829 ( \10515 , \10192 , \10514 );
not \U$9830 ( \10516 , \10192 );
buf \U$9831 ( \10517 , \9099 );
not \U$9832 ( \10518 , \10517 );
buf \U$9833 ( \10519 , \8977 );
nand \U$9834 ( \10520 , \10438 , \10519 );
not \U$9835 ( \10521 , \10520 );
or \U$9836 ( \10522 , \10518 , \10521 );
not \U$9837 ( \10523 , \9192 );
nand \U$9838 ( \10524 , \10522 , \10523 );
nand \U$9839 ( \10525 , \9196 , \9188 );
xor \U$9840 ( \10526 , \10524 , \10525 );
and \U$9841 ( \10527 , \10516 , \10526 );
nor \U$9842 ( \10528 , \10515 , \10527 );
buf \U$9843 ( \10529 , \10528 );
and \U$9844 ( \10530 , \10511 , \4697 );
and \U$9845 ( \10531 , \10530 , \10508 );
not \U$9846 ( \10532 , \10530 );
not \U$9847 ( \10533 , \10508 );
and \U$9848 ( \10534 , \10532 , \10533 );
nor \U$9849 ( \10535 , \10531 , \10534 );
not \U$9850 ( \10536 , \10535 );
and \U$9851 ( \10537 , \10192 , \10536 );
not \U$9852 ( \10538 , \10192 );
nand \U$9853 ( \10539 , \10523 , \10517 );
xor \U$9854 ( \10540 , \10520 , \10539 );
and \U$9855 ( \10541 , \10538 , \10540 );
nor \U$9856 ( \10542 , \10537 , \10541 );
buf \U$9857 ( \10543 , \10542 );
not \U$9858 ( \10544 , \10504 );
buf \U$9859 ( \10545 , \4717 );
nand \U$9860 ( \10546 , \10544 , \10545 );
nand \U$9861 ( \10547 , \4662 , \4718 );
xor \U$9862 ( \10548 , \10546 , \10547 );
and \U$9863 ( \10549 , \10192 , \10548 );
not \U$9864 ( \10550 , \10192 );
not \U$9865 ( \10551 , \10128 );
not \U$9866 ( \10552 , \10125 );
or \U$9867 ( \10553 , \10551 , \10552 );
nand \U$9868 ( \10554 , \10553 , \8975 );
nand \U$9869 ( \10555 , \8857 , \8856 );
xor \U$9870 ( \10556 , \10554 , \10555 );
and \U$9871 ( \10557 , \10550 , \10556 );
nor \U$9872 ( \10558 , \10549 , \10557 );
buf \U$9873 ( \10559 , \10558 );
not \U$9874 ( \10560 , \5948 );
nand \U$9875 ( \10561 , \8975 , \10128 );
not \U$9876 ( \10562 , \10561 );
not \U$9877 ( \10563 , \10125 );
or \U$9878 ( \10564 , \10562 , \10563 );
or \U$9879 ( \10565 , \10125 , \10561 );
nand \U$9880 ( \10566 , \10564 , \10565 );
not \U$9881 ( \10567 , \10566 );
or \U$9882 ( \10568 , \10560 , \10567 );
nand \U$9883 ( \10569 , \10545 , \4674 );
not \U$9884 ( \10570 , \10569 );
buf \U$9885 ( \10571 , \10503 );
not \U$9886 ( \10572 , \10571 );
or \U$9887 ( \10573 , \10570 , \10572 );
or \U$9888 ( \10574 , \10571 , \10569 );
nand \U$9889 ( \10575 , \10573 , \10574 );
nand \U$9890 ( \10576 , \10575 , \10192 );
nand \U$9891 ( \10577 , \10568 , \10576 );
buf \U$9892 ( \10578 , \10577 );
not \U$9893 ( \10579 , \4574 );
not \U$9894 ( \10580 , \10579 );
not \U$9895 ( \10581 , \4571 );
or \U$9896 ( \10582 , \10580 , \10581 );
not \U$9897 ( \10583 , \3988 );
nand \U$9898 ( \10584 , \10582 , \10583 );
not \U$9899 ( \10585 , \4572 );
and \U$9900 ( \10586 , \10584 , \10585 );
not \U$9901 ( \10587 , \4099 );
nor \U$9902 ( \10588 , \10586 , \10587 );
nand \U$9903 ( \10589 , \4184 , \4578 );
xor \U$9904 ( \10590 , \10588 , \10589 );
not \U$9905 ( \10591 , \10590 );
nor \U$9906 ( \10592 , \10591 , \5948 );
not \U$9907 ( \10593 , \10592 );
nand \U$9908 ( \10594 , \9642 , \9645 );
not \U$9909 ( \10595 , \10594 );
buf \U$9910 ( \10596 , \9473 );
not \U$9911 ( \10597 , \10596 );
not \U$9912 ( \10598 , \10123 );
not \U$9913 ( \10599 , \10119 );
or \U$9914 ( \10600 , \10598 , \10599 );
nand \U$9915 ( \10601 , \10600 , \9627 );
not \U$9916 ( \10602 , \10601 );
or \U$9917 ( \10603 , \10597 , \10602 );
buf \U$9918 ( \10604 , \9630 );
nand \U$9919 ( \10605 , \10603 , \10604 );
not \U$9920 ( \10606 , \10605 );
or \U$9921 ( \10607 , \10595 , \10606 );
or \U$9922 ( \10608 , \10605 , \10594 );
nand \U$9923 ( \10609 , \10607 , \10608 );
nand \U$9924 ( \10610 , \10609 , \5948 );
nand \U$9925 ( \10611 , \10593 , \10610 );
buf \U$9926 ( \10612 , \10611 );
nand \U$9927 ( \10613 , \10585 , \4099 );
xnor \U$9928 ( \10614 , \10584 , \10613 );
and \U$9929 ( \10615 , \10192 , \10614 );
not \U$9930 ( \10616 , \10192 );
nand \U$9931 ( \10617 , \10604 , \10596 );
not \U$9932 ( \10618 , \10617 );
not \U$9933 ( \10619 , \10601 );
or \U$9934 ( \10620 , \10618 , \10619 );
or \U$9935 ( \10621 , \10601 , \10617 );
nand \U$9936 ( \10622 , \10620 , \10621 );
and \U$9937 ( \10623 , \10616 , \10622 );
or \U$9938 ( \10624 , \10615 , \10623 );
buf \U$9939 ( \10625 , \10624 );
buf \U$9940 ( \10626 , \4573 );
and \U$9941 ( \10627 , \4571 , \10626 );
buf \U$9942 ( \10628 , \3983 );
nor \U$9943 ( \10629 , \10627 , \10628 );
nand \U$9944 ( \10630 , \3987 , \3927 );
and \U$9945 ( \10631 , \10629 , \10630 );
not \U$9946 ( \10632 , \10629 );
not \U$9947 ( \10633 , \10630 );
and \U$9948 ( \10634 , \10632 , \10633 );
nor \U$9949 ( \10635 , \10631 , \10634 );
not \U$9950 ( \10636 , \10635 );
nor \U$9951 ( \10637 , \10636 , \5948 );
not \U$9952 ( \10638 , \10637 );
nand \U$9953 ( \10639 , \9564 , \9625 );
not \U$9954 ( \10640 , \10639 );
not \U$9955 ( \10641 , \10122 );
not \U$9956 ( \10642 , \10119 );
or \U$9957 ( \10643 , \10641 , \10642 );
nand \U$9958 ( \10644 , \10643 , \9624 );
not \U$9959 ( \10645 , \10644 );
or \U$9960 ( \10646 , \10640 , \10645 );
or \U$9961 ( \10647 , \10644 , \10639 );
nand \U$9962 ( \10648 , \10646 , \10647 );
nand \U$9963 ( \10649 , \10648 , \5948 );
nand \U$9964 ( \10650 , \10638 , \10649 );
buf \U$9965 ( \10651 , \10650 );
not \U$9966 ( \10652 , \10628 );
nand \U$9967 ( \10653 , \10652 , \10626 );
xnor \U$9968 ( \10654 , \4571 , \10653 );
and \U$9969 ( \10655 , \10192 , \10654 );
not \U$9970 ( \10656 , \10192 );
nand \U$9971 ( \10657 , \9624 , \10122 );
not \U$9972 ( \10658 , \10657 );
and \U$9973 ( \10659 , \10119 , \10658 );
not \U$9974 ( \10660 , \10119 );
and \U$9975 ( \10661 , \10660 , \10657 );
nor \U$9976 ( \10662 , \10659 , \10661 );
and \U$9977 ( \10663 , \10656 , \10662 );
or \U$9978 ( \10664 , \10655 , \10663 );
buf \U$9979 ( \10665 , \10664 );
not \U$9980 ( \10666 , \5948 );
nand \U$9981 ( \10667 , \9710 , \10118 );
not \U$9982 ( \10668 , \10667 );
not \U$9983 ( \10669 , \10114 );
not \U$9984 ( \10670 , \10102 );
or \U$9985 ( \10671 , \10669 , \10670 );
not \U$9986 ( \10672 , \10116 );
nand \U$9987 ( \10673 , \10671 , \10672 );
not \U$9988 ( \10674 , \10673 );
or \U$9989 ( \10675 , \10668 , \10674 );
or \U$9990 ( \10676 , \10673 , \10667 );
nand \U$9991 ( \10677 , \10675 , \10676 );
not \U$9992 ( \10678 , \10677 );
or \U$9993 ( \10679 , \10666 , \10678 );
xor \U$9994 ( \10680 , \4252 , \4257 );
xor \U$9995 ( \10681 , \10680 , \4568 );
nand \U$9996 ( \10682 , \10681 , \10192 );
nand \U$9997 ( \10683 , \10679 , \10682 );
buf \U$9998 ( \10684 , \10683 );
not \U$9999 ( \10685 , \5948 );
nand \U$10000 ( \10686 , \10672 , \10114 );
not \U$10001 ( \10687 , \10686 );
xor \U$10002 ( \10688 , \10102 , \10687 );
not \U$10003 ( \10689 , \10688 );
or \U$10004 ( \10690 , \10685 , \10689 );
xor \U$10005 ( \10691 , \4302 , \4304 );
xor \U$10006 ( \10692 , \10691 , \4565 );
nand \U$10007 ( \10693 , \10692 , \10192 );
nand \U$10008 ( \10694 , \10690 , \10693 );
buf \U$10009 ( \10695 , \10694 );
xor \U$10010 ( \10696 , \4340 , \4342 );
xor \U$10011 ( \10697 , \10696 , \4562 );
and \U$10012 ( \10698 , \10192 , \10697 );
not \U$10013 ( \10699 , \10192 );
xor \U$10014 ( \10700 , \9795 , \9829 );
xor \U$10015 ( \10701 , \10700 , \10099 );
and \U$10016 ( \10702 , \10699 , \10701 );
or \U$10017 ( \10703 , \10698 , \10702 );
buf \U$10018 ( \10704 , \10703 );
not \U$10019 ( \10705 , \5948 );
buf \U$10020 ( \10706 , \10094 );
not \U$10021 ( \10707 , \10706 );
nand \U$10022 ( \10708 , \9894 , \10098 );
not \U$10023 ( \10709 , \10708 );
or \U$10024 ( \10710 , \10707 , \10709 );
or \U$10025 ( \10711 , \10706 , \10708 );
nand \U$10026 ( \10712 , \10710 , \10711 );
not \U$10027 ( \10713 , \10712 );
or \U$10028 ( \10714 , \10705 , \10713 );
nand \U$10029 ( \10715 , \4558 , \4561 );
xnor \U$10030 ( \10716 , \10715 , \4546 );
nand \U$10031 ( \10717 , \10716 , \10192 );
nand \U$10032 ( \10718 , \10714 , \10717 );
buf \U$10033 ( \10719 , \10718 );
not \U$10034 ( \10720 , \4416 );
nand \U$10035 ( \10721 , \10720 , \4545 );
xor \U$10036 ( \10722 , \10721 , \4543 );
not \U$10037 ( \10723 , \10722 );
nor \U$10038 ( \10724 , \10723 , \5948 );
not \U$10039 ( \10725 , \10724 );
and \U$10040 ( \10726 , \10093 , \9943 );
and \U$10041 ( \10727 , \10726 , \10088 );
not \U$10042 ( \10728 , \10726 );
not \U$10043 ( \10729 , \10088 );
and \U$10044 ( \10730 , \10728 , \10729 );
nor \U$10045 ( \10731 , \10727 , \10730 );
nand \U$10046 ( \10732 , \10731 , \5948 );
nand \U$10047 ( \10733 , \10725 , \10732 );
buf \U$10048 ( \10734 , \10733 );
nor \U$10049 ( \10735 , RI9921f28_596, RI99222e8_588, RI9922090_593);
nor \U$10050 ( \10736 , RI99221f8_590, RI9922180_591);
nor \U$10051 ( \10737 , RI9922018_594, RI9921fa0_595);
nor \U$10052 ( \10738 , RI9922270_589, RI9922108_592);
nand \U$10053 ( \10739 , \10735 , \10736 , \10737 , \10738 );
not \U$10054 ( \10740 , \10739 );
and \U$10055 ( \10741 , RI9921eb0_597, RI9921e38_598, RI9921dc0_599);
not \U$10056 ( \10742 , RI9921d48_600);
nor \U$10057 ( \10743 , \10741 , \10742 );
and \U$10058 ( \10744 , \10740 , \10743 );
not \U$10059 ( \10745 , \10744 );
not \U$10060 ( \10746 , RI9921dc0_599);
not \U$10061 ( \10747 , \10746 );
and \U$10062 ( \10748 , \10745 , \10747 );
and \U$10063 ( \10749 , \10744 , \10746 );
nor \U$10064 ( \10750 , \10748 , \10749 );
not \U$10065 ( \10751 , \10750 );
not \U$10066 ( \10752 , \10751 );
nand \U$10067 ( \10753 , RI9921eb0_597, RI9921e38_598, RI9921dc0_599, RI9921d48_600);
nand \U$10068 ( \10754 , \10740 , \10753 );
and \U$10069 ( \10755 , \10754 , \10742 );
not \U$10070 ( \10756 , \10754 );
and \U$10071 ( \10757 , \10756 , RI9921d48_600);
nor \U$10072 ( \10758 , \10755 , \10757 );
buf \U$10073 ( \10759 , \10758 );
and \U$10074 ( \10760 , \10752 , \10759 );
not \U$10075 ( \10761 , RI9921e38_598);
not \U$10076 ( \10762 , RI9921dc0_599);
nor \U$10077 ( \10763 , \10762 , RI9921f28_596);
nor \U$10078 ( \10764 , RI9922018_594, RI9921fa0_595);
nor \U$10079 ( \10765 , RI9922108_592, RI9922090_593);
and \U$10080 ( \10766 , \10763 , \10764 , \10765 );
nor \U$10081 ( \10767 , RI99222e8_588, RI9922270_589);
and \U$10082 ( \10768 , \10736 , \10767 );
nand \U$10083 ( \10769 , \10766 , \10753 , \10768 , RI9921d48_600);
not \U$10084 ( \10770 , \10769 );
not \U$10085 ( \10771 , \10770 );
or \U$10086 ( \10772 , \10761 , \10771 );
not \U$10087 ( \10773 , RI9921eb0_597);
nand \U$10088 ( \10774 , \10772 , \10773 );
not \U$10089 ( \10775 , \10774 );
not \U$10090 ( \10776 , \10775 );
not \U$10091 ( \10777 , \10769 );
not \U$10092 ( \10778 , \10777 );
not \U$10093 ( \10779 , RI9921e38_598);
not \U$10094 ( \10780 , \10779 );
and \U$10095 ( \10781 , \10778 , \10780 );
and \U$10096 ( \10782 , \10770 , \10779 );
nor \U$10097 ( \10783 , \10781 , \10782 );
nand \U$10098 ( \10784 , \10776 , \10783 );
not \U$10099 ( \10785 , \10784 );
nand \U$10100 ( \10786 , \10760 , \10785 );
buf \U$10101 ( \10787 , \10786 );
buf \U$10102 ( \10788 , \10787 );
nor \U$10103 ( \10789 , \10788 , \5304 );
not \U$10104 ( \10790 , \10750 );
not \U$10105 ( \10791 , \10759 );
and \U$10106 ( \10792 , \10790 , \10791 );
nand \U$10107 ( \10793 , \10792 , \10785 );
buf \U$10108 ( \10794 , \10793 );
nor \U$10109 ( \10795 , \10794 , \5277 );
nor \U$10110 ( \10796 , \10789 , \10795 );
not \U$10111 ( \10797 , RI9808a98_80);
not \U$10112 ( \10798 , \10783 );
not \U$10113 ( \10799 , \10774 );
nand \U$10114 ( \10800 , \10798 , \10799 );
not \U$10115 ( \10801 , \10800 );
not \U$10116 ( \10802 , \10750 );
nor \U$10117 ( \10803 , \10802 , \10759 );
nand \U$10118 ( \10804 , \10801 , \10803 );
not \U$10119 ( \10805 , \10804 );
not \U$10120 ( \10806 , \10805 );
nor \U$10121 ( \10807 , \10797 , \10806 );
and \U$10122 ( \10808 , \10750 , \10791 );
not \U$10123 ( \10809 , \10784 );
nand \U$10124 ( \10810 , \10808 , \10809 );
not \U$10125 ( \10811 , \10810 );
not \U$10126 ( \10812 , \10811 );
nor \U$10127 ( \10813 , \10812 , \5293 );
nor \U$10128 ( \10814 , \10807 , \10813 );
nand \U$10129 ( \10815 , \10796 , \10814 );
not \U$10130 ( \10816 , \10759 );
nor \U$10131 ( \10817 , \10802 , \10816 );
not \U$10132 ( \10818 , \10774 );
nor \U$10133 ( \10819 , \10818 , \10783 );
buf \U$10134 ( \10820 , \10819 );
nand \U$10135 ( \10821 , \10817 , \10820 );
not \U$10136 ( \10822 , \10821 );
not \U$10137 ( \10823 , \10822 );
nor \U$10138 ( \10824 , \10823 , \815 );
and \U$10139 ( \10825 , \10751 , \10791 );
nand \U$10140 ( \10826 , \10825 , \10820 );
not \U$10141 ( \10827 , \10826 );
not \U$10142 ( \10828 , \10827 );
buf \U$10143 ( \10829 , \10828 );
nor \U$10144 ( \10830 , \10829 , \5301 );
nor \U$10145 ( \10831 , \10824 , \10830 );
and \U$10146 ( \10832 , \10790 , \10759 );
nand \U$10147 ( \10833 , \10832 , \10820 );
not \U$10148 ( \10834 , \10833 );
and \U$10149 ( \10835 , \10834 , RI9967078_223);
and \U$10150 ( \10836 , RI995e450_236, RI9921f28_596);
nor \U$10151 ( \10837 , \10835 , \10836 );
nand \U$10152 ( \10838 , \10799 , \10783 );
not \U$10153 ( \10839 , \10838 );
not \U$10154 ( \10840 , RI9921f28_596);
nand \U$10155 ( \10841 , \10808 , \10839 , \10840 );
not \U$10156 ( \10842 , \10841 );
buf \U$10157 ( \10843 , \10842 );
nand \U$10158 ( \10844 , \10843 , RI994ddd0_28);
nand \U$10159 ( \10845 , \10831 , \10837 , \10844 );
nor \U$10160 ( \10846 , \10815 , \10845 );
nand \U$10161 ( \10847 , \10817 , \10839 );
not \U$10162 ( \10848 , \10847 );
not \U$10163 ( \10849 , \10848 );
not \U$10164 ( \10850 , \10849 );
not \U$10165 ( \10851 , RI98bc8d0_41);
not \U$10166 ( \10852 , \10851 );
and \U$10167 ( \10853 , \10850 , \10852 );
not \U$10168 ( \10854 , \10800 );
nand \U$10169 ( \10855 , \10832 , \10854 );
not \U$10170 ( \10856 , \10855 );
not \U$10171 ( \10857 , \10856 );
not \U$10172 ( \10858 , \10857 );
and \U$10173 ( \10859 , \10858 , RI89ec640_119);
nor \U$10174 ( \10860 , \10853 , \10859 );
nand \U$10175 ( \10861 , \10820 , \10803 );
buf \U$10176 ( \10862 , \10861 );
not \U$10177 ( \10863 , \10862 );
not \U$10178 ( \10864 , \5291 );
and \U$10179 ( \10865 , \10863 , \10864 );
and \U$10180 ( \10866 , \10790 , \10759 );
nand \U$10181 ( \10867 , \10866 , \10785 );
not \U$10182 ( \10868 , \10867 );
and \U$10183 ( \10869 , \10868 , RI89253b0_171);
nor \U$10184 ( \10870 , \10865 , \10869 );
nand \U$10185 ( \10871 , \10860 , \10870 );
nand \U$10186 ( \10872 , \10760 , \10854 );
not \U$10187 ( \10873 , \10872 );
not \U$10188 ( \10874 , \10873 );
not \U$10189 ( \10875 , \10874 );
not \U$10190 ( \10876 , \5317 );
and \U$10191 ( \10877 , \10875 , \10876 );
nand \U$10192 ( \10878 , \10825 , \10854 );
not \U$10193 ( \10879 , \10878 );
not \U$10194 ( \10880 , \10879 );
nor \U$10195 ( \10881 , \10880 , \829 );
nor \U$10196 ( \10882 , \10877 , \10881 );
nand \U$10197 ( \10883 , \10832 , \10839 );
not \U$10198 ( \10884 , \10883 );
not \U$10199 ( \10885 , \10884 );
nor \U$10200 ( \10886 , \10885 , \5311 );
not \U$10201 ( \10887 , RI98abc38_54);
nand \U$10202 ( \10888 , \10792 , \10839 );
buf \U$10203 ( \10889 , \10888 );
nor \U$10204 ( \10890 , \10887 , \10889 );
nor \U$10205 ( \10891 , \10886 , \10890 );
nand \U$10206 ( \10892 , \10882 , \10891 );
nor \U$10207 ( \10893 , \10871 , \10892 );
nand \U$10208 ( \10894 , \10846 , \10893 );
not \U$10209 ( \10895 , RI995ef90_4);
not \U$10210 ( \10896 , RI995ecc0_10);
nand \U$10211 ( \10897 , RI995ec48_11, RI995ebd0_12);
nor \U$10212 ( \10898 , \10896 , \10897 );
nand \U$10213 ( \10899 , \10898 , RI995ed38_9);
not \U$10214 ( \10900 , RI995edb0_8);
nor \U$10215 ( \10901 , \10899 , \10900 );
nand \U$10216 ( \10902 , \10901 , RI995ee28_7);
not \U$10217 ( \10903 , \10902 );
nand \U$10218 ( \10904 , \10903 , RI995eea0_6);
not \U$10219 ( \10905 , \10904 );
nand \U$10220 ( \10906 , \10905 , RI995ef18_5);
nor \U$10221 ( \10907 , \10895 , \10906 );
nand \U$10222 ( \10908 , \10907 , RI995f008_3);
xor \U$10223 ( \10909 , \10908 , RI995f080_2);
nand \U$10224 ( \10910 , \10894 , \10909 );
and \U$10225 ( \10911 , \10834 , RI995e900_226);
and \U$10226 ( \10912 , RI9959f68_239, RI9921f28_596);
nor \U$10227 ( \10913 , \10911 , \10912 );
nand \U$10228 ( \10914 , \10842 , RI994dc68_31);
not \U$10229 ( \10915 , \10828 );
nand \U$10230 ( \10916 , \10915 , RI9967528_213);
buf \U$10231 ( \10917 , \10752 );
buf \U$10232 ( \10918 , \10783 );
and \U$10233 ( \10919 , \10917 , \10918 , \10775 , \10759 );
not \U$10234 ( \10920 , \10919 );
not \U$10235 ( \10921 , \10920 );
nand \U$10236 ( \10922 , \10921 , RI98bc768_44);
and \U$10237 ( \10923 , \10913 , \10914 , \10916 , \10922 );
not \U$10238 ( \10924 , RI8946470_135);
or \U$10239 ( \10925 , \10812 , \10924 );
not \U$10240 ( \10926 , RI9808930_83);
or \U$10241 ( \10927 , \10806 , \10926 );
nand \U$10242 ( \10928 , \10925 , \10927 );
not \U$10243 ( \10929 , RI8939c48_148);
and \U$10244 ( \10930 , \10817 , \10785 );
buf \U$10245 ( \10931 , \10930 );
not \U$10246 ( \10932 , \10931 );
or \U$10247 ( \10933 , \10929 , \10932 );
and \U$10248 ( \10934 , \10792 , \10785 );
not \U$10249 ( \10935 , \10934 );
not \U$10250 ( \10936 , \10935 );
nand \U$10251 ( \10937 , \10936 , RI8930c60_161);
nand \U$10252 ( \10938 , \10933 , \10937 );
nor \U$10253 ( \10939 , \10928 , \10938 );
not \U$10254 ( \10940 , RI9808318_96);
not \U$10255 ( \10941 , \10873 );
or \U$10256 ( \10942 , \10940 , \10941 );
nand \U$10257 ( \10943 , \10879 , RI9776e18_109);
nand \U$10258 ( \10944 , \10942 , \10943 );
not \U$10259 ( \10945 , RI890fa38_200);
not \U$10260 ( \10946 , \10822 );
or \U$10261 ( \10947 , \10945 , \10946 );
nand \U$10262 ( \10948 , \10884 , RI98195c8_70);
nand \U$10263 ( \10949 , \10947 , \10948 );
nor \U$10264 ( \10950 , \10944 , \10949 );
not \U$10265 ( \10951 , RI8925248_174);
not \U$10266 ( \10952 , \10868 );
or \U$10267 ( \10953 , \10951 , \10952 );
and \U$10268 ( \10954 , \10808 , \10820 );
buf \U$10269 ( \10955 , \10954 );
nand \U$10270 ( \10956 , \10955 , RI8918a20_187);
nand \U$10271 ( \10957 , \10953 , \10956 );
not \U$10272 ( \10958 , RI89ec4d8_122);
not \U$10273 ( \10959 , \10856 );
or \U$10274 ( \10960 , \10958 , \10959 );
not \U$10275 ( \10961 , \10792 );
nor \U$10276 ( \10962 , \10961 , \10838 );
buf \U$10277 ( \10963 , \10962 );
nand \U$10278 ( \10964 , \10963 , RI98abad0_57);
nand \U$10279 ( \10965 , \10960 , \10964 );
nor \U$10280 ( \10966 , \10957 , \10965 );
nand \U$10281 ( \10967 , \10923 , \10939 , \10950 , \10966 );
buf \U$10282 ( \10968 , \10967 );
not \U$10283 ( \10969 , \10904 );
not \U$10284 ( \10970 , RI995ef18_5);
and \U$10285 ( \10971 , \10969 , \10970 );
and \U$10286 ( \10972 , \10904 , RI995ef18_5);
nor \U$10287 ( \10973 , \10971 , \10972 );
nand \U$10288 ( \10974 , \10968 , \10973 );
buf \U$10289 ( \10975 , \10826 );
not \U$10290 ( \10976 , \10975 );
not \U$10291 ( \10977 , RI99675a0_212);
not \U$10292 ( \10978 , \10977 );
and \U$10293 ( \10979 , \10976 , \10978 );
and \U$10294 ( \10980 , \10884 , RI9819640_69);
nor \U$10295 ( \10981 , \10979 , \10980 );
and \U$10296 ( \10982 , \10834 , RI995e978_225);
nand \U$10297 ( \10983 , RI9959fe0_238, RI9921f28_596);
not \U$10298 ( \10984 , \10983 );
nor \U$10299 ( \10985 , \10982 , \10984 );
nand \U$10300 ( \10986 , \10842 , RI994dce0_30);
nand \U$10301 ( \10987 , \10981 , \10985 , \10986 );
nand \U$10302 ( \10988 , \10805 , RI98089a8_82);
nand \U$10303 ( \10989 , \10811 , RI89464e8_134);
nand \U$10304 ( \10990 , \10931 , RI8939cc0_147);
nand \U$10305 ( \10991 , \10934 , RI8930cd8_160);
nand \U$10306 ( \10992 , \10988 , \10989 , \10990 , \10991 );
nor \U$10307 ( \10993 , \10987 , \10992 );
nand \U$10308 ( \10994 , \10955 , RI8918a98_186);
nand \U$10309 ( \10995 , \10856 , RI89ec550_121);
nand \U$10310 ( \10996 , \10919 , RI98bc7e0_43);
nand \U$10311 ( \10997 , \10868 , RI89252c0_173);
nand \U$10312 ( \10998 , \10994 , \10995 , \10996 , \10997 );
nand \U$10313 ( \10999 , \10873 , RI9808390_95);
nand \U$10314 ( \11000 , \10822 , RI890fab0_199);
not \U$10315 ( \11001 , \10878 );
nand \U$10316 ( \11002 , \11001 , RI9776e90_108);
nand \U$10317 ( \11003 , \10963 , RI98abb48_56);
nand \U$10318 ( \11004 , \10999 , \11000 , \11002 , \11003 );
nor \U$10319 ( \11005 , \10998 , \11004 );
nand \U$10320 ( \11006 , \10993 , \11005 );
not \U$10321 ( \11007 , \11006 );
not \U$10322 ( \11008 , \10906 );
not \U$10323 ( \11009 , RI995ef90_4);
and \U$10324 ( \11010 , \11008 , \11009 );
and \U$10325 ( \11011 , \10906 , RI995ef90_4);
nor \U$10326 ( \11012 , \11010 , \11011 );
not \U$10327 ( \11013 , \11012 );
nor \U$10328 ( \11014 , \11007 , \11013 );
not \U$10329 ( \11015 , \11014 );
not \U$10330 ( \11016 , \10829 );
not \U$10331 ( \11017 , RI9967618_211);
not \U$10332 ( \11018 , \11017 );
and \U$10333 ( \11019 , \11016 , \11018 );
and \U$10334 ( \11020 , \10856 , RI89ec5c8_120);
nor \U$10335 ( \11021 , \11019 , \11020 );
and \U$10336 ( \11022 , \10834 , RI99669e8_224);
nand \U$10337 ( \11023 , RI995e3d8_237, RI9921f28_596);
not \U$10338 ( \11024 , \11023 );
nor \U$10339 ( \11025 , \11022 , \11024 );
nand \U$10340 ( \11026 , \10843 , RI994dd58_29);
nand \U$10341 ( \11027 , \11021 , \11025 , \11026 );
not \U$10342 ( \11028 , \10812 );
nand \U$10343 ( \11029 , \11028 , RI8946560_133);
buf \U$10344 ( \11030 , \10963 );
nand \U$10345 ( \11031 , \11030 , RI98abbc0_55);
not \U$10346 ( \11032 , \10806 );
nand \U$10347 ( \11033 , \11032 , RI9808a20_81);
nand \U$10348 ( \11034 , \10921 , RI98bc858_42);
nand \U$10349 ( \11035 , \11029 , \11031 , \11033 , \11034 );
nor \U$10350 ( \11036 , \11027 , \11035 );
nand \U$10351 ( \11037 , \10822 , RI890fb28_198);
nand \U$10352 ( \11038 , \10873 , RI9808408_94);
not \U$10353 ( \11039 , \10880 );
nand \U$10354 ( \11040 , \11039 , RI9776f08_107);
nand \U$10355 ( \11041 , \10955 , RI8918b10_185);
nand \U$10356 ( \11042 , \11037 , \11038 , \11040 , \11041 );
nand \U$10357 ( \11043 , \10868 , RI8925338_172);
nand \U$10358 ( \11044 , \10931 , RI8939d38_146);
nand \U$10359 ( \11045 , \10884 , RI98196b8_68);
nand \U$10360 ( \11046 , \10936 , RI8930d50_159);
nand \U$10361 ( \11047 , \11043 , \11044 , \11045 , \11046 );
nor \U$10362 ( \11048 , \11042 , \11047 );
nand \U$10363 ( \11049 , \11036 , \11048 );
xnor \U$10364 ( \11050 , \10907 , RI995f008_3);
nand \U$10365 ( \11051 , \11049 , \11050 );
and \U$10366 ( \11052 , \10910 , \10974 , \11015 , \11051 );
not \U$10367 ( \11053 , \11052 );
not \U$10368 ( \11054 , RI89ec820_115);
not \U$10369 ( \11055 , \11001 );
or \U$10370 ( \11056 , \11054 , \11055 );
not \U$10371 ( \11057 , \10883 );
nand \U$10372 ( \11058 , \11057 , RI98192f8_76);
nand \U$10373 ( \11059 , \11056 , \11058 );
not \U$10374 ( \11060 , RI98ab800_63);
or \U$10375 ( \11061 , \10889 , \11060 );
not \U$10376 ( \11062 , RI98abe18_50);
or \U$10377 ( \11063 , \11062 , \10847 );
nand \U$10378 ( \11064 , \11061 , \11063 );
nor \U$10379 ( \11065 , \11059 , \11064 );
not \U$10380 ( \11066 , RI8939978_154);
not \U$10381 ( \11067 , \10930 );
or \U$10382 ( \11068 , \11066 , \11067 );
nand \U$10383 ( \11069 , \10856 , RI89ec208_128);
nand \U$10384 ( \11070 , \11068 , \11069 );
not \U$10385 ( \11071 , RI8930990_167);
or \U$10386 ( \11072 , \10794 , \11071 );
not \U$10387 ( \11073 , RI9967258_219);
or \U$10388 ( \11074 , \10975 , \11073 );
nand \U$10389 ( \11075 , \11072 , \11074 );
nor \U$10390 ( \11076 , \11070 , \11075 );
not \U$10391 ( \11077 , \10804 );
not \U$10392 ( \11078 , RI9808660_89);
not \U$10393 ( \11079 , \11078 );
and \U$10394 ( \11080 , \11077 , \11079 );
and \U$10395 ( \11081 , \10822 , RI890f768_206);
nor \U$10396 ( \11082 , \11080 , \11081 );
not \U$10397 ( \11083 , \10833 );
and \U$10398 ( \11084 , \11083 , RI995e630_232);
and \U$10399 ( \11085 , RI994d7b8_245, RI9921f28_596);
nor \U$10400 ( \11086 , \11084 , \11085 );
nand \U$10401 ( \11087 , \10842 , RI98bcab0_37);
and \U$10402 ( \11088 , \11082 , \11086 , \11087 );
not \U$10403 ( \11089 , RI9777160_102);
not \U$10404 ( \11090 , \10873 );
or \U$10405 ( \11091 , \11089 , \11090 );
not \U$10406 ( \11092 , \10867 );
nand \U$10407 ( \11093 , \11092 , RI8924f78_180);
nand \U$10408 ( \11094 , \11091 , \11093 );
not \U$10409 ( \11095 , RI8918750_193);
not \U$10410 ( \11096 , \10954 );
or \U$10411 ( \11097 , \11095 , \11096 );
nand \U$10412 ( \11098 , \10811 , RI89461a0_141);
nand \U$10413 ( \11099 , \11097 , \11098 );
nor \U$10414 ( \11100 , \11094 , \11099 );
nand \U$10415 ( \11101 , \11065 , \11076 , \11088 , \11100 );
not \U$10416 ( \11102 , RI995ebd0_12);
and \U$10417 ( \11103 , RI995ec48_11, \11102 );
not \U$10418 ( \11104 , RI995ec48_11);
and \U$10419 ( \11105 , \11104 , RI995ebd0_12);
nor \U$10420 ( \11106 , \11103 , \11105 );
nand \U$10421 ( \11107 , \11101 , \11106 );
not \U$10422 ( \11108 , \11107 );
nand \U$10423 ( \11109 , \10825 , \10820 );
not \U$10424 ( \11110 , \11109 );
not \U$10425 ( \11111 , \1140 );
and \U$10426 ( \11112 , \11110 , \11111 );
not \U$10427 ( \11113 , \10800 );
and \U$10428 ( \11114 , \11113 , \10817 );
and \U$10429 ( \11115 , \11114 , RI97770e8_103);
nor \U$10430 ( \11116 , \11112 , \11115 );
and \U$10431 ( \11117 , \10840 , \10839 , \10803 );
nand \U$10432 ( \11118 , \11117 , RI98bca38_38);
and \U$10433 ( \11119 , \11116 , \11118 );
not \U$10434 ( \11120 , \10786 );
not \U$10435 ( \11121 , RI8939900_155);
not \U$10436 ( \11122 , \11121 );
and \U$10437 ( \11123 , \11120 , \11122 );
nand \U$10438 ( \11124 , \10832 , \11113 );
not \U$10439 ( \11125 , \11124 );
and \U$10440 ( \11126 , \11125 , RI89ec190_129);
nor \U$10441 ( \11127 , \11123 , \11126 );
nand \U$10442 ( \11128 , \10808 , \10809 );
not \U$10443 ( \11129 , \11128 );
not \U$10444 ( \11130 , RI8946128_142);
not \U$10445 ( \11131 , \11130 );
and \U$10446 ( \11132 , \11129 , \11131 );
nand \U$10447 ( \11133 , \10866 , \10839 );
not \U$10448 ( \11134 , \11133 );
and \U$10449 ( \11135 , \11134 , RI9819280_77);
nor \U$10450 ( \11136 , \11132 , \11135 );
and \U$10451 ( \11137 , \11127 , \11136 );
nand \U$10452 ( \11138 , \10760 , \10820 );
not \U$10453 ( \11139 , \11138 );
not \U$10454 ( \11140 , RI890f6f0_207);
not \U$10455 ( \11141 , \11140 );
and \U$10456 ( \11142 , \11139 , \11141 );
nand \U$10457 ( \11143 , \10825 , \11113 );
not \U$10458 ( \11144 , \11143 );
and \U$10459 ( \11145 , \11144 , RI89ec7a8_116);
nor \U$10460 ( \11146 , \11142 , \11145 );
nand \U$10461 ( \11147 , \10866 , \10820 );
not \U$10462 ( \11148 , \11147 );
and \U$10463 ( \11149 , \11148 , RI995e5b8_233);
nand \U$10464 ( \11150 , RI994d740_246, RI9921f28_596);
not \U$10465 ( \11151 , \11150 );
nor \U$10466 ( \11152 , \11149 , \11151 );
not \U$10467 ( \11153 , \10804 );
not \U$10468 ( \11154 , RI98085e8_90);
not \U$10469 ( \11155 , \11154 );
and \U$10470 ( \11156 , \11153 , \11155 );
not \U$10471 ( \11157 , RI89186d8_194);
nor \U$10472 ( \11158 , \11157 , \10861 );
nor \U$10473 ( \11159 , \11156 , \11158 );
and \U$10474 ( \11160 , \11146 , \11152 , \11159 );
nand \U$10475 ( \11161 , \10866 , \10809 );
not \U$10476 ( \11162 , \11161 );
not \U$10477 ( \11163 , RI8924f00_181);
not \U$10478 ( \11164 , \11163 );
and \U$10479 ( \11165 , \11162 , \11164 );
not \U$10480 ( \11166 , RI8930918_168);
nor \U$10481 ( \11167 , \10793 , \11166 );
nor \U$10482 ( \11168 , \11165 , \11167 );
not \U$10483 ( \11169 , \10888 );
not \U$10484 ( \11170 , RI98ab788_64);
not \U$10485 ( \11171 , \11170 );
and \U$10486 ( \11172 , \11169 , \11171 );
not \U$10487 ( \11173 , RI98abda0_51);
nor \U$10488 ( \11174 , \11173 , \10847 );
nor \U$10489 ( \11175 , \11172 , \11174 );
and \U$10490 ( \11176 , \11168 , \11175 );
nand \U$10491 ( \11177 , \11119 , \11137 , \11160 , \11176 );
nand \U$10492 ( \11178 , \11177 , RI995ebd0_12);
not \U$10493 ( \11179 , \11178 );
not \U$10494 ( \11180 , RI995e540_234);
not \U$10495 ( \11181 , \11148 );
or \U$10496 ( \11182 , \11180 , \11181 );
nand \U$10497 ( \11183 , RI994d6c8_247, RI9921f28_596);
nand \U$10498 ( \11184 , \11182 , \11183 );
and \U$10499 ( \11185 , \11117 , RI98bc9c0_39);
nor \U$10500 ( \11186 , \11184 , \11185 );
not \U$10501 ( \11187 , RI8939888_156);
nor \U$10502 ( \11188 , \11187 , \10786 );
not \U$10503 ( \11189 , RI89308a0_169);
nor \U$10504 ( \11190 , \10793 , \11189 );
nor \U$10505 ( \11191 , \11188 , \11190 );
not \U$10506 ( \11192 , \10805 );
not \U$10507 ( \11193 , \11192 );
not \U$10508 ( \11194 , RI9808570_91);
not \U$10509 ( \11195 , \11194 );
and \U$10510 ( \11196 , \11193 , \11195 );
and \U$10511 ( \11197 , \10963 , RI98ab710_65);
nor \U$10512 ( \11198 , \11196 , \11197 );
not \U$10513 ( \11199 , RI9819208_78);
nor \U$10514 ( \11200 , \11199 , \11133 );
not \U$10515 ( \11201 , RI8924e88_182);
nor \U$10516 ( \11202 , \11201 , \11161 );
nor \U$10517 ( \11203 , \11200 , \11202 );
nand \U$10518 ( \11204 , \11186 , \11191 , \11198 , \11203 );
not \U$10519 ( \11205 , \11138 );
not \U$10520 ( \11206 , RI890f678_208);
not \U$10521 ( \11207 , \11206 );
and \U$10522 ( \11208 , \11205 , \11207 );
not \U$10523 ( \11209 , RI8918660_195);
nor \U$10524 ( \11210 , \10861 , \11209 );
nor \U$10525 ( \11211 , \11208 , \11210 );
not \U$10526 ( \11212 , RI89ec118_130);
nor \U$10527 ( \11213 , \11212 , \11124 );
not \U$10528 ( \11214 , RI89ec730_117);
nor \U$10529 ( \11215 , \11214 , \11143 );
nor \U$10530 ( \11216 , \11213 , \11215 );
not \U$10531 ( \11217 , \11128 );
not \U$10532 ( \11218 , RI89460b0_143);
not \U$10533 ( \11219 , \11218 );
and \U$10534 ( \11220 , \11217 , \11219 );
and \U$10535 ( \11221 , \10919 , RI98abd28_52);
nor \U$10536 ( \11222 , \11220 , \11221 );
not \U$10537 ( \11223 , \11109 );
not \U$10538 ( \11224 , RI9967168_221);
not \U$10539 ( \11225 , \11224 );
and \U$10540 ( \11226 , \11223 , \11225 );
and \U$10541 ( \11227 , \11114 , RI9777070_104);
nor \U$10542 ( \11228 , \11226 , \11227 );
nand \U$10543 ( \11229 , \11211 , \11216 , \11222 , \11228 );
or \U$10544 ( \11230 , \11204 , \11229 );
not \U$10545 ( \11231 , RI994e4d8_13);
nand \U$10546 ( \11232 , \11230 , \11231 );
not \U$10547 ( \11233 , \11232 );
or \U$10548 ( \11234 , \11179 , \11233 );
and \U$10549 ( \11235 , \11146 , \11127 );
and \U$10550 ( \11236 , \11116 , \11152 , \11118 );
not \U$10551 ( \11237 , \11136 );
not \U$10552 ( \11238 , \11159 );
nor \U$10553 ( \11239 , \11237 , \11238 );
nand \U$10554 ( \11240 , \11235 , \11176 , \11236 , \11239 );
not \U$10555 ( \11241 , \11240 );
nand \U$10556 ( \11242 , \11241 , \11102 );
nand \U$10557 ( \11243 , \11234 , \11242 );
not \U$10558 ( \11244 , \11243 );
or \U$10559 ( \11245 , \11108 , \11244 );
not \U$10560 ( \11246 , \11101 );
not \U$10561 ( \11247 , \11106 );
and \U$10562 ( \11248 , \11246 , \11247 );
not \U$10563 ( \11249 , \11248 );
nand \U$10564 ( \11250 , \11245 , \11249 );
not \U$10565 ( \11251 , \11250 );
not \U$10566 ( \11252 , RI8939a68_152);
nor \U$10567 ( \11253 , \11252 , \10787 );
nor \U$10568 ( \11254 , \10793 , \5468 );
nor \U$10569 ( \11255 , \11253 , \11254 );
not \U$10570 ( \11256 , \10804 );
not \U$10571 ( \11257 , \5489 );
and \U$10572 ( \11258 , \11256 , \11257 );
not \U$10573 ( \11259 , RI8946290_139);
nor \U$10574 ( \11260 , \11259 , \11128 );
nor \U$10575 ( \11261 , \11258 , \11260 );
nand \U$10576 ( \11262 , \11255 , \11261 );
not \U$10577 ( \11263 , \10826 );
not \U$10578 ( \11264 , RI9967348_217);
not \U$10579 ( \11265 , \11264 );
and \U$10580 ( \11266 , \11263 , \11265 );
and \U$10581 ( \11267 , \10873 , RI9777250_100);
nor \U$10582 ( \11268 , \11266 , \11267 );
not \U$10583 ( \11269 , RI8918840_191);
nor \U$10584 ( \11270 , \11269 , \10862 );
not \U$10585 ( \11271 , RI890f858_204);
nor \U$10586 ( \11272 , \11271 , \10821 );
nor \U$10587 ( \11273 , \11270 , \11272 );
nand \U$10588 ( \11274 , \11268 , \11273 );
nor \U$10589 ( \11275 , \11262 , \11274 );
not \U$10590 ( \11276 , \11275 );
not \U$10591 ( \11277 , \10847 );
not \U$10592 ( \11278 , RI98abf08_48);
not \U$10593 ( \11279 , \11278 );
and \U$10594 ( \11280 , \11277 , \11279 );
and \U$10595 ( \11281 , \10879 , RI89ec910_113);
nor \U$10596 ( \11282 , \11280 , \11281 );
not \U$10597 ( \11283 , RI98ab8f0_61);
nor \U$10598 ( \11284 , \11283 , \10889 );
not \U$10599 ( \11285 , RI89ec2f8_126);
nor \U$10600 ( \11286 , \11285 , \10855 );
nor \U$10601 ( \11287 , \11284 , \11286 );
nand \U$10602 ( \11288 , \11282 , \11287 );
not \U$10603 ( \11289 , RI995e720_230);
not \U$10604 ( \11290 , \11083 );
or \U$10605 ( \11291 , \11289 , \11290 );
nand \U$10606 ( \11292 , RI994d8a8_243, RI9921f28_596);
nand \U$10607 ( \11293 , \11291 , \11292 );
not \U$10608 ( \11294 , \11293 );
nand \U$10609 ( \11295 , \11134 , RI98193e8_74);
not \U$10610 ( \11296 , \10867 );
nand \U$10611 ( \11297 , \11296 , RI8925068_178);
and \U$10612 ( \11298 , \11295 , \11297 );
nand \U$10613 ( \11299 , \10842 , RI98bcba0_35);
nand \U$10614 ( \11300 , \11294 , \11298 , \11299 );
nor \U$10615 ( \11301 , \11288 , \11300 );
not \U$10616 ( \11302 , \11301 );
or \U$10617 ( \11303 , \11276 , \11302 );
not \U$10618 ( \11304 , RI995ed38_9);
and \U$10619 ( \11305 , \10898 , \11304 );
not \U$10620 ( \11306 , \10898 );
and \U$10621 ( \11307 , \11306 , RI995ed38_9);
nor \U$10622 ( \11308 , \11305 , \11307 );
nand \U$10623 ( \11309 , \11303 , \11308 );
nand \U$10624 ( \11310 , \10827 , RI99673c0_216);
nand \U$10625 ( \11311 , \10934 , RI8930af8_164);
nand \U$10626 ( \11312 , \10930 , RI8939ae0_151);
nand \U$10627 ( \11313 , \10822 , RI890f8d0_203);
and \U$10628 ( \11314 , \11310 , \11311 , \11312 , \11313 );
nand \U$10629 ( \11315 , \10811 , RI8946308_138);
nand \U$10630 ( \11316 , \11148 , RI995e798_229);
nand \U$10631 ( \11317 , RI994d920_242, RI9921f28_596);
nand \U$10632 ( \11318 , \11315 , \11316 , \11317 );
not \U$10633 ( \11319 , RI97772c8_99);
not \U$10634 ( \11320 , \10873 );
or \U$10635 ( \11321 , \11319 , \11320 );
nand \U$10636 ( \11322 , \11057 , RI9819460_73);
nand \U$10637 ( \11323 , \11321 , \11322 );
nor \U$10638 ( \11324 , \11318 , \11323 );
not \U$10639 ( \11325 , RI98abf80_47);
not \U$10640 ( \11326 , \10919 );
or \U$10641 ( \11327 , \11325 , \11326 );
nand \U$10642 ( \11328 , \10963 , RI98ab968_60);
nand \U$10643 ( \11329 , \11327 , \11328 );
not \U$10644 ( \11330 , RI89ec370_125);
not \U$10645 ( \11331 , \10856 );
or \U$10646 ( \11332 , \11330 , \11331 );
nand \U$10647 ( \11333 , \10805 , RI98087c8_86);
nand \U$10648 ( \11334 , \11332 , \11333 );
nor \U$10649 ( \11335 , \11329 , \11334 );
not \U$10650 ( \11336 , RI89250e0_177);
not \U$10651 ( \11337 , \10868 );
or \U$10652 ( \11338 , \11336 , \11337 );
nand \U$10653 ( \11339 , \10954 , RI89188b8_190);
nand \U$10654 ( \11340 , \11338 , \11339 );
not \U$10655 ( \11341 , RI89ec988_112);
not \U$10656 ( \11342 , \10879 );
or \U$10657 ( \11343 , \11341 , \11342 );
nand \U$10658 ( \11344 , \11117 , RI98bcc18_34);
nand \U$10659 ( \11345 , \11343 , \11344 );
nor \U$10660 ( \11346 , \11340 , \11345 );
nand \U$10661 ( \11347 , \11314 , \11324 , \11335 , \11346 );
and \U$10662 ( \11348 , \10899 , \10900 );
not \U$10663 ( \11349 , \10899 );
and \U$10664 ( \11350 , \11349 , RI995edb0_8);
or \U$10665 ( \11351 , \11348 , \11350 );
nand \U$10666 ( \11352 , \11347 , \11351 );
and \U$10667 ( \11353 , \11309 , \11352 );
nand \U$10668 ( \11354 , \10842 , RI98bcc90_33);
nand \U$10669 ( \11355 , \11083 , RI995e810_228);
nand \U$10670 ( \11356 , RI994d998_241, RI9921f28_596);
nand \U$10671 ( \11357 , \11354 , \11355 , \11356 );
not \U$10672 ( \11358 , RI9808228_98);
not \U$10673 ( \11359 , \10873 );
or \U$10674 ( \11360 , \11358 , \11359 );
nand \U$10675 ( \11361 , \10827 , RI9967438_215);
nand \U$10676 ( \11362 , \11360 , \11361 );
nor \U$10677 ( \11363 , \11357 , \11362 );
not \U$10678 ( \11364 , RI8925158_176);
not \U$10679 ( \11365 , \11092 );
or \U$10680 ( \11366 , \11364 , \11365 );
nand \U$10681 ( \11367 , \11057 , RI98194d8_72);
nand \U$10682 ( \11368 , \11366 , \11367 );
not \U$10683 ( \11369 , RI8939b58_150);
not \U$10684 ( \11370 , \10930 );
or \U$10685 ( \11371 , \11369 , \11370 );
nand \U$10686 ( \11372 , \11001 , RI9776d28_111);
nand \U$10687 ( \11373 , \11371 , \11372 );
nor \U$10688 ( \11374 , \11368 , \11373 );
not \U$10689 ( \11375 , RI89ec3e8_124);
not \U$10690 ( \11376 , \10856 );
or \U$10691 ( \11377 , \11375 , \11376 );
nand \U$10692 ( \11378 , \10934 , RI8930b70_163);
nand \U$10693 ( \11379 , \11377 , \11378 );
not \U$10694 ( \11380 , RI890f948_202);
not \U$10695 ( \11381 , \10822 );
or \U$10696 ( \11382 , \11380 , \11381 );
nand \U$10697 ( \11383 , \10954 , RI8918930_189);
nand \U$10698 ( \11384 , \11382 , \11383 );
nor \U$10699 ( \11385 , \11379 , \11384 );
not \U$10700 ( \11386 , RI98ab9e0_59);
or \U$10701 ( \11387 , \10889 , \11386 );
not \U$10702 ( \11388 , RI98abff8_46);
or \U$10703 ( \11389 , \10849 , \11388 );
nand \U$10704 ( \11390 , \11387 , \11389 );
not \U$10705 ( \11391 , \10811 );
not \U$10706 ( \11392 , RI8946380_137);
or \U$10707 ( \11393 , \11391 , \11392 );
not \U$10708 ( \11394 , RI9808840_85);
or \U$10709 ( \11395 , \11192 , \11394 );
nand \U$10710 ( \11396 , \11393 , \11395 );
nor \U$10711 ( \11397 , \11390 , \11396 );
nand \U$10712 ( \11398 , \11363 , \11374 , \11385 , \11397 );
xnor \U$10713 ( \11399 , \10901 , RI995ee28_7);
nand \U$10714 ( \11400 , \11398 , \11399 );
not \U$10715 ( \11401 , RI89251d0_175);
not \U$10716 ( \11402 , \11092 );
or \U$10717 ( \11403 , \11401 , \11402 );
nand \U$10718 ( \11404 , \11057 , RI9819550_71);
nand \U$10719 ( \11405 , \11403 , \11404 );
not \U$10720 ( \11406 , RI98082a0_97);
not \U$10721 ( \11407 , \10873 );
or \U$10722 ( \11408 , \11406 , \11407 );
nand \U$10723 ( \11409 , \10934 , RI8930be8_162);
nand \U$10724 ( \11410 , \11408 , \11409 );
nor \U$10725 ( \11411 , \11405 , \11410 );
nand \U$10726 ( \11412 , \11083 , RI995e888_227);
nand \U$10727 ( \11413 , \10842 , RI994dbf0_32);
nand \U$10728 ( \11414 , RI9959860_240, RI9921f28_596);
nand \U$10729 ( \11415 , \11412 , \11413 , \11414 );
not \U$10730 ( \11416 , RI8939bd0_149);
or \U$10731 ( \11417 , \11416 , \10787 );
not \U$10732 ( \11418 , RI99674b0_214);
or \U$10733 ( \11419 , \10828 , \11418 );
nand \U$10734 ( \11420 , \11417 , \11419 );
nor \U$10735 ( \11421 , \11415 , \11420 );
not \U$10736 ( \11422 , RI9776da0_110);
not \U$10737 ( \11423 , \11001 );
or \U$10738 ( \11424 , \11422 , \11423 );
nand \U$10739 ( \11425 , \10856 , RI89ec460_123);
nand \U$10740 ( \11426 , \11424 , \11425 );
not \U$10741 ( \11427 , RI98bc6f0_45);
not \U$10742 ( \11428 , \10919 );
or \U$10743 ( \11429 , \11427 , \11428 );
nand \U$10744 ( \11430 , \10963 , RI98aba58_58);
nand \U$10745 ( \11431 , \11429 , \11430 );
nor \U$10746 ( \11432 , \11426 , \11431 );
not \U$10747 ( \11433 , RI890f9c0_201);
not \U$10748 ( \11434 , \10822 );
or \U$10749 ( \11435 , \11433 , \11434 );
nand \U$10750 ( \11436 , \10954 , RI89189a8_188);
nand \U$10751 ( \11437 , \11435 , \11436 );
not \U$10752 ( \11438 , \10811 );
not \U$10753 ( \11439 , RI89463f8_136);
or \U$10754 ( \11440 , \11438 , \11439 );
not \U$10755 ( \11441 , RI98088b8_84);
or \U$10756 ( \11442 , \11192 , \11441 );
nand \U$10757 ( \11443 , \11440 , \11442 );
nor \U$10758 ( \11444 , \11437 , \11443 );
nand \U$10759 ( \11445 , \11411 , \11421 , \11432 , \11444 );
and \U$10760 ( \11446 , \10902 , RI995eea0_6);
not \U$10761 ( \11447 , \10902 );
not \U$10762 ( \11448 , RI995eea0_6);
and \U$10763 ( \11449 , \11447 , \11448 );
nor \U$10764 ( \11450 , \11446 , \11449 );
nand \U$10765 ( \11451 , \11445 , \11450 );
and \U$10766 ( \11452 , \11400 , \11451 );
not \U$10767 ( \11453 , RI99672d0_218);
or \U$10768 ( \11454 , \10975 , \11453 );
not \U$10769 ( \11455 , \10821 );
nand \U$10770 ( \11456 , \11455 , RI890f7e0_205);
nand \U$10771 ( \11457 , \11454 , \11456 );
not \U$10772 ( \11458 , RI97771d8_101);
not \U$10773 ( \11459 , \10873 );
or \U$10774 ( \11460 , \11458 , \11459 );
nand \U$10775 ( \11461 , \10934 , RI8930a08_166);
nand \U$10776 ( \11462 , \11460 , \11461 );
nor \U$10777 ( \11463 , \11457 , \11462 );
not \U$10778 ( \11464 , \11128 );
not \U$10779 ( \11465 , RI8946218_140);
not \U$10780 ( \11466 , \11465 );
and \U$10781 ( \11467 , \11464 , \11466 );
and \U$10782 ( \11468 , \11001 , RI89ec898_114);
nor \U$10783 ( \11469 , \11467 , \11468 );
and \U$10784 ( \11470 , \11148 , RI995e6a8_231);
and \U$10785 ( \11471 , RI9921f28_596, RI994d830_244);
nor \U$10786 ( \11472 , \11470 , \11471 );
nand \U$10787 ( \11473 , \10842 , RI98bcb28_36);
and \U$10788 ( \11474 , \11469 , \11472 , \11473 );
not \U$10789 ( \11475 , RI8924ff0_179);
not \U$10790 ( \11476 , \11092 );
or \U$10791 ( \11477 , \11475 , \11476 );
nand \U$10792 ( \11478 , \10963 , RI98ab878_62);
nand \U$10793 ( \11479 , \11477 , \11478 );
not \U$10794 ( \11480 , RI98abe90_49);
not \U$10795 ( \11481 , \10919 );
or \U$10796 ( \11482 , \11480 , \11481 );
nand \U$10797 ( \11483 , \11057 , RI9819370_75);
nand \U$10798 ( \11484 , \11482 , \11483 );
nor \U$10799 ( \11485 , \11479 , \11484 );
not \U$10800 ( \11486 , RI89399f0_153);
not \U$10801 ( \11487 , \10930 );
or \U$10802 ( \11488 , \11486 , \11487 );
nand \U$10803 ( \11489 , \11125 , RI89ec280_127);
nand \U$10804 ( \11490 , \11488 , \11489 );
not \U$10805 ( \11491 , RI98086d8_88);
or \U$10806 ( \11492 , \10806 , \11491 );
not \U$10807 ( \11493 , RI89187c8_192);
or \U$10808 ( \11494 , \10862 , \11493 );
nand \U$10809 ( \11495 , \11492 , \11494 );
nor \U$10810 ( \11496 , \11490 , \11495 );
nand \U$10811 ( \11497 , \11463 , \11474 , \11485 , \11496 );
xor \U$10812 ( \11498 , \10897 , RI995ecc0_10);
nand \U$10813 ( \11499 , \11497 , \11498 );
nand \U$10814 ( \11500 , \11353 , \11452 , \11499 );
not \U$10815 ( \11501 , \11500 );
not \U$10816 ( \11502 , \11501 );
or \U$10817 ( \11503 , \11251 , \11502 );
and \U$10818 ( \11504 , \11463 , \11474 , \11485 , \11496 );
not \U$10819 ( \11505 , \11498 );
and \U$10820 ( \11506 , \11504 , \11505 );
not \U$10821 ( \11507 , \11506 );
not \U$10822 ( \11508 , \11309 );
or \U$10823 ( \11509 , \11507 , \11508 );
nor \U$10824 ( \11510 , \11334 , \11318 );
nor \U$10825 ( \11511 , \11323 , \11345 );
nor \U$10826 ( \11512 , \11329 , \11340 );
nand \U$10827 ( \11513 , \11510 , \11314 , \11511 , \11512 );
nor \U$10828 ( \11514 , \11513 , \11351 );
nand \U$10829 ( \11515 , \11294 , \11255 , \11261 );
nor \U$10830 ( \11516 , \11515 , \11288 );
nand \U$10831 ( \11517 , \10842 , RI98bcba0_35);
nand \U$10832 ( \11518 , \11298 , \11517 );
nor \U$10833 ( \11519 , \11518 , \11274 );
nand \U$10834 ( \11520 , \11516 , \11519 );
nor \U$10835 ( \11521 , \11520 , \11308 );
nor \U$10836 ( \11522 , \11514 , \11521 );
nand \U$10837 ( \11523 , \11509 , \11522 );
and \U$10838 ( \11524 , \11400 , \11352 , \11451 );
and \U$10839 ( \11525 , \11523 , \11524 );
not \U$10840 ( \11526 , \11399 );
not \U$10841 ( \11527 , \11398 );
nand \U$10842 ( \11528 , \11526 , \11527 );
not \U$10843 ( \11529 , \11450 );
not \U$10844 ( \11530 , \11445 );
nand \U$10845 ( \11531 , \11529 , \11530 );
and \U$10846 ( \11532 , \11528 , \11531 );
not \U$10847 ( \11533 , \11451 );
nor \U$10848 ( \11534 , \11532 , \11533 );
nor \U$10849 ( \11535 , \11525 , \11534 );
nand \U$10850 ( \11536 , \11503 , \11535 );
not \U$10851 ( \11537 , \11536 );
or \U$10852 ( \11538 , \11053 , \11537 );
not \U$10853 ( \11539 , \11051 );
not \U$10854 ( \11540 , \10967 );
not \U$10855 ( \11541 , \10973 );
nand \U$10856 ( \11542 , \11540 , \11541 );
not \U$10857 ( \11543 , \11006 );
nand \U$10858 ( \11544 , \11543 , \11013 );
and \U$10859 ( \11545 , \11542 , \11544 );
nor \U$10860 ( \11546 , \11545 , \11014 );
not \U$10861 ( \11547 , \11546 );
or \U$10862 ( \11548 , \11539 , \11547 );
not \U$10863 ( \11549 , \11049 );
not \U$10864 ( \11550 , \11050 );
nand \U$10865 ( \11551 , \11549 , \11550 );
nand \U$10866 ( \11552 , \11548 , \11551 );
nor \U$10867 ( \11553 , \10894 , \10909 );
or \U$10868 ( \11554 , \11552 , \11553 );
buf \U$10869 ( \11555 , \10910 );
nand \U$10870 ( \11556 , \11554 , \11555 );
nand \U$10871 ( \11557 , \11538 , \11556 );
not \U$10872 ( \11558 , RI8946038_144);
buf \U$10873 ( \11559 , \10788 );
nor \U$10874 ( \11560 , \11558 , \11559 );
nor \U$10875 ( \11561 , \10794 , \5840 );
nor \U$10876 ( \11562 , \11560 , \11561 );
buf \U$10877 ( \11563 , \10812 );
not \U$10878 ( \11564 , \11563 );
not \U$10879 ( \11565 , RI89ec0a0_131);
not \U$10880 ( \11566 , \11565 );
and \U$10881 ( \11567 , \11564 , \11566 );
buf \U$10882 ( \11568 , \10857 );
not \U$10883 ( \11569 , \11568 );
and \U$10884 ( \11570 , \11569 , RI89ec6b8_118);
nor \U$10885 ( \11571 , \11567 , \11570 );
nand \U$10886 ( \11572 , \11562 , \11571 );
buf \U$10887 ( \11573 , \10880 );
not \U$10888 ( \11574 , \11573 );
nand \U$10889 ( \11575 , \11574 , RI9776ff8_105);
not \U$10890 ( \11576 , \10874 );
nand \U$10891 ( \11577 , \11576 , RI98084f8_92);
and \U$10892 ( \11578 , \10834 , RI99670f0_222);
nand \U$10893 ( \11579 , RI995e4c8_235, RI9921f28_596);
not \U$10894 ( \11580 , \11579 );
nor \U$10895 ( \11581 , \11578 , \11580 );
buf \U$10896 ( \11582 , \10805 );
nand \U$10897 ( \11583 , \11582 , RI9808b10_79);
nand \U$10898 ( \11584 , \11575 , \11577 , \11581 , \11583 );
nor \U$10899 ( \11585 , \11572 , \11584 );
buf \U$10900 ( \11586 , \10829 );
not \U$10901 ( \11587 , \11586 );
not \U$10902 ( \11588 , \5825 );
and \U$10903 ( \11589 , \11587 , \11588 );
and \U$10904 ( \11590 , \10843 , RI994de48_27);
nor \U$10905 ( \11591 , \11589 , \11590 );
not \U$10906 ( \11592 , RI89185e8_196);
nor \U$10907 ( \11593 , \11592 , \10823 );
not \U$10908 ( \11594 , RI8924e10_183);
nor \U$10909 ( \11595 , \11594 , \10862 );
nor \U$10910 ( \11596 , \11593 , \11595 );
nand \U$10911 ( \11597 , \11591 , \11596 );
not \U$10912 ( \11598 , \10889 );
not \U$10913 ( \11599 , \11598 );
not \U$10914 ( \11600 , \11599 );
not \U$10915 ( \11601 , \5855 );
and \U$10916 ( \11602 , \11600 , \11601 );
not \U$10917 ( \11603 , \10868 );
not \U$10918 ( \11604 , \11603 );
and \U$10919 ( \11605 , \11604 , RI8930828_170);
nor \U$10920 ( \11606 , \11602 , \11605 );
not \U$10921 ( \11607 , \10848 );
nor \U$10922 ( \11608 , \11607 , \714 );
nor \U$10923 ( \11609 , \10885 , \5833 );
nor \U$10924 ( \11610 , \11608 , \11609 );
nand \U$10925 ( \11611 , \11606 , \11610 );
nor \U$10926 ( \11612 , \11597 , \11611 );
nand \U$10927 ( \11613 , \11585 , \11612 );
nand \U$10928 ( \11614 , RI995f080_2, RI995ef90_4, RI995f008_3, RI995ef18_5);
nor \U$10929 ( \11615 , \10904 , \11614 );
xor \U$10930 ( \11616 , RI995f0f8_1, \11615 );
not \U$10931 ( \11617 , \11616 );
and \U$10932 ( \11618 , \11613 , \11617 );
not \U$10933 ( \11619 , \11618 );
and \U$10934 ( \11620 , \11557 , \11619 );
not \U$10935 ( \11621 , \11613 );
nand \U$10936 ( \11622 , \11621 , \11616 );
not \U$10937 ( \11623 , \11622 );
nor \U$10938 ( \11624 , \11620 , \11623 );
and \U$10939 ( \11625 , RI995f0f8_1, \11615 );
not \U$10940 ( \11626 , \11625 );
nor \U$10941 ( \11627 , \11624 , \11626 );
not \U$10942 ( \11628 , \11627 );
not \U$10943 ( \11629 , \11625 );
nand \U$10944 ( \11630 , \11629 , \11624 );
nand \U$10945 ( \11631 , \11628 , \11630 );
not \U$10946 ( \11632 , \11631 );
not \U$10947 ( \11633 , \11632 );
not \U$10948 ( \11634 , \11630 );
not \U$10949 ( \11635 , \11634 );
and \U$10950 ( \11636 , \11633 , \11635 );
buf \U$10951 ( \11637 , \11636 );
buf \U$10952 ( \11638 , \11637 );
buf \U$10953 ( \11639 , \11635 );
buf \U$10954 ( \11640 , \10740 );
nand \U$10955 ( \11641 , \10832 , \11640 );
not \U$10956 ( \11642 , \11641 );
and \U$10957 ( \11643 , \11642 , \10918 );
not \U$10958 ( \11644 , \11642 );
not \U$10959 ( \11645 , \10918 );
and \U$10960 ( \11646 , \11644 , \11645 );
nor \U$10961 ( \11647 , \11643 , \11646 );
not \U$10962 ( \11648 , \11640 );
not \U$10963 ( \11649 , \11648 );
not \U$10964 ( \11650 , \10759 );
or \U$10965 ( \11651 , \11649 , \11650 );
not \U$10966 ( \11652 , \10744 );
nand \U$10967 ( \11653 , \11651 , \11652 );
not \U$10968 ( \11654 , \11653 );
nand \U$10969 ( \11655 , \11647 , \11654 );
not \U$10970 ( \11656 , \11655 );
nor \U$10971 ( \11657 , \11641 , \10800 );
not \U$10972 ( \11658 , \11657 );
not \U$10973 ( \11659 , \10775 );
nand \U$10974 ( \11660 , \11659 , \11641 );
not \U$10975 ( \11661 , \10809 );
nand \U$10976 ( \11662 , \11658 , \11660 , \11661 );
not \U$10977 ( \11663 , \10825 );
not \U$10978 ( \11664 , \11663 );
not \U$10979 ( \11665 , \10917 );
and \U$10980 ( \11666 , \11648 , \11665 );
not \U$10981 ( \11667 , \11648 );
and \U$10982 ( \11668 , \11667 , \10760 );
or \U$10983 ( \11669 , \11666 , \11668 );
nor \U$10984 ( \11670 , \11664 , \11669 );
not \U$10985 ( \11671 , \11670 );
and \U$10986 ( \11672 , \11662 , \11671 );
nand \U$10987 ( \11673 , \11656 , \11672 );
buf \U$10988 ( \11674 , \11673 );
not \U$10989 ( \11675 , \11674 );
not \U$10990 ( \11676 , \1650 );
and \U$10991 ( \11677 , \11675 , \11676 );
not \U$10992 ( \11678 , \11647 );
nor \U$10993 ( \11679 , \11678 , \11654 );
nand \U$10994 ( \11680 , \11672 , \11679 );
buf \U$10995 ( \11681 , \11680 );
nor \U$10996 ( \11682 , \11681 , \1654 );
nor \U$10997 ( \11683 , \11677 , \11682 );
and \U$10998 ( \11684 , \11662 , \11670 );
buf \U$10999 ( \11685 , \11684 );
nand \U$11000 ( \11686 , \11685 , \11679 );
not \U$11001 ( \11687 , \11686 );
not \U$11002 ( \11688 , \11687 );
not \U$11003 ( \11689 , \11688 );
not \U$11004 ( \11690 , \6128 );
and \U$11005 ( \11691 , \11689 , \11690 );
nand \U$11006 ( \11692 , \11685 , \11656 );
nor \U$11007 ( \11693 , \11692 , \6133 );
nor \U$11008 ( \11694 , \11691 , \11693 );
nand \U$11009 ( \11695 , \11683 , \11694 );
nor \U$11010 ( \11696 , \11647 , \11653 );
buf \U$11011 ( \11697 , \11696 );
nand \U$11012 ( \11698 , \11672 , \11697 );
buf \U$11013 ( \11699 , \11698 );
not \U$11014 ( \11700 , \11699 );
not \U$11015 ( \11701 , \1673 );
and \U$11016 ( \11702 , \11700 , \11701 );
nor \U$11017 ( \11703 , \11654 , \11647 );
nand \U$11018 ( \11704 , \11672 , \11703 );
buf \U$11019 ( \11705 , \11704 );
nor \U$11020 ( \11706 , \11705 , \1644 );
nor \U$11021 ( \11707 , \11702 , \11706 );
nand \U$11022 ( \11708 , \11685 , \11703 );
not \U$11023 ( \11709 , \11708 );
not \U$11024 ( \11710 , \11709 );
not \U$11025 ( \11711 , \11710 );
not \U$11026 ( \11712 , \6088 );
and \U$11027 ( \11713 , \11711 , \11712 );
nand \U$11028 ( \11714 , \11685 , \11697 );
buf \U$11029 ( \11715 , \11714 );
nor \U$11030 ( \11716 , \11715 , \6096 );
nor \U$11031 ( \11717 , \11713 , \11716 );
nand \U$11032 ( \11718 , \11707 , \11717 );
nor \U$11033 ( \11719 , \11695 , \11718 );
not \U$11034 ( \11720 , \11654 );
nand \U$11035 ( \11721 , \11720 , \11678 );
not \U$11036 ( \11722 , \11662 );
not \U$11037 ( \11723 , \11670 );
nand \U$11038 ( \11724 , \11722 , \11723 );
nor \U$11039 ( \11725 , \11721 , \11724 );
buf \U$11040 ( \11726 , \11725 );
nand \U$11041 ( \11727 , \11726 , RI992a1f0_389);
nand \U$11042 ( \11728 , \11647 , \11653 );
or \U$11043 ( \11729 , \11724 , \11728 );
not \U$11044 ( \11730 , \11729 );
nand \U$11045 ( \11731 , \11730 , RI992eed0_309);
not \U$11046 ( \11732 , \11696 );
nor \U$11047 ( \11733 , \11724 , \11732 );
buf \U$11048 ( \11734 , \11733 );
nand \U$11049 ( \11735 , \11734 , RI992ab50_369);
nor \U$11050 ( \11736 , \11724 , \11655 );
buf \U$11051 ( \11737 , \11736 );
nand \U$11052 ( \11738 , \11737 , RI992f830_289);
nand \U$11053 ( \11739 , \11727 , \11731 , \11735 , \11738 );
not \U$11054 ( \11740 , \11723 );
nand \U$11055 ( \11741 , \11740 , \11722 );
nor \U$11056 ( \11742 , \11741 , \11732 );
buf \U$11057 ( \11743 , \11742 );
and \U$11058 ( \11744 , \11743 , RI992cfe0_329);
not \U$11059 ( \11745 , RI9922bd0_569);
not \U$11060 ( \11746 , \10820 );
not \U$11061 ( \11747 , \11642 );
or \U$11062 ( \11748 , \11746 , \11747 );
nand \U$11063 ( \11749 , \11748 , \10840 );
not \U$11064 ( \11750 , \11749 );
or \U$11065 ( \11751 , \11745 , \11750 );
nand \U$11066 ( \11752 , \10843 , RI994d5d8_249);
nand \U$11067 ( \11753 , \11751 , \11752 );
nor \U$11068 ( \11754 , \11744 , \11753 );
nor \U$11069 ( \11755 , \11741 , \11728 );
buf \U$11070 ( \11756 , \11755 );
nand \U$11071 ( \11757 , \11756 , RI9931ae0_269);
nor \U$11072 ( \11758 , \11741 , \11721 );
buf \U$11073 ( \11759 , \11758 );
nand \U$11074 ( \11760 , \11759 , RI992b4b0_349);
nand \U$11075 ( \11761 , \11754 , \11757 , \11760 );
nor \U$11076 ( \11762 , \11739 , \11761 );
nand \U$11077 ( \11763 , \11719 , \11762 );
buf \U$11078 ( \11764 , \11763 );
not \U$11079 ( \11765 , \11764 );
and \U$11080 ( \11766 , \11639 , \11765 );
not \U$11081 ( \11767 , \11639 );
and \U$11082 ( \11768 , \11767 , \11764 );
nor \U$11083 ( \11769 , \11766 , \11768 );
nand \U$11084 ( \11770 , \11638 , \11769 );
not \U$11085 ( \11771 , \11770 );
not \U$11086 ( \11772 , RI9923878_548);
not \U$11087 ( \11773 , \11672 );
nor \U$11088 ( \11774 , \11773 , \11721 );
buf \U$11089 ( \11775 , \11774 );
not \U$11090 ( \11776 , \11775 );
or \U$11091 ( \11777 , \11772 , \11776 );
not \U$11092 ( \11778 , \11699 );
nand \U$11093 ( \11779 , \11778 , RI99241d8_528);
nand \U$11094 ( \11780 , \11777 , \11779 );
not \U$11095 ( \11781 , RI9924b38_508);
and \U$11096 ( \11782 , \11684 , \11703 );
not \U$11097 ( \11783 , \11782 );
or \U$11098 ( \11784 , \11781 , \11783 );
and \U$11099 ( \11785 , \11684 , \11697 );
buf \U$11100 ( \11786 , \11785 );
nand \U$11101 ( \11787 , \11786 , RI9925b28_488);
nand \U$11102 ( \11788 , \11784 , \11787 );
nor \U$11103 ( \11789 , \11780 , \11788 );
not \U$11104 ( \11790 , RI9926488_468);
not \U$11105 ( \11791 , \11681 );
not \U$11106 ( \11792 , \11791 );
or \U$11107 ( \11793 , \11790 , \11792 );
not \U$11108 ( \11794 , \11672 );
nor \U$11109 ( \11795 , \11794 , \11655 );
buf \U$11110 ( \11796 , \11795 );
nand \U$11111 ( \11797 , \11796 , RI9926de8_448);
nand \U$11112 ( \11798 , \11793 , \11797 );
not \U$11113 ( \11799 , RI9928198_428);
nand \U$11114 ( \11800 , \11685 , \11679 );
not \U$11115 ( \11801 , \11800 );
not \U$11116 ( \11802 , \11801 );
or \U$11117 ( \11803 , \11799 , \11802 );
nand \U$11118 ( \11804 , \11685 , \11656 );
not \U$11119 ( \11805 , \11804 );
nand \U$11120 ( \11806 , \11805 , RI9928af8_408);
nand \U$11121 ( \11807 , \11803 , \11806 );
nor \U$11122 ( \11808 , \11798 , \11807 );
not \U$11123 ( \11809 , RI992a268_388);
not \U$11124 ( \11810 , \11726 );
or \U$11125 ( \11811 , \11809 , \11810 );
nand \U$11126 ( \11812 , \11734 , RI992abc8_368);
nand \U$11127 ( \11813 , \11811 , \11812 );
not \U$11128 ( \11814 , RI992ef48_308);
or \U$11129 ( \11815 , \11724 , \11728 );
not \U$11130 ( \11816 , \11815 );
not \U$11131 ( \11817 , \11816 );
or \U$11132 ( \11818 , \11814 , \11817 );
nand \U$11133 ( \11819 , \11737 , RI992f8a8_288);
nand \U$11134 ( \11820 , \11818 , \11819 );
nor \U$11135 ( \11821 , \11813 , \11820 );
not \U$11136 ( \11822 , RI9931b58_268);
not \U$11137 ( \11823 , \11756 );
or \U$11138 ( \11824 , \11822 , \11823 );
nor \U$11139 ( \11825 , \11721 , \11741 );
buf \U$11140 ( \11826 , \11825 );
nand \U$11141 ( \11827 , \11826 , RI992c6f8_348);
nand \U$11142 ( \11828 , \11824 , \11827 );
not \U$11143 ( \11829 , RI992d058_328);
not \U$11144 ( \11830 , \11743 );
or \U$11145 ( \11831 , \11829 , \11830 );
and \U$11146 ( \11832 , \11749 , RI9922f18_568);
nand \U$11147 ( \11833 , \10843 , RI994d650_248);
not \U$11148 ( \11834 , \11833 );
nor \U$11149 ( \11835 , \11832 , \11834 );
nand \U$11150 ( \11836 , \11831 , \11835 );
nor \U$11151 ( \11837 , \11828 , \11836 );
nand \U$11152 ( \11838 , \11789 , \11808 , \11821 , \11837 );
buf \U$11153 ( \11839 , \11838 );
not \U$11154 ( \11840 , \11839 );
and \U$11155 ( \11841 , \11840 , \11639 );
not \U$11156 ( \11842 , \11840 );
and \U$11157 ( \11843 , \11842 , \11767 );
nor \U$11158 ( \11844 , \11841 , \11843 );
nand \U$11159 ( \11845 , \11638 , \11844 );
not \U$11160 ( \11846 , \11845 );
not \U$11161 ( \11847 , \11618 );
nand \U$11162 ( \11848 , \11847 , \11622 );
xnor \U$11163 ( \11849 , \11557 , \11848 );
not \U$11164 ( \11850 , \11849 );
not \U$11165 ( \11851 , \11850 );
not \U$11166 ( \11852 , \11051 );
nand \U$11167 ( \11853 , \10974 , \11015 );
nor \U$11168 ( \11854 , \11852 , \11853 );
not \U$11169 ( \11855 , \11854 );
not \U$11170 ( \11856 , \11536 );
or \U$11171 ( \11857 , \11855 , \11856 );
not \U$11172 ( \11858 , \11552 );
nand \U$11173 ( \11859 , \11857 , \11858 );
nor \U$11174 ( \11860 , \10894 , \10909 );
not \U$11175 ( \11861 , \11860 );
nand \U$11176 ( \11862 , \11861 , \11555 );
not \U$11177 ( \11863 , \11862 );
and \U$11178 ( \11864 , \11859 , \11863 );
not \U$11179 ( \11865 , \11859 );
and \U$11180 ( \11866 , \11865 , \11862 );
nor \U$11181 ( \11867 , \11864 , \11866 );
not \U$11182 ( \11868 , \11867 );
or \U$11183 ( \11869 , \11851 , \11868 );
not \U$11184 ( \11870 , \11867 );
nand \U$11185 ( \11871 , \11870 , \11849 );
nand \U$11186 ( \11872 , \11869 , \11871 );
buf \U$11187 ( \11873 , \11872 );
not \U$11188 ( \11874 , \11873 );
not \U$11189 ( \11875 , \11874 );
not \U$11190 ( \11876 , \11850 );
not \U$11191 ( \11877 , \11876 );
not \U$11192 ( \11878 , \11632 );
or \U$11193 ( \11879 , \11877 , \11878 );
nand \U$11194 ( \11880 , \11631 , \11850 );
nand \U$11195 ( \11881 , \11879 , \11880 );
not \U$11196 ( \11882 , \11872 );
nand \U$11197 ( \11883 , \11881 , \11882 );
not \U$11198 ( \11884 , \11883 );
buf \U$11199 ( \11885 , \11884 );
not \U$11200 ( \11886 , \11885 );
not \U$11201 ( \11887 , \11886 );
or \U$11202 ( \11888 , \11875 , \11887 );
buf \U$11203 ( \11889 , \11632 );
not \U$11204 ( \11890 , \11889 );
not \U$11205 ( \11891 , \11890 );
not \U$11206 ( \11892 , \11891 );
nand \U$11207 ( \11893 , \11888 , \11892 );
not \U$11208 ( \11894 , \11893 );
or \U$11209 ( \11895 , \11846 , \11894 );
or \U$11210 ( \11896 , \11893 , \11845 );
nand \U$11211 ( \11897 , \11895 , \11896 );
not \U$11212 ( \11898 , \11897 );
or \U$11213 ( \11899 , \11771 , \11898 );
or \U$11214 ( \11900 , \11897 , \11770 );
nand \U$11215 ( \11901 , \11899 , \11900 );
and \U$11216 ( \11902 , \11839 , \11891 );
not \U$11217 ( \11903 , \11839 );
and \U$11218 ( \11904 , \11903 , \11892 );
nor \U$11219 ( \11905 , \11902 , \11904 );
or \U$11220 ( \11906 , \11886 , \11905 );
or \U$11221 ( \11907 , \11874 , \11891 );
nand \U$11222 ( \11908 , \11906 , \11907 );
xor \U$11223 ( \11909 , \11908 , \11770 );
not \U$11224 ( \11910 , \11692 );
and \U$11225 ( \11911 , \11910 , RI9928a08_410);
buf \U$11226 ( \11912 , \11686 );
not \U$11227 ( \11913 , \11912 );
and \U$11228 ( \11914 , \11913 , RI99280a8_430);
nor \U$11229 ( \11915 , \11911 , \11914 );
and \U$11230 ( \11916 , \11796 , RI9926cf8_450);
not \U$11231 ( \11917 , \11681 );
and \U$11232 ( \11918 , \11917 , RI9926398_470);
nor \U$11233 ( \11919 , \11916 , \11918 );
nand \U$11234 ( \11920 , \11915 , \11919 );
and \U$11235 ( \11921 , \11786 , RI9925a38_490);
not \U$11236 ( \11922 , \11782 );
not \U$11237 ( \11923 , \11922 );
and \U$11238 ( \11924 , \11923 , RI9924a48_510);
nor \U$11239 ( \11925 , \11921 , \11924 );
not \U$11240 ( \11926 , \11699 );
and \U$11241 ( \11927 , \11926 , RI99240e8_530);
and \U$11242 ( \11928 , \11775 , RI9923788_550);
nor \U$11243 ( \11929 , \11927 , \11928 );
nand \U$11244 ( \11930 , \11925 , \11929 );
nor \U$11245 ( \11931 , \11920 , \11930 );
nand \U$11246 ( \11932 , \11726 , RI992a178_390);
nand \U$11247 ( \11933 , \11734 , RI992aad8_370);
nand \U$11248 ( \11934 , \11730 , RI992ee58_310);
nand \U$11249 ( \11935 , \11737 , RI992f7b8_290);
nand \U$11250 ( \11936 , \11932 , \11933 , \11934 , \11935 );
nand \U$11251 ( \11937 , \11743 , RI992cf68_330);
nand \U$11252 ( \11938 , \11826 , RI992b438_350);
nand \U$11253 ( \11939 , \11756 , RI9931a68_270);
and \U$11254 ( \11940 , \11749 , RI9922b58_570);
nand \U$11255 ( \11941 , \10843 , RI994d560_250);
not \U$11256 ( \11942 , \11941 );
nor \U$11257 ( \11943 , \11940 , \11942 );
nand \U$11258 ( \11944 , \11937 , \11938 , \11939 , \11943 );
nor \U$11259 ( \11945 , \11936 , \11944 );
nand \U$11260 ( \11946 , \11931 , \11945 );
not \U$11261 ( \11947 , \11946 );
and \U$11262 ( \11948 , \11639 , \11947 );
not \U$11263 ( \11949 , \11947 );
and \U$11264 ( \11950 , \11767 , \11949 );
nor \U$11265 ( \11951 , \11948 , \11950 );
nand \U$11266 ( \11952 , \11638 , \11951 );
not \U$11267 ( \11953 , \11952 );
not \U$11268 ( \11954 , \11953 );
not \U$11269 ( \11955 , \11886 );
not \U$11270 ( \11956 , \11764 );
not \U$11271 ( \11957 , \11891 );
or \U$11272 ( \11958 , \11956 , \11957 );
nand \U$11273 ( \11959 , \11892 , \11765 );
nand \U$11274 ( \11960 , \11958 , \11959 );
not \U$11275 ( \11961 , \11960 );
not \U$11276 ( \11962 , \11961 );
and \U$11277 ( \11963 , \11955 , \11962 );
nor \U$11278 ( \11964 , \11905 , \11874 );
nor \U$11279 ( \11965 , \11963 , \11964 );
not \U$11280 ( \11966 , \11965 );
not \U$11281 ( \11967 , \11966 );
or \U$11282 ( \11968 , \11954 , \11967 );
or \U$11283 ( \11969 , \11966 , \11953 );
buf \U$11284 ( \11970 , \10974 );
not \U$11285 ( \11971 , \11970 );
not \U$11286 ( \11972 , \11536 );
or \U$11287 ( \11973 , \11971 , \11972 );
buf \U$11288 ( \11974 , \11542 );
nand \U$11289 ( \11975 , \11973 , \11974 );
nand \U$11290 ( \11976 , \11544 , \11015 );
not \U$11291 ( \11977 , \11976 );
and \U$11292 ( \11978 , \11975 , \11977 );
not \U$11293 ( \11979 , \11975 );
and \U$11294 ( \11980 , \11979 , \11976 );
nor \U$11295 ( \11981 , \11978 , \11980 );
buf \U$11296 ( \11982 , \11981 );
not \U$11297 ( \11983 , \11853 );
not \U$11298 ( \11984 , \11983 );
buf \U$11299 ( \11985 , \11536 );
not \U$11300 ( \11986 , \11985 );
or \U$11301 ( \11987 , \11984 , \11986 );
not \U$11302 ( \11988 , \11546 );
nand \U$11303 ( \11989 , \11987 , \11988 );
not \U$11304 ( \11990 , \11852 );
nand \U$11305 ( \11991 , \11990 , \11551 );
not \U$11306 ( \11992 , \11991 );
and \U$11307 ( \11993 , \11989 , \11992 );
not \U$11308 ( \11994 , \11989 );
and \U$11309 ( \11995 , \11994 , \11991 );
nor \U$11310 ( \11996 , \11993 , \11995 );
and \U$11311 ( \11997 , \11982 , \11996 );
not \U$11312 ( \11998 , \11982 );
not \U$11313 ( \11999 , \11996 );
and \U$11314 ( \12000 , \11998 , \11999 );
nor \U$11315 ( \12001 , \11997 , \12000 );
buf \U$11316 ( \12002 , \12001 );
buf \U$11317 ( \12003 , \12002 );
not \U$11318 ( \12004 , \12003 );
not \U$11319 ( \12005 , \12004 );
not \U$11320 ( \12006 , \12001 );
not \U$11321 ( \12007 , \11867 );
not \U$11322 ( \12008 , \12007 );
not \U$11323 ( \12009 , \11996 );
or \U$11324 ( \12010 , \12008 , \12009 );
not \U$11325 ( \12011 , \11999 );
buf \U$11326 ( \12012 , \12007 );
or \U$11327 ( \12013 , \12011 , \12012 );
nand \U$11328 ( \12014 , \12010 , \12013 );
nand \U$11329 ( \12015 , \12006 , \12014 );
not \U$11330 ( \12016 , \12015 );
not \U$11331 ( \12017 , \12016 );
not \U$11332 ( \12018 , \12017 );
or \U$11333 ( \12019 , \12005 , \12018 );
not \U$11334 ( \12020 , \12012 );
nand \U$11335 ( \12021 , \12019 , \12020 );
nand \U$11336 ( \12022 , \11969 , \12021 );
nand \U$11337 ( \12023 , \11968 , \12022 );
and \U$11338 ( \12024 , \11909 , \12023 );
and \U$11339 ( \12025 , \11908 , \11770 );
or \U$11340 ( \12026 , \12024 , \12025 );
xnor \U$11341 ( \12027 , \11901 , \12026 );
not \U$11342 ( \12028 , \12027 );
not \U$11343 ( \12029 , \12012 );
and \U$11344 ( \12030 , \11840 , \12029 );
not \U$11345 ( \12031 , \11840 );
not \U$11346 ( \12032 , \12012 );
not \U$11347 ( \12033 , \12032 );
and \U$11348 ( \12034 , \12031 , \12033 );
nor \U$11349 ( \12035 , \12030 , \12034 );
not \U$11350 ( \12036 , \12035 );
not \U$11351 ( \12037 , \12036 );
not \U$11352 ( \12038 , \12017 );
not \U$11353 ( \12039 , \12038 );
or \U$11354 ( \12040 , \12037 , \12039 );
nand \U$11355 ( \12041 , \12003 , \12020 );
nand \U$11356 ( \12042 , \12040 , \12041 );
not \U$11357 ( \12043 , \12042 );
and \U$11358 ( \12044 , \12021 , \11952 );
not \U$11359 ( \12045 , \12021 );
and \U$11360 ( \12046 , \12045 , \11953 );
or \U$11361 ( \12047 , \12044 , \12046 );
and \U$11362 ( \12048 , \12047 , \11965 );
not \U$11363 ( \12049 , \12047 );
and \U$11364 ( \12050 , \12049 , \11966 );
nor \U$11365 ( \12051 , \12048 , \12050 );
not \U$11366 ( \12052 , \12051 );
not \U$11367 ( \12053 , \12052 );
or \U$11368 ( \12054 , \12043 , \12053 );
not \U$11369 ( \12055 , \12042 );
nand \U$11370 ( \12056 , \12051 , \12055 );
not \U$11371 ( \12057 , RI99249d0_511);
not \U$11372 ( \12058 , \11923 );
or \U$11373 ( \12059 , \12057 , \12058 );
nand \U$11374 ( \12060 , \11786 , RI99259c0_491);
nand \U$11375 ( \12061 , \12059 , \12060 );
not \U$11376 ( \12062 , RI9926320_471);
not \U$11377 ( \12063 , \11791 );
or \U$11378 ( \12064 , \12062 , \12063 );
nand \U$11379 ( \12065 , \11796 , RI9926c80_451);
nand \U$11380 ( \12066 , \12064 , \12065 );
nor \U$11381 ( \12067 , \12061 , \12066 );
not \U$11382 ( \12068 , RI9923710_551);
not \U$11383 ( \12069 , \11775 );
or \U$11384 ( \12070 , \12068 , \12069 );
nand \U$11385 ( \12071 , \11778 , RI9924070_531);
nand \U$11386 ( \12072 , \12070 , \12071 );
not \U$11387 ( \12073 , RI9928030_431);
not \U$11388 ( \12074 , \11801 );
or \U$11389 ( \12075 , \12073 , \12074 );
nand \U$11390 ( \12076 , \11805 , RI9928990_411);
nand \U$11391 ( \12077 , \12075 , \12076 );
nor \U$11392 ( \12078 , \12072 , \12077 );
not \U$11393 ( \12079 , RI992ede0_311);
not \U$11394 ( \12080 , \11816 );
or \U$11395 ( \12081 , \12079 , \12080 );
nand \U$11396 ( \12082 , \11737 , RI992f740_291);
nand \U$11397 ( \12083 , \12081 , \12082 );
not \U$11398 ( \12084 , RI992a100_391);
not \U$11399 ( \12085 , \11726 );
or \U$11400 ( \12086 , \12084 , \12085 );
nand \U$11401 ( \12087 , \11734 , RI992aa60_371);
nand \U$11402 ( \12088 , \12086 , \12087 );
nor \U$11403 ( \12089 , \12083 , \12088 );
not \U$11404 ( \12090 , RI99319f0_271);
not \U$11405 ( \12091 , \11756 );
or \U$11406 ( \12092 , \12090 , \12091 );
nand \U$11407 ( \12093 , \11826 , RI992b3c0_351);
nand \U$11408 ( \12094 , \12092 , \12093 );
not \U$11409 ( \12095 , RI992cef0_331);
not \U$11410 ( \12096 , \11743 );
or \U$11411 ( \12097 , \12095 , \12096 );
and \U$11412 ( \12098 , \11749 , RI9922ae0_571);
nand \U$11413 ( \12099 , \10843 , RI994d4e8_251);
not \U$11414 ( \12100 , \12099 );
nor \U$11415 ( \12101 , \12098 , \12100 );
nand \U$11416 ( \12102 , \12097 , \12101 );
nor \U$11417 ( \12103 , \12094 , \12102 );
nand \U$11418 ( \12104 , \12067 , \12078 , \12089 , \12103 );
not \U$11419 ( \12105 , \12104 );
not \U$11420 ( \12106 , \12105 );
not \U$11421 ( \12107 , \12106 );
not \U$11422 ( \12108 , \12107 );
and \U$11423 ( \12109 , \12108 , \11767 );
not \U$11424 ( \12110 , \12108 );
and \U$11425 ( \12111 , \12110 , \11639 );
nor \U$11426 ( \12112 , \12109 , \12111 );
and \U$11427 ( \12113 , \11638 , \12112 );
xor \U$11428 ( \12114 , \12113 , \12055 );
not \U$11429 ( \12115 , \11949 );
not \U$11430 ( \12116 , \11891 );
or \U$11431 ( \12117 , \12115 , \12116 );
buf \U$11432 ( \12118 , \11889 );
not \U$11433 ( \12119 , \12118 );
nand \U$11434 ( \12120 , \12119 , \11947 );
nand \U$11435 ( \12121 , \12117 , \12120 );
not \U$11436 ( \12122 , \12121 );
not \U$11437 ( \12123 , \11885 );
or \U$11438 ( \12124 , \12122 , \12123 );
nand \U$11439 ( \12125 , \11960 , \11873 );
nand \U$11440 ( \12126 , \12124 , \12125 );
and \U$11441 ( \12127 , \12114 , \12126 );
and \U$11442 ( \12128 , \12113 , \12055 );
or \U$11443 ( \12129 , \12127 , \12128 );
nand \U$11444 ( \12130 , \12056 , \12129 );
nand \U$11445 ( \12131 , \12054 , \12130 );
xor \U$11446 ( \12132 , \11908 , \11770 );
xor \U$11447 ( \12133 , \12132 , \12023 );
or \U$11448 ( \12134 , \12131 , \12133 );
not \U$11449 ( \12135 , \12134 );
not \U$11450 ( \12136 , \11839 );
buf \U$11451 ( \12137 , \11982 );
not \U$11452 ( \12138 , \12137 );
not \U$11453 ( \12139 , \12138 );
or \U$11454 ( \12140 , \12136 , \12139 );
nand \U$11455 ( \12141 , \12137 , \11840 );
nand \U$11456 ( \12142 , \12140 , \12141 );
not \U$11457 ( \12143 , \12142 );
nand \U$11458 ( \12144 , \11974 , \11970 );
not \U$11459 ( \12145 , \12144 );
not \U$11460 ( \12146 , \12145 );
not \U$11461 ( \12147 , \11985 );
not \U$11462 ( \12148 , \12147 );
or \U$11463 ( \12149 , \12146 , \12148 );
not \U$11464 ( \12150 , \12147 );
nand \U$11465 ( \12151 , \12150 , \12144 );
nand \U$11466 ( \12152 , \12149 , \12151 );
not \U$11467 ( \12153 , \12152 );
not \U$11468 ( \12154 , \11982 );
not \U$11469 ( \12155 , \12154 );
or \U$11470 ( \12156 , \12153 , \12155 );
not \U$11471 ( \12157 , \12152 );
nand \U$11472 ( \12158 , \12157 , \11982 );
nand \U$11473 ( \12159 , \12156 , \12158 );
not \U$11474 ( \12160 , \12152 );
and \U$11475 ( \12161 , \11451 , \11531 );
not \U$11476 ( \12162 , \12161 );
not \U$11477 ( \12163 , \12162 );
not \U$11478 ( \12164 , \11522 );
not \U$11479 ( \12165 , \11352 );
not \U$11480 ( \12166 , \12165 );
and \U$11481 ( \12167 , \12164 , \12166 );
nor \U$11482 ( \12168 , \11101 , \11106 );
and \U$11483 ( \12169 , \12168 , \11499 );
nor \U$11484 ( \12170 , \11497 , \11498 );
nor \U$11485 ( \12171 , \12169 , \12170 );
nand \U$11486 ( \12172 , \11243 , \11499 , \11107 );
nand \U$11487 ( \12173 , \12171 , \12172 );
buf \U$11488 ( \12174 , \11353 );
and \U$11489 ( \12175 , \12173 , \12174 );
nor \U$11490 ( \12176 , \12167 , \12175 );
buf \U$11491 ( \12177 , \11400 );
not \U$11492 ( \12178 , \12177 );
or \U$11493 ( \12179 , \12176 , \12178 );
nand \U$11494 ( \12180 , \12179 , \11528 );
not \U$11495 ( \12181 , \12180 );
or \U$11496 ( \12182 , \12163 , \12181 );
or \U$11497 ( \12183 , \12176 , \12178 );
nand \U$11498 ( \12184 , \12183 , \12161 , \11528 );
nand \U$11499 ( \12185 , \12182 , \12184 );
not \U$11500 ( \12186 , \12185 );
not \U$11501 ( \12187 , \12186 );
or \U$11502 ( \12188 , \12160 , \12187 );
not \U$11503 ( \12189 , \12186 );
nand \U$11504 ( \12190 , \12157 , \12189 );
nand \U$11505 ( \12191 , \12188 , \12190 );
not \U$11506 ( \12192 , \12191 );
nand \U$11507 ( \12193 , \12159 , \12192 );
not \U$11508 ( \12194 , \12193 );
not \U$11509 ( \12195 , \12194 );
or \U$11510 ( \12196 , \12143 , \12195 );
not \U$11511 ( \12197 , \12192 );
buf \U$11512 ( \12198 , \12154 );
not \U$11513 ( \12199 , \12198 );
nand \U$11514 ( \12200 , \12197 , \12199 );
nand \U$11515 ( \12201 , \12196 , \12200 );
not \U$11516 ( \12202 , \11674 );
not \U$11517 ( \12203 , \6571 );
and \U$11518 ( \12204 , \12202 , \12203 );
nor \U$11519 ( \12205 , \11681 , \2129 );
nor \U$11520 ( \12206 , \12204 , \12205 );
not \U$11521 ( \12207 , \11688 );
not \U$11522 ( \12208 , RI9927f40_433);
not \U$11523 ( \12209 , \12208 );
and \U$11524 ( \12210 , \12207 , \12209 );
buf \U$11525 ( \12211 , \11804 );
not \U$11526 ( \12212 , RI99288a0_413);
nor \U$11527 ( \12213 , \12211 , \12212 );
nor \U$11528 ( \12214 , \12210 , \12213 );
nand \U$11529 ( \12215 , \12206 , \12214 );
not \U$11530 ( \12216 , \11705 );
not \U$11531 ( \12217 , \2108 );
and \U$11532 ( \12218 , \12216 , \12217 );
nor \U$11533 ( \12219 , \11699 , \2136 );
nor \U$11534 ( \12220 , \12218 , \12219 );
not \U$11535 ( \12221 , \11710 );
not \U$11536 ( \12222 , RI99248e0_513);
not \U$11537 ( \12223 , \12222 );
and \U$11538 ( \12224 , \12221 , \12223 );
not \U$11539 ( \12225 , RI99258d0_493);
nor \U$11540 ( \12226 , \11715 , \12225 );
nor \U$11541 ( \12227 , \12224 , \12226 );
nand \U$11542 ( \12228 , \12220 , \12227 );
nor \U$11543 ( \12229 , \12215 , \12228 );
nand \U$11544 ( \12230 , \11737 , RI992f650_293);
nand \U$11545 ( \12231 , \11816 , RI992ecf0_313);
nand \U$11546 ( \12232 , \11734 , RI992a970_373);
nand \U$11547 ( \12233 , \11726 , RI9929200_393);
nand \U$11548 ( \12234 , \12230 , \12231 , \12232 , \12233 );
and \U$11549 ( \12235 , \11743 , RI992ce00_333);
not \U$11550 ( \12236 , RI99229f0_573);
not \U$11551 ( \12237 , \11749 );
or \U$11552 ( \12238 , \12236 , \12237 );
nand \U$11553 ( \12239 , \10843 , RI994d3f8_253);
nand \U$11554 ( \12240 , \12238 , \12239 );
nor \U$11555 ( \12241 , \12235 , \12240 );
nand \U$11556 ( \12242 , \11756 , RI9931900_273);
nand \U$11557 ( \12243 , \11759 , RI992b2d0_353);
nand \U$11558 ( \12244 , \12241 , \12242 , \12243 );
nor \U$11559 ( \12245 , \12234 , \12244 );
nand \U$11560 ( \12246 , \12229 , \12245 );
buf \U$11561 ( \12247 , \12246 );
and \U$11562 ( \12248 , \12247 , \11767 );
not \U$11563 ( \12249 , \12247 );
and \U$11564 ( \12250 , \12249 , \11639 );
nor \U$11565 ( \12251 , \12248 , \12250 );
and \U$11566 ( \12252 , \11638 , \12251 );
xor \U$11567 ( \12253 , \12201 , \12252 );
not \U$11568 ( \12254 , RI9923698_552);
not \U$11569 ( \12255 , \11775 );
or \U$11570 ( \12256 , \12254 , \12255 );
nand \U$11571 ( \12257 , \11926 , RI9923ff8_532);
nand \U$11572 ( \12258 , \12256 , \12257 );
not \U$11573 ( \12259 , RI9924958_512);
not \U$11574 ( \12260 , \11923 );
or \U$11575 ( \12261 , \12259 , \12260 );
nand \U$11576 ( \12262 , \11786 , RI9925948_492);
nand \U$11577 ( \12263 , \12261 , \12262 );
nor \U$11578 ( \12264 , \12258 , \12263 );
not \U$11579 ( \12265 , RI99262a8_472);
not \U$11580 ( \12266 , \11791 );
or \U$11581 ( \12267 , \12265 , \12266 );
nand \U$11582 ( \12268 , \11796 , RI9926c08_452);
nand \U$11583 ( \12269 , \12267 , \12268 );
not \U$11584 ( \12270 , RI9927fb8_432);
not \U$11585 ( \12271 , \11801 );
or \U$11586 ( \12272 , \12270 , \12271 );
nand \U$11587 ( \12273 , \11805 , RI9928918_412);
nand \U$11588 ( \12274 , \12272 , \12273 );
nor \U$11589 ( \12275 , \12269 , \12274 );
not \U$11590 ( \12276 , RI9929278_392);
not \U$11591 ( \12277 , \11726 );
or \U$11592 ( \12278 , \12276 , \12277 );
nand \U$11593 ( \12279 , \11734 , RI992a9e8_372);
nand \U$11594 ( \12280 , \12278 , \12279 );
not \U$11595 ( \12281 , RI992ed68_312);
not \U$11596 ( \12282 , \11816 );
or \U$11597 ( \12283 , \12281 , \12282 );
nand \U$11598 ( \12284 , \11737 , RI992f6c8_292);
nand \U$11599 ( \12285 , \12283 , \12284 );
nor \U$11600 ( \12286 , \12280 , \12285 );
not \U$11601 ( \12287 , RI9931978_272);
not \U$11602 ( \12288 , \11756 );
or \U$11603 ( \12289 , \12287 , \12288 );
nand \U$11604 ( \12290 , \11826 , RI992b348_352);
nand \U$11605 ( \12291 , \12289 , \12290 );
not \U$11606 ( \12292 , RI992ce78_332);
not \U$11607 ( \12293 , \11743 );
or \U$11608 ( \12294 , \12292 , \12293 );
and \U$11609 ( \12295 , \11749 , RI9922a68_572);
nand \U$11610 ( \12296 , \10843 , RI994d470_252);
not \U$11611 ( \12297 , \12296 );
nor \U$11612 ( \12298 , \12295 , \12297 );
nand \U$11613 ( \12299 , \12294 , \12298 );
nor \U$11614 ( \12300 , \12291 , \12299 );
nand \U$11615 ( \12301 , \12264 , \12275 , \12286 , \12300 );
buf \U$11616 ( \12302 , \12301 );
not \U$11617 ( \12303 , \12302 );
not \U$11618 ( \12304 , \11891 );
or \U$11619 ( \12305 , \12303 , \12304 );
not \U$11620 ( \12306 , \12302 );
nand \U$11621 ( \12307 , \12119 , \12306 );
nand \U$11622 ( \12308 , \12305 , \12307 );
not \U$11623 ( \12309 , \12308 );
not \U$11624 ( \12310 , \11885 );
or \U$11625 ( \12311 , \12309 , \12310 );
not \U$11626 ( \12312 , \12108 );
not \U$11627 ( \12313 , \11891 );
or \U$11628 ( \12314 , \12312 , \12313 );
nand \U$11629 ( \12315 , \12119 , \12107 );
nand \U$11630 ( \12316 , \12314 , \12315 );
nand \U$11631 ( \12317 , \12316 , \11873 );
nand \U$11632 ( \12318 , \12311 , \12317 );
xor \U$11633 ( \12319 , \12253 , \12318 );
not \U$11634 ( \12320 , \12319 );
not \U$11635 ( \12321 , \11949 );
buf \U$11636 ( \12322 , \11867 );
not \U$11637 ( \12323 , \12322 );
not \U$11638 ( \12324 , \12323 );
or \U$11639 ( \12325 , \12321 , \12324 );
not \U$11640 ( \12326 , \12012 );
not \U$11641 ( \12327 , \12326 );
not \U$11642 ( \12328 , \12327 );
nand \U$11643 ( \12329 , \12328 , \11947 );
nand \U$11644 ( \12330 , \12325 , \12329 );
not \U$11645 ( \12331 , \12330 );
not \U$11646 ( \12332 , \12038 );
or \U$11647 ( \12333 , \12331 , \12332 );
and \U$11648 ( \12334 , \11764 , \12033 );
not \U$11649 ( \12335 , \11764 );
and \U$11650 ( \12336 , \12335 , \12020 );
nor \U$11651 ( \12337 , \12334 , \12336 );
not \U$11652 ( \12338 , \12337 );
nand \U$11653 ( \12339 , \12338 , \12003 );
nand \U$11654 ( \12340 , \12333 , \12339 );
not \U$11655 ( \12341 , \12340 );
not \U$11656 ( \12342 , \12178 );
nand \U$11657 ( \12343 , \12342 , \11528 );
xor \U$11658 ( \12344 , \12176 , \12343 );
buf \U$11659 ( \12345 , \11309 );
not \U$11660 ( \12346 , \12345 );
not \U$11661 ( \12347 , \12173 );
or \U$11662 ( \12348 , \12346 , \12347 );
not \U$11663 ( \12349 , \11521 );
nand \U$11664 ( \12350 , \12348 , \12349 );
nor \U$11665 ( \12351 , \12165 , \11514 );
and \U$11666 ( \12352 , \12350 , \12351 );
not \U$11667 ( \12353 , \12350 );
not \U$11668 ( \12354 , \12351 );
and \U$11669 ( \12355 , \12353 , \12354 );
nor \U$11670 ( \12356 , \12352 , \12355 );
buf \U$11671 ( \12357 , \12356 );
not \U$11672 ( \12358 , \12357 );
and \U$11673 ( \12359 , \12344 , \12358 );
not \U$11674 ( \12360 , \12344 );
and \U$11675 ( \12361 , \12360 , \12357 );
nor \U$11676 ( \12362 , \12359 , \12361 );
buf \U$11677 ( \12363 , \12362 );
not \U$11678 ( \12364 , \12363 );
buf \U$11679 ( \12365 , \12364 );
not \U$11680 ( \12366 , \12365 );
not \U$11681 ( \12367 , \12366 );
not \U$11682 ( \12368 , \12185 );
not \U$11683 ( \12369 , \12344 );
nand \U$11684 ( \12370 , \12368 , \12369 );
buf \U$11685 ( \12371 , \12185 );
not \U$11686 ( \12372 , \12369 );
nand \U$11687 ( \12373 , \12371 , \12372 );
nand \U$11688 ( \12374 , \12362 , \12370 , \12373 );
not \U$11689 ( \12375 , \12374 );
not \U$11690 ( \12376 , \12375 );
not \U$11691 ( \12377 , \12376 );
or \U$11692 ( \12378 , \12367 , \12377 );
nand \U$11693 ( \12379 , \12378 , \12371 );
not \U$11694 ( \12380 , \11764 );
not \U$11695 ( \12381 , \12138 );
or \U$11696 ( \12382 , \12380 , \12381 );
not \U$11697 ( \12383 , \12154 );
nand \U$11698 ( \12384 , \12383 , \11765 );
nand \U$11699 ( \12385 , \12382 , \12384 );
not \U$11700 ( \12386 , \12385 );
not \U$11701 ( \12387 , \12194 );
or \U$11702 ( \12388 , \12386 , \12387 );
nand \U$11703 ( \12389 , \12142 , \12197 );
nand \U$11704 ( \12390 , \12388 , \12389 );
xor \U$11705 ( \12391 , \12379 , \12390 );
not \U$11706 ( \12392 , \12108 );
not \U$11707 ( \12393 , \12020 );
not \U$11708 ( \12394 , \12393 );
or \U$11709 ( \12395 , \12392 , \12394 );
nand \U$11710 ( \12396 , \12322 , \12107 );
nand \U$11711 ( \12397 , \12395 , \12396 );
not \U$11712 ( \12398 , \12397 );
buf \U$11713 ( \12399 , \12016 );
not \U$11714 ( \12400 , \12399 );
or \U$11715 ( \12401 , \12398 , \12400 );
nand \U$11716 ( \12402 , \12003 , \12330 );
nand \U$11717 ( \12403 , \12401 , \12402 );
and \U$11718 ( \12404 , \12391 , \12403 );
and \U$11719 ( \12405 , \12379 , \12390 );
or \U$11720 ( \12406 , \12404 , \12405 );
xor \U$11721 ( \12407 , \12341 , \12406 );
not \U$11722 ( \12408 , \12247 );
not \U$11723 ( \12409 , \12118 );
or \U$11724 ( \12410 , \12408 , \12409 );
not \U$11725 ( \12411 , \12247 );
nand \U$11726 ( \12412 , \11890 , \12411 );
nand \U$11727 ( \12413 , \12410 , \12412 );
not \U$11728 ( \12414 , \12413 );
not \U$11729 ( \12415 , \11885 );
or \U$11730 ( \12416 , \12414 , \12415 );
nand \U$11731 ( \12417 , \12308 , \11873 );
nand \U$11732 ( \12418 , \12416 , \12417 );
not \U$11733 ( \12419 , \12418 );
not \U$11734 ( \12420 , \11709 );
not \U$11735 ( \12421 , \12420 );
not \U$11736 ( \12422 , \6761 );
and \U$11737 ( \12423 , \12421 , \12422 );
not \U$11738 ( \12424 , RI9925858_494);
nor \U$11739 ( \12425 , \11715 , \12424 );
nor \U$11740 ( \12426 , \12423 , \12425 );
not \U$11741 ( \12427 , \11801 );
not \U$11742 ( \12428 , \12427 );
not \U$11743 ( \12429 , \6783 );
and \U$11744 ( \12430 , \12428 , \12429 );
nor \U$11745 ( \12431 , \11692 , \6787 );
nor \U$11746 ( \12432 , \12430 , \12431 );
nand \U$11747 ( \12433 , \12426 , \12432 );
not \U$11748 ( \12434 , \11674 );
not \U$11749 ( \12435 , \6775 );
and \U$11750 ( \12436 , \12434 , \12435 );
nor \U$11751 ( \12437 , \11681 , \2057 );
nor \U$11752 ( \12438 , \12436 , \12437 );
not \U$11753 ( \12439 , \11705 );
not \U$11754 ( \12440 , \2036 );
and \U$11755 ( \12441 , \12439 , \12440 );
nor \U$11756 ( \12442 , \11699 , \2064 );
nor \U$11757 ( \12443 , \12441 , \12442 );
nand \U$11758 ( \12444 , \12438 , \12443 );
nor \U$11759 ( \12445 , \12433 , \12444 );
nand \U$11760 ( \12446 , \11737 , RI992f5d8_294);
nand \U$11761 ( \12447 , \11816 , RI992d6e8_314);
nand \U$11762 ( \12448 , \11734 , RI992a8f8_374);
nand \U$11763 ( \12449 , \11726 , RI9929188_394);
nand \U$11764 ( \12450 , \12446 , \12447 , \12448 , \12449 );
nand \U$11765 ( \12451 , \11759 , RI992b258_354);
nand \U$11766 ( \12452 , \11756 , RI9931888_274);
and \U$11767 ( \12453 , \11743 , RI992cd88_334);
not \U$11768 ( \12454 , RI9922978_574);
not \U$11769 ( \12455 , \11749 );
or \U$11770 ( \12456 , \12454 , \12455 );
nand \U$11771 ( \12457 , \10843 , RI9935fc8_254);
nand \U$11772 ( \12458 , \12456 , \12457 );
nor \U$11773 ( \12459 , \12453 , \12458 );
nand \U$11774 ( \12460 , \12451 , \12452 , \12459 );
nor \U$11775 ( \12461 , \12450 , \12460 );
nand \U$11776 ( \12462 , \12445 , \12461 );
buf \U$11777 ( \12463 , \12462 );
not \U$11778 ( \12464 , \12463 );
and \U$11779 ( \12465 , \12464 , \11635 );
not \U$11780 ( \12466 , \12464 );
not \U$11781 ( \12467 , \11635 );
and \U$11782 ( \12468 , \12466 , \12467 );
nor \U$11783 ( \12469 , \12465 , \12468 );
nand \U$11784 ( \12470 , \11638 , \12469 );
not \U$11785 ( \12471 , \12376 );
not \U$11786 ( \12472 , \11839 );
not \U$11787 ( \12473 , \12189 );
not \U$11788 ( \12474 , \12473 );
or \U$11789 ( \12475 , \12472 , \12474 );
nand \U$11790 ( \12476 , \12371 , \11840 );
nand \U$11791 ( \12477 , \12475 , \12476 );
not \U$11792 ( \12478 , \12477 );
not \U$11793 ( \12479 , \12478 );
and \U$11794 ( \12480 , \12471 , \12479 );
not \U$11795 ( \12481 , \12371 );
nor \U$11796 ( \12482 , \12366 , \12481 );
nor \U$11797 ( \12483 , \12480 , \12482 );
buf \U$11798 ( \12484 , \12483 );
nand \U$11799 ( \12485 , \12470 , \12484 );
not \U$11800 ( \12486 , \12485 );
or \U$11801 ( \12487 , \12419 , \12486 );
not \U$11802 ( \12488 , \12470 );
not \U$11803 ( \12489 , \12484 );
nand \U$11804 ( \12490 , \12488 , \12489 );
nand \U$11805 ( \12491 , \12487 , \12490 );
xor \U$11806 ( \12492 , \12407 , \12491 );
not \U$11807 ( \12493 , \12492 );
or \U$11808 ( \12494 , \12320 , \12493 );
or \U$11809 ( \12495 , \12492 , \12319 );
xor \U$11810 ( \12496 , \12483 , \12488 );
xor \U$11811 ( \12497 , \12496 , \12418 );
not \U$11812 ( \12498 , \12497 );
xor \U$11813 ( \12499 , \12379 , \12390 );
xor \U$11814 ( \12500 , \12499 , \12403 );
not \U$11815 ( \12501 , \12500 );
not \U$11816 ( \12502 , \12501 );
or \U$11817 ( \12503 , \12498 , \12502 );
not \U$11818 ( \12504 , \11949 );
not \U$11819 ( \12505 , \12138 );
or \U$11820 ( \12506 , \12504 , \12505 );
nand \U$11821 ( \12507 , \12137 , \11947 );
nand \U$11822 ( \12508 , \12506 , \12507 );
not \U$11823 ( \12509 , \12508 );
not \U$11824 ( \12510 , \12194 );
or \U$11825 ( \12511 , \12509 , \12510 );
nand \U$11826 ( \12512 , \12385 , \12197 );
nand \U$11827 ( \12513 , \12511 , \12512 );
not \U$11828 ( \12514 , \12302 );
not \U$11829 ( \12515 , \12323 );
or \U$11830 ( \12516 , \12514 , \12515 );
nand \U$11831 ( \12517 , \12020 , \12306 );
nand \U$11832 ( \12518 , \12516 , \12517 );
not \U$11833 ( \12519 , \12518 );
buf \U$11834 ( \12520 , \12015 );
not \U$11835 ( \12521 , \12520 );
not \U$11836 ( \12522 , \12521 );
or \U$11837 ( \12523 , \12519 , \12522 );
not \U$11838 ( \12524 , \12002 );
not \U$11839 ( \12525 , \12524 );
nand \U$11840 ( \12526 , \12525 , \12397 );
nand \U$11841 ( \12527 , \12523 , \12526 );
xor \U$11842 ( \12528 , \12513 , \12527 );
not \U$11843 ( \12529 , \12463 );
not \U$11844 ( \12530 , \12118 );
or \U$11845 ( \12531 , \12529 , \12530 );
buf \U$11846 ( \12532 , \11631 );
not \U$11847 ( \12533 , \12532 );
not \U$11848 ( \12534 , \12533 );
nand \U$11849 ( \12535 , \12534 , \12464 );
nand \U$11850 ( \12536 , \12531 , \12535 );
not \U$11851 ( \12537 , \12536 );
not \U$11852 ( \12538 , \11884 );
or \U$11853 ( \12539 , \12537 , \12538 );
not \U$11854 ( \12540 , \11882 );
nand \U$11855 ( \12541 , \12413 , \12540 );
nand \U$11856 ( \12542 , \12539 , \12541 );
and \U$11857 ( \12543 , \12528 , \12542 );
and \U$11858 ( \12544 , \12513 , \12527 );
or \U$11859 ( \12545 , \12543 , \12544 );
nand \U$11860 ( \12546 , \12503 , \12545 );
not \U$11861 ( \12547 , \12497 );
nand \U$11862 ( \12548 , \12547 , \12500 );
nand \U$11863 ( \12549 , \12546 , \12548 );
nand \U$11864 ( \12550 , \12495 , \12549 );
nand \U$11865 ( \12551 , \12494 , \12550 );
xor \U$11866 ( \12552 , \12201 , \12252 );
and \U$11867 ( \12553 , \12552 , \12318 );
and \U$11868 ( \12554 , \12201 , \12252 );
or \U$11869 ( \12555 , \12553 , \12554 );
xor \U$11870 ( \12556 , \12341 , \12406 );
and \U$11871 ( \12557 , \12556 , \12491 );
and \U$11872 ( \12558 , \12341 , \12406 );
or \U$11873 ( \12559 , \12557 , \12558 );
xor \U$11874 ( \12560 , \12555 , \12559 );
and \U$11875 ( \12561 , \11767 , \12302 );
not \U$11876 ( \12562 , \11767 );
and \U$11877 ( \12563 , \12562 , \12306 );
nor \U$11878 ( \12564 , \12561 , \12563 );
nand \U$11879 ( \12565 , \11638 , \12564 );
and \U$11880 ( \12566 , \12565 , \12340 );
not \U$11881 ( \12567 , \12565 );
and \U$11882 ( \12568 , \12567 , \12341 );
or \U$11883 ( \12569 , \12566 , \12568 );
not \U$11884 ( \12570 , \12399 );
not \U$11885 ( \12571 , \12570 );
not \U$11886 ( \12572 , \12337 );
and \U$11887 ( \12573 , \12571 , \12572 );
nor \U$11888 ( \12574 , \12004 , \12035 );
nor \U$11889 ( \12575 , \12573 , \12574 );
not \U$11890 ( \12576 , \12192 );
not \U$11891 ( \12577 , \12193 );
or \U$11892 ( \12578 , \12576 , \12577 );
nand \U$11893 ( \12579 , \12578 , \12199 );
not \U$11894 ( \12580 , \12579 );
and \U$11895 ( \12581 , \12575 , \12580 );
not \U$11896 ( \12582 , \12575 );
and \U$11897 ( \12583 , \12582 , \12579 );
nor \U$11898 ( \12584 , \12581 , \12583 );
not \U$11899 ( \12585 , \12316 );
not \U$11900 ( \12586 , \11885 );
or \U$11901 ( \12587 , \12585 , \12586 );
nand \U$11902 ( \12588 , \12121 , \11873 );
nand \U$11903 ( \12589 , \12587 , \12588 );
not \U$11904 ( \12590 , \12589 );
and \U$11905 ( \12591 , \12584 , \12590 );
not \U$11906 ( \12592 , \12584 );
and \U$11907 ( \12593 , \12592 , \12589 );
nor \U$11908 ( \12594 , \12591 , \12593 );
xnor \U$11909 ( \12595 , \12569 , \12594 );
xor \U$11910 ( \12596 , \12560 , \12595 );
nor \U$11911 ( \12597 , \12551 , \12596 );
not \U$11912 ( \12598 , \12597 );
not \U$11913 ( \12599 , \11767 );
nand \U$11914 ( \12600 , \11791 , RI9926140_475);
nand \U$11915 ( \12601 , \11795 , RI9926aa0_455);
nand \U$11916 ( \12602 , \11782 , RI99247f0_515);
nand \U$11917 ( \12603 , \11785 , RI99257e0_495);
nand \U$11918 ( \12604 , \12600 , \12601 , \12602 , \12603 );
nand \U$11919 ( \12605 , \11775 , RI9923530_555);
nand \U$11920 ( \12606 , \11778 , RI9923e90_535);
nand \U$11921 ( \12607 , \11687 , RI9927e50_435);
nand \U$11922 ( \12608 , \11805 , RI99287b0_415);
nand \U$11923 ( \12609 , \12605 , \12606 , \12607 , \12608 );
nor \U$11924 ( \12610 , \12604 , \12609 );
nand \U$11925 ( \12611 , \11726 , RI9929110_395);
nand \U$11926 ( \12612 , \11734 , RI992a880_375);
nand \U$11927 ( \12613 , \11737 , RI992f560_295);
nand \U$11928 ( \12614 , \11730 , RI992d670_315);
nand \U$11929 ( \12615 , \12611 , \12612 , \12613 , \12614 );
nand \U$11930 ( \12616 , \11743 , RI992cd10_335);
nand \U$11931 ( \12617 , \11756 , RI9931810_275);
nand \U$11932 ( \12618 , \11825 , RI992b1e0_355);
and \U$11933 ( \12619 , \11749 , RI9922900_575);
nand \U$11934 ( \12620 , \10843 , RI9935f50_255);
not \U$11935 ( \12621 , \12620 );
nor \U$11936 ( \12622 , \12619 , \12621 );
nand \U$11937 ( \12623 , \12616 , \12617 , \12618 , \12622 );
nor \U$11938 ( \12624 , \12615 , \12623 );
nand \U$11939 ( \12625 , \12610 , \12624 );
not \U$11940 ( \12626 , \12625 );
not \U$11941 ( \12627 , \12626 );
not \U$11942 ( \12628 , \12627 );
and \U$11943 ( \12629 , \12599 , \12628 );
and \U$11944 ( \12630 , \11767 , \12627 );
nor \U$11945 ( \12631 , \12629 , \12630 );
nand \U$11946 ( \12632 , \11638 , \12631 );
not \U$11947 ( \12633 , \12632 );
not \U$11948 ( \12634 , \12489 );
and \U$11949 ( \12635 , \12633 , \12634 );
not \U$11950 ( \12636 , \11763 );
buf \U$11951 ( \12637 , \12186 );
not \U$11952 ( \12638 , \12637 );
or \U$11953 ( \12639 , \12636 , \12638 );
not \U$11954 ( \12640 , \11763 );
nand \U$11955 ( \12641 , \12189 , \12640 );
nand \U$11956 ( \12642 , \12639 , \12641 );
not \U$11957 ( \12643 , \12642 );
and \U$11958 ( \12644 , \12373 , \12370 , \12362 );
not \U$11959 ( \12645 , \12644 );
or \U$11960 ( \12646 , \12643 , \12645 );
nand \U$11961 ( \12647 , \12477 , \12364 );
nand \U$11962 ( \12648 , \12646 , \12647 );
not \U$11963 ( \12649 , \12648 );
nand \U$11964 ( \12650 , \12345 , \12349 );
xnor \U$11965 ( \12651 , \12650 , \12173 );
not \U$11966 ( \12652 , \12651 );
not \U$11967 ( \12653 , \12652 );
not \U$11968 ( \12654 , \11506 );
nand \U$11969 ( \12655 , \12654 , \11499 );
not \U$11970 ( \12656 , \12655 );
and \U$11971 ( \12657 , \11250 , \12656 );
not \U$11972 ( \12658 , \11250 );
and \U$11973 ( \12659 , \12658 , \12655 );
nor \U$11974 ( \12660 , \12657 , \12659 );
not \U$11975 ( \12661 , \12660 );
not \U$11976 ( \12662 , \12661 );
not \U$11977 ( \12663 , \12662 );
or \U$11978 ( \12664 , \12653 , \12663 );
nand \U$11979 ( \12665 , \12651 , \12661 );
nand \U$11980 ( \12666 , \12664 , \12665 );
buf \U$11981 ( \12667 , \12666 );
not \U$11982 ( \12668 , \12667 );
not \U$11983 ( \12669 , \12668 );
not \U$11984 ( \12670 , \12357 );
not \U$11985 ( \12671 , \12652 );
not \U$11986 ( \12672 , \12671 );
nand \U$11987 ( \12673 , \12670 , \12672 );
nand \U$11988 ( \12674 , \12357 , \12671 );
not \U$11989 ( \12675 , \12652 );
not \U$11990 ( \12676 , \12662 );
or \U$11991 ( \12677 , \12675 , \12676 );
nand \U$11992 ( \12678 , \12677 , \12665 );
not \U$11993 ( \12679 , \12678 );
and \U$11994 ( \12680 , \12673 , \12674 , \12679 );
buf \U$11995 ( \12681 , \12680 );
not \U$11996 ( \12682 , \12681 );
not \U$11997 ( \12683 , \12682 );
or \U$11998 ( \12684 , \12669 , \12683 );
not \U$11999 ( \12685 , \12357 );
buf \U$12000 ( \12686 , \12685 );
not \U$12001 ( \12687 , \12686 );
nand \U$12002 ( \12688 , \12684 , \12687 );
not \U$12003 ( \12689 , \12688 );
nand \U$12004 ( \12690 , \12649 , \12689 );
not \U$12005 ( \12691 , \12690 );
not \U$12006 ( \12692 , \12247 );
not \U$12007 ( \12693 , \12327 );
or \U$12008 ( \12694 , \12692 , \12693 );
nand \U$12009 ( \12695 , \12322 , \12411 );
nand \U$12010 ( \12696 , \12694 , \12695 );
not \U$12011 ( \12697 , \12696 );
not \U$12012 ( \12698 , \12520 );
not \U$12013 ( \12699 , \12698 );
or \U$12014 ( \12700 , \12697 , \12699 );
nand \U$12015 ( \12701 , \12002 , \12518 );
nand \U$12016 ( \12702 , \12700 , \12701 );
not \U$12017 ( \12703 , \12702 );
or \U$12018 ( \12704 , \12691 , \12703 );
not \U$12019 ( \12705 , \12689 );
nand \U$12020 ( \12706 , \12705 , \12648 );
nand \U$12021 ( \12707 , \12704 , \12706 );
nand \U$12022 ( \12708 , \12632 , \12489 );
and \U$12023 ( \12709 , \12707 , \12708 );
nor \U$12024 ( \12710 , \12635 , \12709 );
xor \U$12025 ( \12711 , \12500 , \12545 );
xor \U$12026 ( \12712 , \12711 , \12497 );
xor \U$12027 ( \12713 , \12710 , \12712 );
not \U$12028 ( \12714 , \11884 );
not \U$12029 ( \12715 , \12627 );
not \U$12030 ( \12716 , \12118 );
or \U$12031 ( \12717 , \12715 , \12716 );
nand \U$12032 ( \12718 , \12534 , \12626 );
nand \U$12033 ( \12719 , \12717 , \12718 );
not \U$12034 ( \12720 , \12719 );
or \U$12035 ( \12721 , \12714 , \12720 );
nand \U$12036 ( \12722 , \12536 , \12540 );
nand \U$12037 ( \12723 , \12721 , \12722 );
not \U$12038 ( \12724 , \12723 );
and \U$12039 ( \12725 , \12648 , \12689 );
not \U$12040 ( \12726 , \12648 );
and \U$12041 ( \12727 , \12726 , \12688 );
nor \U$12042 ( \12728 , \12725 , \12727 );
not \U$12043 ( \12729 , \12728 );
not \U$12044 ( \12730 , \12702 );
or \U$12045 ( \12731 , \12729 , \12730 );
not \U$12046 ( \12732 , \12702 );
not \U$12047 ( \12733 , \12728 );
nand \U$12048 ( \12734 , \12732 , \12733 );
nand \U$12049 ( \12735 , \12731 , \12734 );
not \U$12050 ( \12736 , \12735 );
or \U$12051 ( \12737 , \12724 , \12736 );
not \U$12052 ( \12738 , \12735 );
not \U$12053 ( \12739 , \12738 );
not \U$12054 ( \12740 , \12723 );
not \U$12055 ( \12741 , \12740 );
or \U$12056 ( \12742 , \12739 , \12741 );
not \U$12057 ( \12743 , \11949 );
not \U$12058 ( \12744 , \12637 );
or \U$12059 ( \12745 , \12743 , \12744 );
not \U$12060 ( \12746 , \12637 );
nand \U$12061 ( \12747 , \12746 , \11947 );
nand \U$12062 ( \12748 , \12745 , \12747 );
not \U$12063 ( \12749 , \12748 );
not \U$12064 ( \12750 , \12644 );
or \U$12065 ( \12751 , \12749 , \12750 );
nand \U$12066 ( \12752 , \12642 , \12364 );
nand \U$12067 ( \12753 , \12751 , \12752 );
not \U$12068 ( \12754 , \12198 );
not \U$12069 ( \12755 , \12302 );
or \U$12070 ( \12756 , \12754 , \12755 );
nand \U$12071 ( \12757 , \12137 , \12306 );
nand \U$12072 ( \12758 , \12756 , \12757 );
not \U$12073 ( \12759 , \12758 );
nand \U$12074 ( \12760 , \12159 , \12192 );
not \U$12075 ( \12761 , \12760 );
not \U$12076 ( \12762 , \12761 );
or \U$12077 ( \12763 , \12759 , \12762 );
not \U$12078 ( \12764 , \12106 );
not \U$12079 ( \12765 , \12198 );
or \U$12080 ( \12766 , \12764 , \12765 );
nand \U$12081 ( \12767 , \12383 , \12107 );
nand \U$12082 ( \12768 , \12766 , \12767 );
nand \U$12083 ( \12769 , \12768 , \12197 );
nand \U$12084 ( \12770 , \12763 , \12769 );
xor \U$12085 ( \12771 , \12753 , \12770 );
not \U$12086 ( \12772 , \12463 );
not \U$12087 ( \12773 , \12327 );
or \U$12088 ( \12774 , \12772 , \12773 );
nand \U$12089 ( \12775 , \12029 , \12464 );
nand \U$12090 ( \12776 , \12774 , \12775 );
not \U$12091 ( \12777 , \12776 );
not \U$12092 ( \12778 , \12520 );
not \U$12093 ( \12779 , \12778 );
or \U$12094 ( \12780 , \12777 , \12779 );
nand \U$12095 ( \12781 , \12002 , \12696 );
nand \U$12096 ( \12782 , \12780 , \12781 );
and \U$12097 ( \12783 , \12771 , \12782 );
and \U$12098 ( \12784 , \12753 , \12770 );
or \U$12099 ( \12785 , \12783 , \12784 );
buf \U$12100 ( \12786 , \12785 );
nand \U$12101 ( \12787 , \12742 , \12786 );
nand \U$12102 ( \12788 , \12737 , \12787 );
xor \U$12103 ( \12789 , \12513 , \12527 );
xor \U$12104 ( \12790 , \12789 , \12542 );
not \U$12105 ( \12791 , \12790 );
and \U$12106 ( \12792 , \11910 , RI9928738_416);
and \U$12107 ( \12793 , \11913 , RI9927dd8_436);
nor \U$12108 ( \12794 , \12792 , \12793 );
and \U$12109 ( \12795 , \11786 , RI9925768_496);
and \U$12110 ( \12796 , \11923 , RI9924778_516);
nor \U$12111 ( \12797 , \12795 , \12796 );
nand \U$12112 ( \12798 , \12794 , \12797 );
and \U$12113 ( \12799 , \11796 , RI9926a28_456);
and \U$12114 ( \12800 , \11917 , RI99260c8_476);
nor \U$12115 ( \12801 , \12799 , \12800 );
and \U$12116 ( \12802 , \11778 , RI9923e18_536);
and \U$12117 ( \12803 , \11775 , RI99234b8_556);
nor \U$12118 ( \12804 , \12802 , \12803 );
nand \U$12119 ( \12805 , \12801 , \12804 );
nor \U$12120 ( \12806 , \12798 , \12805 );
nand \U$12121 ( \12807 , \11743 , RI992cc98_336);
nand \U$12122 ( \12808 , \11826 , RI992b168_356);
nand \U$12123 ( \12809 , \11756 , RI9931798_276);
and \U$12124 ( \12810 , \11749 , RI9922888_576);
nand \U$12125 ( \12811 , \10843 , RI9935ed8_256);
not \U$12126 ( \12812 , \12811 );
nor \U$12127 ( \12813 , \12810 , \12812 );
nand \U$12128 ( \12814 , \12807 , \12808 , \12809 , \12813 );
nand \U$12129 ( \12815 , \11737 , RI992f4e8_296);
nand \U$12130 ( \12816 , \11734 , RI992a808_376);
nand \U$12131 ( \12817 , \11730 , RI992d5f8_316);
nand \U$12132 ( \12818 , \11726 , RI9929098_396);
nand \U$12133 ( \12819 , \12815 , \12816 , \12817 , \12818 );
nor \U$12134 ( \12820 , \12814 , \12819 );
nand \U$12135 ( \12821 , \12806 , \12820 );
not \U$12136 ( \12822 , \12821 );
not \U$12137 ( \12823 , \12822 );
not \U$12138 ( \12824 , \11639 );
and \U$12139 ( \12825 , \12823 , \12824 );
not \U$12140 ( \12826 , \12823 );
buf \U$12141 ( \12827 , \11634 );
not \U$12142 ( \12828 , \12827 );
and \U$12143 ( \12829 , \12826 , \12828 );
nor \U$12144 ( \12830 , \12825 , \12829 );
nand \U$12145 ( \12831 , \11638 , \12830 );
not \U$12146 ( \12832 , \12831 );
not \U$12147 ( \12833 , \12768 );
not \U$12148 ( \12834 , \12194 );
or \U$12149 ( \12835 , \12833 , \12834 );
buf \U$12150 ( \12836 , \12192 );
not \U$12151 ( \12837 , \12836 );
nand \U$12152 ( \12838 , \12837 , \12508 );
nand \U$12153 ( \12839 , \12835 , \12838 );
not \U$12154 ( \12840 , \12839 );
not \U$12155 ( \12841 , \12840 );
or \U$12156 ( \12842 , \12832 , \12841 );
not \U$12157 ( \12843 , \11839 );
not \U$12158 ( \12844 , \12686 );
or \U$12159 ( \12845 , \12843 , \12844 );
not \U$12160 ( \12846 , \12686 );
nand \U$12161 ( \12847 , \12846 , \11840 );
nand \U$12162 ( \12848 , \12845 , \12847 );
not \U$12163 ( \12849 , \12848 );
buf \U$12164 ( \12850 , \12681 );
not \U$12165 ( \12851 , \12850 );
or \U$12166 ( \12852 , \12849 , \12851 );
nand \U$12167 ( \12853 , \12667 , \12687 );
nand \U$12168 ( \12854 , \12852 , \12853 );
buf \U$12169 ( \12855 , \12854 );
nand \U$12170 ( \12856 , \12842 , \12855 );
not \U$12171 ( \12857 , \12831 );
nand \U$12172 ( \12858 , \12857 , \12839 );
and \U$12173 ( \12859 , \12856 , \12858 );
nand \U$12174 ( \12860 , \12791 , \12859 );
and \U$12175 ( \12861 , \12788 , \12860 );
nor \U$12176 ( \12862 , \12791 , \12859 );
nor \U$12177 ( \12863 , \12861 , \12862 );
and \U$12178 ( \12864 , \12713 , \12863 );
and \U$12179 ( \12865 , \12710 , \12712 );
or \U$12180 ( \12866 , \12864 , \12865 );
xor \U$12181 ( \12867 , \12319 , \12492 );
xnor \U$12182 ( \12868 , \12867 , \12549 );
nand \U$12183 ( \12869 , \12866 , \12868 );
nand \U$12184 ( \12870 , \12598 , \12869 );
xor \U$12185 ( \12871 , \12555 , \12559 );
and \U$12186 ( \12872 , \12871 , \12595 );
and \U$12187 ( \12873 , \12555 , \12559 );
or \U$12188 ( \12874 , \12872 , \12873 );
not \U$12189 ( \12875 , \12579 );
not \U$12190 ( \12876 , \12589 );
or \U$12191 ( \12877 , \12875 , \12876 );
or \U$12192 ( \12878 , \12589 , \12579 );
not \U$12193 ( \12879 , \12575 );
nand \U$12194 ( \12880 , \12878 , \12879 );
nand \U$12195 ( \12881 , \12877 , \12880 );
not \U$12196 ( \12882 , \12881 );
xor \U$12197 ( \12883 , \12113 , \12055 );
xor \U$12198 ( \12884 , \12883 , \12126 );
not \U$12199 ( \12885 , \12884 );
not \U$12200 ( \12886 , \12885 );
or \U$12201 ( \12887 , \12882 , \12886 );
not \U$12202 ( \12888 , \12881 );
nand \U$12203 ( \12889 , \12884 , \12888 );
nand \U$12204 ( \12890 , \12887 , \12889 );
nand \U$12205 ( \12891 , \12341 , \12565 );
not \U$12206 ( \12892 , \12891 );
not \U$12207 ( \12893 , \12594 );
not \U$12208 ( \12894 , \12893 );
or \U$12209 ( \12895 , \12892 , \12894 );
not \U$12210 ( \12896 , \12565 );
nand \U$12211 ( \12897 , \12896 , \12340 );
nand \U$12212 ( \12898 , \12895 , \12897 );
xor \U$12213 ( \12899 , \12890 , \12898 );
nor \U$12214 ( \12900 , \12874 , \12899 );
nor \U$12215 ( \12901 , \12870 , \12900 );
nand \U$12216 ( \12902 , \12885 , \12888 );
nand \U$12217 ( \12903 , \12898 , \12902 );
nand \U$12218 ( \12904 , \12884 , \12881 );
and \U$12219 ( \12905 , \12903 , \12904 );
not \U$12220 ( \12906 , \12055 );
not \U$12221 ( \12907 , \12052 );
or \U$12222 ( \12908 , \12906 , \12907 );
nand \U$12223 ( \12909 , \12051 , \12042 );
nand \U$12224 ( \12910 , \12908 , \12909 );
xnor \U$12225 ( \12911 , \12910 , \12129 );
nand \U$12226 ( \12912 , \12905 , \12911 );
nand \U$12227 ( \12913 , \12901 , \12912 );
buf \U$12228 ( \12914 , \11241 );
or \U$12229 ( \12915 , \12914 , \11102 );
buf \U$12230 ( \12916 , \11242 );
nand \U$12231 ( \12917 , \12915 , \12916 );
and \U$12232 ( \12918 , \11186 , \11191 , \11222 , \11211 );
and \U$12233 ( \12919 , \11228 , \11198 , \11216 , \11203 );
nand \U$12234 ( \12920 , \12918 , \12919 );
nand \U$12235 ( \12921 , \12920 , \11231 );
not \U$12236 ( \12922 , \12921 );
and \U$12237 ( \12923 , \12917 , \12922 );
not \U$12238 ( \12924 , \12917 );
and \U$12239 ( \12925 , \12924 , \12921 );
nor \U$12240 ( \12926 , \12923 , \12925 );
not \U$12241 ( \12927 , \11248 );
nand \U$12242 ( \12928 , \12927 , \11107 );
buf \U$12243 ( \12929 , \11243 );
not \U$12244 ( \12930 , \12929 );
and \U$12245 ( \12931 , \12928 , \12930 );
not \U$12246 ( \12932 , \12928 );
and \U$12247 ( \12933 , \12932 , \12929 );
nor \U$12248 ( \12934 , \12931 , \12933 );
xnor \U$12249 ( \12935 , \12926 , \12934 );
not \U$12250 ( \12936 , \12935 );
not \U$12251 ( \12937 , \12936 );
not \U$12252 ( \12938 , \12937 );
not \U$12253 ( \12939 , \12934 );
not \U$12254 ( \12940 , \12939 );
not \U$12255 ( \12941 , \12940 );
not \U$12256 ( \12942 , \12660 );
not \U$12257 ( \12943 , \12942 );
or \U$12258 ( \12944 , \12941 , \12943 );
nand \U$12259 ( \12945 , \12939 , \12660 );
nand \U$12260 ( \12946 , \12944 , \12945 );
nand \U$12261 ( \12947 , \12946 , \12935 );
not \U$12262 ( \12948 , \12947 );
or \U$12263 ( \12949 , \12938 , \12948 );
buf \U$12264 ( \12950 , \12942 );
not \U$12265 ( \12951 , \12950 );
nand \U$12266 ( \12952 , \12949 , \12951 );
not \U$12267 ( \12953 , \11763 );
not \U$12268 ( \12954 , \12686 );
or \U$12269 ( \12955 , \12953 , \12954 );
buf \U$12270 ( \12956 , \12357 );
nand \U$12271 ( \12957 , \12956 , \12640 );
nand \U$12272 ( \12958 , \12955 , \12957 );
not \U$12273 ( \12959 , \12958 );
not \U$12274 ( \12960 , \12850 );
or \U$12275 ( \12961 , \12959 , \12960 );
nand \U$12276 ( \12962 , \12848 , \12667 );
nand \U$12277 ( \12963 , \12961 , \12962 );
xor \U$12278 ( \12964 , \12952 , \12963 );
not \U$12279 ( \12965 , \12108 );
not \U$12280 ( \12966 , \12637 );
or \U$12281 ( \12967 , \12965 , \12966 );
not \U$12282 ( \12968 , \12186 );
nand \U$12283 ( \12969 , \12968 , \12107 );
nand \U$12284 ( \12970 , \12967 , \12969 );
not \U$12285 ( \12971 , \12970 );
not \U$12286 ( \12972 , \12375 );
or \U$12287 ( \12973 , \12971 , \12972 );
nand \U$12288 ( \12974 , \12365 , \12748 );
nand \U$12289 ( \12975 , \12973 , \12974 );
xor \U$12290 ( \12976 , \12964 , \12975 );
not \U$12291 ( \12977 , \12937 );
not \U$12292 ( \12978 , \12950 );
and \U$12293 ( \12979 , \12977 , \12978 );
not \U$12294 ( \12980 , \12947 );
not \U$12295 ( \12981 , \11839 );
not \U$12296 ( \12982 , \12950 );
or \U$12297 ( \12983 , \12981 , \12982 );
nand \U$12298 ( \12984 , \11840 , \12951 );
nand \U$12299 ( \12985 , \12983 , \12984 );
and \U$12300 ( \12986 , \12980 , \12985 );
nor \U$12301 ( \12987 , \12979 , \12986 );
not \U$12302 ( \12988 , \12197 );
not \U$12303 ( \12989 , \12758 );
or \U$12304 ( \12990 , \12988 , \12989 );
not \U$12305 ( \12991 , \12247 );
not \U$12306 ( \12992 , \12383 );
not \U$12307 ( \12993 , \12992 );
or \U$12308 ( \12994 , \12991 , \12993 );
nand \U$12309 ( \12995 , \12137 , \12411 );
nand \U$12310 ( \12996 , \12994 , \12995 );
nand \U$12311 ( \12997 , \12996 , \12159 , \12836 );
nand \U$12312 ( \12998 , \12990 , \12997 );
xor \U$12313 ( \12999 , \12987 , \12998 );
not \U$12314 ( \13000 , \12627 );
not \U$12315 ( \13001 , \12323 );
or \U$12316 ( \13002 , \13000 , \13001 );
nand \U$12317 ( \13003 , \12326 , \12626 );
nand \U$12318 ( \13004 , \13002 , \13003 );
not \U$12319 ( \13005 , \13004 );
not \U$12320 ( \13006 , \12399 );
or \U$12321 ( \13007 , \13005 , \13006 );
nand \U$12322 ( \13008 , \12003 , \12776 );
nand \U$12323 ( \13009 , \13007 , \13008 );
xnor \U$12324 ( \13010 , \12999 , \13009 );
or \U$12325 ( \13011 , \12976 , \13010 );
not \U$12326 ( \13012 , \12823 );
not \U$12327 ( \13013 , \12327 );
or \U$12328 ( \13014 , \13012 , \13013 );
nand \U$12329 ( \13015 , \12322 , \12822 );
nand \U$12330 ( \13016 , \13014 , \13015 );
not \U$12331 ( \13017 , \13016 );
not \U$12332 ( \13018 , \12016 );
or \U$12333 ( \13019 , \13017 , \13018 );
nand \U$12334 ( \13020 , \12002 , \13004 );
nand \U$12335 ( \13021 , \13019 , \13020 );
not \U$12336 ( \13022 , \13021 );
not \U$12337 ( \13023 , \12463 );
not \U$12338 ( \13024 , \12154 );
or \U$12339 ( \13025 , \13023 , \13024 );
nand \U$12340 ( \13026 , \12137 , \12464 );
nand \U$12341 ( \13027 , \13025 , \13026 );
not \U$12342 ( \13028 , \13027 );
not \U$12343 ( \13029 , \12194 );
or \U$12344 ( \13030 , \13028 , \13029 );
nand \U$12345 ( \13031 , \12837 , \12996 );
nand \U$12346 ( \13032 , \13030 , \13031 );
not \U$12347 ( \13033 , \13032 );
or \U$12348 ( \13034 , \13022 , \13033 );
or \U$12349 ( \13035 , \13032 , \13021 );
not \U$12350 ( \13036 , \11763 );
not \U$12351 ( \13037 , \12662 );
not \U$12352 ( \13038 , \13037 );
or \U$12353 ( \13039 , \13036 , \13038 );
nand \U$12354 ( \13040 , \12951 , \12640 );
nand \U$12355 ( \13041 , \13039 , \13040 );
not \U$12356 ( \13042 , \13041 );
not \U$12357 ( \13043 , \12980 );
or \U$12358 ( \13044 , \13042 , \13043 );
buf \U$12359 ( \13045 , \12936 );
nand \U$12360 ( \13046 , \12985 , \13045 );
nand \U$12361 ( \13047 , \13044 , \13046 );
buf \U$12362 ( \13048 , \12926 );
not \U$12363 ( \13049 , \13048 );
buf \U$12364 ( \13050 , \13049 );
or \U$12365 ( \13051 , \13047 , \13050 );
nand \U$12366 ( \13052 , \13035 , \13051 );
nand \U$12367 ( \13053 , \13034 , \13052 );
nand \U$12368 ( \13054 , \13011 , \13053 );
nand \U$12369 ( \13055 , \13010 , \12976 );
nand \U$12370 ( \13056 , \13054 , \13055 );
not \U$12371 ( \13057 , \11705 );
not \U$12372 ( \13058 , \2302 );
and \U$12373 ( \13059 , \13057 , \13058 );
nor \U$12374 ( \13060 , \11699 , \2327 );
nor \U$12375 ( \13061 , \13059 , \13060 );
not \U$12376 ( \13062 , \11801 );
not \U$12377 ( \13063 , \13062 );
not \U$12378 ( \13064 , \2285 );
and \U$12379 ( \13065 , \13063 , \13064 );
nor \U$12380 ( \13066 , \12211 , \7477 );
nor \U$12381 ( \13067 , \13065 , \13066 );
nand \U$12382 ( \13068 , \13061 , \13067 );
not \U$12383 ( \13069 , \11674 );
not \U$12384 ( \13070 , \2317 );
and \U$12385 ( \13071 , \13069 , \13070 );
nor \U$12386 ( \13072 , \11681 , \2320 );
nor \U$12387 ( \13073 , \13071 , \13072 );
not \U$12388 ( \13074 , \11710 );
not \U$12389 ( \13075 , \7448 );
and \U$12390 ( \13076 , \13074 , \13075 );
nor \U$12391 ( \13077 , \11715 , \7451 );
nor \U$12392 ( \13078 , \13076 , \13077 );
nand \U$12393 ( \13079 , \13073 , \13078 );
nor \U$12394 ( \13080 , \13068 , \13079 );
nand \U$12395 ( \13081 , \11726 , RI9928fa8_398);
nand \U$12396 ( \13082 , \11730 , RI992d508_318);
nand \U$12397 ( \13083 , \11734 , RI992a718_378);
nand \U$12398 ( \13084 , \11737 , RI992f3f8_298);
nand \U$12399 ( \13085 , \13081 , \13082 , \13083 , \13084 );
and \U$12400 ( \13086 , \11743 , RI992cba8_338);
not \U$12401 ( \13087 , RI9922798_578);
not \U$12402 ( \13088 , \11749 );
or \U$12403 ( \13089 , \13087 , \13088 );
nand \U$12404 ( \13090 , \10843 , RI9933d18_258);
nand \U$12405 ( \13091 , \13089 , \13090 );
nor \U$12406 ( \13092 , \13086 , \13091 );
nand \U$12407 ( \13093 , \11756 , RI99316a8_278);
nand \U$12408 ( \13094 , \11826 , RI992b078_358);
nand \U$12409 ( \13095 , \13092 , \13093 , \13094 );
nor \U$12410 ( \13096 , \13085 , \13095 );
nand \U$12411 ( \13097 , \13080 , \13096 );
buf \U$12412 ( \13098 , \13097 );
not \U$12413 ( \13099 , \13098 );
not \U$12414 ( \13100 , \11889 );
or \U$12415 ( \13101 , \13099 , \13100 );
not \U$12416 ( \13102 , \13098 );
nand \U$12417 ( \13103 , \12532 , \13102 );
nand \U$12418 ( \13104 , \13101 , \13103 );
not \U$12419 ( \13105 , \13104 );
not \U$12420 ( \13106 , \11884 );
or \U$12421 ( \13107 , \13105 , \13106 );
not \U$12422 ( \13108 , \11705 );
not \U$12423 ( \13109 , \2391 );
and \U$12424 ( \13110 , \13108 , \13109 );
nor \U$12425 ( \13111 , \11699 , \2365 );
nor \U$12426 ( \13112 , \13110 , \13111 );
not \U$12427 ( \13113 , \13062 );
not \U$12428 ( \13114 , \2376 );
and \U$12429 ( \13115 , \13113 , \13114 );
nor \U$12430 ( \13116 , \11692 , \7268 );
nor \U$12431 ( \13117 , \13115 , \13116 );
nand \U$12432 ( \13118 , \13112 , \13117 );
not \U$12433 ( \13119 , \11681 );
not \U$12434 ( \13120 , \2349 );
and \U$12435 ( \13121 , \13119 , \13120 );
nor \U$12436 ( \13122 , \11674 , \2346 );
nor \U$12437 ( \13123 , \13121 , \13122 );
not \U$12438 ( \13124 , \11710 );
not \U$12439 ( \13125 , \7283 );
and \U$12440 ( \13126 , \13124 , \13125 );
nor \U$12441 ( \13127 , \11715 , \7285 );
nor \U$12442 ( \13128 , \13126 , \13127 );
nand \U$12443 ( \13129 , \13123 , \13128 );
nor \U$12444 ( \13130 , \13118 , \13129 );
nand \U$12445 ( \13131 , \11737 , RI992f470_297);
nand \U$12446 ( \13132 , \11730 , RI992d580_317);
nand \U$12447 ( \13133 , \11734 , RI992a790_377);
nand \U$12448 ( \13134 , \11726 , RI9929020_397);
nand \U$12449 ( \13135 , \13131 , \13132 , \13133 , \13134 );
and \U$12450 ( \13136 , \11743 , RI992cc20_337);
not \U$12451 ( \13137 , RI9922810_577);
not \U$12452 ( \13138 , \11749 );
or \U$12453 ( \13139 , \13137 , \13138 );
nand \U$12454 ( \13140 , \10843 , RI9933d90_257);
nand \U$12455 ( \13141 , \13139 , \13140 );
nor \U$12456 ( \13142 , \13136 , \13141 );
nand \U$12457 ( \13143 , \11756 , RI9931720_277);
nand \U$12458 ( \13144 , \11759 , RI992b0f0_357);
nand \U$12459 ( \13145 , \13142 , \13143 , \13144 );
nor \U$12460 ( \13146 , \13135 , \13145 );
nand \U$12461 ( \13147 , \13130 , \13146 );
not \U$12462 ( \13148 , \13147 );
not \U$12463 ( \13149 , \13148 );
not \U$12464 ( \13150 , \13149 );
not \U$12465 ( \13151 , \12118 );
or \U$12466 ( \13152 , \13150 , \13151 );
nand \U$12467 ( \13153 , \11890 , \13148 );
nand \U$12468 ( \13154 , \13152 , \13153 );
nand \U$12469 ( \13155 , \13154 , \12540 );
nand \U$12470 ( \13156 , \13107 , \13155 );
not \U$12471 ( \13157 , \11705 );
not \U$12472 ( \13158 , \2424 );
and \U$12473 ( \13159 , \13157 , \13158 );
not \U$12474 ( \13160 , RI9923cb0_539);
nor \U$12475 ( \13161 , \11699 , \13160 );
nor \U$12476 ( \13162 , \13159 , \13161 );
not \U$12477 ( \13163 , RI9927c70_439);
nor \U$12478 ( \13164 , \13163 , \12427 );
not \U$12479 ( \13165 , RI99285d0_419);
nor \U$12480 ( \13166 , \13165 , \11692 );
nor \U$12481 ( \13167 , \13164 , \13166 );
nand \U$12482 ( \13168 , \13162 , \13167 );
not \U$12483 ( \13169 , \11681 );
not \U$12484 ( \13170 , \7628 );
and \U$12485 ( \13171 , \13169 , \13170 );
not \U$12486 ( \13172 , RI99268c0_459);
nor \U$12487 ( \13173 , \11674 , \13172 );
nor \U$12488 ( \13174 , \13171 , \13173 );
not \U$12489 ( \13175 , \11710 );
not \U$12490 ( \13176 , RI9924610_519);
not \U$12491 ( \13177 , \13176 );
and \U$12492 ( \13178 , \13175 , \13177 );
not \U$12493 ( \13179 , RI9925600_499);
nor \U$12494 ( \13180 , \11715 , \13179 );
nor \U$12495 ( \13181 , \13178 , \13180 );
nand \U$12496 ( \13182 , \13174 , \13181 );
nor \U$12497 ( \13183 , \13168 , \13182 );
nand \U$12498 ( \13184 , \11737 , RI992f380_299);
nand \U$12499 ( \13185 , \11816 , RI992d490_319);
nand \U$12500 ( \13186 , \11734 , RI992a6a0_379);
nand \U$12501 ( \13187 , \11726 , RI9928f30_399);
nand \U$12502 ( \13188 , \13184 , \13185 , \13186 , \13187 );
and \U$12503 ( \13189 , \11743 , RI992cb30_339);
nand \U$12504 ( \13190 , \11749 , RI9922720_579);
nand \U$12505 ( \13191 , \10843 , RI9933ca0_259);
nand \U$12506 ( \13192 , \13190 , \13191 );
nor \U$12507 ( \13193 , \13189 , \13192 );
nand \U$12508 ( \13194 , \11756 , RI9931630_279);
nand \U$12509 ( \13195 , \11759 , RI992b000_359);
nand \U$12510 ( \13196 , \13193 , \13194 , \13195 );
nor \U$12511 ( \13197 , \13188 , \13196 );
nand \U$12512 ( \13198 , \13183 , \13197 );
buf \U$12513 ( \13199 , \13198 );
and \U$12514 ( \13200 , \13199 , \12467 );
not \U$12515 ( \13201 , \13199 );
and \U$12516 ( \13202 , \13201 , \12828 );
nor \U$12517 ( \13203 , \13200 , \13202 );
nand \U$12518 ( \13204 , \11637 , \13203 );
not \U$12519 ( \13205 , \13204 );
or \U$12520 ( \13206 , \13156 , \13205 );
not \U$12521 ( \13207 , \12247 );
not \U$12522 ( \13208 , \12637 );
or \U$12523 ( \13209 , \13207 , \13208 );
nand \U$12524 ( \13210 , \12189 , \12411 );
nand \U$12525 ( \13211 , \13209 , \13210 );
not \U$12526 ( \13212 , \13211 );
not \U$12527 ( \13213 , \12644 );
or \U$12528 ( \13214 , \13212 , \13213 );
not \U$12529 ( \13215 , \12302 );
not \U$12530 ( \13216 , \12637 );
or \U$12531 ( \13217 , \13215 , \13216 );
nand \U$12532 ( \13218 , \12968 , \12306 );
nand \U$12533 ( \13219 , \13217 , \13218 );
nand \U$12534 ( \13220 , \13219 , \12364 );
nand \U$12535 ( \13221 , \13214 , \13220 );
not \U$12536 ( \13222 , \13221 );
not \U$12537 ( \13223 , \12106 );
not \U$12538 ( \13224 , \12956 );
not \U$12539 ( \13225 , \13224 );
or \U$12540 ( \13226 , \13223 , \13225 );
nand \U$12541 ( \13227 , \12107 , \12956 );
nand \U$12542 ( \13228 , \13226 , \13227 );
not \U$12543 ( \13229 , \13228 );
not \U$12544 ( \13230 , \12681 );
or \U$12545 ( \13231 , \13229 , \13230 );
not \U$12546 ( \13232 , \11949 );
not \U$12547 ( \13233 , \13224 );
or \U$12548 ( \13234 , \13232 , \13233 );
nand \U$12549 ( \13235 , \12956 , \11947 );
nand \U$12550 ( \13236 , \13234 , \13235 );
nand \U$12551 ( \13237 , \13236 , \12667 );
nand \U$12552 ( \13238 , \13231 , \13237 );
not \U$12553 ( \13239 , \13238 );
nand \U$12554 ( \13240 , \13222 , \13239 );
buf \U$12555 ( \13241 , \12661 );
and \U$12556 ( \13242 , \11946 , \13241 );
not \U$12557 ( \13243 , \11946 );
not \U$12558 ( \13244 , \13241 );
and \U$12559 ( \13245 , \13243 , \13244 );
or \U$12560 ( \13246 , \13242 , \13245 );
not \U$12561 ( \13247 , \13246 );
and \U$12562 ( \13248 , \12946 , \12935 );
not \U$12563 ( \13249 , \13248 );
or \U$12564 ( \13250 , \13247 , \13249 );
not \U$12565 ( \13251 , \12935 );
nand \U$12566 ( \13252 , \13041 , \13251 );
nand \U$12567 ( \13253 , \13250 , \13252 );
nor \U$12568 ( \13254 , \12920 , \11231 );
not \U$12569 ( \13255 , \13254 );
nand \U$12570 ( \13256 , \13255 , \12921 );
not \U$12571 ( \13257 , \13256 );
nand \U$12572 ( \13258 , \13257 , \13048 );
not \U$12573 ( \13259 , \13258 );
not \U$12574 ( \13260 , \13259 );
not \U$12575 ( \13261 , \13048 );
and \U$12576 ( \13262 , \11838 , \13261 );
not \U$12577 ( \13263 , \11838 );
not \U$12578 ( \13264 , \13049 );
and \U$12579 ( \13265 , \13263 , \13264 );
or \U$12580 ( \13266 , \13262 , \13265 );
not \U$12581 ( \13267 , \13266 );
or \U$12582 ( \13268 , \13260 , \13267 );
not \U$12583 ( \13269 , \13050 );
buf \U$12584 ( \13270 , \13256 );
nand \U$12585 ( \13271 , \13269 , \13270 );
nand \U$12586 ( \13272 , \13268 , \13271 );
nand \U$12587 ( \13273 , \13253 , \13272 );
not \U$12588 ( \13274 , \13273 );
and \U$12589 ( \13275 , \13240 , \13274 );
and \U$12590 ( \13276 , \13221 , \13238 );
nor \U$12591 ( \13277 , \13275 , \13276 );
not \U$12592 ( \13278 , \13277 );
nand \U$12593 ( \13279 , \13206 , \13278 );
nand \U$12594 ( \13280 , \13156 , \13205 );
nand \U$12595 ( \13281 , \13279 , \13280 );
and \U$12596 ( \13282 , \13098 , \12824 );
not \U$12597 ( \13283 , \13098 );
and \U$12598 ( \13284 , \13283 , \11639 );
nor \U$12599 ( \13285 , \13282 , \13284 );
nand \U$12600 ( \13286 , \11637 , \13285 );
not \U$12601 ( \13287 , \13154 );
not \U$12602 ( \13288 , \11884 );
or \U$12603 ( \13289 , \13287 , \13288 );
not \U$12604 ( \13290 , \12823 );
not \U$12605 ( \13291 , \12533 );
or \U$12606 ( \13292 , \13290 , \13291 );
nand \U$12607 ( \13293 , \11890 , \12822 );
nand \U$12608 ( \13294 , \13292 , \13293 );
nand \U$12609 ( \13295 , \13294 , \12540 );
nand \U$12610 ( \13296 , \13289 , \13295 );
xor \U$12611 ( \13297 , \13286 , \13296 );
not \U$12612 ( \13298 , \13236 );
not \U$12613 ( \13299 , \12850 );
or \U$12614 ( \13300 , \13298 , \13299 );
nand \U$12615 ( \13301 , \12958 , \12667 );
nand \U$12616 ( \13302 , \13300 , \13301 );
xor \U$12617 ( \13303 , \12987 , \13302 );
not \U$12618 ( \13304 , \13219 );
not \U$12619 ( \13305 , \12375 );
or \U$12620 ( \13306 , \13304 , \13305 );
buf \U$12621 ( \13307 , \12363 );
not \U$12622 ( \13308 , \13307 );
nand \U$12623 ( \13309 , \12970 , \13308 );
nand \U$12624 ( \13310 , \13306 , \13309 );
and \U$12625 ( \13311 , \13303 , \13310 );
and \U$12626 ( \13312 , \12987 , \13302 );
or \U$12627 ( \13313 , \13311 , \13312 );
xnor \U$12628 ( \13314 , \13297 , \13313 );
xor \U$12629 ( \13315 , \13281 , \13314 );
xor \U$12630 ( \13316 , \13051 , \13021 );
xnor \U$12631 ( \13317 , \13316 , \13032 );
xor \U$12632 ( \13318 , \12987 , \13302 );
xor \U$12633 ( \13319 , \13318 , \13310 );
not \U$12634 ( \13320 , \13319 );
nand \U$12635 ( \13321 , \13317 , \13320 );
not \U$12636 ( \13322 , \13321 );
not \U$12637 ( \13323 , \13047 );
not \U$12638 ( \13324 , \13050 );
or \U$12639 ( \13325 , \13323 , \13324 );
nand \U$12640 ( \13326 , \13325 , \13051 );
not \U$12641 ( \13327 , \12627 );
not \U$12642 ( \13328 , \12198 );
or \U$12643 ( \13329 , \13327 , \13328 );
nand \U$12644 ( \13330 , \12383 , \12626 );
nand \U$12645 ( \13331 , \13329 , \13330 );
not \U$12646 ( \13332 , \13331 );
not \U$12647 ( \13333 , \12194 );
or \U$12648 ( \13334 , \13332 , \13333 );
nand \U$12649 ( \13335 , \13027 , \12197 );
nand \U$12650 ( \13336 , \13334 , \13335 );
xor \U$12651 ( \13337 , \13326 , \13336 );
not \U$12652 ( \13338 , \13149 );
not \U$12653 ( \13339 , \12323 );
or \U$12654 ( \13340 , \13338 , \13339 );
nand \U$12655 ( \13341 , \12322 , \13148 );
nand \U$12656 ( \13342 , \13340 , \13341 );
not \U$12657 ( \13343 , \13342 );
not \U$12658 ( \13344 , \12038 );
or \U$12659 ( \13345 , \13343 , \13344 );
nand \U$12660 ( \13346 , \12003 , \13016 );
nand \U$12661 ( \13347 , \13345 , \13346 );
and \U$12662 ( \13348 , \13337 , \13347 );
and \U$12663 ( \13349 , \13326 , \13336 );
or \U$12664 ( \13350 , \13348 , \13349 );
not \U$12665 ( \13351 , \13350 );
or \U$12666 ( \13352 , \13322 , \13351 );
not \U$12667 ( \13353 , \13320 );
not \U$12668 ( \13354 , \13317 );
nand \U$12669 ( \13355 , \13353 , \13354 );
nand \U$12670 ( \13356 , \13352 , \13355 );
and \U$12671 ( \13357 , \13315 , \13356 );
and \U$12672 ( \13358 , \13281 , \13314 );
or \U$12673 ( \13359 , \13357 , \13358 );
xor \U$12674 ( \13360 , \13056 , \13359 );
xor \U$12675 ( \13361 , \12952 , \12963 );
and \U$12676 ( \13362 , \13361 , \12975 );
and \U$12677 ( \13363 , \12952 , \12963 );
or \U$12678 ( \13364 , \13362 , \13363 );
xor \U$12679 ( \13365 , \12753 , \12770 );
xor \U$12680 ( \13366 , \13365 , \12782 );
xor \U$12681 ( \13367 , \13364 , \13366 );
not \U$12682 ( \13368 , \12998 );
nand \U$12683 ( \13369 , \13368 , \12987 );
not \U$12684 ( \13370 , \13369 );
not \U$12685 ( \13371 , \13009 );
or \U$12686 ( \13372 , \13370 , \13371 );
not \U$12687 ( \13373 , \12987 );
nand \U$12688 ( \13374 , \13373 , \12998 );
nand \U$12689 ( \13375 , \13372 , \13374 );
xor \U$12690 ( \13376 , \13367 , \13375 );
not \U$12691 ( \13377 , \13376 );
not \U$12692 ( \13378 , \13294 );
not \U$12693 ( \13379 , \11884 );
or \U$12694 ( \13380 , \13378 , \13379 );
nand \U$12695 ( \13381 , \12719 , \12540 );
nand \U$12696 ( \13382 , \13380 , \13381 );
xor \U$12697 ( \13383 , \12854 , \13382 );
and \U$12698 ( \13384 , \13149 , \12824 );
not \U$12699 ( \13385 , \13149 );
and \U$12700 ( \13386 , \13385 , \11639 );
nor \U$12701 ( \13387 , \13384 , \13386 );
nand \U$12702 ( \13388 , \11638 , \13387 );
xnor \U$12703 ( \13389 , \13383 , \13388 );
not \U$12704 ( \13390 , \13389 );
not \U$12705 ( \13391 , \13286 );
not \U$12706 ( \13392 , \13391 );
not \U$12707 ( \13393 , \13296 );
or \U$12708 ( \13394 , \13392 , \13393 );
not \U$12709 ( \13395 , \13286 );
not \U$12710 ( \13396 , \13296 );
not \U$12711 ( \13397 , \13396 );
or \U$12712 ( \13398 , \13395 , \13397 );
nand \U$12713 ( \13399 , \13398 , \13313 );
nand \U$12714 ( \13400 , \13394 , \13399 );
not \U$12715 ( \13401 , \13400 );
and \U$12716 ( \13402 , \13390 , \13401 );
and \U$12717 ( \13403 , \13389 , \13400 );
nor \U$12718 ( \13404 , \13402 , \13403 );
not \U$12719 ( \13405 , \13404 );
or \U$12720 ( \13406 , \13377 , \13405 );
or \U$12721 ( \13407 , \13404 , \13376 );
nand \U$12722 ( \13408 , \13406 , \13407 );
and \U$12723 ( \13409 , \13360 , \13408 );
and \U$12724 ( \13410 , \13056 , \13359 );
or \U$12725 ( \13411 , \13409 , \13410 );
xor \U$12726 ( \13412 , \13364 , \13366 );
and \U$12727 ( \13413 , \13412 , \13375 );
and \U$12728 ( \13414 , \13364 , \13366 );
or \U$12729 ( \13415 , \13413 , \13414 );
not \U$12730 ( \13416 , \12855 );
not \U$12731 ( \13417 , \13388 );
or \U$12732 ( \13418 , \13416 , \13417 );
nand \U$12733 ( \13419 , \13418 , \13382 );
or \U$12734 ( \13420 , \13388 , \12855 );
nand \U$12735 ( \13421 , \13419 , \13420 );
xor \U$12736 ( \13422 , \12854 , \12839 );
xnor \U$12737 ( \13423 , \13422 , \12831 );
xor \U$12738 ( \13424 , \13421 , \13423 );
not \U$12739 ( \13425 , \13424 );
not \U$12740 ( \13426 , \13425 );
xor \U$12741 ( \13427 , \12723 , \12785 );
xnor \U$12742 ( \13428 , \13427 , \12735 );
not \U$12743 ( \13429 , \13428 );
not \U$12744 ( \13430 , \13429 );
or \U$12745 ( \13431 , \13426 , \13430 );
nand \U$12746 ( \13432 , \13428 , \13424 );
nand \U$12747 ( \13433 , \13431 , \13432 );
xor \U$12748 ( \13434 , \13415 , \13433 );
not \U$12749 ( \13435 , \13400 );
nand \U$12750 ( \13436 , \13435 , \13389 );
not \U$12751 ( \13437 , \13436 );
not \U$12752 ( \13438 , \13376 );
or \U$12753 ( \13439 , \13437 , \13438 );
not \U$12754 ( \13440 , \13389 );
nand \U$12755 ( \13441 , \13440 , \13400 );
nand \U$12756 ( \13442 , \13439 , \13441 );
not \U$12757 ( \13443 , \13442 );
xnor \U$12758 ( \13444 , \13434 , \13443 );
nor \U$12759 ( \13445 , \13411 , \13444 );
xor \U$12760 ( \13446 , \13281 , \13314 );
xor \U$12761 ( \13447 , \13446 , \13356 );
xor \U$12762 ( \13448 , \12976 , \13053 );
xnor \U$12763 ( \13449 , \13448 , \13010 );
not \U$12764 ( \13450 , \13449 );
or \U$12765 ( \13451 , \13447 , \13450 );
and \U$12766 ( \13452 , \11881 , \11882 );
not \U$12767 ( \13453 , \13452 );
not \U$12768 ( \13454 , \13199 );
not \U$12769 ( \13455 , \12533 );
or \U$12770 ( \13456 , \13454 , \13455 );
not \U$12771 ( \13457 , \13199 );
nand \U$12772 ( \13458 , \12532 , \13457 );
nand \U$12773 ( \13459 , \13456 , \13458 );
not \U$12774 ( \13460 , \13459 );
or \U$12775 ( \13461 , \13453 , \13460 );
nand \U$12776 ( \13462 , \13104 , \11873 );
nand \U$12777 ( \13463 , \13461 , \13462 );
not \U$12778 ( \13464 , \13463 );
and \U$12779 ( \13465 , \11910 , RI9928558_420);
not \U$12780 ( \13466 , \11912 );
and \U$12781 ( \13467 , \13466 , RI9927bf8_440);
nor \U$12782 ( \13468 , \13465 , \13467 );
and \U$12783 ( \13469 , \11786 , RI9925588_500);
and \U$12784 ( \13470 , \11782 , RI9924598_520);
nor \U$12785 ( \13471 , \13469 , \13470 );
nand \U$12786 ( \13472 , \13468 , \13471 );
and \U$12787 ( \13473 , \11796 , RI9926848_460);
not \U$12788 ( \13474 , \11681 );
and \U$12789 ( \13475 , \13474 , RI9925ee8_480);
nor \U$12790 ( \13476 , \13473 , \13475 );
not \U$12791 ( \13477 , \11699 );
and \U$12792 ( \13478 , \13477 , RI9923c38_540);
and \U$12793 ( \13479 , \11775 , RI99232d8_560);
nor \U$12794 ( \13480 , \13478 , \13479 );
nand \U$12795 ( \13481 , \13476 , \13480 );
nor \U$12796 ( \13482 , \13472 , \13481 );
and \U$12797 ( \13483 , \11734 , RI992a628_380);
and \U$12798 ( \13484 , \11726 , RI9928eb8_400);
nor \U$12799 ( \13485 , \13483 , \13484 );
and \U$12800 ( \13486 , \11737 , RI992f308_300);
and \U$12801 ( \13487 , \11730 , RI992d418_320);
nor \U$12802 ( \13488 , \13486 , \13487 );
nand \U$12803 ( \13489 , \13485 , \13488 );
and \U$12804 ( \13490 , \11743 , RI992cab8_340);
not \U$12805 ( \13491 , RI99226a8_580);
not \U$12806 ( \13492 , \11749 );
or \U$12807 ( \13493 , \13491 , \13492 );
nand \U$12808 ( \13494 , \10843 , RI9933c28_260);
nand \U$12809 ( \13495 , \13493 , \13494 );
nor \U$12810 ( \13496 , \13490 , \13495 );
nand \U$12811 ( \13497 , \11759 , RI992af88_360);
nand \U$12812 ( \13498 , \11756 , RI99315b8_280);
nand \U$12813 ( \13499 , \13496 , \13497 , \13498 );
nor \U$12814 ( \13500 , \13489 , \13499 );
nand \U$12815 ( \13501 , \13482 , \13500 );
not \U$12816 ( \13502 , \13501 );
buf \U$12817 ( \13503 , \13502 );
and \U$12818 ( \13504 , \13503 , \11635 );
not \U$12819 ( \13505 , \13503 );
and \U$12820 ( \13506 , \13505 , \11634 );
nor \U$12821 ( \13507 , \13504 , \13506 );
nand \U$12822 ( \13508 , \11636 , \13507 );
nand \U$12823 ( \13509 , \13464 , \13508 );
and \U$12824 ( \13510 , \12104 , \12950 );
not \U$12825 ( \13511 , \12104 );
and \U$12826 ( \13512 , \13511 , \12662 );
or \U$12827 ( \13513 , \13510 , \13512 );
not \U$12828 ( \13514 , \13513 );
not \U$12829 ( \13515 , \13248 );
or \U$12830 ( \13516 , \13514 , \13515 );
nand \U$12831 ( \13517 , \13246 , \12936 );
nand \U$12832 ( \13518 , \13516 , \13517 );
not \U$12833 ( \13519 , \13259 );
buf \U$12834 ( \13520 , \12926 );
not \U$12835 ( \13521 , \13520 );
and \U$12836 ( \13522 , \11763 , \13521 );
not \U$12837 ( \13523 , \11763 );
and \U$12838 ( \13524 , \13523 , \13264 );
or \U$12839 ( \13525 , \13522 , \13524 );
not \U$12840 ( \13526 , \13525 );
or \U$12841 ( \13527 , \13519 , \13526 );
nand \U$12842 ( \13528 , \13266 , \13270 );
nand \U$12843 ( \13529 , \13527 , \13528 );
and \U$12844 ( \13530 , \13518 , \13529 );
not \U$12845 ( \13531 , \12302 );
not \U$12846 ( \13532 , \13224 );
or \U$12847 ( \13533 , \13531 , \13532 );
nand \U$12848 ( \13534 , \12956 , \12306 );
nand \U$12849 ( \13535 , \13533 , \13534 );
not \U$12850 ( \13536 , \13535 );
not \U$12851 ( \13537 , \12681 );
or \U$12852 ( \13538 , \13536 , \13537 );
nand \U$12853 ( \13539 , \13228 , \12667 );
nand \U$12854 ( \13540 , \13538 , \13539 );
xor \U$12855 ( \13541 , \13530 , \13540 );
and \U$12856 ( \13542 , \12463 , \12481 );
not \U$12857 ( \13543 , \12463 );
not \U$12858 ( \13544 , \12637 );
and \U$12859 ( \13545 , \13543 , \13544 );
or \U$12860 ( \13546 , \13542 , \13545 );
not \U$12861 ( \13547 , \13546 );
not \U$12862 ( \13548 , \12644 );
or \U$12863 ( \13549 , \13547 , \13548 );
nand \U$12864 ( \13550 , \13211 , \12364 );
nand \U$12865 ( \13551 , \13549 , \13550 );
and \U$12866 ( \13552 , \13541 , \13551 );
and \U$12867 ( \13553 , \13530 , \13540 );
or \U$12868 ( \13554 , \13552 , \13553 );
and \U$12869 ( \13555 , \13509 , \13554 );
not \U$12870 ( \13556 , \13463 );
nor \U$12871 ( \13557 , \13556 , \13508 );
nor \U$12872 ( \13558 , \13555 , \13557 );
not \U$12873 ( \13559 , \13558 );
xor \U$12874 ( \13560 , \13204 , \13156 );
xnor \U$12875 ( \13561 , \13560 , \13277 );
not \U$12876 ( \13562 , \13561 );
or \U$12877 ( \13563 , \13559 , \13562 );
xor \U$12878 ( \13564 , \13273 , \13238 );
xnor \U$12879 ( \13565 , \13564 , \13221 );
not \U$12880 ( \13566 , \13565 );
not \U$12881 ( \13567 , \13272 );
not \U$12882 ( \13568 , \13567 );
not \U$12883 ( \13569 , \13253 );
or \U$12884 ( \13570 , \13568 , \13569 );
or \U$12885 ( \13571 , \13253 , \13567 );
nand \U$12886 ( \13572 , \13570 , \13571 );
not \U$12887 ( \13573 , \12823 );
not \U$12888 ( \13574 , \12138 );
or \U$12889 ( \13575 , \13573 , \13574 );
nand \U$12890 ( \13576 , \12383 , \12822 );
nand \U$12891 ( \13577 , \13575 , \13576 );
not \U$12892 ( \13578 , \13577 );
not \U$12893 ( \13579 , \12761 );
or \U$12894 ( \13580 , \13578 , \13579 );
nand \U$12895 ( \13581 , \13331 , \12197 );
nand \U$12896 ( \13582 , \13580 , \13581 );
xor \U$12897 ( \13583 , \13572 , \13582 );
not \U$12898 ( \13584 , \13098 );
not \U$12899 ( \13585 , \12012 );
or \U$12900 ( \13586 , \13584 , \13585 );
nand \U$12901 ( \13587 , \12322 , \13102 );
nand \U$12902 ( \13588 , \13586 , \13587 );
not \U$12903 ( \13589 , \13588 );
not \U$12904 ( \13590 , \12521 );
or \U$12905 ( \13591 , \13589 , \13590 );
nand \U$12906 ( \13592 , \12002 , \13342 );
nand \U$12907 ( \13593 , \13591 , \13592 );
and \U$12908 ( \13594 , \13583 , \13593 );
and \U$12909 ( \13595 , \13572 , \13582 );
or \U$12910 ( \13596 , \13594 , \13595 );
not \U$12911 ( \13597 , \13596 );
or \U$12912 ( \13598 , \13566 , \13597 );
or \U$12913 ( \13599 , \13565 , \13596 );
xor \U$12914 ( \13600 , \13326 , \13336 );
xor \U$12915 ( \13601 , \13600 , \13347 );
nand \U$12916 ( \13602 , \13599 , \13601 );
nand \U$12917 ( \13603 , \13598 , \13602 );
nand \U$12918 ( \13604 , \13563 , \13603 );
not \U$12919 ( \13605 , \13561 );
not \U$12920 ( \13606 , \13558 );
nand \U$12921 ( \13607 , \13605 , \13606 );
nand \U$12922 ( \13608 , \13604 , \13607 );
not \U$12923 ( \13609 , \13608 );
not \U$12924 ( \13610 , \13609 );
nand \U$12925 ( \13611 , \13451 , \13610 );
nand \U$12926 ( \13612 , \13447 , \13450 );
nand \U$12927 ( \13613 , \13611 , \13612 );
xor \U$12928 ( \13614 , \13056 , \13359 );
xor \U$12929 ( \13615 , \13614 , \13408 );
nor \U$12930 ( \13616 , \13613 , \13615 );
nor \U$12931 ( \13617 , \13445 , \13616 );
xor \U$12932 ( \13618 , \12632 , \12484 );
xor \U$12933 ( \13619 , \13618 , \12707 );
and \U$12934 ( \13620 , \12859 , \12790 );
not \U$12935 ( \13621 , \12859 );
and \U$12936 ( \13622 , \13621 , \12791 );
nor \U$12937 ( \13623 , \13620 , \13622 );
not \U$12938 ( \13624 , \13623 );
not \U$12939 ( \13625 , \12788 );
and \U$12940 ( \13626 , \13624 , \13625 );
and \U$12941 ( \13627 , \13623 , \12788 );
nor \U$12942 ( \13628 , \13626 , \13627 );
xor \U$12943 ( \13629 , \13619 , \13628 );
buf \U$12944 ( \13630 , \13429 );
or \U$12945 ( \13631 , \13421 , \13423 );
and \U$12946 ( \13632 , \13630 , \13631 );
and \U$12947 ( \13633 , \13421 , \13423 );
nor \U$12948 ( \13634 , \13632 , \13633 );
xor \U$12949 ( \13635 , \13629 , \13634 );
not \U$12950 ( \13636 , \13415 );
not \U$12951 ( \13637 , \13433 );
nand \U$12952 ( \13638 , \13636 , \13637 );
and \U$12953 ( \13639 , \13638 , \13442 );
and \U$12954 ( \13640 , \13433 , \13415 );
nor \U$12955 ( \13641 , \13639 , \13640 );
nand \U$12956 ( \13642 , \13635 , \13641 );
xor \U$12957 ( \13643 , \12710 , \12712 );
xor \U$12958 ( \13644 , \13643 , \12863 );
xor \U$12959 ( \13645 , \13619 , \13628 );
and \U$12960 ( \13646 , \13645 , \13634 );
and \U$12961 ( \13647 , \13619 , \13628 );
or \U$12962 ( \13648 , \13646 , \13647 );
nand \U$12963 ( \13649 , \13644 , \13648 );
and \U$12964 ( \13650 , \13642 , \13649 );
nand \U$12965 ( \13651 , \13617 , \13650 );
not \U$12966 ( \13652 , \13651 );
not \U$12967 ( \13653 , \13652 );
nor \U$12968 ( \13654 , \12913 , \13653 );
not \U$12969 ( \13655 , \13654 );
not \U$12970 ( \13656 , \12980 );
and \U$12971 ( \13657 , \12462 , \13037 );
not \U$12972 ( \13658 , \12462 );
and \U$12973 ( \13659 , \13658 , \12662 );
or \U$12974 ( \13660 , \13657 , \13659 );
not \U$12975 ( \13661 , \13660 );
or \U$12976 ( \13662 , \13656 , \13661 );
and \U$12977 ( \13663 , \12246 , \13241 );
not \U$12978 ( \13664 , \12246 );
and \U$12979 ( \13665 , \13664 , \12662 );
or \U$12980 ( \13666 , \13663 , \13665 );
nand \U$12981 ( \13667 , \13666 , \13045 );
nand \U$12982 ( \13668 , \13662 , \13667 );
not \U$12983 ( \13669 , \13270 );
and \U$12984 ( \13670 , \13520 , \12106 );
not \U$12985 ( \13671 , \13520 );
and \U$12986 ( \13672 , \13671 , \12105 );
nor \U$12987 ( \13673 , \13670 , \13672 );
not \U$12988 ( \13674 , \13673 );
or \U$12989 ( \13675 , \13669 , \13674 );
and \U$12990 ( \13676 , \13521 , \12301 );
not \U$12991 ( \13677 , \13521 );
not \U$12992 ( \13678 , \12301 );
and \U$12993 ( \13679 , \13677 , \13678 );
nor \U$12994 ( \13680 , \13676 , \13679 );
not \U$12995 ( \13681 , \13680 );
nand \U$12996 ( \13682 , \13681 , \13259 );
nand \U$12997 ( \13683 , \13675 , \13682 );
nand \U$12998 ( \13684 , \13668 , \13683 );
not \U$12999 ( \13685 , \12627 );
not \U$13000 ( \13686 , \12686 );
or \U$13001 ( \13687 , \13685 , \13686 );
nand \U$13002 ( \13688 , \12956 , \12626 );
nand \U$13003 ( \13689 , \13687 , \13688 );
not \U$13004 ( \13690 , \13689 );
not \U$13005 ( \13691 , \12681 );
or \U$13006 ( \13692 , \13690 , \13691 );
and \U$13007 ( \13693 , \12463 , \12686 );
not \U$13008 ( \13694 , \12463 );
and \U$13009 ( \13695 , \13694 , \12956 );
or \U$13010 ( \13696 , \13693 , \13695 );
nand \U$13011 ( \13697 , \13696 , \12667 );
nand \U$13012 ( \13698 , \13692 , \13697 );
xor \U$13013 ( \13699 , \13684 , \13698 );
not \U$13014 ( \13700 , \13149 );
not \U$13015 ( \13701 , \12481 );
or \U$13016 ( \13702 , \13700 , \13701 );
nand \U$13017 ( \13703 , \12746 , \13148 );
nand \U$13018 ( \13704 , \13702 , \13703 );
not \U$13019 ( \13705 , \13704 );
not \U$13020 ( \13706 , \12375 );
or \U$13021 ( \13707 , \13705 , \13706 );
not \U$13022 ( \13708 , \12823 );
not \U$13023 ( \13709 , \12637 );
or \U$13024 ( \13710 , \13708 , \13709 );
nand \U$13025 ( \13711 , \13544 , \12822 );
nand \U$13026 ( \13712 , \13710 , \13711 );
nand \U$13027 ( \13713 , \13712 , \12364 );
nand \U$13028 ( \13714 , \13707 , \13713 );
xor \U$13029 ( \13715 , \13699 , \13714 );
and \U$13030 ( \13716 , \11796 , RI9926758_462);
and \U$13031 ( \13717 , \11917 , RI9925df8_482);
nor \U$13032 ( \13718 , \13716 , \13717 );
and \U$13033 ( \13719 , \11926 , RI9923b48_542);
and \U$13034 ( \13720 , \11775 , RI99231e8_562);
nor \U$13035 ( \13721 , \13719 , \13720 );
nand \U$13036 ( \13722 , \13718 , \13721 );
and \U$13037 ( \13723 , \11910 , RI9928468_422);
and \U$13038 ( \13724 , \11913 , RI9927b08_442);
nor \U$13039 ( \13725 , \13723 , \13724 );
and \U$13040 ( \13726 , \11786 , RI9924e08_502);
and \U$13041 ( \13727 , \11923 , RI99244a8_522);
nor \U$13042 ( \13728 , \13726 , \13727 );
nand \U$13043 ( \13729 , \13725 , \13728 );
nor \U$13044 ( \13730 , \13722 , \13729 );
and \U$13045 ( \13731 , \11734 , RI992a538_382);
and \U$13046 ( \13732 , \11726 , RI9928dc8_402);
nor \U$13047 ( \13733 , \13731 , \13732 );
and \U$13048 ( \13734 , \11737 , RI992f218_302);
and \U$13049 ( \13735 , \11730 , RI992d328_322);
nor \U$13050 ( \13736 , \13734 , \13735 );
nand \U$13051 ( \13737 , \13733 , \13736 );
and \U$13052 ( \13738 , \11743 , RI992c9c8_342);
not \U$13053 ( \13739 , RI99225b8_582);
not \U$13054 ( \13740 , \11749 );
or \U$13055 ( \13741 , \13739 , \13740 );
nand \U$13056 ( \13742 , \10843 , RI9933b38_262);
nand \U$13057 ( \13743 , \13741 , \13742 );
nor \U$13058 ( \13744 , \13738 , \13743 );
nand \U$13059 ( \13745 , \11759 , RI992ae98_362);
nand \U$13060 ( \13746 , \11756 , RI99314c8_282);
nand \U$13061 ( \13747 , \13744 , \13745 , \13746 );
nor \U$13062 ( \13748 , \13737 , \13747 );
nand \U$13063 ( \13749 , \13730 , \13748 );
not \U$13064 ( \13750 , \13749 );
not \U$13065 ( \13751 , \13750 );
and \U$13066 ( \13752 , \13751 , \12323 );
not \U$13067 ( \13753 , \13751 );
and \U$13068 ( \13754 , \13753 , \12020 );
nor \U$13069 ( \13755 , \13752 , \13754 );
not \U$13070 ( \13756 , \13755 );
not \U$13071 ( \13757 , \13756 );
not \U$13072 ( \13758 , \12016 );
or \U$13073 ( \13759 , \13757 , \13758 );
and \U$13074 ( \13760 , \11805 , RI99284e0_421);
and \U$13075 ( \13761 , \13466 , RI9927b80_441);
nor \U$13076 ( \13762 , \13760 , \13761 );
not \U$13077 ( \13763 , \11795 );
not \U$13078 ( \13764 , \13763 );
and \U$13079 ( \13765 , \13764 , RI99267d0_461);
and \U$13080 ( \13766 , \13474 , RI9925e70_481);
nor \U$13081 ( \13767 , \13765 , \13766 );
nand \U$13082 ( \13768 , \13762 , \13767 );
and \U$13083 ( \13769 , \11786 , RI9925510_501);
and \U$13084 ( \13770 , \11923 , RI9924520_521);
nor \U$13085 ( \13771 , \13769 , \13770 );
and \U$13086 ( \13772 , \13477 , RI9923bc0_541);
and \U$13087 ( \13773 , \11775 , RI9923260_561);
nor \U$13088 ( \13774 , \13772 , \13773 );
nand \U$13089 ( \13775 , \13771 , \13774 );
nor \U$13090 ( \13776 , \13768 , \13775 );
nand \U$13091 ( \13777 , \11726 , RI9928e40_401);
nand \U$13092 ( \13778 , \11734 , RI992a5b0_381);
nand \U$13093 ( \13779 , \11730 , RI992d3a0_321);
nand \U$13094 ( \13780 , \11737 , RI992f290_301);
nand \U$13095 ( \13781 , \13777 , \13778 , \13779 , \13780 );
nand \U$13096 ( \13782 , \11743 , RI992ca40_341);
nand \U$13097 ( \13783 , \11825 , RI992af10_361);
nand \U$13098 ( \13784 , \11756 , RI9931540_281);
and \U$13099 ( \13785 , \11749 , RI9922630_581);
nand \U$13100 ( \13786 , \10843 , RI9933bb0_261);
not \U$13101 ( \13787 , \13786 );
nor \U$13102 ( \13788 , \13785 , \13787 );
nand \U$13103 ( \13789 , \13782 , \13783 , \13784 , \13788 );
nor \U$13104 ( \13790 , \13781 , \13789 );
nand \U$13105 ( \13791 , \13776 , \13790 );
buf \U$13106 ( \13792 , \13791 );
not \U$13107 ( \13793 , \13792 );
and \U$13108 ( \13794 , \12032 , \13793 );
not \U$13109 ( \13795 , \12032 );
and \U$13110 ( \13796 , \13795 , \13792 );
or \U$13111 ( \13797 , \13794 , \13796 );
nand \U$13112 ( \13798 , \12002 , \13797 );
nand \U$13113 ( \13799 , \13759 , \13798 );
not \U$13114 ( \13800 , \13799 );
not \U$13115 ( \13801 , \13503 );
not \U$13116 ( \13802 , \13801 );
not \U$13117 ( \13803 , \12198 );
or \U$13118 ( \13804 , \13802 , \13803 );
nand \U$13119 ( \13805 , \12383 , \13503 );
nand \U$13120 ( \13806 , \13804 , \13805 );
not \U$13121 ( \13807 , \13806 );
not \U$13122 ( \13808 , \12194 );
or \U$13123 ( \13809 , \13807 , \13808 );
not \U$13124 ( \13810 , \13199 );
not \U$13125 ( \13811 , \12138 );
or \U$13126 ( \13812 , \13810 , \13811 );
nand \U$13127 ( \13813 , \12137 , \13457 );
nand \U$13128 ( \13814 , \13812 , \13813 );
nand \U$13129 ( \13815 , \13814 , \12837 );
nand \U$13130 ( \13816 , \13809 , \13815 );
not \U$13131 ( \13817 , \13816 );
nand \U$13132 ( \13818 , \13800 , \13817 );
xor \U$13133 ( \13819 , \13668 , \13683 );
and \U$13134 ( \13820 , \13818 , \13819 );
and \U$13135 ( \13821 , \13799 , \13816 );
nor \U$13136 ( \13822 , \13820 , \13821 );
not \U$13137 ( \13823 , \13822 );
xor \U$13138 ( \13824 , \13715 , \13823 );
not \U$13139 ( \13825 , \13259 );
not \U$13140 ( \13826 , \13673 );
or \U$13141 ( \13827 , \13825 , \13826 );
not \U$13142 ( \13828 , \13520 );
not \U$13143 ( \13829 , \11947 );
or \U$13144 ( \13830 , \13828 , \13829 );
nand \U$13145 ( \13831 , \11946 , \13261 );
nand \U$13146 ( \13832 , \13830 , \13831 );
nand \U$13147 ( \13833 , \13832 , \13270 );
nand \U$13148 ( \13834 , \13827 , \13833 );
not \U$13149 ( \13835 , \13666 );
not \U$13150 ( \13836 , \12980 );
or \U$13151 ( \13837 , \13835 , \13836 );
not \U$13152 ( \13838 , \13037 );
not \U$13153 ( \13839 , \12301 );
or \U$13154 ( \13840 , \13838 , \13839 );
nand \U$13155 ( \13841 , \13244 , \13678 );
nand \U$13156 ( \13842 , \13840 , \13841 );
nand \U$13157 ( \13843 , \13842 , \12936 );
nand \U$13158 ( \13844 , \13837 , \13843 );
xor \U$13159 ( \13845 , \13834 , \13844 );
not \U$13160 ( \13846 , \13814 );
not \U$13161 ( \13847 , \12194 );
or \U$13162 ( \13848 , \13846 , \13847 );
not \U$13163 ( \13849 , \13098 );
not \U$13164 ( \13850 , \12154 );
or \U$13165 ( \13851 , \13849 , \13850 );
nand \U$13166 ( \13852 , \12199 , \13102 );
nand \U$13167 ( \13853 , \13851 , \13852 );
nand \U$13168 ( \13854 , \13853 , \12837 );
nand \U$13169 ( \13855 , \13848 , \13854 );
xor \U$13170 ( \13856 , \13845 , \13855 );
not \U$13171 ( \13857 , \13797 );
not \U$13172 ( \13858 , \12016 );
or \U$13173 ( \13859 , \13857 , \13858 );
not \U$13174 ( \13860 , \13801 );
not \U$13175 ( \13861 , \12323 );
or \U$13176 ( \13862 , \13860 , \13861 );
nand \U$13177 ( \13863 , \12029 , \13503 );
nand \U$13178 ( \13864 , \13862 , \13863 );
nand \U$13179 ( \13865 , \12002 , \13864 );
nand \U$13180 ( \13866 , \13859 , \13865 );
xor \U$13181 ( \13867 , \13856 , \13866 );
xnor \U$13182 ( \13868 , \13824 , \13867 );
nor \U$13183 ( \13869 , \11681 , \3487 );
nor \U$13184 ( \13870 , \11674 , \3485 );
nor \U$13185 ( \13871 , \13869 , \13870 );
nor \U$13186 ( \13872 , \12427 , \8237 );
nor \U$13187 ( \13873 , \11692 , \8240 );
nor \U$13188 ( \13874 , \13872 , \13873 );
nand \U$13189 ( \13875 , \13871 , \13874 );
nor \U$13190 ( \13876 , \11705 , \3465 );
nor \U$13191 ( \13877 , \11699 , \3490 );
nor \U$13192 ( \13878 , \13876 , \13877 );
not \U$13193 ( \13879 , \12420 );
not \U$13194 ( \13880 , \8262 );
and \U$13195 ( \13881 , \13879 , \13880 );
nor \U$13196 ( \13882 , \11715 , \8265 );
nor \U$13197 ( \13883 , \13881 , \13882 );
nand \U$13198 ( \13884 , \13878 , \13883 );
nor \U$13199 ( \13885 , \13875 , \13884 );
nand \U$13200 ( \13886 , \11737 , RI992f0b0_305);
nand \U$13201 ( \13887 , \11816 , RI992d1c0_325);
nand \U$13202 ( \13888 , \11734 , RI992a3d0_385);
nand \U$13203 ( \13889 , RI9928c60_405, \11726 );
nand \U$13204 ( \13890 , \13886 , \13887 , \13888 , \13889 );
and \U$13205 ( \13891 , \11743 , RI992c860_345);
nand \U$13206 ( \13892 , \11749 , RI9922450_585);
nand \U$13207 ( \13893 , \10843 , RI99339d0_265);
nand \U$13208 ( \13894 , \13892 , \13893 );
nor \U$13209 ( \13895 , \13891 , \13894 );
nand \U$13210 ( \13896 , \11756 , RI9931360_285);
nand \U$13211 ( \13897 , \11759 , RI992ad30_365);
nand \U$13212 ( \13898 , \13895 , \13896 , \13897 );
nor \U$13213 ( \13899 , \13890 , \13898 );
nand \U$13214 ( \13900 , \13885 , \13899 );
buf \U$13215 ( \13901 , \13900 );
not \U$13216 ( \13902 , \13901 );
and \U$13217 ( \13903 , \11639 , \13902 );
and \U$13218 ( \13904 , \12827 , \13901 );
nor \U$13219 ( \13905 , \13903 , \13904 );
nand \U$13220 ( \13906 , \11637 , \13905 );
not \U$13221 ( \13907 , \13906 );
not \U$13222 ( \13908 , \11884 );
and \U$13223 ( \13909 , \11910 , RI9928378_424);
and \U$13224 ( \13910 , \11913 , RI9926fc8_444);
nor \U$13225 ( \13911 , \13909 , \13910 );
and \U$13226 ( \13912 , \11796 , RI9926668_464);
and \U$13227 ( \13913 , \11917 , RI9925d08_484);
nor \U$13228 ( \13914 , \13912 , \13913 );
nand \U$13229 ( \13915 , \13911 , \13914 );
and \U$13230 ( \13916 , \11786 , RI9924d18_504);
and \U$13231 ( \13917 , \11923 , RI99243b8_524);
nor \U$13232 ( \13918 , \13916 , \13917 );
and \U$13233 ( \13919 , \11926 , RI9923a58_544);
and \U$13234 ( \13920 , \11775 , RI99230f8_564);
nor \U$13235 ( \13921 , \13919 , \13920 );
nand \U$13236 ( \13922 , \13918 , \13921 );
nor \U$13237 ( \13923 , \13915 , \13922 );
nand \U$13238 ( \13924 , \11737 , RI992f128_304);
nand \U$13239 ( \13925 , \11816 , RI992d238_324);
nand \U$13240 ( \13926 , \11726 , RI9928cd8_404);
nand \U$13241 ( \13927 , \11734 , RI992a448_384);
nand \U$13242 ( \13928 , \13924 , \13925 , \13926 , \13927 );
and \U$13243 ( \13929 , \11743 , RI992c8d8_344);
not \U$13244 ( \13930 , RI99224c8_584);
not \U$13245 ( \13931 , \11749 );
or \U$13246 ( \13932 , \13930 , \13931 );
nand \U$13247 ( \13933 , \10843 , RI9933a48_264);
nand \U$13248 ( \13934 , \13932 , \13933 );
nor \U$13249 ( \13935 , \13929 , \13934 );
nand \U$13250 ( \13936 , \11759 , RI992ada8_364);
nand \U$13251 ( \13937 , \11756 , RI99313d8_284);
nand \U$13252 ( \13938 , \13935 , \13936 , \13937 );
nor \U$13253 ( \13939 , \13928 , \13938 );
nand \U$13254 ( \13940 , \13923 , \13939 );
not \U$13255 ( \13941 , \13940 );
not \U$13256 ( \13942 , \13941 );
not \U$13257 ( \13943 , \13942 );
not \U$13258 ( \13944 , \12118 );
or \U$13259 ( \13945 , \13943 , \13944 );
nand \U$13260 ( \13946 , \12534 , \13941 );
nand \U$13261 ( \13947 , \13945 , \13946 );
not \U$13262 ( \13948 , \13947 );
or \U$13263 ( \13949 , \13908 , \13948 );
nor \U$13264 ( \13950 , \11912 , \8359 );
not \U$13265 ( \13951 , \13950 );
not \U$13266 ( \13952 , \8362 );
nand \U$13267 ( \13953 , \13952 , \11805 );
not \U$13268 ( \13954 , \11705 );
not \U$13269 ( \13955 , \2616 );
and \U$13270 ( \13956 , \13954 , \13955 );
nor \U$13271 ( \13957 , \11699 , \8339 );
nor \U$13272 ( \13958 , \13956 , \13957 );
nand \U$13273 ( \13959 , \13951 , \13953 , \13958 );
not \U$13274 ( \13960 , \11715 );
not \U$13275 ( \13961 , \8327 );
and \U$13276 ( \13962 , \13960 , \13961 );
nor \U$13277 ( \13963 , \12420 , \8324 );
nor \U$13278 ( \13964 , \13962 , \13963 );
not \U$13279 ( \13965 , \11681 );
not \U$13280 ( \13966 , \8368 );
and \U$13281 ( \13967 , \13965 , \13966 );
nor \U$13282 ( \13968 , \11674 , \8352 );
nor \U$13283 ( \13969 , \13967 , \13968 );
nand \U$13284 ( \13970 , \13964 , \13969 );
nor \U$13285 ( \13971 , \13959 , \13970 );
and \U$13286 ( \13972 , \11743 , RI992c950_343);
not \U$13287 ( \13973 , RI9922540_583);
not \U$13288 ( \13974 , \11749 );
or \U$13289 ( \13975 , \13973 , \13974 );
nand \U$13290 ( \13976 , \10843 , RI9933ac0_263);
nand \U$13291 ( \13977 , \13975 , \13976 );
nor \U$13292 ( \13978 , \13972 , \13977 );
nand \U$13293 ( \13979 , \11756 , RI9931450_283);
nand \U$13294 ( \13980 , \11826 , RI992ae20_363);
nand \U$13295 ( \13981 , \13978 , \13979 , \13980 );
nand \U$13296 ( \13982 , \11737 , RI992f1a0_303);
nand \U$13297 ( \13983 , \11816 , RI992d2b0_323);
nand \U$13298 ( \13984 , \11734 , RI992a4c0_383);
nand \U$13299 ( \13985 , \11726 , RI9928d50_403);
nand \U$13300 ( \13986 , \13982 , \13983 , \13984 , \13985 );
nor \U$13301 ( \13987 , \13981 , \13986 );
nand \U$13302 ( \13988 , \13971 , \13987 );
buf \U$13303 ( \13989 , \13988 );
not \U$13304 ( \13990 , \13989 );
not \U$13305 ( \13991 , \12533 );
or \U$13306 ( \13992 , \13990 , \13991 );
not \U$13307 ( \13993 , \13989 );
nand \U$13308 ( \13994 , \11890 , \13993 );
nand \U$13309 ( \13995 , \13992 , \13994 );
nand \U$13310 ( \13996 , \13995 , \12540 );
nand \U$13311 ( \13997 , \13949 , \13996 );
not \U$13312 ( \13998 , \13997 );
not \U$13313 ( \13999 , \13998 );
or \U$13314 ( \14000 , \13907 , \13999 );
buf \U$13315 ( \14001 , \13147 );
not \U$13316 ( \14002 , \14001 );
not \U$13317 ( \14003 , \13224 );
or \U$13318 ( \14004 , \14002 , \14003 );
not \U$13319 ( \14005 , \14001 );
nand \U$13320 ( \14006 , \14005 , \12956 );
nand \U$13321 ( \14007 , \14004 , \14006 );
not \U$13322 ( \14008 , \14007 );
not \U$13323 ( \14009 , \12681 );
or \U$13324 ( \14010 , \14008 , \14009 );
not \U$13325 ( \14011 , \12823 );
not \U$13326 ( \14012 , \12686 );
or \U$13327 ( \14013 , \14011 , \14012 );
nand \U$13328 ( \14014 , \12956 , \12822 );
nand \U$13329 ( \14015 , \14013 , \14014 );
nand \U$13330 ( \14016 , \14015 , \12667 );
nand \U$13331 ( \14017 , \14010 , \14016 );
xor \U$13333 ( \14018 , \14017 , 1'b0 );
not \U$13334 ( \14019 , \13199 );
not \U$13335 ( \14020 , \12481 );
or \U$13336 ( \14021 , \14019 , \14020 );
nand \U$13337 ( \14022 , \12746 , \13457 );
nand \U$13338 ( \14023 , \14021 , \14022 );
not \U$13339 ( \14024 , \14023 );
not \U$13340 ( \14025 , \12375 );
or \U$13341 ( \14026 , \14024 , \14025 );
and \U$13342 ( \14027 , \13102 , \13544 );
not \U$13343 ( \14028 , \13102 );
and \U$13344 ( \14029 , \14028 , \12637 );
or \U$13345 ( \14030 , \14027 , \14029 );
nand \U$13346 ( \14031 , \14030 , \12365 );
nand \U$13347 ( \14032 , \14026 , \14031 );
and \U$13348 ( \14033 , \14018 , \14032 );
or \U$13350 ( \14034 , \14033 , 1'b0 );
nand \U$13351 ( \14035 , \14000 , \14034 );
not \U$13352 ( \14036 , \13906 );
nand \U$13353 ( \14037 , \14036 , \13997 );
nand \U$13354 ( \14038 , \14035 , \14037 );
and \U$13355 ( \14039 , \13941 , \11639 );
not \U$13356 ( \14040 , \13941 );
and \U$13357 ( \14041 , \14040 , \12467 );
nor \U$13358 ( \14042 , \14039 , \14041 );
and \U$13359 ( \14043 , \11637 , \14042 );
not \U$13360 ( \14044 , \13751 );
not \U$13361 ( \14045 , \12533 );
or \U$13362 ( \14046 , \14044 , \14045 );
nand \U$13363 ( \14047 , \11890 , \13750 );
nand \U$13364 ( \14048 , \14046 , \14047 );
not \U$13365 ( \14049 , \14048 );
not \U$13366 ( \14050 , \11873 );
or \U$13367 ( \14051 , \14049 , \14050 );
buf \U$13368 ( \14052 , \11881 );
nand \U$13369 ( \14053 , \13995 , \14052 , \11882 );
nand \U$13370 ( \14054 , \14051 , \14053 );
xor \U$13371 ( \14055 , \14043 , \14054 );
not \U$13372 ( \14056 , \14015 );
not \U$13373 ( \14057 , \12681 );
or \U$13374 ( \14058 , \14056 , \14057 );
nand \U$13375 ( \14059 , \13689 , \12667 );
nand \U$13376 ( \14060 , \14058 , \14059 );
and \U$13377 ( \14061 , \12625 , \13037 );
not \U$13378 ( \14062 , \12625 );
and \U$13379 ( \14063 , \14062 , \13244 );
or \U$13380 ( \14064 , \14061 , \14063 );
not \U$13381 ( \14065 , \14064 );
not \U$13382 ( \14066 , \13248 );
or \U$13383 ( \14067 , \14065 , \14066 );
nand \U$13384 ( \14068 , \13251 , \13660 );
nand \U$13385 ( \14069 , \14067 , \14068 );
not \U$13386 ( \14070 , \14069 );
and \U$13387 ( \14071 , \12246 , \13050 );
not \U$13388 ( \14072 , \12246 );
and \U$13389 ( \14073 , \14072 , \13264 );
or \U$13390 ( \14074 , \14071 , \14073 );
and \U$13391 ( \14075 , \14074 , \13259 );
not \U$13392 ( \14076 , \13270 );
nor \U$13393 ( \14077 , \14076 , \13680 );
nor \U$13394 ( \14078 , \14075 , \14077 );
nor \U$13395 ( \14079 , \14070 , \14078 );
xor \U$13396 ( \14080 , \14060 , \14079 );
not \U$13397 ( \14081 , \14030 );
not \U$13398 ( \14082 , \12644 );
or \U$13399 ( \14083 , \14081 , \14082 );
not \U$13400 ( \14084 , \12363 );
nand \U$13401 ( \14085 , \14084 , \13704 );
nand \U$13402 ( \14086 , \14083 , \14085 );
and \U$13403 ( \14087 , \14080 , \14086 );
and \U$13404 ( \14088 , \14060 , \14079 );
or \U$13405 ( \14089 , \14087 , \14088 );
xor \U$13406 ( \14090 , \14055 , \14089 );
xor \U$13407 ( \14091 , \14038 , \14090 );
xor \U$13408 ( \14092 , \14060 , \14079 );
xor \U$13409 ( \14093 , \14092 , \14086 );
xnor \U$13410 ( \14094 , \14078 , \14069 );
not \U$13411 ( \14095 , \13793 );
not \U$13412 ( \14096 , \12383 );
or \U$13413 ( \14097 , \14095 , \14096 );
not \U$13414 ( \14098 , \12137 );
nand \U$13415 ( \14099 , \14098 , \13792 );
nand \U$13416 ( \14100 , \14097 , \14099 );
not \U$13417 ( \14101 , \14100 );
not \U$13418 ( \14102 , \12761 );
or \U$13419 ( \14103 , \14101 , \14102 );
nand \U$13420 ( \14104 , \13806 , \12197 );
nand \U$13421 ( \14105 , \14103 , \14104 );
xor \U$13422 ( \14106 , \14094 , \14105 );
and \U$13423 ( \14107 , \13993 , \12322 );
not \U$13424 ( \14108 , \13993 );
and \U$13425 ( \14109 , \14108 , \12327 );
nor \U$13426 ( \14110 , \14107 , \14109 );
or \U$13427 ( \14111 , \12520 , \14110 );
or \U$13428 ( \14112 , \12524 , \13755 );
nand \U$13429 ( \14113 , \14111 , \14112 );
and \U$13430 ( \14114 , \14106 , \14113 );
and \U$13431 ( \14115 , \14094 , \14105 );
or \U$13432 ( \14116 , \14114 , \14115 );
xor \U$13433 ( \14117 , \14093 , \14116 );
not \U$13434 ( \14118 , \11873 );
not \U$13435 ( \14119 , \13947 );
or \U$13436 ( \14120 , \14118 , \14119 );
not \U$13437 ( \14121 , \13901 );
not \U$13438 ( \14122 , \12533 );
or \U$13439 ( \14123 , \14121 , \14122 );
nand \U$13440 ( \14124 , \11890 , \13902 );
nand \U$13441 ( \14125 , \14123 , \14124 );
nand \U$13442 ( \14126 , \14125 , \14052 , \11882 );
nand \U$13443 ( \14127 , \14120 , \14126 );
not \U$13444 ( \14128 , RI99242c8_526);
nor \U$13445 ( \14129 , \14128 , \11710 );
not \U$13446 ( \14130 , RI9924c28_506);
nor \U$13447 ( \14131 , \11715 , \14130 );
nor \U$13448 ( \14132 , \14129 , \14131 );
not \U$13449 ( \14133 , \12211 );
not \U$13450 ( \14134 , \8542 );
and \U$13451 ( \14135 , \14133 , \14134 );
nor \U$13452 ( \14136 , \12427 , \8539 );
nor \U$13453 ( \14137 , \14135 , \14136 );
nand \U$13454 ( \14138 , \14132 , \14137 );
not \U$13455 ( \14139 , \11705 );
not \U$13456 ( \14140 , \3683 );
and \U$13457 ( \14141 , \14139 , \14140 );
nor \U$13458 ( \14142 , \11699 , \8535 );
nor \U$13459 ( \14143 , \14141 , \14142 );
not \U$13460 ( \14144 , \11674 );
not \U$13461 ( \14145 , \8523 );
and \U$13462 ( \14146 , \14144 , \14145 );
nor \U$13463 ( \14147 , \11681 , \8520 );
nor \U$13464 ( \14148 , \14146 , \14147 );
nand \U$13465 ( \14149 , \14143 , \14148 );
nor \U$13466 ( \14150 , \14138 , \14149 );
nand \U$13467 ( \14151 , \11737 , RI992f038_306);
nand \U$13468 ( \14152 , \11816 , RI992d148_326);
nand \U$13469 ( \14153 , \11734 , RI992a358_386);
nand \U$13470 ( \14154 , \11726 , RI9928be8_406);
nand \U$13471 ( \14155 , \14151 , \14152 , \14153 , \14154 );
and \U$13472 ( \14156 , \11743 , RI992c7e8_346);
not \U$13473 ( \14157 , RI99223d8_586);
not \U$13474 ( \14158 , \11749 );
or \U$13475 ( \14159 , \14157 , \14158 );
nand \U$13476 ( \14160 , \10843 , RI9933958_266);
nand \U$13477 ( \14161 , \14159 , \14160 );
nor \U$13478 ( \14162 , \14156 , \14161 );
nand \U$13479 ( \14163 , \11756 , RI99312e8_286);
nand \U$13480 ( \14164 , \11759 , RI992acb8_366);
nand \U$13481 ( \14165 , \14162 , \14163 , \14164 );
nor \U$13482 ( \14166 , \14155 , \14165 );
nand \U$13483 ( \14167 , \14150 , \14166 );
buf \U$13484 ( \14168 , \14167 );
and \U$13485 ( \14169 , \14168 , \12827 );
not \U$13486 ( \14170 , \14168 );
and \U$13487 ( \14171 , \14170 , \11635 );
nor \U$13488 ( \14172 , \14169 , \14171 );
and \U$13489 ( \14173 , \11637 , \14172 );
or \U$13490 ( \14174 , \14127 , \14173 );
and \U$13491 ( \14175 , \12821 , \13241 );
not \U$13492 ( \14176 , \12821 );
and \U$13493 ( \14177 , \14176 , \13244 );
or \U$13494 ( \14178 , \14175 , \14177 );
not \U$13495 ( \14179 , \14178 );
not \U$13496 ( \14180 , \12980 );
or \U$13497 ( \14181 , \14179 , \14180 );
not \U$13498 ( \14182 , \12937 );
nand \U$13499 ( \14183 , \14064 , \14182 );
nand \U$13500 ( \14184 , \14181 , \14183 );
not \U$13501 ( \14185 , \14184 );
not \U$13502 ( \14186 , \13259 );
xor \U$13503 ( \14187 , \13264 , \12462 );
not \U$13504 ( \14188 , \14187 );
or \U$13505 ( \14189 , \14186 , \14188 );
nand \U$13506 ( \14190 , \14074 , \13270 );
nand \U$13507 ( \14191 , \14189 , \14190 );
not \U$13508 ( \14192 , \14191 );
or \U$13509 ( \14193 , \14185 , \14192 );
not \U$13510 ( \14194 , \14191 );
not \U$13511 ( \14195 , \14194 );
not \U$13512 ( \14196 , \14184 );
not \U$13513 ( \14197 , \14196 );
or \U$13514 ( \14198 , \14195 , \14197 );
not \U$13515 ( \14199 , \13098 );
not \U$13516 ( \14200 , \12686 );
or \U$13517 ( \14201 , \14199 , \14200 );
nand \U$13518 ( \14202 , \12956 , \13102 );
nand \U$13519 ( \14203 , \14201 , \14202 );
not \U$13520 ( \14204 , \14203 );
not \U$13521 ( \14205 , \12681 );
or \U$13522 ( \14206 , \14204 , \14205 );
nand \U$13523 ( \14207 , \14007 , \12667 );
nand \U$13524 ( \14208 , \14206 , \14207 );
nand \U$13525 ( \14209 , \14198 , \14208 );
nand \U$13526 ( \14210 , \14193 , \14209 );
nand \U$13527 ( \14211 , \14174 , \14210 );
nand \U$13528 ( \14212 , \14127 , \14173 );
nand \U$13529 ( \14213 , \14211 , \14212 );
and \U$13530 ( \14214 , \14117 , \14213 );
and \U$13531 ( \14215 , \14093 , \14116 );
or \U$13532 ( \14216 , \14214 , \14215 );
xor \U$13533 ( \14217 , \14091 , \14216 );
xor \U$13534 ( \14218 , \13868 , \14217 );
xor \U$13535 ( \14219 , \13819 , \13799 );
xnor \U$13536 ( \14220 , \14219 , \13817 );
xor \U$13537 ( \14221 , \13906 , \14034 );
xor \U$13538 ( \14222 , \14221 , \13998 );
xor \U$13539 ( \14223 , \14220 , \14222 );
xor \U$13540 ( \14224 , \14093 , \14116 );
xor \U$13541 ( \14225 , \14224 , \14213 );
and \U$13542 ( \14226 , \14223 , \14225 );
and \U$13543 ( \14227 , \14220 , \14222 );
or \U$13544 ( \14228 , \14226 , \14227 );
and \U$13545 ( \14229 , \14218 , \14228 );
not \U$13546 ( \14230 , \14218 );
not \U$13547 ( \14231 , \14228 );
and \U$13548 ( \14232 , \14230 , \14231 );
nor \U$13549 ( \14233 , \14229 , \14232 );
not \U$13550 ( \14234 , \14233 );
xor \U$13551 ( \14235 , \14017 , 1'b0 );
xor \U$13552 ( \14236 , \14235 , \14032 );
not \U$13553 ( \14237 , \11705 );
not \U$13554 ( \14238 , \8659 );
and \U$13555 ( \14239 , \14237 , \14238 );
nor \U$13556 ( \14240 , \11699 , \8682 );
nor \U$13557 ( \14241 , \14239 , \14240 );
nor \U$13558 ( \14242 , \11800 , \8651 );
nor \U$13559 ( \14243 , \12211 , \8655 );
nor \U$13560 ( \14244 , \14242 , \14243 );
not \U$13561 ( \14245 , \12420 );
not \U$13562 ( \14246 , \8666 );
and \U$13563 ( \14247 , \14245 , \14246 );
nor \U$13564 ( \14248 , \11715 , \8668 );
nor \U$13565 ( \14249 , \14247 , \14248 );
and \U$13566 ( \14250 , \13764 , RI9926500_467);
and \U$13567 ( \14251 , \11791 , RI9925ba0_487);
nor \U$13568 ( \14252 , \14250 , \14251 );
nand \U$13569 ( \14253 , \14241 , \14244 , \14249 , \14252 );
and \U$13570 ( \14254 , \11737 , RI992efc0_307);
and \U$13571 ( \14255 , \11816 , RI992d0d0_327);
nor \U$13572 ( \14256 , \14254 , \14255 );
and \U$13573 ( \14257 , \11734 , RI992a2e0_387);
and \U$13574 ( \14258 , \11726 , RI9928b70_407);
nor \U$13575 ( \14259 , \14257 , \14258 );
and \U$13576 ( \14260 , \11743 , RI992c770_347);
and \U$13577 ( \14261 , \11826 , RI992ac40_367);
nor \U$13578 ( \14262 , \14260 , \14261 );
and \U$13579 ( \14263 , \11756 , RI992f920_287);
not \U$13580 ( \14264 , RI9922360_587);
not \U$13581 ( \14265 , \11749 );
or \U$13582 ( \14266 , \14264 , \14265 );
nand \U$13583 ( \14267 , \10843 , RI99338e0_267);
nand \U$13584 ( \14268 , \14266 , \14267 );
nor \U$13585 ( \14269 , \14263 , \14268 );
nand \U$13586 ( \14270 , \14256 , \14259 , \14262 , \14269 );
nor \U$13587 ( \14271 , \14253 , \14270 );
not \U$13588 ( \14272 , \14271 );
buf \U$13589 ( \14273 , \14272 );
nand \U$13590 ( \14274 , \11637 , \14273 );
not \U$13591 ( \14275 , \14274 );
not \U$13592 ( \14276 , \13801 );
not \U$13593 ( \14277 , \12968 );
not \U$13594 ( \14278 , \14277 );
or \U$13595 ( \14279 , \14276 , \14278 );
nand \U$13596 ( \14280 , \12371 , \13503 );
nand \U$13597 ( \14281 , \14279 , \14280 );
not \U$13598 ( \14282 , \14281 );
not \U$13599 ( \14283 , \12375 );
or \U$13600 ( \14284 , \14282 , \14283 );
nand \U$13601 ( \14285 , \14023 , \13308 );
nand \U$13602 ( \14286 , \14284 , \14285 );
not \U$13603 ( \14287 , \14286 );
not \U$13604 ( \14288 , \14287 );
or \U$13605 ( \14289 , \14275 , \14288 );
and \U$13606 ( \14290 , \13147 , \12950 );
not \U$13607 ( \14291 , \13147 );
and \U$13608 ( \14292 , \14291 , \12662 );
or \U$13609 ( \14293 , \14290 , \14292 );
not \U$13610 ( \14294 , \14293 );
not \U$13611 ( \14295 , \13248 );
or \U$13612 ( \14296 , \14294 , \14295 );
nand \U$13613 ( \14297 , \14178 , \13251 );
nand \U$13614 ( \14298 , \14296 , \14297 );
not \U$13615 ( \14299 , \13270 );
not \U$13616 ( \14300 , \14187 );
or \U$13617 ( \14301 , \14299 , \14300 );
not \U$13618 ( \14302 , \13264 );
not \U$13619 ( \14303 , \12625 );
not \U$13620 ( \14304 , \14303 );
or \U$13621 ( \14305 , \14302 , \14304 );
nand \U$13622 ( \14306 , \12625 , \13521 );
nand \U$13623 ( \14307 , \14305 , \14306 );
nand \U$13624 ( \14308 , \14307 , \13259 );
nand \U$13625 ( \14309 , \14301 , \14308 );
nand \U$13626 ( \14310 , \14298 , \14309 );
not \U$13627 ( \14311 , \14310 );
nand \U$13628 ( \14312 , \14289 , \14311 );
not \U$13629 ( \14313 , \14274 );
nand \U$13630 ( \14314 , \14313 , \14286 );
nand \U$13631 ( \14315 , \14312 , \14314 );
xor \U$13632 ( \14316 , \14236 , \14315 );
not \U$13633 ( \14317 , \13751 );
not \U$13634 ( \14318 , \12992 );
or \U$13635 ( \14319 , \14317 , \14318 );
nand \U$13636 ( \14320 , \12199 , \13750 );
nand \U$13637 ( \14321 , \14319 , \14320 );
not \U$13638 ( \14322 , \14321 );
not \U$13639 ( \14323 , \12761 );
or \U$13640 ( \14324 , \14322 , \14323 );
nand \U$13641 ( \14325 , \14100 , \12837 );
nand \U$13642 ( \14326 , \14324 , \14325 );
not \U$13643 ( \14327 , \13942 );
not \U$13644 ( \14328 , \12012 );
or \U$13645 ( \14329 , \14327 , \14328 );
nand \U$13646 ( \14330 , \12322 , \13941 );
nand \U$13647 ( \14331 , \14329 , \14330 );
not \U$13648 ( \14332 , \14331 );
not \U$13649 ( \14333 , \12698 );
or \U$13650 ( \14334 , \14332 , \14333 );
not \U$13651 ( \14335 , \14110 );
nand \U$13652 ( \14336 , \14335 , \12002 );
nand \U$13653 ( \14337 , \14334 , \14336 );
xor \U$13654 ( \14338 , \14326 , \14337 );
not \U$13655 ( \14339 , \14168 );
not \U$13656 ( \14340 , \12533 );
or \U$13657 ( \14341 , \14339 , \14340 );
not \U$13658 ( \14342 , \14168 );
nand \U$13659 ( \14343 , \11890 , \14342 );
nand \U$13660 ( \14344 , \14341 , \14343 );
not \U$13661 ( \14345 , \14344 );
not \U$13662 ( \14346 , \11884 );
or \U$13663 ( \14347 , \14345 , \14346 );
nand \U$13664 ( \14348 , \14125 , \11873 );
nand \U$13665 ( \14349 , \14347 , \14348 );
and \U$13666 ( \14350 , \14338 , \14349 );
and \U$13667 ( \14351 , \14326 , \14337 );
or \U$13668 ( \14352 , \14350 , \14351 );
and \U$13669 ( \14353 , \14316 , \14352 );
and \U$13670 ( \14354 , \14236 , \14315 );
or \U$13671 ( \14355 , \14353 , \14354 );
not \U$13672 ( \14356 , \14355 );
xor \U$13673 ( \14357 , \14210 , \14173 );
xnor \U$13674 ( \14358 , \14357 , \14127 );
not \U$13675 ( \14359 , \14358 );
not \U$13676 ( \14360 , \14359 );
xor \U$13677 ( \14361 , \14094 , \14105 );
xor \U$13678 ( \14362 , \14361 , \14113 );
not \U$13679 ( \14363 , \14362 );
or \U$13680 ( \14364 , \14360 , \14363 );
not \U$13681 ( \14365 , \14362 );
not \U$13682 ( \14366 , \14365 );
not \U$13683 ( \14367 , \14358 );
or \U$13684 ( \14368 , \14366 , \14367 );
not \U$13685 ( \14369 , \13199 );
not \U$13686 ( \14370 , \13224 );
or \U$13687 ( \14371 , \14369 , \14370 );
not \U$13688 ( \14372 , \13198 );
nand \U$13689 ( \14373 , \12956 , \14372 );
nand \U$13690 ( \14374 , \14371 , \14373 );
not \U$13691 ( \14375 , \14374 );
not \U$13692 ( \14376 , \12681 );
or \U$13693 ( \14377 , \14375 , \14376 );
nand \U$13694 ( \14378 , \14203 , \12667 );
nand \U$13695 ( \14379 , \14377 , \14378 );
buf \U$13696 ( \14380 , \11633 );
not \U$13697 ( \14381 , \11850 );
not \U$13698 ( \14382 , \12323 );
or \U$13699 ( \14383 , \14381 , \14382 );
nand \U$13700 ( \14384 , \14383 , \14273 );
nand \U$13701 ( \14385 , \12032 , \11876 );
and \U$13702 ( \14386 , \14380 , \14384 , \14385 );
xor \U$13703 ( \14387 , \14379 , \14386 );
not \U$13704 ( \14388 , \13792 );
not \U$13705 ( \14389 , \12473 );
or \U$13706 ( \14390 , \14388 , \14389 );
nand \U$13707 ( \14391 , \12746 , \13793 );
nand \U$13708 ( \14392 , \14390 , \14391 );
not \U$13709 ( \14393 , \14392 );
not \U$13710 ( \14394 , \12375 );
or \U$13711 ( \14395 , \14393 , \14394 );
nand \U$13712 ( \14396 , \14281 , \13308 );
nand \U$13713 ( \14397 , \14395 , \14396 );
and \U$13714 ( \14398 , \14387 , \14397 );
and \U$13715 ( \14399 , \14379 , \14386 );
or \U$13716 ( \14400 , \14398 , \14399 );
not \U$13717 ( \14401 , \14400 );
xor \U$13718 ( \14402 , \14184 , \14191 );
xnor \U$13719 ( \14403 , \14402 , \14208 );
nand \U$13720 ( \14404 , \14401 , \14403 );
not \U$13721 ( \14405 , \14404 );
xor \U$13722 ( \14406 , \14309 , \14298 );
not \U$13723 ( \14407 , \13989 );
not \U$13724 ( \14408 , \12138 );
or \U$13725 ( \14409 , \14407 , \14408 );
nand \U$13726 ( \14410 , \12383 , \13993 );
nand \U$13727 ( \14411 , \14409 , \14410 );
not \U$13728 ( \14412 , \14411 );
not \U$13729 ( \14413 , \12761 );
or \U$13730 ( \14414 , \14412 , \14413 );
nand \U$13731 ( \14415 , \14321 , \12197 );
nand \U$13732 ( \14416 , \14414 , \14415 );
xor \U$13733 ( \14417 , \14406 , \14416 );
not \U$13734 ( \14418 , \13901 );
not \U$13735 ( \14419 , \12323 );
or \U$13736 ( \14420 , \14418 , \14419 );
nand \U$13737 ( \14421 , \12322 , \13902 );
nand \U$13738 ( \14422 , \14420 , \14421 );
not \U$13739 ( \14423 , \14422 );
not \U$13740 ( \14424 , \12016 );
or \U$13741 ( \14425 , \14423 , \14424 );
nand \U$13742 ( \14426 , \12002 , \14331 );
nand \U$13743 ( \14427 , \14425 , \14426 );
and \U$13744 ( \14428 , \14417 , \14427 );
and \U$13745 ( \14429 , \14406 , \14416 );
or \U$13746 ( \14430 , \14428 , \14429 );
not \U$13747 ( \14431 , \14430 );
or \U$13748 ( \14432 , \14405 , \14431 );
not \U$13749 ( \14433 , \14403 );
nand \U$13750 ( \14434 , \14433 , \14400 );
nand \U$13751 ( \14435 , \14432 , \14434 );
nand \U$13752 ( \14436 , \14368 , \14435 );
nand \U$13753 ( \14437 , \14364 , \14436 );
not \U$13754 ( \14438 , \14437 );
nand \U$13755 ( \14439 , \14356 , \14438 );
not \U$13756 ( \14440 , \14439 );
xor \U$13757 ( \14441 , \14220 , \14222 );
xor \U$13758 ( \14442 , \14441 , \14225 );
not \U$13759 ( \14443 , \14442 );
or \U$13760 ( \14444 , \14440 , \14443 );
not \U$13761 ( \14445 , \14438 );
nand \U$13762 ( \14446 , \14445 , \14355 );
nand \U$13763 ( \14447 , \14444 , \14446 );
not \U$13764 ( \14448 , \14447 );
nand \U$13765 ( \14449 , \14234 , \14448 );
nand \U$13766 ( \14450 , \14233 , \14447 );
and \U$13767 ( \14451 , \14355 , \14438 );
not \U$13768 ( \14452 , \14355 );
and \U$13769 ( \14453 , \14452 , \14437 );
nor \U$13770 ( \14454 , \14451 , \14453 );
not \U$13771 ( \14455 , \14454 );
not \U$13772 ( \14456 , \14442 );
or \U$13773 ( \14457 , \14455 , \14456 );
or \U$13774 ( \14458 , \14454 , \14442 );
nand \U$13775 ( \14459 , \14457 , \14458 );
xor \U$13776 ( \14460 , \14236 , \14315 );
xor \U$13777 ( \14461 , \14460 , \14352 );
xor \U$13778 ( \14462 , \14310 , \14286 );
xnor \U$13779 ( \14463 , \14462 , \14274 );
not \U$13780 ( \14464 , \14463 );
not \U$13781 ( \14465 , \14464 );
xor \U$13782 ( \14466 , \14326 , \14337 );
xor \U$13783 ( \14467 , \14466 , \14349 );
not \U$13784 ( \14468 , \14467 );
or \U$13785 ( \14469 , \14465 , \14468 );
or \U$13786 ( \14470 , \14467 , \14464 );
not \U$13787 ( \14471 , \13259 );
not \U$13788 ( \14472 , \13048 );
not \U$13789 ( \14473 , \12821 );
not \U$13790 ( \14474 , \14473 );
or \U$13791 ( \14475 , \14472 , \14474 );
nand \U$13792 ( \14476 , \12821 , \13261 );
nand \U$13793 ( \14477 , \14475 , \14476 );
not \U$13794 ( \14478 , \14477 );
or \U$13795 ( \14479 , \14471 , \14478 );
nand \U$13796 ( \14480 , \14307 , \13270 );
nand \U$13797 ( \14481 , \14479 , \14480 );
not \U$13798 ( \14482 , \14481 );
not \U$13799 ( \14483 , \14482 );
nand \U$13800 ( \14484 , \11872 , \14273 );
not \U$13801 ( \14485 , \14484 );
or \U$13802 ( \14486 , \14483 , \14485 );
and \U$13803 ( \14487 , \13097 , \13241 );
not \U$13804 ( \14488 , \13097 );
and \U$13805 ( \14489 , \14488 , \12662 );
or \U$13806 ( \14490 , \14487 , \14489 );
not \U$13807 ( \14491 , \14490 );
not \U$13808 ( \14492 , \13248 );
or \U$13809 ( \14493 , \14491 , \14492 );
nand \U$13810 ( \14494 , \14293 , \12936 );
nand \U$13811 ( \14495 , \14493 , \14494 );
nand \U$13812 ( \14496 , \14486 , \14495 );
or \U$13813 ( \14497 , \14484 , \14482 );
nand \U$13814 ( \14498 , \14496 , \14497 );
not \U$13815 ( \14499 , \14273 );
and \U$13816 ( \14500 , \14499 , \11891 );
not \U$13817 ( \14501 , \14499 );
and \U$13818 ( \14502 , \14501 , \12119 );
nor \U$13819 ( \14503 , \14500 , \14502 );
not \U$13820 ( \14504 , \14503 );
not \U$13821 ( \14505 , \11884 );
or \U$13822 ( \14506 , \14504 , \14505 );
nand \U$13823 ( \14507 , \14344 , \11873 );
nand \U$13824 ( \14508 , \14506 , \14507 );
xor \U$13825 ( \14509 , \14498 , \14508 );
not \U$13826 ( \14510 , \13801 );
not \U$13827 ( \14511 , \13224 );
or \U$13828 ( \14512 , \14510 , \14511 );
nand \U$13829 ( \14513 , \12956 , \13503 );
nand \U$13830 ( \14514 , \14512 , \14513 );
not \U$13831 ( \14515 , \14514 );
not \U$13832 ( \14516 , \12681 );
or \U$13833 ( \14517 , \14515 , \14516 );
nand \U$13834 ( \14518 , \14374 , \12667 );
nand \U$13835 ( \14519 , \14517 , \14518 );
not \U$13836 ( \14520 , \13199 );
not \U$13837 ( \14521 , \13241 );
or \U$13838 ( \14522 , \14520 , \14521 );
nand \U$13839 ( \14523 , \13244 , \14372 );
nand \U$13840 ( \14524 , \14522 , \14523 );
not \U$13841 ( \14525 , \14524 );
not \U$13842 ( \14526 , \12980 );
or \U$13843 ( \14527 , \14525 , \14526 );
nand \U$13844 ( \14528 , \14182 , \14490 );
nand \U$13845 ( \14529 , \14527 , \14528 );
not \U$13846 ( \14530 , \13259 );
not \U$13847 ( \14531 , \13264 );
not \U$13848 ( \14532 , \14531 );
not \U$13849 ( \14533 , \14532 );
not \U$13850 ( \14534 , \13148 );
or \U$13851 ( \14535 , \14533 , \14534 );
nand \U$13852 ( \14536 , \14001 , \14531 );
nand \U$13853 ( \14537 , \14535 , \14536 );
not \U$13854 ( \14538 , \14537 );
or \U$13855 ( \14539 , \14530 , \14538 );
nand \U$13856 ( \14540 , \14477 , \13270 );
nand \U$13857 ( \14541 , \14539 , \14540 );
and \U$13858 ( \14542 , \14529 , \14541 );
xor \U$13859 ( \14543 , \14519 , \14542 );
not \U$13860 ( \14544 , \13751 );
not \U$13861 ( \14545 , \14277 );
or \U$13862 ( \14546 , \14544 , \14545 );
nand \U$13863 ( \14547 , \13544 , \13750 );
nand \U$13864 ( \14548 , \14546 , \14547 );
not \U$13865 ( \14549 , \14548 );
not \U$13866 ( \14550 , \12375 );
or \U$13867 ( \14551 , \14549 , \14550 );
nand \U$13868 ( \14552 , \14392 , \12365 );
nand \U$13869 ( \14553 , \14551 , \14552 );
and \U$13870 ( \14554 , \14543 , \14553 );
and \U$13871 ( \14555 , \14519 , \14542 );
or \U$13872 ( \14556 , \14554 , \14555 );
and \U$13873 ( \14557 , \14509 , \14556 );
and \U$13874 ( \14558 , \14498 , \14508 );
or \U$13875 ( \14559 , \14557 , \14558 );
nand \U$13876 ( \14560 , \14470 , \14559 );
nand \U$13877 ( \14561 , \14469 , \14560 );
xor \U$13878 ( \14562 , \14461 , \14561 );
xor \U$13879 ( \14563 , \14362 , \14359 );
xor \U$13880 ( \14564 , \14563 , \14435 );
and \U$13881 ( \14565 , \14562 , \14564 );
and \U$13882 ( \14566 , \14461 , \14561 );
or \U$13883 ( \14567 , \14565 , \14566 );
nand \U$13884 ( \14568 , \14459 , \14567 );
nand \U$13885 ( \14569 , \14450 , \14568 );
nand \U$13886 ( \14570 , \14449 , \14569 );
and \U$13887 ( \14571 , \13844 , \13834 );
not \U$13888 ( \14572 , \13696 );
not \U$13889 ( \14573 , \12850 );
or \U$13890 ( \14574 , \14572 , \14573 );
not \U$13891 ( \14575 , \12247 );
not \U$13892 ( \14576 , \13224 );
or \U$13893 ( \14577 , \14575 , \14576 );
not \U$13894 ( \14578 , \12686 );
nand \U$13895 ( \14579 , \14578 , \12411 );
nand \U$13896 ( \14580 , \14577 , \14579 );
nand \U$13897 ( \14581 , \14580 , \12667 );
nand \U$13898 ( \14582 , \14574 , \14581 );
xor \U$13899 ( \14583 , \14571 , \14582 );
not \U$13900 ( \14584 , \13712 );
not \U$13901 ( \14585 , \12375 );
or \U$13902 ( \14586 , \14584 , \14585 );
not \U$13903 ( \14587 , \12627 );
not \U$13904 ( \14588 , \12637 );
or \U$13905 ( \14589 , \14587 , \14588 );
nand \U$13906 ( \14590 , \13544 , \12626 );
nand \U$13907 ( \14591 , \14589 , \14590 );
nand \U$13908 ( \14592 , \14591 , \12365 );
nand \U$13909 ( \14593 , \14586 , \14592 );
xor \U$13910 ( \14594 , \14583 , \14593 );
or \U$13911 ( \14595 , \13866 , \13855 );
nand \U$13912 ( \14596 , \14595 , \13845 );
nand \U$13913 ( \14597 , \13866 , \13855 );
and \U$13914 ( \14598 , \14596 , \14597 );
not \U$13915 ( \14599 , \14598 );
xor \U$13916 ( \14600 , \14594 , \14599 );
not \U$13917 ( \14601 , \13270 );
not \U$13918 ( \14602 , \13525 );
or \U$13919 ( \14603 , \14601 , \14602 );
nand \U$13920 ( \14604 , \13832 , \13259 );
nand \U$13921 ( \14605 , \14603 , \14604 );
not \U$13922 ( \14606 , \13842 );
not \U$13923 ( \14607 , \12980 );
or \U$13924 ( \14608 , \14606 , \14607 );
nand \U$13925 ( \14609 , \13513 , \13045 );
nand \U$13926 ( \14610 , \14608 , \14609 );
xor \U$13927 ( \14611 , \14605 , \14610 );
not \U$13928 ( \14612 , \13853 );
not \U$13929 ( \14613 , \12194 );
or \U$13930 ( \14614 , \14612 , \14613 );
not \U$13931 ( \14615 , \13149 );
not \U$13932 ( \14616 , \12992 );
or \U$13933 ( \14617 , \14615 , \14616 );
nand \U$13934 ( \14618 , \12137 , \13148 );
nand \U$13935 ( \14619 , \14617 , \14618 );
nand \U$13936 ( \14620 , \14619 , \12197 );
nand \U$13937 ( \14621 , \14614 , \14620 );
xor \U$13938 ( \14622 , \14611 , \14621 );
not \U$13939 ( \14623 , \13864 );
or \U$13940 ( \14624 , \12017 , \14623 );
and \U$13941 ( \14625 , \13457 , \12029 );
not \U$13942 ( \14626 , \13457 );
and \U$13943 ( \14627 , \14626 , \12323 );
nor \U$13944 ( \14628 , \14625 , \14627 );
or \U$13945 ( \14629 , \12524 , \14628 );
nand \U$13946 ( \14630 , \14624 , \14629 );
xor \U$13947 ( \14631 , \14622 , \14630 );
xnor \U$13948 ( \14632 , \14600 , \14631 );
xor \U$13949 ( \14633 , \14038 , \14090 );
and \U$13950 ( \14634 , \14633 , \14216 );
and \U$13951 ( \14635 , \14038 , \14090 );
or \U$13952 ( \14636 , \14634 , \14635 );
not \U$13953 ( \14637 , \14636 );
xor \U$13954 ( \14638 , \14632 , \14637 );
xor \U$13955 ( \14639 , \14043 , \14054 );
and \U$13956 ( \14640 , \14639 , \14089 );
and \U$13957 ( \14641 , \14043 , \14054 );
or \U$13958 ( \14642 , \14640 , \14641 );
not \U$13959 ( \14643 , \14642 );
and \U$13960 ( \14644 , \13993 , \11639 );
not \U$13961 ( \14645 , \13993 );
and \U$13962 ( \14646 , \14645 , \12827 );
nor \U$13963 ( \14647 , \14644 , \14646 );
and \U$13964 ( \14648 , \11637 , \14647 );
not \U$13965 ( \14649 , \14048 );
not \U$13966 ( \14650 , \11884 );
or \U$13967 ( \14651 , \14649 , \14650 );
and \U$13968 ( \14652 , \13792 , \12118 );
not \U$13969 ( \14653 , \13792 );
and \U$13970 ( \14654 , \14653 , \12534 );
or \U$13971 ( \14655 , \14652 , \14654 );
nand \U$13972 ( \14656 , \14655 , \12540 );
nand \U$13973 ( \14657 , \14651 , \14656 );
xor \U$13974 ( \14658 , \14648 , \14657 );
nor \U$13975 ( \14659 , \13714 , \13698 );
or \U$13976 ( \14660 , \14659 , \13684 );
nand \U$13977 ( \14661 , \13714 , \13698 );
nand \U$13978 ( \14662 , \14660 , \14661 );
xor \U$13979 ( \14663 , \14658 , \14662 );
not \U$13980 ( \14664 , \14663 );
not \U$13981 ( \14665 , \14664 );
or \U$13982 ( \14666 , \14643 , \14665 );
not \U$13983 ( \14667 , \14642 );
nand \U$13984 ( \14668 , \14663 , \14667 );
nand \U$13985 ( \14669 , \14666 , \14668 );
not \U$13986 ( \14670 , \13715 );
not \U$13987 ( \14671 , \14670 );
not \U$13988 ( \14672 , \13823 );
or \U$13989 ( \14673 , \14671 , \14672 );
not \U$13990 ( \14674 , \13715 );
not \U$13991 ( \14675 , \13822 );
or \U$13992 ( \14676 , \14674 , \14675 );
nand \U$13993 ( \14677 , \14676 , \13867 );
nand \U$13994 ( \14678 , \14673 , \14677 );
not \U$13995 ( \14679 , \14678 );
and \U$13996 ( \14680 , \14669 , \14679 );
not \U$13997 ( \14681 , \14669 );
and \U$13998 ( \14682 , \14681 , \14678 );
nor \U$13999 ( \14683 , \14680 , \14682 );
xor \U$14000 ( \14684 , \14638 , \14683 );
or \U$14001 ( \14685 , \14217 , \13868 );
and \U$14002 ( \14686 , \14685 , \14228 );
and \U$14003 ( \14687 , \13868 , \14217 );
nor \U$14004 ( \14688 , \14686 , \14687 );
nand \U$14005 ( \14689 , \14684 , \14688 );
nand \U$14006 ( \14690 , \14610 , \14605 );
not \U$14007 ( \14691 , \14580 );
not \U$14008 ( \14692 , \12681 );
or \U$14009 ( \14693 , \14691 , \14692 );
nand \U$14010 ( \14694 , \13535 , \12667 );
nand \U$14011 ( \14695 , \14693 , \14694 );
xor \U$14012 ( \14696 , \14690 , \14695 );
not \U$14013 ( \14697 , \14591 );
not \U$14014 ( \14698 , \12644 );
or \U$14015 ( \14699 , \14697 , \14698 );
nand \U$14016 ( \14700 , \13546 , \12364 );
nand \U$14017 ( \14701 , \14699 , \14700 );
xnor \U$14018 ( \14702 , \14696 , \14701 );
xor \U$14019 ( \14703 , \14611 , \14621 );
and \U$14020 ( \14704 , \14703 , \14630 );
and \U$14021 ( \14705 , \14611 , \14621 );
or \U$14022 ( \14706 , \14704 , \14705 );
xor \U$14023 ( \14707 , \14702 , \14706 );
xor \U$14024 ( \14708 , \13529 , \13518 );
not \U$14025 ( \14709 , \14619 );
not \U$14026 ( \14710 , \12761 );
or \U$14027 ( \14711 , \14709 , \14710 );
nand \U$14028 ( \14712 , \12197 , \13577 );
nand \U$14029 ( \14713 , \14711 , \14712 );
xor \U$14030 ( \14714 , \14708 , \14713 );
not \U$14031 ( \14715 , \14628 );
not \U$14032 ( \14716 , \14715 );
not \U$14033 ( \14717 , \12521 );
or \U$14034 ( \14718 , \14716 , \14717 );
nand \U$14035 ( \14719 , \12002 , \13588 );
nand \U$14036 ( \14720 , \14718 , \14719 );
xor \U$14037 ( \14721 , \14714 , \14720 );
xnor \U$14038 ( \14722 , \14707 , \14721 );
not \U$14039 ( \14723 , \14678 );
nand \U$14040 ( \14724 , \14664 , \14667 );
not \U$14041 ( \14725 , \14724 );
or \U$14042 ( \14726 , \14723 , \14725 );
nand \U$14043 ( \14727 , \14663 , \14642 );
nand \U$14044 ( \14728 , \14726 , \14727 );
not \U$14045 ( \14729 , \14728 );
xor \U$14046 ( \14730 , \14722 , \14729 );
and \U$14047 ( \14731 , \13751 , \12827 );
not \U$14048 ( \14732 , \13751 );
and \U$14049 ( \14733 , \14732 , \11639 );
nor \U$14050 ( \14734 , \14731 , \14733 );
and \U$14051 ( \14735 , \11637 , \14734 );
not \U$14052 ( \14736 , \14655 );
not \U$14053 ( \14737 , \11884 );
or \U$14054 ( \14738 , \14736 , \14737 );
not \U$14055 ( \14739 , \13801 );
not \U$14056 ( \14740 , \11889 );
or \U$14057 ( \14741 , \14739 , \14740 );
nand \U$14058 ( \14742 , \14380 , \13503 );
nand \U$14059 ( \14743 , \14741 , \14742 );
nand \U$14060 ( \14744 , \14743 , \12540 );
nand \U$14061 ( \14745 , \14738 , \14744 );
xor \U$14062 ( \14746 , \14735 , \14745 );
xor \U$14063 ( \14747 , \14571 , \14582 );
and \U$14064 ( \14748 , \14747 , \14593 );
and \U$14065 ( \14749 , \14571 , \14582 );
or \U$14066 ( \14750 , \14748 , \14749 );
xor \U$14067 ( \14751 , \14746 , \14750 );
xor \U$14068 ( \14752 , \14648 , \14657 );
and \U$14069 ( \14753 , \14752 , \14662 );
and \U$14070 ( \14754 , \14648 , \14657 );
or \U$14071 ( \14755 , \14753 , \14754 );
and \U$14072 ( \14756 , \14751 , \14755 );
not \U$14073 ( \14757 , \14751 );
not \U$14074 ( \14758 , \14755 );
and \U$14075 ( \14759 , \14757 , \14758 );
nor \U$14076 ( \14760 , \14756 , \14759 );
not \U$14077 ( \14761 , \14594 );
nand \U$14078 ( \14762 , \14761 , \14598 );
not \U$14079 ( \14763 , \14762 );
not \U$14080 ( \14764 , \14631 );
or \U$14081 ( \14765 , \14763 , \14764 );
nand \U$14082 ( \14766 , \14599 , \14594 );
nand \U$14083 ( \14767 , \14765 , \14766 );
not \U$14084 ( \14768 , \14767 );
and \U$14085 ( \14769 , \14760 , \14768 );
not \U$14086 ( \14770 , \14760 );
and \U$14087 ( \14771 , \14770 , \14767 );
nor \U$14088 ( \14772 , \14769 , \14771 );
xor \U$14089 ( \14773 , \14730 , \14772 );
xor \U$14090 ( \14774 , \14632 , \14637 );
and \U$14091 ( \14775 , \14774 , \14683 );
and \U$14092 ( \14776 , \14632 , \14637 );
or \U$14093 ( \14777 , \14775 , \14776 );
nand \U$14094 ( \14778 , \14773 , \14777 );
nand \U$14095 ( \14779 , \14689 , \14778 );
nor \U$14096 ( \14780 , \14570 , \14779 );
not \U$14097 ( \14781 , \14780 );
nor \U$14098 ( \14782 , \14684 , \14688 );
not \U$14099 ( \14783 , \14782 );
not \U$14100 ( \14784 , \14778 );
or \U$14101 ( \14785 , \14783 , \14784 );
or \U$14102 ( \14786 , \14773 , \14777 );
nand \U$14103 ( \14787 , \14785 , \14786 );
not \U$14104 ( \14788 , \14787 );
nand \U$14105 ( \14789 , \14781 , \14788 );
xor \U$14106 ( \14790 , \13565 , \13596 );
xnor \U$14107 ( \14791 , \14790 , \13601 );
xor \U$14108 ( \14792 , \13530 , \13540 );
xor \U$14109 ( \14793 , \14792 , \13551 );
not \U$14110 ( \14794 , \14793 );
not \U$14111 ( \14795 , \14794 );
xor \U$14112 ( \14796 , \14708 , \14713 );
and \U$14113 ( \14797 , \14796 , \14720 );
and \U$14114 ( \14798 , \14708 , \14713 );
or \U$14115 ( \14799 , \14797 , \14798 );
not \U$14116 ( \14800 , \14799 );
not \U$14117 ( \14801 , \14800 );
or \U$14118 ( \14802 , \14795 , \14801 );
xor \U$14119 ( \14803 , \13572 , \13582 );
xor \U$14120 ( \14804 , \14803 , \13593 );
nand \U$14121 ( \14805 , \14802 , \14804 );
nand \U$14122 ( \14806 , \14799 , \14793 );
nand \U$14123 ( \14807 , \14805 , \14806 );
not \U$14124 ( \14808 , \14807 );
xor \U$14125 ( \14809 , \13508 , \13463 );
xnor \U$14126 ( \14810 , \14809 , \13554 );
not \U$14127 ( \14811 , \14810 );
and \U$14128 ( \14812 , \13792 , \11634 );
not \U$14129 ( \14813 , \13792 );
and \U$14130 ( \14814 , \14813 , \11635 );
nor \U$14131 ( \14815 , \14812 , \14814 );
and \U$14132 ( \14816 , \11636 , \14815 );
not \U$14133 ( \14817 , \14743 );
not \U$14134 ( \14818 , \13452 );
or \U$14135 ( \14819 , \14817 , \14818 );
nand \U$14136 ( \14820 , \13459 , \11873 );
nand \U$14137 ( \14821 , \14819 , \14820 );
xor \U$14138 ( \14822 , \14816 , \14821 );
nor \U$14139 ( \14823 , \14701 , \14695 );
or \U$14140 ( \14824 , \14823 , \14690 );
nand \U$14141 ( \14825 , \14701 , \14695 );
nand \U$14142 ( \14826 , \14824 , \14825 );
and \U$14143 ( \14827 , \14822 , \14826 );
and \U$14144 ( \14828 , \14816 , \14821 );
or \U$14145 ( \14829 , \14827 , \14828 );
not \U$14146 ( \14830 , \14829 );
not \U$14147 ( \14831 , \14830 );
and \U$14148 ( \14832 , \14811 , \14831 );
and \U$14149 ( \14833 , \14810 , \14830 );
nor \U$14150 ( \14834 , \14832 , \14833 );
not \U$14151 ( \14835 , \14834 );
or \U$14152 ( \14836 , \14808 , \14835 );
not \U$14153 ( \14837 , \14834 );
not \U$14154 ( \14838 , \14807 );
nand \U$14155 ( \14839 , \14837 , \14838 );
nand \U$14156 ( \14840 , \14836 , \14839 );
xor \U$14157 ( \14841 , \14791 , \14840 );
xor \U$14158 ( \14842 , \14735 , \14745 );
and \U$14159 ( \14843 , \14842 , \14750 );
and \U$14160 ( \14844 , \14735 , \14745 );
or \U$14161 ( \14845 , \14843 , \14844 );
not \U$14162 ( \14846 , \14845 );
xor \U$14163 ( \14847 , \14816 , \14821 );
xor \U$14164 ( \14848 , \14847 , \14826 );
not \U$14165 ( \14849 , \14848 );
or \U$14166 ( \14850 , \14846 , \14849 );
or \U$14167 ( \14851 , \14706 , \14702 );
nand \U$14168 ( \14852 , \14851 , \14721 );
nand \U$14169 ( \14853 , \14706 , \14702 );
nand \U$14170 ( \14854 , \14852 , \14853 );
not \U$14171 ( \14855 , \14848 );
not \U$14172 ( \14856 , \14845 );
nand \U$14173 ( \14857 , \14855 , \14856 );
nand \U$14174 ( \14858 , \14854 , \14857 );
nand \U$14175 ( \14859 , \14850 , \14858 );
xor \U$14176 ( \14860 , \14841 , \14859 );
buf \U$14177 ( \14861 , \14799 );
xor \U$14178 ( \14862 , \14793 , \14861 );
xnor \U$14179 ( \14863 , \14862 , \14804 );
not \U$14180 ( \14864 , \14767 );
not \U$14181 ( \14865 , \14751 );
nand \U$14182 ( \14866 , \14865 , \14758 );
not \U$14183 ( \14867 , \14866 );
or \U$14184 ( \14868 , \14864 , \14867 );
not \U$14185 ( \14869 , \14865 );
nand \U$14186 ( \14870 , \14869 , \14755 );
nand \U$14187 ( \14871 , \14868 , \14870 );
not \U$14188 ( \14872 , \14871 );
xor \U$14189 ( \14873 , \14863 , \14872 );
not \U$14190 ( \14874 , \14845 );
not \U$14191 ( \14875 , \14855 );
or \U$14192 ( \14876 , \14874 , \14875 );
nand \U$14193 ( \14877 , \14848 , \14856 );
nand \U$14194 ( \14878 , \14876 , \14877 );
not \U$14195 ( \14879 , \14854 );
and \U$14196 ( \14880 , \14878 , \14879 );
not \U$14197 ( \14881 , \14878 );
and \U$14198 ( \14882 , \14881 , \14854 );
nor \U$14199 ( \14883 , \14880 , \14882 );
and \U$14200 ( \14884 , \14873 , \14883 );
and \U$14201 ( \14885 , \14863 , \14872 );
or \U$14202 ( \14886 , \14884 , \14885 );
nand \U$14203 ( \14887 , \14860 , \14886 );
xor \U$14204 ( \14888 , \13319 , \13350 );
xnor \U$14205 ( \14889 , \14888 , \13354 );
not \U$14206 ( \14890 , \14810 );
nand \U$14207 ( \14891 , \14890 , \14830 );
and \U$14208 ( \14892 , \14891 , \14807 );
nor \U$14209 ( \14893 , \14890 , \14830 );
nor \U$14210 ( \14894 , \14892 , \14893 );
xor \U$14211 ( \14895 , \14889 , \14894 );
not \U$14212 ( \14896 , \13606 );
not \U$14213 ( \14897 , \13561 );
or \U$14214 ( \14898 , \14896 , \14897 );
nand \U$14215 ( \14899 , \13605 , \13558 );
nand \U$14216 ( \14900 , \14898 , \14899 );
not \U$14217 ( \14901 , \13603 );
and \U$14218 ( \14902 , \14900 , \14901 );
not \U$14219 ( \14903 , \14900 );
and \U$14220 ( \14904 , \14903 , \13603 );
nor \U$14221 ( \14905 , \14902 , \14904 );
xor \U$14222 ( \14906 , \14895 , \14905 );
not \U$14223 ( \14907 , \14840 );
nand \U$14224 ( \14908 , \14907 , \14791 );
and \U$14225 ( \14909 , \14908 , \14859 );
nor \U$14226 ( \14910 , \14907 , \14791 );
nor \U$14227 ( \14911 , \14909 , \14910 );
nand \U$14228 ( \14912 , \14906 , \14911 );
xor \U$14229 ( \14913 , \14863 , \14872 );
xor \U$14230 ( \14914 , \14913 , \14883 );
xor \U$14231 ( \14915 , \14722 , \14729 );
and \U$14232 ( \14916 , \14915 , \14772 );
and \U$14233 ( \14917 , \14722 , \14729 );
or \U$14234 ( \14918 , \14916 , \14917 );
nand \U$14235 ( \14919 , \14914 , \14918 );
xor \U$14236 ( \14920 , \13449 , \13609 );
xnor \U$14237 ( \14921 , \14920 , \13447 );
xor \U$14238 ( \14922 , \14889 , \14894 );
and \U$14239 ( \14923 , \14922 , \14905 );
and \U$14240 ( \14924 , \14889 , \14894 );
or \U$14241 ( \14925 , \14923 , \14924 );
nand \U$14242 ( \14926 , \14921 , \14925 );
nand \U$14243 ( \14927 , \14887 , \14912 , \14919 , \14926 );
not \U$14244 ( \14928 , \14927 );
buf \U$14245 ( \14929 , \14928 );
nand \U$14246 ( \14930 , \14789 , \14929 );
xor \U$14247 ( \14931 , \14379 , \14386 );
xor \U$14248 ( \14932 , \14931 , \14397 );
xor \U$14249 ( \14933 , \14406 , \14416 );
xor \U$14250 ( \14934 , \14933 , \14427 );
xor \U$14251 ( \14935 , \14932 , \14934 );
not \U$14252 ( \14936 , \14484 );
and \U$14253 ( \14937 , \14495 , \14481 );
not \U$14254 ( \14938 , \14495 );
and \U$14255 ( \14939 , \14938 , \14482 );
nor \U$14256 ( \14940 , \14937 , \14939 );
not \U$14257 ( \14941 , \14940 );
or \U$14258 ( \14942 , \14936 , \14941 );
or \U$14259 ( \14943 , \14484 , \14940 );
nand \U$14260 ( \14944 , \14942 , \14943 );
not \U$14261 ( \14945 , \13942 );
not \U$14262 ( \14946 , \12138 );
or \U$14263 ( \14947 , \14945 , \14946 );
nand \U$14264 ( \14948 , \12383 , \13941 );
nand \U$14265 ( \14949 , \14947 , \14948 );
not \U$14266 ( \14950 , \14949 );
not \U$14267 ( \14951 , \12194 );
or \U$14268 ( \14952 , \14950 , \14951 );
nand \U$14269 ( \14953 , \14411 , \12837 );
nand \U$14270 ( \14954 , \14952 , \14953 );
xor \U$14271 ( \14955 , \14944 , \14954 );
not \U$14272 ( \14956 , \14168 );
not \U$14273 ( \14957 , \12029 );
not \U$14274 ( \14958 , \14957 );
or \U$14275 ( \14959 , \14956 , \14958 );
nand \U$14276 ( \14960 , \12032 , \14342 );
nand \U$14277 ( \14961 , \14959 , \14960 );
not \U$14278 ( \14962 , \14961 );
not \U$14279 ( \14963 , \12399 );
or \U$14280 ( \14964 , \14962 , \14963 );
nand \U$14281 ( \14965 , \12003 , \14422 );
nand \U$14282 ( \14966 , \14964 , \14965 );
and \U$14283 ( \14967 , \14955 , \14966 );
and \U$14284 ( \14968 , \14944 , \14954 );
or \U$14285 ( \14969 , \14967 , \14968 );
and \U$14286 ( \14970 , \14935 , \14969 );
and \U$14287 ( \14971 , \14932 , \14934 );
or \U$14288 ( \14972 , \14970 , \14971 );
not \U$14289 ( \14973 , \14972 );
xor \U$14290 ( \14974 , \14400 , \14403 );
xor \U$14291 ( \14975 , \14974 , \14430 );
not \U$14292 ( \14976 , \14975 );
and \U$14293 ( \14977 , \14973 , \14976 );
and \U$14294 ( \14978 , \14972 , \14975 );
nor \U$14295 ( \14979 , \14977 , \14978 );
not \U$14296 ( \14980 , \14979 );
xor \U$14297 ( \14981 , \14463 , \14467 );
xor \U$14298 ( \14982 , \14981 , \14559 );
not \U$14299 ( \14983 , \14982 );
not \U$14300 ( \14984 , \14983 );
and \U$14301 ( \14985 , \14980 , \14984 );
and \U$14302 ( \14986 , \14983 , \14979 );
nor \U$14303 ( \14987 , \14985 , \14986 );
xor \U$14304 ( \14988 , \14498 , \14508 );
xor \U$14305 ( \14989 , \14988 , \14556 );
not \U$14306 ( \14990 , \13792 );
not \U$14307 ( \14991 , \12686 );
or \U$14308 ( \14992 , \14990 , \14991 );
nand \U$14309 ( \14993 , \12956 , \13793 );
nand \U$14310 ( \14994 , \14992 , \14993 );
not \U$14311 ( \14995 , \14994 );
not \U$14312 ( \14996 , \12681 );
or \U$14313 ( \14997 , \14995 , \14996 );
nand \U$14314 ( \14998 , \14514 , \12667 );
nand \U$14315 ( \14999 , \14997 , \14998 );
not \U$14316 ( \15000 , \12383 );
buf \U$14317 ( \15001 , \12011 );
not \U$14318 ( \15002 , \15001 );
nand \U$14319 ( \15003 , \15000 , \15002 );
and \U$14320 ( \15004 , \15003 , \14273 );
not \U$14321 ( \15005 , \12383 );
not \U$14322 ( \15006 , \15001 );
or \U$14323 ( \15007 , \15005 , \15006 );
nand \U$14324 ( \15008 , \15007 , \12326 );
nor \U$14325 ( \15009 , \15004 , \15008 );
xor \U$14326 ( \15010 , \14999 , \15009 );
and \U$14327 ( \15011 , \12637 , \13989 );
not \U$14328 ( \15012 , \12637 );
and \U$14329 ( \15013 , \15012 , \13993 );
or \U$14330 ( \15014 , \15011 , \15013 );
not \U$14331 ( \15015 , \15014 );
not \U$14332 ( \15016 , \12375 );
or \U$14333 ( \15017 , \15015 , \15016 );
nand \U$14334 ( \15018 , \12365 , \14548 );
nand \U$14335 ( \15019 , \15017 , \15018 );
and \U$14336 ( \15020 , \15010 , \15019 );
and \U$14337 ( \15021 , \14999 , \15009 );
or \U$14338 ( \15022 , \15020 , \15021 );
xor \U$14339 ( \15023 , \14519 , \14542 );
xor \U$14340 ( \15024 , \15023 , \14553 );
xor \U$14341 ( \15025 , \15022 , \15024 );
xor \U$14342 ( \15026 , \14541 , \14529 );
not \U$14343 ( \15027 , \13902 );
not \U$14344 ( \15028 , \12199 );
or \U$14345 ( \15029 , \15027 , \15028 );
not \U$14346 ( \15030 , \12383 );
nand \U$14347 ( \15031 , \15030 , \13901 );
nand \U$14348 ( \15032 , \15029 , \15031 );
not \U$14349 ( \15033 , \15032 );
not \U$14350 ( \15034 , \12194 );
or \U$14351 ( \15035 , \15033 , \15034 );
nand \U$14352 ( \15036 , \14949 , \12197 );
nand \U$14353 ( \15037 , \15035 , \15036 );
xor \U$14354 ( \15038 , \15026 , \15037 );
not \U$14355 ( \15039 , \14273 );
not \U$14356 ( \15040 , \12323 );
or \U$14357 ( \15041 , \15039 , \15040 );
nand \U$14358 ( \15042 , \12029 , \14499 );
nand \U$14359 ( \15043 , \15041 , \15042 );
not \U$14360 ( \15044 , \15043 );
not \U$14361 ( \15045 , \12521 );
or \U$14362 ( \15046 , \15044 , \15045 );
nand \U$14363 ( \15047 , \12003 , \14961 );
nand \U$14364 ( \15048 , \15046 , \15047 );
and \U$14365 ( \15049 , \15038 , \15048 );
and \U$14366 ( \15050 , \15026 , \15037 );
or \U$14367 ( \15051 , \15049 , \15050 );
and \U$14368 ( \15052 , \15025 , \15051 );
and \U$14369 ( \15053 , \15022 , \15024 );
or \U$14370 ( \15054 , \15052 , \15053 );
xor \U$14371 ( \15055 , \14989 , \15054 );
xor \U$14372 ( \15056 , \14932 , \14934 );
xor \U$14373 ( \15057 , \15056 , \14969 );
and \U$14374 ( \15058 , \15055 , \15057 );
and \U$14375 ( \15059 , \14989 , \15054 );
or \U$14376 ( \15060 , \15058 , \15059 );
not \U$14377 ( \15061 , \15060 );
nand \U$14378 ( \15062 , \14987 , \15061 );
not \U$14379 ( \15063 , \15062 );
xor \U$14380 ( \15064 , \14989 , \15054 );
xor \U$14381 ( \15065 , \15064 , \15057 );
xor \U$14382 ( \15066 , \15022 , \15024 );
xor \U$14383 ( \15067 , \15066 , \15051 );
not \U$14384 ( \15068 , \15067 );
not \U$14385 ( \15069 , \13259 );
and \U$14386 ( \15070 , \14532 , \13098 );
not \U$14387 ( \15071 , \14532 );
and \U$14388 ( \15072 , \15071 , \13102 );
nor \U$14389 ( \15073 , \15070 , \15072 );
not \U$14390 ( \15074 , \15073 );
or \U$14391 ( \15075 , \15069 , \15074 );
nand \U$14392 ( \15076 , \14537 , \13270 );
nand \U$14393 ( \15077 , \15075 , \15076 );
not \U$14394 ( \15078 , \13801 );
not \U$14395 ( \15079 , \13241 );
or \U$14396 ( \15080 , \15078 , \15079 );
nand \U$14397 ( \15081 , \13244 , \13503 );
nand \U$14398 ( \15082 , \15080 , \15081 );
not \U$14399 ( \15083 , \15082 );
not \U$14400 ( \15084 , \12980 );
or \U$14401 ( \15085 , \15083 , \15084 );
nand \U$14402 ( \15086 , \14524 , \14182 );
nand \U$14403 ( \15087 , \15085 , \15086 );
xor \U$14404 ( \15088 , \15077 , \15087 );
and \U$14405 ( \15089 , \12002 , \14273 );
and \U$14406 ( \15090 , \15088 , \15089 );
and \U$14407 ( \15091 , \15077 , \15087 );
or \U$14408 ( \15092 , \15090 , \15091 );
xor \U$14409 ( \15093 , \14999 , \15009 );
xor \U$14410 ( \15094 , \15093 , \15019 );
xor \U$14411 ( \15095 , \15092 , \15094 );
not \U$14412 ( \15096 , \13792 );
not \U$14413 ( \15097 , \12950 );
or \U$14414 ( \15098 , \15096 , \15097 );
nand \U$14415 ( \15099 , \13244 , \13793 );
nand \U$14416 ( \15100 , \15098 , \15099 );
not \U$14417 ( \15101 , \15100 );
not \U$14418 ( \15102 , \12980 );
or \U$14419 ( \15103 , \15101 , \15102 );
nand \U$14420 ( \15104 , \15082 , \14182 );
nand \U$14421 ( \15105 , \15103 , \15104 );
not \U$14422 ( \15106 , \13270 );
not \U$14423 ( \15107 , \15073 );
or \U$14424 ( \15108 , \15106 , \15107 );
not \U$14425 ( \15109 , \13269 );
not \U$14426 ( \15110 , \14372 );
or \U$14427 ( \15111 , \15109 , \15110 );
nand \U$14428 ( \15112 , \13198 , \14531 );
nand \U$14429 ( \15113 , \15111 , \15112 );
nand \U$14430 ( \15114 , \15113 , \13259 );
nand \U$14431 ( \15115 , \15108 , \15114 );
and \U$14432 ( \15116 , \15105 , \15115 );
not \U$14433 ( \15117 , \13751 );
not \U$14434 ( \15118 , \13224 );
or \U$14435 ( \15119 , \15117 , \15118 );
nand \U$14436 ( \15120 , \12956 , \13750 );
nand \U$14437 ( \15121 , \15119 , \15120 );
not \U$14438 ( \15122 , \15121 );
not \U$14439 ( \15123 , \12682 );
not \U$14440 ( \15124 , \15123 );
or \U$14441 ( \15125 , \15122 , \15124 );
nand \U$14442 ( \15126 , \14994 , \12667 );
nand \U$14443 ( \15127 , \15125 , \15126 );
xor \U$14444 ( \15128 , \15116 , \15127 );
not \U$14445 ( \15129 , \13942 );
not \U$14446 ( \15130 , \12481 );
or \U$14447 ( \15131 , \15129 , \15130 );
nand \U$14448 ( \15132 , \12371 , \13941 );
nand \U$14449 ( \15133 , \15131 , \15132 );
not \U$14450 ( \15134 , \15133 );
or \U$14451 ( \15135 , \12376 , \15134 );
not \U$14452 ( \15136 , \15014 );
or \U$14453 ( \15137 , \12366 , \15136 );
nand \U$14454 ( \15138 , \15135 , \15137 );
and \U$14455 ( \15139 , \15128 , \15138 );
and \U$14456 ( \15140 , \15116 , \15127 );
or \U$14457 ( \15141 , \15139 , \15140 );
and \U$14458 ( \15142 , \15095 , \15141 );
and \U$14459 ( \15143 , \15092 , \15094 );
or \U$14460 ( \15144 , \15142 , \15143 );
not \U$14461 ( \15145 , \15144 );
xor \U$14462 ( \15146 , \14944 , \14954 );
xor \U$14463 ( \15147 , \15146 , \14966 );
not \U$14464 ( \15148 , \15147 );
nand \U$14465 ( \15149 , \15145 , \15148 );
not \U$14466 ( \15150 , \15149 );
or \U$14467 ( \15151 , \15068 , \15150 );
nand \U$14468 ( \15152 , \15144 , \15147 );
nand \U$14469 ( \15153 , \15151 , \15152 );
nand \U$14470 ( \15154 , \15065 , \15153 );
not \U$14471 ( \15155 , \15154 );
and \U$14472 ( \15156 , \15144 , \15147 );
not \U$14473 ( \15157 , \15144 );
and \U$14474 ( \15158 , \15157 , \15148 );
nor \U$14475 ( \15159 , \15156 , \15158 );
and \U$14476 ( \15160 , \15159 , \15067 );
not \U$14477 ( \15161 , \15159 );
not \U$14478 ( \15162 , \15067 );
and \U$14479 ( \15163 , \15161 , \15162 );
nor \U$14480 ( \15164 , \15160 , \15163 );
xor \U$14481 ( \15165 , \15026 , \15037 );
xor \U$14482 ( \15166 , \15165 , \15048 );
not \U$14483 ( \15167 , \14168 );
not \U$14484 ( \15168 , \12138 );
or \U$14485 ( \15169 , \15167 , \15168 );
nand \U$14486 ( \15170 , \12137 , \14342 );
nand \U$14487 ( \15171 , \15169 , \15170 );
not \U$14488 ( \15172 , \15171 );
not \U$14489 ( \15173 , \12194 );
or \U$14490 ( \15174 , \15172 , \15173 );
nand \U$14491 ( \15175 , \15032 , \12197 );
nand \U$14492 ( \15176 , \15174 , \15175 );
not \U$14493 ( \15177 , \12198 );
not \U$14494 ( \15178 , \12157 );
not \U$14495 ( \15179 , \12637 );
or \U$14496 ( \15180 , \15178 , \15179 );
nand \U$14497 ( \15181 , \15180 , \14273 );
nand \U$14498 ( \15182 , \12968 , \12152 );
nand \U$14499 ( \15183 , \15177 , \15181 , \15182 );
not \U$14500 ( \15184 , \15183 );
not \U$14501 ( \15185 , \12681 );
not \U$14502 ( \15186 , \13989 );
not \U$14503 ( \15187 , \12686 );
or \U$14504 ( \15188 , \15186 , \15187 );
nand \U$14505 ( \15189 , \12846 , \13993 );
nand \U$14506 ( \15190 , \15188 , \15189 );
not \U$14507 ( \15191 , \15190 );
or \U$14508 ( \15192 , \15185 , \15191 );
nand \U$14509 ( \15193 , \15121 , \12667 );
nand \U$14510 ( \15194 , \15192 , \15193 );
not \U$14511 ( \15195 , \15194 );
not \U$14512 ( \15196 , \15195 );
or \U$14513 ( \15197 , \15184 , \15196 );
xor \U$14514 ( \15198 , \15115 , \15105 );
nand \U$14515 ( \15199 , \15197 , \15198 );
not \U$14516 ( \15200 , \15195 );
not \U$14517 ( \15201 , \15183 );
nand \U$14518 ( \15202 , \15200 , \15201 );
nand \U$14519 ( \15203 , \15199 , \15202 );
xor \U$14520 ( \15204 , \15176 , \15203 );
xor \U$14521 ( \15205 , \15077 , \15087 );
xor \U$14522 ( \15206 , \15205 , \15089 );
and \U$14523 ( \15207 , \15204 , \15206 );
and \U$14524 ( \15208 , \15176 , \15203 );
or \U$14525 ( \15209 , \15207 , \15208 );
xor \U$14526 ( \15210 , \15166 , \15209 );
xor \U$14527 ( \15211 , \15092 , \15094 );
xor \U$14528 ( \15212 , \15211 , \15141 );
and \U$14529 ( \15213 , \15210 , \15212 );
and \U$14530 ( \15214 , \15166 , \15209 );
or \U$14531 ( \15215 , \15213 , \15214 );
nand \U$14532 ( \15216 , \15164 , \15215 );
not \U$14533 ( \15217 , \15216 );
or \U$14534 ( \15218 , \15155 , \15217 );
or \U$14535 ( \15219 , \15065 , \15153 );
nand \U$14536 ( \15220 , \15218 , \15219 );
nor \U$14537 ( \15221 , \15063 , \15220 );
not \U$14538 ( \15222 , \14987 );
nand \U$14539 ( \15223 , \15222 , \15060 );
xor \U$14540 ( \15224 , \14461 , \14561 );
xor \U$14541 ( \15225 , \15224 , \14564 );
not \U$14542 ( \15226 , \14975 );
not \U$14543 ( \15227 , \15226 );
not \U$14544 ( \15228 , \14983 );
or \U$14545 ( \15229 , \15227 , \15228 );
not \U$14546 ( \15230 , \14975 );
not \U$14547 ( \15231 , \14982 );
or \U$14548 ( \15232 , \15230 , \15231 );
buf \U$14549 ( \15233 , \14972 );
nand \U$14550 ( \15234 , \15232 , \15233 );
nand \U$14551 ( \15235 , \15229 , \15234 );
nand \U$14552 ( \15236 , \15225 , \15235 );
nand \U$14553 ( \15237 , \15223 , \15236 );
or \U$14554 ( \15238 , \15221 , \15237 );
nor \U$14555 ( \15239 , \15225 , \15235 );
not \U$14556 ( \15240 , \15239 );
nand \U$14557 ( \15241 , \15238 , \15240 );
not \U$14558 ( \15242 , \15239 );
xor \U$14559 ( \15243 , \15166 , \15209 );
xor \U$14560 ( \15244 , \15243 , \15212 );
xor \U$14561 ( \15245 , \15116 , \15127 );
xor \U$14562 ( \15246 , \15245 , \15138 );
not \U$14563 ( \15247 , \12481 );
not \U$14564 ( \15248 , \13901 );
or \U$14565 ( \15249 , \15247 , \15248 );
nand \U$14566 ( \15250 , \12371 , \13902 );
nand \U$14567 ( \15251 , \15249 , \15250 );
not \U$14568 ( \15252 , \15251 );
not \U$14569 ( \15253 , \12375 );
or \U$14570 ( \15254 , \15252 , \15253 );
nand \U$14571 ( \15255 , \15133 , \12365 );
nand \U$14572 ( \15256 , \15254 , \15255 );
not \U$14573 ( \15257 , \15256 );
not \U$14574 ( \15258 , \15257 );
and \U$14575 ( \15259 , \14499 , \12198 );
not \U$14576 ( \15260 , \14499 );
and \U$14577 ( \15261 , \15260 , \12199 );
nor \U$14578 ( \15262 , \15259 , \15261 );
not \U$14579 ( \15263 , \15262 );
not \U$14580 ( \15264 , \12194 );
or \U$14581 ( \15265 , \15263 , \15264 );
nand \U$14582 ( \15266 , \15171 , \12197 );
nand \U$14583 ( \15267 , \15265 , \15266 );
not \U$14584 ( \15268 , \15267 );
not \U$14585 ( \15269 , \15268 );
or \U$14586 ( \15270 , \15258 , \15269 );
not \U$14587 ( \15271 , \13270 );
not \U$14588 ( \15272 , \15113 );
or \U$14589 ( \15273 , \15271 , \15272 );
not \U$14590 ( \15274 , \13048 );
not \U$14591 ( \15275 , \13502 );
or \U$14592 ( \15276 , \15274 , \15275 );
nand \U$14593 ( \15277 , \13501 , \13049 );
nand \U$14594 ( \15278 , \15276 , \15277 );
nand \U$14595 ( \15279 , \15278 , \13259 );
nand \U$14596 ( \15280 , \15273 , \15279 );
not \U$14597 ( \15281 , \13751 );
not \U$14598 ( \15282 , \12950 );
or \U$14599 ( \15283 , \15281 , \15282 );
nand \U$14600 ( \15284 , \13244 , \13750 );
nand \U$14601 ( \15285 , \15283 , \15284 );
not \U$14602 ( \15286 , \15285 );
not \U$14603 ( \15287 , \12980 );
or \U$14604 ( \15288 , \15286 , \15287 );
nand \U$14605 ( \15289 , \15100 , \13045 );
nand \U$14606 ( \15290 , \15288 , \15289 );
xor \U$14607 ( \15291 , \15280 , \15290 );
nor \U$14608 ( \15292 , \12836 , \14499 );
and \U$14609 ( \15293 , \15291 , \15292 );
and \U$14610 ( \15294 , \15280 , \15290 );
or \U$14611 ( \15295 , \15293 , \15294 );
nand \U$14612 ( \15296 , \15270 , \15295 );
nand \U$14613 ( \15297 , \15267 , \15256 );
nand \U$14614 ( \15298 , \15296 , \15297 );
xor \U$14615 ( \15299 , \15246 , \15298 );
xor \U$14616 ( \15300 , \15176 , \15203 );
xor \U$14617 ( \15301 , \15300 , \15206 );
and \U$14618 ( \15302 , \15299 , \15301 );
and \U$14619 ( \15303 , \15246 , \15298 );
or \U$14620 ( \15304 , \15302 , \15303 );
nor \U$14621 ( \15305 , \15244 , \15304 );
not \U$14622 ( \15306 , \15305 );
not \U$14623 ( \15307 , \13942 );
not \U$14624 ( \15308 , \12686 );
or \U$14625 ( \15309 , \15307 , \15308 );
nand \U$14626 ( \15310 , \12956 , \13941 );
nand \U$14627 ( \15311 , \15309 , \15310 );
not \U$14628 ( \15312 , \15311 );
not \U$14629 ( \15313 , \12681 );
or \U$14630 ( \15314 , \15312 , \15313 );
nand \U$14631 ( \15315 , \15190 , \12667 );
nand \U$14632 ( \15316 , \15314 , \15315 );
not \U$14633 ( \15317 , \12685 );
not \U$14634 ( \15318 , \12369 );
or \U$14635 ( \15319 , \15317 , \15318 );
nand \U$14636 ( \15320 , \15319 , \14272 );
not \U$14637 ( \15321 , \12685 );
nand \U$14638 ( \15322 , \15321 , \12372 );
and \U$14639 ( \15323 , \15320 , \12189 , \15322 );
not \U$14640 ( \15324 , \13259 );
and \U$14641 ( \15325 , \13791 , \13261 );
not \U$14642 ( \15326 , \13791 );
and \U$14643 ( \15327 , \15326 , \13520 );
or \U$14644 ( \15328 , \15325 , \15327 );
not \U$14645 ( \15329 , \15328 );
or \U$14646 ( \15330 , \15324 , \15329 );
nand \U$14647 ( \15331 , \15278 , \13270 );
nand \U$14648 ( \15332 , \15330 , \15331 );
nand \U$14649 ( \15333 , \15323 , \15332 );
xor \U$14650 ( \15334 , \15316 , \15333 );
not \U$14651 ( \15335 , \14168 );
not \U$14652 ( \15336 , \12481 );
or \U$14653 ( \15337 , \15335 , \15336 );
nand \U$14654 ( \15338 , \13544 , \14342 );
nand \U$14655 ( \15339 , \15337 , \15338 );
not \U$14656 ( \15340 , \15339 );
not \U$14657 ( \15341 , \12375 );
or \U$14658 ( \15342 , \15340 , \15341 );
nand \U$14659 ( \15343 , \15251 , \12365 );
nand \U$14660 ( \15344 , \15342 , \15343 );
xor \U$14661 ( \15345 , \15334 , \15344 );
not \U$14662 ( \15346 , \15345 );
not \U$14663 ( \15347 , \15346 );
xor \U$14664 ( \15348 , \15280 , \15290 );
xor \U$14665 ( \15349 , \15348 , \15292 );
not \U$14666 ( \15350 , \15349 );
or \U$14667 ( \15351 , \15347 , \15350 );
not \U$14668 ( \15352 , \15349 );
not \U$14669 ( \15353 , \15352 );
not \U$14670 ( \15354 , \15345 );
or \U$14671 ( \15355 , \15353 , \15354 );
not \U$14672 ( \15356 , \12980 );
not \U$14673 ( \15357 , \13989 );
not \U$14674 ( \15358 , \12950 );
or \U$14675 ( \15359 , \15357 , \15358 );
nand \U$14676 ( \15360 , \13993 , \12662 );
nand \U$14677 ( \15361 , \15359 , \15360 );
not \U$14678 ( \15362 , \15361 );
or \U$14679 ( \15363 , \15356 , \15362 );
nand \U$14680 ( \15364 , \15285 , \14182 );
nand \U$14681 ( \15365 , \15363 , \15364 );
not \U$14682 ( \15366 , \15365 );
not \U$14683 ( \15367 , \15332 );
and \U$14684 ( \15368 , \15323 , \15367 );
not \U$14685 ( \15369 , \15323 );
and \U$14686 ( \15370 , \15369 , \15332 );
nor \U$14687 ( \15371 , \15368 , \15370 );
nand \U$14688 ( \15372 , \15366 , \15371 );
not \U$14689 ( \15373 , \12686 );
not \U$14690 ( \15374 , \15373 );
not \U$14691 ( \15375 , \13902 );
or \U$14692 ( \15376 , \15374 , \15375 );
not \U$14693 ( \15377 , \12846 );
nand \U$14694 ( \15378 , \15377 , \13901 );
nand \U$14695 ( \15379 , \15376 , \15378 );
not \U$14696 ( \15380 , \15379 );
not \U$14697 ( \15381 , \15123 );
or \U$14698 ( \15382 , \15380 , \15381 );
nand \U$14699 ( \15383 , \15311 , \12667 );
nand \U$14700 ( \15384 , \15382 , \15383 );
and \U$14701 ( \15385 , \15372 , \15384 );
nor \U$14702 ( \15386 , \15371 , \15366 );
nor \U$14703 ( \15387 , \15385 , \15386 );
not \U$14704 ( \15388 , \15387 );
nand \U$14705 ( \15389 , \15355 , \15388 );
nand \U$14706 ( \15390 , \15351 , \15389 );
not \U$14707 ( \15391 , \15316 );
nand \U$14708 ( \15392 , \15391 , \15333 );
not \U$14709 ( \15393 , \15392 );
not \U$14710 ( \15394 , \15344 );
or \U$14711 ( \15395 , \15393 , \15394 );
or \U$14712 ( \15396 , \15333 , \15391 );
nand \U$14713 ( \15397 , \15395 , \15396 );
not \U$14714 ( \15398 , \15397 );
not \U$14715 ( \15399 , \15195 );
not \U$14716 ( \15400 , \15201 );
or \U$14717 ( \15401 , \15399 , \15400 );
nand \U$14718 ( \15402 , \15194 , \15183 );
nand \U$14719 ( \15403 , \15401 , \15402 );
not \U$14720 ( \15404 , \15198 );
and \U$14721 ( \15405 , \15403 , \15404 );
not \U$14722 ( \15406 , \15403 );
and \U$14723 ( \15407 , \15406 , \15198 );
nor \U$14724 ( \15408 , \15405 , \15407 );
not \U$14725 ( \15409 , \15408 );
or \U$14726 ( \15410 , \15398 , \15409 );
or \U$14727 ( \15411 , \15397 , \15408 );
nand \U$14728 ( \15412 , \15410 , \15411 );
not \U$14729 ( \15413 , \15412 );
not \U$14730 ( \15414 , \15295 );
not \U$14731 ( \15415 , \15257 );
or \U$14732 ( \15416 , \15414 , \15415 );
or \U$14733 ( \15417 , \15257 , \15295 );
nand \U$14734 ( \15418 , \15416 , \15417 );
xor \U$14735 ( \15419 , \15418 , \15268 );
not \U$14736 ( \15420 , \15419 );
or \U$14737 ( \15421 , \15413 , \15420 );
or \U$14738 ( \15422 , \15419 , \15412 );
nand \U$14739 ( \15423 , \15421 , \15422 );
xor \U$14740 ( \15424 , \15390 , \15423 );
not \U$14741 ( \15425 , \14273 );
not \U$14742 ( \15426 , \12481 );
or \U$14743 ( \15427 , \15425 , \15426 );
nand \U$14744 ( \15428 , \13544 , \14499 );
nand \U$14745 ( \15429 , \15427 , \15428 );
not \U$14746 ( \15430 , \15429 );
not \U$14747 ( \15431 , \12375 );
or \U$14748 ( \15432 , \15430 , \15431 );
nand \U$14749 ( \15433 , \15339 , \13308 );
nand \U$14750 ( \15434 , \15432 , \15433 );
not \U$14751 ( \15435 , \15434 );
not \U$14752 ( \15436 , \14272 );
or \U$14753 ( \15437 , \12362 , \15436 );
not \U$14754 ( \15438 , \13259 );
not \U$14755 ( \15439 , \13520 );
not \U$14756 ( \15440 , \13750 );
or \U$14757 ( \15441 , \15439 , \15440 );
nand \U$14758 ( \15442 , \13749 , \13521 );
nand \U$14759 ( \15443 , \15441 , \15442 );
not \U$14760 ( \15444 , \15443 );
or \U$14761 ( \15445 , \15438 , \15444 );
nand \U$14762 ( \15446 , \15328 , \13270 );
nand \U$14763 ( \15447 , \15445 , \15446 );
not \U$14764 ( \15448 , \15447 );
nand \U$14765 ( \15449 , \15437 , \15448 );
not \U$14766 ( \15450 , \12980 );
not \U$14767 ( \15451 , \13241 );
not \U$14768 ( \15452 , \13942 );
or \U$14769 ( \15453 , \15451 , \15452 );
nand \U$14770 ( \15454 , \12951 , \13941 );
nand \U$14771 ( \15455 , \15453 , \15454 );
not \U$14772 ( \15456 , \15455 );
or \U$14773 ( \15457 , \15450 , \15456 );
nand \U$14774 ( \15458 , \15361 , \14182 );
nand \U$14775 ( \15459 , \15457 , \15458 );
and \U$14776 ( \15460 , \15449 , \15459 );
nor \U$14777 ( \15461 , \15437 , \15448 );
nor \U$14778 ( \15462 , \15460 , \15461 );
nand \U$14779 ( \15463 , \15435 , \15462 );
not \U$14780 ( \15464 , \15463 );
not \U$14781 ( \15465 , \15384 );
not \U$14782 ( \15466 , \15371 );
and \U$14783 ( \15467 , \15366 , \15466 );
not \U$14784 ( \15468 , \15366 );
and \U$14785 ( \15469 , \15468 , \15371 );
nor \U$14786 ( \15470 , \15467 , \15469 );
not \U$14787 ( \15471 , \15470 );
or \U$14788 ( \15472 , \15465 , \15471 );
or \U$14789 ( \15473 , \15470 , \15384 );
nand \U$14790 ( \15474 , \15472 , \15473 );
not \U$14791 ( \15475 , \15474 );
or \U$14792 ( \15476 , \15464 , \15475 );
not \U$14793 ( \15477 , \15462 );
nand \U$14794 ( \15478 , \15477 , \15434 );
nand \U$14795 ( \15479 , \15476 , \15478 );
not \U$14796 ( \15480 , \15479 );
and \U$14797 ( \15481 , \15387 , \15352 );
not \U$14798 ( \15482 , \15387 );
and \U$14799 ( \15483 , \15482 , \15349 );
nor \U$14800 ( \15484 , \15481 , \15483 );
and \U$14801 ( \15485 , \15484 , \15345 );
not \U$14802 ( \15486 , \15484 );
and \U$14803 ( \15487 , \15486 , \15346 );
nor \U$14804 ( \15488 , \15485 , \15487 );
nand \U$14805 ( \15489 , \15480 , \15488 );
not \U$14806 ( \15490 , \15489 );
nand \U$14807 ( \15491 , \12666 , \14273 );
not \U$14808 ( \15492 , \15491 );
not \U$14809 ( \15493 , \13259 );
not \U$14810 ( \15494 , \13264 );
not \U$14811 ( \15495 , \13940 );
not \U$14812 ( \15496 , \15495 );
or \U$14813 ( \15497 , \15494 , \15496 );
nand \U$14814 ( \15498 , \13940 , \13521 );
nand \U$14815 ( \15499 , \15497 , \15498 );
not \U$14816 ( \15500 , \15499 );
or \U$14817 ( \15501 , \15493 , \15500 );
and \U$14818 ( \15502 , \13988 , \13261 );
not \U$14819 ( \15503 , \13988 );
and \U$14820 ( \15504 , \15503 , \13520 );
or \U$14821 ( \15505 , \15502 , \15504 );
nand \U$14822 ( \15506 , \15505 , \13270 );
nand \U$14823 ( \15507 , \15501 , \15506 );
not \U$14824 ( \15508 , \15507 );
not \U$14825 ( \15509 , \15508 );
or \U$14826 ( \15510 , \15492 , \15509 );
and \U$14827 ( \15511 , \14167 , \12661 );
not \U$14828 ( \15512 , \14167 );
and \U$14829 ( \15513 , \15512 , \12951 );
or \U$14830 ( \15514 , \15511 , \15513 );
and \U$14831 ( \15515 , \12980 , \15514 );
and \U$14832 ( \15516 , \13900 , \13241 );
not \U$14833 ( \15517 , \13900 );
and \U$14834 ( \15518 , \15517 , \12662 );
or \U$14835 ( \15519 , \15516 , \15518 );
and \U$14836 ( \15520 , \15519 , \13251 );
nor \U$14837 ( \15521 , \15515 , \15520 );
not \U$14838 ( \15522 , \15521 );
nand \U$14839 ( \15523 , \15510 , \15522 );
not \U$14840 ( \15524 , \15491 );
nand \U$14841 ( \15525 , \15524 , \15507 );
nand \U$14842 ( \15526 , \15523 , \15525 );
not \U$14843 ( \15527 , \15526 );
and \U$14844 ( \15528 , \12980 , \15519 );
and \U$14845 ( \15529 , \15455 , \13045 );
nor \U$14846 ( \15530 , \15528 , \15529 );
not \U$14847 ( \15531 , \13270 );
not \U$14848 ( \15532 , \15443 );
or \U$14849 ( \15533 , \15531 , \15532 );
nand \U$14850 ( \15534 , \15505 , \13259 );
nand \U$14851 ( \15535 , \15533 , \15534 );
not \U$14852 ( \15536 , \15535 );
not \U$14853 ( \15537 , \13241 );
not \U$14854 ( \15538 , \12652 );
or \U$14855 ( \15539 , \15537 , \15538 );
nand \U$14856 ( \15540 , \15539 , \14272 );
nand \U$14857 ( \15541 , \12662 , \12671 );
nand \U$14858 ( \15542 , \12956 , \15540 , \15541 );
not \U$14859 ( \15543 , \15542 );
and \U$14860 ( \15544 , \15536 , \15543 );
and \U$14861 ( \15545 , \15542 , \15535 );
nor \U$14862 ( \15546 , \15544 , \15545 );
xor \U$14863 ( \15547 , \15530 , \15546 );
not \U$14864 ( \15548 , \12681 );
not \U$14865 ( \15549 , \14273 );
not \U$14866 ( \15550 , \13224 );
or \U$14867 ( \15551 , \15549 , \15550 );
nand \U$14868 ( \15552 , \12846 , \15436 );
nand \U$14869 ( \15553 , \15551 , \15552 );
not \U$14870 ( \15554 , \15553 );
or \U$14871 ( \15555 , \15548 , \15554 );
not \U$14872 ( \15556 , \14168 );
not \U$14873 ( \15557 , \13224 );
or \U$14874 ( \15558 , \15556 , \15557 );
not \U$14875 ( \15559 , \14167 );
nand \U$14876 ( \15560 , \15559 , \15373 );
nand \U$14877 ( \15561 , \15558 , \15560 );
nand \U$14878 ( \15562 , \15561 , \12667 );
nand \U$14879 ( \15563 , \15555 , \15562 );
not \U$14880 ( \15564 , \15563 );
xor \U$14881 ( \15565 , \15547 , \15564 );
nand \U$14882 ( \15566 , \15527 , \15565 );
not \U$14883 ( \15567 , \15566 );
not \U$14884 ( \15568 , \13270 );
or \U$14885 ( \15569 , \14531 , \13900 );
nand \U$14886 ( \15570 , \13900 , \13050 );
nand \U$14887 ( \15571 , \15569 , \15570 );
not \U$14888 ( \15572 , \15571 );
or \U$14889 ( \15573 , \15568 , \15572 );
and \U$14890 ( \15574 , \14167 , \13049 );
not \U$14891 ( \15575 , \14167 );
and \U$14892 ( \15576 , \15575 , \13269 );
or \U$14893 ( \15577 , \15574 , \15576 );
nand \U$14894 ( \15578 , \15577 , \13259 );
nand \U$14895 ( \15579 , \15573 , \15578 );
not \U$14896 ( \15580 , \15579 );
nor \U$14897 ( \15581 , \14499 , \12937 );
not \U$14898 ( \15582 , \15581 );
nand \U$14899 ( \15583 , \15580 , \15582 );
not \U$14900 ( \15584 , \14273 );
not \U$14901 ( \15585 , \13258 );
and \U$14902 ( \15586 , \15584 , \15585 );
and \U$14903 ( \15587 , \15577 , \13270 );
nor \U$14904 ( \15588 , \15586 , \15587 );
nand \U$14905 ( \15589 , \14273 , \13270 );
nand \U$14906 ( \15590 , \15589 , \13269 );
nor \U$14907 ( \15591 , \15588 , \15590 );
and \U$14908 ( \15592 , \15583 , \15591 );
and \U$14909 ( \15593 , \15581 , \15579 );
nor \U$14910 ( \15594 , \15592 , \15593 );
not \U$14911 ( \15595 , \13049 );
not \U$14912 ( \15596 , \12939 );
or \U$14913 ( \15597 , \15595 , \15596 );
nand \U$14914 ( \15598 , \15597 , \14272 );
nand \U$14915 ( \15599 , \12940 , \13048 );
and \U$14916 ( \15600 , \13244 , \15598 , \15599 );
not \U$14917 ( \15601 , \13270 );
not \U$14918 ( \15602 , \15499 );
or \U$14919 ( \15603 , \15601 , \15602 );
nand \U$14920 ( \15604 , \15571 , \13259 );
nand \U$14921 ( \15605 , \15603 , \15604 );
xor \U$14922 ( \15606 , \15600 , \15605 );
and \U$14923 ( \15607 , \15436 , \12950 );
not \U$14924 ( \15608 , \15436 );
and \U$14925 ( \15609 , \15608 , \12951 );
nor \U$14926 ( \15610 , \15607 , \15609 );
not \U$14927 ( \15611 , \15610 );
not \U$14928 ( \15612 , \12980 );
or \U$14929 ( \15613 , \15611 , \15612 );
nand \U$14930 ( \15614 , \15514 , \14182 );
nand \U$14931 ( \15615 , \15613 , \15614 );
nor \U$14932 ( \15616 , \15606 , \15615 );
or \U$14933 ( \15617 , \15594 , \15616 );
nand \U$14934 ( \15618 , \15606 , \15615 );
nand \U$14935 ( \15619 , \15617 , \15618 );
not \U$14936 ( \15620 , \15619 );
and \U$14937 ( \15621 , \15600 , \15605 );
not \U$14938 ( \15622 , \15621 );
not \U$14939 ( \15623 , \15491 );
not \U$14940 ( \15624 , \15507 );
or \U$14941 ( \15625 , \15623 , \15624 );
or \U$14942 ( \15626 , \15491 , \15507 );
nand \U$14943 ( \15627 , \15625 , \15626 );
not \U$14944 ( \15628 , \15627 );
not \U$14945 ( \15629 , \15521 );
and \U$14946 ( \15630 , \15628 , \15629 );
and \U$14947 ( \15631 , \15627 , \15521 );
nor \U$14948 ( \15632 , \15630 , \15631 );
nand \U$14949 ( \15633 , \15622 , \15632 );
not \U$14950 ( \15634 , \15633 );
or \U$14951 ( \15635 , \15620 , \15634 );
not \U$14952 ( \15636 , \15632 );
nand \U$14953 ( \15637 , \15636 , \15621 );
nand \U$14954 ( \15638 , \15635 , \15637 );
not \U$14955 ( \15639 , \15638 );
or \U$14956 ( \15640 , \15567 , \15639 );
not \U$14957 ( \15641 , \15565 );
nand \U$14958 ( \15642 , \15641 , \15526 );
nand \U$14959 ( \15643 , \15640 , \15642 );
not \U$14960 ( \15644 , \15643 );
not \U$14961 ( \15645 , \15561 );
not \U$14962 ( \15646 , \12681 );
or \U$14963 ( \15647 , \15645 , \15646 );
nand \U$14964 ( \15648 , \15379 , \12667 );
nand \U$14965 ( \15649 , \15647 , \15648 );
not \U$14966 ( \15650 , \15649 );
not \U$14967 ( \15651 , \15542 );
nand \U$14968 ( \15652 , \15651 , \15535 );
not \U$14969 ( \15653 , \15652 );
and \U$14970 ( \15654 , \15650 , \15653 );
and \U$14971 ( \15655 , \15649 , \15652 );
nor \U$14972 ( \15656 , \15654 , \15655 );
not \U$14973 ( \15657 , \15656 );
xor \U$14974 ( \15658 , \15447 , \15437 );
xnor \U$14975 ( \15659 , \15658 , \15459 );
not \U$14976 ( \15660 , \15659 );
and \U$14977 ( \15661 , \15657 , \15660 );
and \U$14978 ( \15662 , \15659 , \15656 );
nor \U$14979 ( \15663 , \15661 , \15662 );
xor \U$14980 ( \15664 , \15530 , \15546 );
and \U$14981 ( \15665 , \15664 , \15564 );
and \U$14982 ( \15666 , \15530 , \15546 );
or \U$14983 ( \15667 , \15665 , \15666 );
nand \U$14984 ( \15668 , \15663 , \15667 );
not \U$14985 ( \15669 , \15668 );
or \U$14986 ( \15670 , \15644 , \15669 );
not \U$14987 ( \15671 , \15663 );
not \U$14988 ( \15672 , \15667 );
nand \U$14989 ( \15673 , \15671 , \15672 );
nand \U$14990 ( \15674 , \15670 , \15673 );
not \U$14991 ( \15675 , \15474 );
not \U$14992 ( \15676 , \15434 );
not \U$14993 ( \15677 , \15462 );
and \U$14994 ( \15678 , \15676 , \15677 );
and \U$14995 ( \15679 , \15434 , \15462 );
nor \U$14996 ( \15680 , \15678 , \15679 );
not \U$14997 ( \15681 , \15680 );
and \U$14998 ( \15682 , \15675 , \15681 );
and \U$14999 ( \15683 , \15474 , \15680 );
nor \U$15000 ( \15684 , \15682 , \15683 );
not \U$15001 ( \15685 , \15649 );
nand \U$15002 ( \15686 , \15685 , \15652 );
and \U$15003 ( \15687 , \15686 , \15659 );
nor \U$15004 ( \15688 , \15685 , \15652 );
nor \U$15005 ( \15689 , \15687 , \15688 );
nand \U$15006 ( \15690 , \15684 , \15689 );
nand \U$15007 ( \15691 , \15674 , \15690 );
not \U$15008 ( \15692 , \15684 );
not \U$15009 ( \15693 , \15689 );
nand \U$15010 ( \15694 , \15692 , \15693 );
nand \U$15011 ( \15695 , \15691 , \15694 );
not \U$15012 ( \15696 , \15695 );
or \U$15013 ( \15697 , \15490 , \15696 );
not \U$15014 ( \15698 , \15488 );
nand \U$15015 ( \15699 , \15698 , \15479 );
nand \U$15016 ( \15700 , \15697 , \15699 );
and \U$15017 ( \15701 , \15424 , \15700 );
and \U$15018 ( \15702 , \15390 , \15423 );
or \U$15019 ( \15703 , \15701 , \15702 );
xor \U$15020 ( \15704 , \15246 , \15298 );
xor \U$15021 ( \15705 , \15704 , \15301 );
not \U$15022 ( \15706 , \15397 );
nand \U$15023 ( \15707 , \15706 , \15408 );
not \U$15024 ( \15708 , \15707 );
not \U$15025 ( \15709 , \15419 );
not \U$15026 ( \15710 , \15709 );
or \U$15027 ( \15711 , \15708 , \15710 );
not \U$15028 ( \15712 , \15408 );
nand \U$15029 ( \15713 , \15712 , \15397 );
nand \U$15030 ( \15714 , \15711 , \15713 );
or \U$15031 ( \15715 , \15705 , \15714 );
nand \U$15032 ( \15716 , \15306 , \15703 , \15715 );
and \U$15033 ( \15717 , \15705 , \15714 );
nand \U$15034 ( \15718 , \15306 , \15717 );
nand \U$15035 ( \15719 , \15244 , \15304 );
nand \U$15036 ( \15720 , \15716 , \15718 , \15719 );
not \U$15037 ( \15721 , \15164 );
not \U$15038 ( \15722 , \15215 );
nand \U$15039 ( \15723 , \15721 , \15722 );
and \U$15040 ( \15724 , \15219 , \15723 );
nand \U$15041 ( \15725 , \15242 , \15720 , \15724 , \15062 );
nand \U$15042 ( \15726 , \15241 , \15725 );
not \U$15043 ( \15727 , \14459 );
not \U$15044 ( \15728 , \14567 );
nand \U$15045 ( \15729 , \15727 , \15728 );
nand \U$15046 ( \15730 , \14449 , \15729 );
nor \U$15047 ( \15731 , \15730 , \14779 );
nand \U$15048 ( \15732 , \15726 , \14928 , \15731 );
not \U$15049 ( \15733 , \14886 );
not \U$15050 ( \15734 , \14860 );
or \U$15051 ( \15735 , \15733 , \15734 );
nor \U$15052 ( \15736 , \14914 , \14918 );
nand \U$15053 ( \15737 , \15735 , \15736 );
nor \U$15054 ( \15738 , \14906 , \14911 );
nor \U$15055 ( \15739 , \14860 , \14886 );
nor \U$15056 ( \15740 , \15738 , \15739 );
nand \U$15057 ( \15741 , \15737 , \15740 );
buf \U$15058 ( \15742 , \14926 );
and \U$15059 ( \15743 , \14912 , \15742 );
nand \U$15060 ( \15744 , \15741 , \15743 );
nor \U$15061 ( \15745 , \14921 , \14925 );
not \U$15062 ( \15746 , \15745 );
nand \U$15063 ( \15747 , \14930 , \15732 , \15744 , \15746 );
not \U$15064 ( \15748 , \15747 );
or \U$15065 ( \15749 , \13655 , \15748 );
not \U$15066 ( \15750 , \12913 );
not \U$15067 ( \15751 , \15750 );
buf \U$15068 ( \15752 , \13649 );
not \U$15069 ( \15753 , \15752 );
and \U$15070 ( \15754 , \13444 , \13411 );
and \U$15071 ( \15755 , \13615 , \13613 );
or \U$15072 ( \15756 , \15754 , \15755 );
not \U$15073 ( \15757 , \13445 );
nand \U$15074 ( \15758 , \15756 , \15757 );
not \U$15075 ( \15759 , \13642 );
or \U$15076 ( \15760 , \15758 , \15759 );
or \U$15077 ( \15761 , \13635 , \13641 );
nand \U$15078 ( \15762 , \15760 , \15761 );
not \U$15079 ( \15763 , \15762 );
or \U$15080 ( \15764 , \15753 , \15763 );
or \U$15081 ( \15765 , \13644 , \13648 );
nand \U$15082 ( \15766 , \15764 , \15765 );
not \U$15083 ( \15767 , \15766 );
or \U$15084 ( \15768 , \15751 , \15767 );
not \U$15085 ( \15769 , \12900 );
not \U$15086 ( \15770 , \15769 );
not \U$15087 ( \15771 , \12866 );
not \U$15088 ( \15772 , \12868 );
nand \U$15089 ( \15773 , \15771 , \15772 );
buf \U$15090 ( \15774 , \12597 );
or \U$15091 ( \15775 , \15773 , \15774 );
nand \U$15092 ( \15776 , \12596 , \12551 );
nand \U$15093 ( \15777 , \15775 , \15776 );
not \U$15094 ( \15778 , \15777 );
or \U$15095 ( \15779 , \15770 , \15778 );
nand \U$15096 ( \15780 , \12874 , \12899 );
nand \U$15097 ( \15781 , \15779 , \15780 );
and \U$15098 ( \15782 , \15781 , \12912 );
nor \U$15099 ( \15783 , \12905 , \12911 );
nor \U$15100 ( \15784 , \15782 , \15783 );
nand \U$15101 ( \15785 , \15768 , \15784 );
not \U$15102 ( \15786 , \15785 );
nand \U$15103 ( \15787 , \15749 , \15786 );
not \U$15104 ( \15788 , \15787 );
or \U$15105 ( \15789 , \12135 , \15788 );
nand \U$15106 ( \15790 , \12131 , \12133 );
nand \U$15107 ( \15791 , \15789 , \15790 );
not \U$15108 ( \15792 , \15791 );
or \U$15109 ( \15793 , \12028 , \15792 );
or \U$15110 ( \15794 , \12027 , \15791 );
nand \U$15111 ( \15795 , \15793 , \15794 );
not \U$15112 ( \15796 , RI9921eb0_597);
nor \U$15113 ( \15797 , \15796 , RI9921d48_600);
not \U$15114 ( \15798 , RI9921e38_598);
nor \U$15115 ( \15799 , \15798 , RI9921dc0_599);
nand \U$15116 ( \15800 , \15797 , \15799 );
buf \U$15117 ( \15801 , \15800 );
not \U$15118 ( \15802 , \15801 );
nand \U$15119 ( \15803 , \15802 , RI8918a20_187);
nor \U$15120 ( \15804 , RI9921e38_598, RI9921dc0_599);
nor \U$15121 ( \15805 , RI9921eb0_597, RI9921d48_600);
and \U$15122 ( \15806 , \15804 , \15805 , \10840 );
not \U$15123 ( \15807 , \15806 );
not \U$15124 ( \15808 , \15807 );
nand \U$15125 ( \15809 , \15808 , RI994dc68_31);
nand \U$15126 ( \15810 , RI9921e38_598, RI9921dc0_599);
not \U$15127 ( \15811 , \15810 );
nand \U$15128 ( \15812 , \15811 , \15797 );
buf \U$15129 ( \15813 , \15812 );
not \U$15130 ( \15814 , \15813 );
nand \U$15131 ( \15815 , \15814 , RI9967528_213);
not \U$15132 ( \15816 , \10753 );
buf \U$15133 ( \15817 , \15816 );
and \U$15134 ( \15818 , \15817 , RI995e900_226);
nor \U$15135 ( \15819 , \15818 , \10912 );
nand \U$15136 ( \15820 , \15803 , \15809 , \15815 , \15819 );
not \U$15137 ( \15821 , \15804 );
not \U$15138 ( \15822 , \15821 );
nand \U$15139 ( \15823 , \15822 , \15797 );
not \U$15140 ( \15824 , \15823 );
nand \U$15141 ( \15825 , \15824 , RI8946470_135);
nand \U$15142 ( \15826 , \10779 , RI9921dc0_599);
not \U$15143 ( \15827 , \15826 );
nand \U$15144 ( \15828 , \15827 , \15797 );
not \U$15145 ( \15829 , \15828 );
nand \U$15146 ( \15830 , \15829 , RI8930c60_161);
nand \U$15147 ( \15831 , \10773 , \10742 );
not \U$15148 ( \15832 , \15831 );
nand \U$15149 ( \15833 , \15832 , \15799 );
not \U$15150 ( \15834 , \15833 );
nand \U$15151 ( \15835 , \15834 , RI9808930_83);
nand \U$15152 ( \15836 , RI9921eb0_597, RI9921d48_600);
not \U$15153 ( \15837 , \15836 );
nand \U$15154 ( \15838 , \15799 , \15837 );
not \U$15155 ( \15839 , \15838 );
nand \U$15156 ( \15840 , \15839 , RI890fa38_200);
nand \U$15157 ( \15841 , \15825 , \15830 , \15835 , \15840 );
nor \U$15158 ( \15842 , \15820 , \15841 );
not \U$15159 ( \15843 , \15826 );
not \U$15160 ( \15844 , RI9921d48_600);
nor \U$15161 ( \15845 , \15844 , RI9921eb0_597);
nand \U$15162 ( \15846 , \15843 , \15845 );
not \U$15163 ( \15847 , \15846 );
buf \U$15164 ( \15848 , \15847 );
nand \U$15165 ( \15849 , \15848 , RI98195c8_70);
nand \U$15166 ( \15850 , \15845 , \15799 );
not \U$15167 ( \15851 , \15850 );
nand \U$15168 ( \15852 , \15851 , RI9808318_96);
not \U$15169 ( \15853 , \15810 );
nand \U$15170 ( \15854 , \15853 , \15845 );
not \U$15171 ( \15855 , \15854 );
nand \U$15172 ( \15856 , \15855 , RI89ec4d8_122);
not \U$15173 ( \15857 , RI9921eb0_597);
not \U$15174 ( \15858 , RI9921d48_600);
nand \U$15175 ( \15859 , \15857 , \15858 , RI9921e38_598, RI9921dc0_599);
not \U$15176 ( \15860 , \15859 );
nand \U$15177 ( \15861 , \15860 , RI9776e18_109);
nand \U$15178 ( \15862 , \15849 , \15852 , \15856 , \15861 );
not \U$15179 ( \15863 , \15826 );
nand \U$15180 ( \15864 , \15863 , \15805 );
not \U$15181 ( \15865 , \15864 );
nand \U$15182 ( \15866 , \15865 , RI98abad0_57);
and \U$15183 ( \15867 , \15845 , \15804 );
buf \U$15184 ( \15868 , \15867 );
nand \U$15185 ( \15869 , \15868 , RI98bc768_44);
not \U$15186 ( \15870 , \15826 );
nand \U$15187 ( \15871 , \15870 , \15837 );
not \U$15188 ( \15872 , \15871 );
buf \U$15189 ( \15873 , \15872 );
nand \U$15190 ( \15874 , \15873 , RI8925248_174);
not \U$15191 ( \15875 , \15836 );
nand \U$15192 ( \15876 , \15875 , \15804 );
not \U$15193 ( \15877 , \15876 );
nand \U$15194 ( \15878 , \15877 , RI8939c48_148);
nand \U$15195 ( \15879 , \15866 , \15869 , \15874 , \15878 );
nor \U$15196 ( \15880 , \15862 , \15879 );
nand \U$15197 ( \15881 , \15842 , \15880 );
not \U$15198 ( \15882 , \15881 );
nor \U$15199 ( \15883 , \10968 , \15882 );
not \U$15200 ( \15884 , \15883 );
buf \U$15201 ( \15885 , \11543 );
not \U$15202 ( \15886 , \15885 );
not \U$15203 ( \15887 , \15813 );
not \U$15204 ( \15888 , \10977 );
and \U$15205 ( \15889 , \15887 , \15888 );
and \U$15206 ( \15890 , RI8918a98_186, \15802 );
nor \U$15207 ( \15891 , \15889 , \15890 );
not \U$15208 ( \15892 , RI89464e8_134);
nor \U$15209 ( \15893 , \15892 , \15823 );
not \U$15210 ( \15894 , RI8930cd8_160);
nor \U$15211 ( \15895 , \15894 , \15828 );
nor \U$15212 ( \15896 , \15893 , \15895 );
and \U$15213 ( \15897 , \15834 , RI98089a8_82);
and \U$15214 ( \15898 , \15839 , RI890fab0_199);
nor \U$15215 ( \15899 , \15897 , \15898 );
and \U$15216 ( \15900 , \15808 , RI994dce0_30);
not \U$15217 ( \15901 , RI995e978_225);
not \U$15218 ( \15902 , \15817 );
or \U$15219 ( \15903 , \15901 , \15902 );
nand \U$15220 ( \15904 , \15903 , \10983 );
nor \U$15221 ( \15905 , \15900 , \15904 );
nand \U$15222 ( \15906 , \15891 , \15896 , \15899 , \15905 );
and \U$15223 ( \15907 , \15865 , RI98abb48_56);
and \U$15224 ( \15908 , \15868 , RI98bc7e0_43);
nor \U$15225 ( \15909 , \15907 , \15908 );
and \U$15226 ( \15910 , \15851 , RI9808390_95);
and \U$15227 ( \15911 , \15848 , RI9819640_69);
nor \U$15228 ( \15912 , \15910 , \15911 );
and \U$15229 ( \15913 , \15860 , RI9776e90_108);
and \U$15230 ( \15914 , \15855 , RI89ec550_121);
nor \U$15231 ( \15915 , \15913 , \15914 );
and \U$15232 ( \15916 , \15877 , RI8939cc0_147);
and \U$15233 ( \15917 , \15873 , RI89252c0_173);
nor \U$15234 ( \15918 , \15916 , \15917 );
nand \U$15235 ( \15919 , \15909 , \15912 , \15915 , \15918 );
nor \U$15236 ( \15920 , \15906 , \15919 );
and \U$15237 ( \15921 , \15886 , \15920 );
and \U$15238 ( \15922 , \15824 , RI8946560_133);
and \U$15239 ( \15923 , \15829 , RI8930d50_159);
nor \U$15240 ( \15924 , \15922 , \15923 );
and \U$15241 ( \15925 , \15802 , RI8918b10_185);
and \U$15242 ( \15926 , \15814 , RI9967618_211);
nor \U$15243 ( \15927 , \15925 , \15926 );
and \U$15244 ( \15928 , \15834 , RI9808a20_81);
and \U$15245 ( \15929 , \15839 , RI890fb28_198);
nor \U$15246 ( \15930 , \15928 , \15929 );
and \U$15247 ( \15931 , \15808 , RI994dd58_29);
not \U$15248 ( \15932 , RI99669e8_224);
not \U$15249 ( \15933 , \15817 );
or \U$15250 ( \15934 , \15932 , \15933 );
nand \U$15251 ( \15935 , \15934 , \11023 );
nor \U$15252 ( \15936 , \15931 , \15935 );
nand \U$15253 ( \15937 , \15924 , \15927 , \15930 , \15936 );
and \U$15254 ( \15938 , \15865 , RI98abbc0_55);
and \U$15255 ( \15939 , \15851 , RI9808408_94);
nor \U$15256 ( \15940 , \15938 , \15939 );
and \U$15257 ( \15941 , \15860 , RI9776f08_107);
and \U$15258 ( \15942 , \15855 , RI89ec5c8_120);
nor \U$15259 ( \15943 , \15941 , \15942 );
and \U$15260 ( \15944 , \15868 , RI98bc858_42);
and \U$15261 ( \15945 , \15873 , RI8925338_172);
nor \U$15262 ( \15946 , \15944 , \15945 );
and \U$15263 ( \15947 , \15877 , RI8939d38_146);
and \U$15264 ( \15948 , \15848 , RI98196b8_68);
nor \U$15265 ( \15949 , \15947 , \15948 );
nand \U$15266 ( \15950 , \15940 , \15943 , \15946 , \15949 );
nor \U$15267 ( \15951 , \15937 , \15950 );
not \U$15268 ( \15952 , \15951 );
not \U$15269 ( \15953 , \11549 );
not \U$15270 ( \15954 , \15953 );
or \U$15271 ( \15955 , \15952 , \15954 );
buf \U$15272 ( \15956 , \10894 );
and \U$15273 ( \15957 , \15865 , RI98abc38_54);
and \U$15274 ( \15958 , \15868 , RI98bc8d0_41);
nor \U$15275 ( \15959 , \15957 , \15958 );
and \U$15276 ( \15960 , \15860 , RI9776f80_106);
and \U$15277 ( \15961 , \15855 , RI89ec640_119);
nor \U$15278 ( \15962 , \15960 , \15961 );
and \U$15279 ( \15963 , \15851 , RI9808480_93);
and \U$15280 ( \15964 , \15873 , RI89253b0_171);
nor \U$15281 ( \15965 , \15963 , \15964 );
and \U$15282 ( \15966 , \15877 , RI8939db0_145);
and \U$15283 ( \15967 , \15848 , RI9819730_67);
nor \U$15284 ( \15968 , \15966 , \15967 );
nand \U$15285 ( \15969 , \15959 , \15962 , \15965 , \15968 );
and \U$15286 ( \15970 , \15824 , RI89465d8_132);
and \U$15287 ( \15971 , \15829 , RI8930dc8_158);
nor \U$15288 ( \15972 , \15970 , \15971 );
and \U$15289 ( \15973 , \15802 , RI8918b88_184);
and \U$15290 ( \15974 , \15814 , RI9967690_210);
nor \U$15291 ( \15975 , \15973 , \15974 );
and \U$15292 ( \15976 , \15834 , RI9808a98_80);
and \U$15293 ( \15977 , \15839 , RI890fba0_197);
nor \U$15294 ( \15978 , \15976 , \15977 );
and \U$15295 ( \15979 , \15808 , RI994ddd0_28);
and \U$15296 ( \15980 , \15817 , RI9967078_223);
nor \U$15297 ( \15981 , \15979 , \15980 , \10836 );
nand \U$15298 ( \15982 , \15972 , \15975 , \15978 , \15981 );
or \U$15299 ( \15983 , \15969 , \15982 );
not \U$15300 ( \15984 , \15983 );
nand \U$15301 ( \15985 , \15956 , \15984 );
nand \U$15302 ( \15986 , \15955 , \15985 );
nor \U$15303 ( \15987 , \15921 , \15986 );
not \U$15304 ( \15988 , \15987 );
or \U$15305 ( \15989 , \15884 , \15988 );
nor \U$15306 ( \15990 , \15986 , \15886 , \15920 );
not \U$15307 ( \15991 , \15951 );
nand \U$15308 ( \15992 , \15991 , \15985 , \11549 );
not \U$15309 ( \15993 , \11613 );
and \U$15310 ( \15994 , \15802 , RI8924e10_183);
and \U$15311 ( \15995 , \15814 , RI890f600_209);
nor \U$15312 ( \15996 , \15994 , \15995 );
and \U$15313 ( \15997 , \15824 , RI89ec0a0_131);
and \U$15314 ( \15998 , \15829 , RI8939810_157);
nor \U$15315 ( \15999 , \15997 , \15998 );
and \U$15316 ( \16000 , \15834 , RI9808b10_79);
and \U$15317 ( \16001 , \15839 , RI89185e8_196);
nor \U$15318 ( \16002 , \16000 , \16001 );
and \U$15319 ( \16003 , \15808 , RI994de48_27);
not \U$15320 ( \16004 , RI99670f0_222);
not \U$15321 ( \16005 , \15817 );
or \U$15322 ( \16006 , \16004 , \16005 );
nand \U$15323 ( \16007 , \16006 , \11579 );
nor \U$15324 ( \16008 , \16003 , \16007 );
nand \U$15325 ( \16009 , \15996 , \15999 , \16002 , \16008 );
and \U$15326 ( \16010 , \15865 , RI98abcb0_53);
and \U$15327 ( \16011 , \15868 , RI98bc948_40);
nor \U$15328 ( \16012 , \16010 , \16011 );
and \U$15329 ( \16013 , \15848 , RI98197a8_66);
and \U$15330 ( \16014 , \15873 , RI8930828_170);
nor \U$15331 ( \16015 , \16013 , \16014 );
and \U$15332 ( \16016 , \15860 , RI9776ff8_105);
and \U$15333 ( \16017 , \15855 , RI89ec6b8_118);
nor \U$15334 ( \16018 , \16016 , \16017 );
and \U$15335 ( \16019 , \15877 , RI8946038_144);
and \U$15336 ( \16020 , \15851 , RI98084f8_92);
nor \U$15337 ( \16021 , \16019 , \16020 );
nand \U$15338 ( \16022 , \16012 , \16015 , \16018 , \16021 );
nor \U$15339 ( \16023 , \16009 , \16022 );
not \U$15340 ( \16024 , \16023 );
and \U$15341 ( \16025 , \15993 , \16024 );
not \U$15342 ( \16026 , \15956 );
and \U$15343 ( \16027 , \16026 , \15983 );
nor \U$15344 ( \16028 , \16025 , \16027 );
nand \U$15345 ( \16029 , \15992 , \16028 );
nor \U$15346 ( \16030 , \15990 , \16029 );
nand \U$15347 ( \16031 , \15989 , \16030 );
nor \U$15348 ( \16032 , \11102 , RI99216b8_614);
and \U$15349 ( \16033 , \16032 , RI995ec48_11);
nand \U$15350 ( \16034 , \16033 , RI995ecc0_10);
nor \U$15351 ( \16035 , \16034 , \11304 );
nand \U$15352 ( \16036 , \16035 , RI995edb0_8);
not \U$15353 ( \16037 , \16036 );
nand \U$15354 ( \16038 , \16037 , RI995ee28_7);
nor \U$15355 ( \16039 , \16038 , \11448 );
not \U$15356 ( \16040 , \16039 );
nor \U$15357 ( \16041 , \16040 , \11614 );
xor \U$15358 ( \16042 , \16041 , RI995f0f8_1);
nor \U$15359 ( \16043 , \11621 , \16042 );
nor \U$15360 ( \16044 , \16031 , \16043 );
not \U$15361 ( \16045 , \16044 );
not \U$15362 ( \16046 , \15812 );
not \U$15363 ( \16047 , \11224 );
and \U$15364 ( \16048 , \16046 , \16047 );
and \U$15365 ( \16049 , \15806 , RI98bc9c0_39);
nor \U$15366 ( \16050 , \16048 , \16049 );
nor \U$15367 ( \16051 , \15828 , \11189 );
nor \U$15368 ( \16052 , \15800 , \11209 );
nor \U$15369 ( \16053 , \16051 , \16052 );
not \U$15370 ( \16054 , \15833 );
not \U$15371 ( \16055 , \11194 );
and \U$15372 ( \16056 , \16054 , \16055 );
nor \U$15373 ( \16057 , \15838 , \11206 );
nor \U$15374 ( \16058 , \16056 , \16057 );
and \U$15375 ( \16059 , \15824 , RI89460b0_143);
not \U$15376 ( \16060 , RI995e540_234);
not \U$15377 ( \16061 , \15816 );
or \U$15378 ( \16062 , \16060 , \16061 );
nand \U$15379 ( \16063 , \16062 , \11183 );
nor \U$15380 ( \16064 , \16059 , \16063 );
nand \U$15381 ( \16065 , \16050 , \16053 , \16058 , \16064 );
not \U$15382 ( \16066 , RI9777070_104);
nor \U$15383 ( \16067 , \16066 , \15850 );
nor \U$15384 ( \16068 , \15846 , \11199 );
nor \U$15385 ( \16069 , \16067 , \16068 );
not \U$15386 ( \16070 , \15864 );
not \U$15387 ( \16071 , RI98ab710_65);
not \U$15388 ( \16072 , \16071 );
and \U$15389 ( \16073 , \16070 , \16072 );
and \U$15390 ( \16074 , \15867 , RI98abd28_52);
nor \U$15391 ( \16075 , \16073 , \16074 );
and \U$15392 ( \16076 , \15872 , RI8924e88_182);
not \U$15393 ( \16077 , RI8939888_156);
nor \U$15394 ( \16078 , \16077 , \15876 );
nor \U$15395 ( \16079 , \16076 , \16078 );
and \U$15396 ( \16080 , \15860 , RI89ec730_117);
not \U$15397 ( \16081 , RI89ec118_130);
nor \U$15398 ( \16082 , \16081 , \15854 );
nor \U$15399 ( \16083 , \16080 , \16082 );
nand \U$15400 ( \16084 , \16069 , \16075 , \16079 , \16083 );
nor \U$15401 ( \16085 , \16065 , \16084 );
buf \U$15402 ( \16086 , \16085 );
not \U$15403 ( \16087 , \16086 );
not \U$15404 ( \16088 , \12920 );
or \U$15405 ( \16089 , \16087 , \16088 );
not \U$15406 ( \16090 , \15828 );
not \U$15407 ( \16091 , \11166 );
and \U$15408 ( \16092 , \16090 , \16091 );
and \U$15409 ( \16093 , \15806 , RI98bca38_38);
nor \U$15410 ( \16094 , \16092 , \16093 );
not \U$15411 ( \16095 , \15823 );
not \U$15412 ( \16096 , \11130 );
and \U$15413 ( \16097 , \16095 , \16096 );
not \U$15414 ( \16098 , RI99671e0_220);
nor \U$15415 ( \16099 , \16098 , \15812 );
nor \U$15416 ( \16100 , \16097 , \16099 );
not \U$15417 ( \16101 , \15833 );
not \U$15418 ( \16102 , \11154 );
and \U$15419 ( \16103 , \16101 , \16102 );
not \U$15420 ( \16104 , RI890f6f0_207);
nor \U$15421 ( \16105 , \16104 , \15838 );
nor \U$15422 ( \16106 , \16103 , \16105 );
not \U$15423 ( \16107 , \15800 );
not \U$15424 ( \16108 , RI89186d8_194);
not \U$15425 ( \16109 , \16108 );
and \U$15426 ( \16110 , \16107 , \16109 );
not \U$15427 ( \16111 , RI995e5b8_233);
not \U$15428 ( \16112 , \15816 );
or \U$15429 ( \16113 , \16111 , \16112 );
nand \U$15430 ( \16114 , \16113 , \11150 );
nor \U$15431 ( \16115 , \16110 , \16114 );
nand \U$15432 ( \16116 , \16094 , \16100 , \16106 , \16115 );
not \U$15433 ( \16117 , \15850 );
not \U$15434 ( \16118 , RI97770e8_103);
not \U$15435 ( \16119 , \16118 );
and \U$15436 ( \16120 , \16117 , \16119 );
and \U$15437 ( \16121 , \15877 , RI8939900_155);
nor \U$15438 ( \16122 , \16120 , \16121 );
not \U$15439 ( \16123 , \15864 );
not \U$15440 ( \16124 , \11170 );
and \U$15441 ( \16125 , \16123 , \16124 );
and \U$15442 ( \16126 , \15867 , RI98abda0_51);
nor \U$15443 ( \16127 , \16125 , \16126 );
not \U$15444 ( \16128 , \15871 );
not \U$15445 ( \16129 , \11163 );
and \U$15446 ( \16130 , \16128 , \16129 );
not \U$15447 ( \16131 , RI9819280_77);
nor \U$15448 ( \16132 , \16131 , \15846 );
nor \U$15449 ( \16133 , \16130 , \16132 );
not \U$15450 ( \16134 , RI89ec7a8_116);
nor \U$15451 ( \16135 , \16134 , \15859 );
not \U$15452 ( \16136 , RI89ec190_129);
nor \U$15453 ( \16137 , \16136 , \15854 );
nor \U$15454 ( \16138 , \16135 , \16137 );
nand \U$15455 ( \16139 , \16122 , \16127 , \16133 , \16138 );
nor \U$15456 ( \16140 , \16116 , \16139 );
not \U$15457 ( \16141 , \16140 );
nand \U$15458 ( \16142 , \16089 , \16141 );
not \U$15459 ( \16143 , \16086 );
nor \U$15460 ( \16144 , \16143 , \16141 );
not \U$15461 ( \16145 , \16144 );
not \U$15462 ( \16146 , \12920 );
or \U$15463 ( \16147 , \16145 , \16146 );
nand \U$15464 ( \16148 , \16147 , \12914 );
nand \U$15465 ( \16149 , \16142 , \16148 );
buf \U$15466 ( \16150 , \11246 );
or \U$15467 ( \16151 , \16149 , \16150 );
nand \U$15468 ( \16152 , \15806 , RI98bcab0_37);
not \U$15469 ( \16153 , \15800 );
nand \U$15470 ( \16154 , \16153 , RI8918750_193);
not \U$15471 ( \16155 , \15812 );
nand \U$15472 ( \16156 , \16155 , RI9967258_219);
and \U$15473 ( \16157 , \15816 , RI995e630_232);
nor \U$15474 ( \16158 , \16157 , \11085 );
nand \U$15475 ( \16159 , \16152 , \16154 , \16156 , \16158 );
nand \U$15476 ( \16160 , \15824 , RI89461a0_141);
nand \U$15477 ( \16161 , \15829 , RI8930990_167);
nand \U$15478 ( \16162 , \15834 , RI9808660_89);
nand \U$15479 ( \16163 , \15839 , RI890f768_206);
nand \U$15480 ( \16164 , \16160 , \16161 , \16162 , \16163 );
nor \U$15481 ( \16165 , \16159 , \16164 );
nand \U$15482 ( \16166 , \15847 , RI98192f8_76);
nand \U$15483 ( \16167 , RI9777160_102, \15851 );
nand \U$15484 ( \16168 , \15855 , RI89ec208_128);
nand \U$15485 ( \16169 , \15860 , RI89ec820_115);
nand \U$15486 ( \16170 , \16166 , \16167 , \16168 , \16169 );
not \U$15487 ( \16171 , \15864 );
nand \U$15488 ( \16172 , \16171 , RI98ab800_63);
nand \U$15489 ( \16173 , \15867 , RI98abe18_50);
nand \U$15490 ( \16174 , \15872 , RI8924f78_180);
nand \U$15491 ( \16175 , \15877 , RI8939978_154);
nand \U$15492 ( \16176 , \16172 , \16173 , \16174 , \16175 );
nor \U$15493 ( \16177 , \16170 , \16176 );
nand \U$15494 ( \16178 , \16165 , \16177 );
not \U$15495 ( \16179 , \16178 );
not \U$15496 ( \16180 , \16179 );
nand \U$15497 ( \16181 , \16151 , \16180 );
nand \U$15498 ( \16182 , \16149 , \16150 );
not \U$15499 ( \16183 , \15801 );
nand \U$15500 ( \16184 , \16183 , RI89187c8_192);
nand \U$15501 ( \16185 , \15806 , RI98bcb28_36);
not \U$15502 ( \16186 , \15813 );
nand \U$15503 ( \16187 , \16186 , RI99672d0_218);
and \U$15504 ( \16188 , \15817 , RI995e6a8_231);
nor \U$15505 ( \16189 , \16188 , \11471 );
nand \U$15506 ( \16190 , \16184 , \16185 , \16187 , \16189 );
nand \U$15507 ( \16191 , \15824 , RI8946218_140);
nand \U$15508 ( \16192 , \15829 , RI8930a08_166);
nand \U$15509 ( \16193 , \15834 , RI98086d8_88);
nand \U$15510 ( \16194 , \15839 , RI890f7e0_205);
nand \U$15511 ( \16195 , \16191 , \16192 , \16193 , \16194 );
nor \U$15512 ( \16196 , \16190 , \16195 );
nand \U$15513 ( \16197 , \15868 , RI98abe90_49);
nand \U$15514 ( \16198 , \15848 , RI9819370_75);
nand \U$15515 ( \16199 , \15873 , RI8924ff0_179);
nand \U$15516 ( \16200 , \15877 , RI89399f0_153);
nand \U$15517 ( \16201 , \16197 , \16198 , \16199 , \16200 );
nand \U$15518 ( \16202 , \15865 , RI98ab878_62);
nand \U$15519 ( \16203 , \15851 , RI97771d8_101);
nand \U$15520 ( \16204 , \15855 , RI89ec280_127);
nand \U$15521 ( \16205 , \15860 , RI89ec898_114);
nand \U$15522 ( \16206 , \16202 , \16203 , \16204 , \16205 );
nor \U$15523 ( \16207 , \16201 , \16206 );
nand \U$15524 ( \16208 , \16196 , \16207 );
not \U$15525 ( \16209 , \16208 );
nand \U$15526 ( \16210 , \16181 , \16182 , \16209 );
buf \U$15527 ( \16211 , \11504 );
and \U$15528 ( \16212 , \16210 , \16211 );
and \U$15529 ( \16213 , \16181 , \16182 );
nor \U$15530 ( \16214 , \16213 , \16209 );
nor \U$15531 ( \16215 , \16212 , \16214 );
nand \U$15532 ( \16216 , \15860 , RI89ec910_113);
nand \U$15533 ( \16217 , \15851 , RI9777250_100);
nand \U$15534 ( \16218 , \15855 , RI89ec2f8_126);
nand \U$15535 ( \16219 , \15873 , RI8925068_178);
nand \U$15536 ( \16220 , \16216 , \16217 , \16218 , \16219 );
nand \U$15537 ( \16221 , \15865 , RI98ab8f0_61);
nand \U$15538 ( \16222 , \15868 , RI98abf08_48);
nand \U$15539 ( \16223 , \15848 , RI98193e8_74);
nand \U$15540 ( \16224 , \15877 , RI8939a68_152);
nand \U$15541 ( \16225 , \16221 , \16222 , \16223 , \16224 );
nor \U$15542 ( \16226 , \16220 , \16225 );
nand \U$15543 ( \16227 , \15808 , RI98bcba0_35);
nand \U$15544 ( \16228 , \15802 , RI8918840_191);
nand \U$15545 ( \16229 , \15814 , RI9967348_217);
and \U$15546 ( \16230 , \15817 , RI995e720_230);
and \U$15547 ( \16231 , RI994d8a8_243, RI9921f28_596);
nor \U$15548 ( \16232 , \16230 , \16231 );
nand \U$15549 ( \16233 , \16227 , \16228 , \16229 , \16232 );
nand \U$15550 ( \16234 , \15824 , RI8946290_139);
nand \U$15551 ( \16235 , \15829 , RI8930a80_165);
nand \U$15552 ( \16236 , \15834 , RI9808750_87);
nand \U$15553 ( \16237 , \15839 , RI890f858_204);
nand \U$15554 ( \16238 , \16234 , \16235 , \16236 , \16237 );
nor \U$15555 ( \16239 , \16233 , \16238 );
nand \U$15556 ( \16240 , \16226 , \16239 );
not \U$15557 ( \16241 , \16240 );
not \U$15558 ( \16242 , \16241 );
buf \U$15559 ( \16243 , \11520 );
not \U$15560 ( \16244 , \16243 );
or \U$15561 ( \16245 , \16242 , \16244 );
buf \U$15562 ( \16246 , \11513 );
not \U$15563 ( \16247 , \16246 );
nand \U$15564 ( \16248 , \15814 , RI99673c0_216);
nand \U$15565 ( \16249 , \15802 , RI89188b8_190);
nand \U$15566 ( \16250 , \15808 , RI98bcc18_34);
and \U$15567 ( \16251 , \15817 , RI995e798_229);
not \U$15568 ( \16252 , \11317 );
nor \U$15569 ( \16253 , \16251 , \16252 );
nand \U$15570 ( \16254 , \16248 , \16249 , \16250 , \16253 );
nand \U$15571 ( \16255 , \15824 , RI8946308_138);
nand \U$15572 ( \16256 , \15829 , RI8930af8_164);
nand \U$15573 ( \16257 , \15834 , RI98087c8_86);
nand \U$15574 ( \16258 , \15839 , RI890f8d0_203);
nand \U$15575 ( \16259 , \16255 , \16256 , \16257 , \16258 );
nor \U$15576 ( \16260 , \16254 , \16259 );
nand \U$15577 ( \16261 , \15868 , RI98abf80_47);
nand \U$15578 ( \16262 , \15848 , RI9819460_73);
nand \U$15579 ( \16263 , \15873 , RI89250e0_177);
nand \U$15580 ( \16264 , \15877 , RI8939ae0_151);
nand \U$15581 ( \16265 , \16261 , \16262 , \16263 , \16264 );
nand \U$15582 ( \16266 , \15865 , RI98ab968_60);
nand \U$15583 ( \16267 , \15851 , RI97772c8_99);
nand \U$15584 ( \16268 , \15855 , RI89ec370_125);
nand \U$15585 ( \16269 , \15860 , RI89ec988_112);
nand \U$15586 ( \16270 , \16266 , \16267 , \16268 , \16269 );
nor \U$15587 ( \16271 , \16265 , \16270 );
nand \U$15588 ( \16272 , \16260 , \16271 );
or \U$15589 ( \16273 , \16247 , \16272 );
not \U$15590 ( \16274 , \11530 );
nand \U$15591 ( \16275 , \15808 , RI994dbf0_32);
nand \U$15592 ( \16276 , \16183 , RI89189a8_188);
nand \U$15593 ( \16277 , \16186 , RI99674b0_214);
and \U$15594 ( \16278 , \15817 , RI995e888_227);
not \U$15595 ( \16279 , \11414 );
nor \U$15596 ( \16280 , \16278 , \16279 );
nand \U$15597 ( \16281 , \16275 , \16276 , \16277 , \16280 );
nand \U$15598 ( \16282 , \15824 , RI89463f8_136);
nand \U$15599 ( \16283 , \15829 , RI8930be8_162);
nand \U$15600 ( \16284 , \15834 , RI98088b8_84);
nand \U$15601 ( \16285 , \15839 , RI890f9c0_201);
nand \U$15602 ( \16286 , \16282 , \16283 , \16284 , \16285 );
nor \U$15603 ( \16287 , \16281 , \16286 );
nand \U$15604 ( \16288 , \15865 , RI98aba58_58);
nand \U$15605 ( \16289 , \15851 , RI98082a0_97);
nand \U$15606 ( \16290 , \15860 , RI9776da0_110);
nand \U$15607 ( \16291 , \15855 , RI89ec460_123);
nand \U$15608 ( \16292 , \16288 , \16289 , \16290 , \16291 );
nand \U$15609 ( \16293 , \15868 , RI98bc6f0_45);
nand \U$15610 ( \16294 , \15847 , RI9819550_71);
nand \U$15611 ( \16295 , \15872 , RI89251d0_175);
nand \U$15612 ( \16296 , \15877 , RI8939bd0_149);
nand \U$15613 ( \16297 , \16293 , \16294 , \16295 , \16296 );
nor \U$15614 ( \16298 , \16292 , \16297 );
nand \U$15615 ( \16299 , \16287 , \16298 );
not \U$15616 ( \16300 , \16299 );
nand \U$15617 ( \16301 , \16274 , \16300 );
nand \U$15618 ( \16302 , \15808 , RI98bcc90_33);
nand \U$15619 ( \16303 , \16183 , RI8918930_189);
nand \U$15620 ( \16304 , \16186 , RI9967438_215);
and \U$15621 ( \16305 , \15817 , RI995e810_228);
not \U$15622 ( \16306 , \11356 );
nor \U$15623 ( \16307 , \16305 , \16306 );
nand \U$15624 ( \16308 , \16302 , \16303 , \16304 , \16307 );
nand \U$15625 ( \16309 , \15824 , RI8946380_137);
nand \U$15626 ( \16310 , \15829 , RI8930b70_163);
nand \U$15627 ( \16311 , \15834 , RI9808840_85);
nand \U$15628 ( \16312 , \15839 , RI890f948_202);
nand \U$15629 ( \16313 , \16309 , \16310 , \16311 , \16312 );
nor \U$15630 ( \16314 , \16308 , \16313 );
nand \U$15631 ( \16315 , \15851 , RI9808228_98);
nand \U$15632 ( \16316 , \15847 , RI98194d8_72);
nand \U$15633 ( \16317 , \15855 , RI89ec3e8_124);
nand \U$15634 ( \16318 , \15860 , RI9776d28_111);
nand \U$15635 ( \16319 , \16315 , \16316 , \16317 , \16318 );
nand \U$15636 ( \16320 , \15865 , RI98ab9e0_59);
nand \U$15637 ( \16321 , \15868 , RI98abff8_46);
nand \U$15638 ( \16322 , \15872 , RI8925158_176);
nand \U$15639 ( \16323 , \15877 , RI8939b58_150);
nand \U$15640 ( \16324 , \16320 , \16321 , \16322 , \16323 );
nor \U$15641 ( \16325 , \16319 , \16324 );
nand \U$15642 ( \16326 , \16314 , \16325 );
not \U$15643 ( \16327 , \16326 );
buf \U$15644 ( \16328 , \11527 );
not \U$15645 ( \16329 , \16328 );
nand \U$15646 ( \16330 , \16327 , \16329 );
nand \U$15647 ( \16331 , \16273 , \16301 , \16330 );
not \U$15648 ( \16332 , \16331 );
nand \U$15649 ( \16333 , \16245 , \16332 );
or \U$15650 ( \16334 , \16215 , \16333 );
nor \U$15651 ( \16335 , \16243 , \16241 );
and \U$15652 ( \16336 , \16332 , \16335 );
nand \U$15653 ( \16337 , \16301 , \16330 , \16247 , \16272 );
and \U$15654 ( \16338 , \16301 , \16328 , \16326 );
nor \U$15655 ( \16339 , \16274 , \16300 );
nor \U$15656 ( \16340 , \16338 , \16339 );
nand \U$15657 ( \16341 , \16337 , \16340 );
nor \U$15658 ( \16342 , \16336 , \16341 );
nand \U$15659 ( \16343 , \16334 , \16342 );
nand \U$15660 ( \16344 , \10968 , \15882 );
and \U$15661 ( \16345 , \15987 , \16344 );
nand \U$15662 ( \16346 , \16343 , \16345 );
not \U$15663 ( \16347 , \16346 );
or \U$15664 ( \16348 , \16045 , \16347 );
nand \U$15665 ( \16349 , \11613 , \16042 , \16023 );
nand \U$15666 ( \16350 , \16348 , \16349 );
not \U$15667 ( \16351 , \15885 );
not \U$15668 ( \16352 , RI995ef90_4);
nand \U$15669 ( \16353 , \16039 , RI995ef18_5);
not \U$15670 ( \16354 , \16353 );
or \U$15671 ( \16355 , \16352 , \16354 );
or \U$15672 ( \16356 , \16353 , RI995ef90_4);
nand \U$15673 ( \16357 , \16355 , \16356 );
not \U$15674 ( \16358 , \16357 );
and \U$15675 ( \16359 , \16351 , \16358 );
not \U$15676 ( \16360 , \16353 );
nand \U$15677 ( \16361 , \16360 , RI995ef90_4);
and \U$15678 ( \16362 , \16361 , RI995f008_3);
nor \U$15679 ( \16363 , \16361 , RI995f008_3);
nor \U$15680 ( \16364 , \16362 , \16363 );
not \U$15681 ( \16365 , \16364 );
not \U$15682 ( \16366 , \15953 );
or \U$15683 ( \16367 , \16365 , \16366 );
not \U$15684 ( \16368 , \16361 );
nand \U$15685 ( \16369 , \16368 , RI995f008_3);
and \U$15686 ( \16370 , \16369 , RI995f080_2);
nor \U$15687 ( \16371 , \16369 , RI995f080_2);
nor \U$15688 ( \16372 , \16370 , \16371 );
nand \U$15689 ( \16373 , \16372 , \15956 );
nand \U$15690 ( \16374 , \16367 , \16373 );
nor \U$15691 ( \16375 , \16359 , \16374 );
not \U$15692 ( \16376 , RI995ef18_5);
not \U$15693 ( \16377 , \16040 );
or \U$15694 ( \16378 , \16376 , \16377 );
or \U$15695 ( \16379 , \16040 , RI995ef18_5);
nand \U$15696 ( \16380 , \16378 , \16379 );
nand \U$15697 ( \16381 , \16375 , \16380 );
not \U$15698 ( \16382 , \16381 );
not \U$15699 ( \16383 , \10968 );
nand \U$15700 ( \16384 , \16383 , \16375 );
not \U$15701 ( \16385 , \16384 );
or \U$15702 ( \16386 , \16382 , \16385 );
and \U$15703 ( \16387 , \11102 , RI99216b8_614);
nor \U$15704 ( \16388 , \16387 , \16032 );
not \U$15705 ( \16389 , \16388 );
not \U$15706 ( \16390 , \12914 );
or \U$15707 ( \16391 , \16389 , \16390 );
nand \U$15708 ( \16392 , \16391 , \12922 );
not \U$15709 ( \16393 , \16150 );
not \U$15710 ( \16394 , RI995ec48_11);
not \U$15711 ( \16395 , \16032 );
not \U$15712 ( \16396 , \16395 );
or \U$15713 ( \16397 , \16394 , \16396 );
or \U$15714 ( \16398 , \16395 , RI995ec48_11);
nand \U$15715 ( \16399 , \16397 , \16398 );
not \U$15716 ( \16400 , \16399 );
and \U$15717 ( \16401 , \16393 , \16400 );
not \U$15718 ( \16402 , \12914 );
not \U$15719 ( \16403 , \16388 );
and \U$15720 ( \16404 , \16402 , \16403 );
nor \U$15721 ( \16405 , \16401 , \16404 );
not \U$15722 ( \16406 , \16211 );
not \U$15723 ( \16407 , \16033 );
not \U$15724 ( \16408 , \16407 );
not \U$15725 ( \16409 , RI995ecc0_10);
and \U$15726 ( \16410 , \16408 , \16409 );
and \U$15727 ( \16411 , \16407 , RI995ecc0_10);
nor \U$15728 ( \16412 , \16410 , \16411 );
nand \U$15729 ( \16413 , \16406 , \16412 );
nand \U$15730 ( \16414 , \16392 , \16405 , \16413 );
and \U$15731 ( \16415 , \16413 , \16150 , \16399 );
nor \U$15732 ( \16416 , \16406 , \16412 );
nor \U$15733 ( \16417 , \16415 , \16416 );
nand \U$15734 ( \16418 , \16414 , \16417 );
not \U$15735 ( \16419 , \16038 );
not \U$15736 ( \16420 , RI995eea0_6);
and \U$15737 ( \16421 , \16419 , \16420 );
and \U$15738 ( \16422 , \16038 , RI995eea0_6);
nor \U$15739 ( \16423 , \16421 , \16422 );
nand \U$15740 ( \16424 , \16274 , \16423 );
not \U$15741 ( \16425 , RI995ee28_7);
not \U$15742 ( \16426 , \16036 );
or \U$15743 ( \16427 , \16425 , \16426 );
or \U$15744 ( \16428 , \16036 , RI995ee28_7);
nand \U$15745 ( \16429 , \16427 , \16428 );
not \U$15746 ( \16430 , \16429 );
nand \U$15747 ( \16431 , \16430 , \16329 );
and \U$15748 ( \16432 , \16424 , \16431 );
not \U$15749 ( \16433 , RI995edb0_8);
not \U$15750 ( \16434 , \16035 );
not \U$15751 ( \16435 , \16434 );
or \U$15752 ( \16436 , \16433 , \16435 );
or \U$15753 ( \16437 , \16434 , RI995edb0_8);
nand \U$15754 ( \16438 , \16436 , \16437 );
not \U$15755 ( \16439 , \16438 );
nand \U$15756 ( \16440 , \16439 , \16246 );
and \U$15757 ( \16441 , \16432 , \16440 );
not \U$15758 ( \16442 , RI995ed38_9);
not \U$15759 ( \16443 , \16034 );
or \U$15760 ( \16444 , \16442 , \16443 );
or \U$15761 ( \16445 , \16034 , RI995ed38_9);
nand \U$15762 ( \16446 , \16444 , \16445 );
not \U$15763 ( \16447 , \16446 );
nand \U$15764 ( \16448 , \16447 , \16243 );
nand \U$15765 ( \16449 , \16418 , \16441 , \16448 );
not \U$15766 ( \16450 , \16243 );
nand \U$15767 ( \16451 , \16450 , \16441 , \16446 );
and \U$15768 ( \16452 , \16432 , \16247 , \16438 );
or \U$15769 ( \16453 , \16274 , \16423 );
nand \U$15770 ( \16454 , \16424 , \16328 , \16429 );
nand \U$15771 ( \16455 , \16453 , \16454 );
nor \U$15772 ( \16456 , \16452 , \16455 );
nand \U$15773 ( \16457 , \16449 , \16451 , \16456 );
nand \U$15774 ( \16458 , \16386 , \16457 );
not \U$15775 ( \16459 , \16384 );
nand \U$15776 ( \16460 , \16459 , \16380 );
not \U$15777 ( \16461 , \16374 );
and \U$15778 ( \16462 , \16461 , \15885 , \16357 );
or \U$15779 ( \16463 , \15956 , \16372 );
not \U$15780 ( \16464 , \16364 );
nand \U$15781 ( \16465 , \16464 , \16373 , \11549 );
nand \U$15782 ( \16466 , \16463 , \16465 );
nor \U$15783 ( \16467 , \16462 , \16466 );
nand \U$15784 ( \16468 , \16458 , \16460 , \16467 );
nand \U$15785 ( \16469 , \16350 , \16468 );
nand \U$15786 ( \16470 , \11621 , \16042 );
nor \U$15787 ( \16471 , \16031 , \16470 );
nand \U$15788 ( \16472 , \16346 , \16471 );
nand \U$15789 ( \16473 , \16469 , \16472 );
not \U$15790 ( \16474 , \16473 );
not \U$15791 ( \16475 , \16474 );
not \U$15792 ( \16476 , \16475 );
not \U$15793 ( \16477 , \16476 );
nand \U$15794 ( \16478 , \15795 , \16477 );
not \U$15795 ( \16479 , \16475 );
or \U$15796 ( \16480 , \11616 , \16023 );
not \U$15797 ( \16481 , \16480 );
nand \U$15798 ( \16482 , \10909 , \15983 );
not \U$15799 ( \16483 , \16482 );
not \U$15800 ( \16484 , \15951 );
nand \U$15801 ( \16485 , \16484 , \11050 );
not \U$15802 ( \16486 , \16485 );
not \U$15803 ( \16487 , \15920 );
nand \U$15804 ( \16488 , \16487 , \11012 );
not \U$15805 ( \16489 , \16488 );
nand \U$15806 ( \16490 , \10973 , \15881 );
nand \U$15807 ( \16491 , \16299 , \11450 );
nand \U$15808 ( \16492 , \16490 , \16491 );
nand \U$15809 ( \16493 , \16326 , \11399 );
nand \U$15810 ( \16494 , \16272 , \11351 );
nand \U$15811 ( \16495 , \16493 , \16494 );
nor \U$15812 ( \16496 , \16492 , \16495 );
not \U$15813 ( \16497 , \16496 );
nand \U$15814 ( \16498 , \16178 , \11106 );
not \U$15815 ( \16499 , \16498 );
nor \U$15816 ( \16500 , \16140 , \11102 );
nor \U$15817 ( \16501 , \16085 , RI994e4d8_13);
or \U$15818 ( \16502 , \16500 , \16501 );
nand \U$15819 ( \16503 , \16140 , \11102 );
nand \U$15820 ( \16504 , \16502 , \16503 );
not \U$15821 ( \16505 , \16504 );
or \U$15822 ( \16506 , \16499 , \16505 );
nand \U$15823 ( \16507 , \16179 , \11247 );
nand \U$15824 ( \16508 , \16506 , \16507 );
nand \U$15825 ( \16509 , \16208 , \11498 );
and \U$15826 ( \16510 , \16508 , \16509 );
nor \U$15827 ( \16511 , \16208 , \11498 );
nor \U$15828 ( \16512 , \16510 , \16511 );
nand \U$15829 ( \16513 , \16240 , \11308 );
not \U$15830 ( \16514 , \16513 );
nor \U$15831 ( \16515 , \16512 , \16514 );
not \U$15832 ( \16516 , \16515 );
or \U$15833 ( \16517 , \16497 , \16516 );
not \U$15834 ( \16518 , \16493 );
nor \U$15835 ( \16519 , \16518 , \16492 );
nor \U$15836 ( \16520 , \16240 , \11308 );
not \U$15837 ( \16521 , \16520 );
not \U$15838 ( \16522 , \16494 );
or \U$15839 ( \16523 , \16521 , \16522 );
or \U$15840 ( \16524 , \16272 , \11351 );
nand \U$15841 ( \16525 , \16523 , \16524 );
and \U$15842 ( \16526 , \16519 , \16525 );
nor \U$15843 ( \16527 , \16326 , \11399 );
and \U$15844 ( \16528 , \16527 , \16491 );
nor \U$15845 ( \16529 , \16299 , \11450 );
nor \U$15846 ( \16530 , \16528 , \16529 );
not \U$15847 ( \16531 , \16490 );
or \U$15848 ( \16532 , \16530 , \16531 );
nand \U$15849 ( \16533 , \11541 , \15882 );
nand \U$15850 ( \16534 , \16532 , \16533 );
nor \U$15851 ( \16535 , \16526 , \16534 );
nand \U$15852 ( \16536 , \16517 , \16535 );
not \U$15853 ( \16537 , \16536 );
or \U$15854 ( \16538 , \16489 , \16537 );
nand \U$15855 ( \16539 , \11013 , \15920 );
nand \U$15856 ( \16540 , \16538 , \16539 );
not \U$15857 ( \16541 , \16540 );
or \U$15858 ( \16542 , \16486 , \16541 );
nand \U$15859 ( \16543 , \11550 , \15951 );
nand \U$15860 ( \16544 , \16542 , \16543 );
not \U$15861 ( \16545 , \16544 );
or \U$15862 ( \16546 , \16483 , \16545 );
not \U$15863 ( \16547 , \10909 );
nand \U$15864 ( \16548 , \16547 , \15984 );
nand \U$15865 ( \16549 , \16546 , \16548 );
not \U$15866 ( \16550 , \16549 );
or \U$15867 ( \16551 , \16481 , \16550 );
nand \U$15868 ( \16552 , \11616 , \16023 );
nand \U$15869 ( \16553 , \16551 , \16552 );
nor \U$15870 ( \16554 , \16553 , \11625 );
not \U$15871 ( \16555 , \16554 );
nand \U$15872 ( \16556 , \16553 , \11625 );
nand \U$15873 ( \16557 , \16555 , \16556 );
not \U$15874 ( \16558 , \16557 );
nand \U$15875 ( \16559 , \16480 , \16552 );
nor \U$15876 ( \16560 , \16549 , \16559 );
not \U$15877 ( \16561 , \16560 );
nand \U$15878 ( \16562 , \16549 , \16559 );
nand \U$15879 ( \16563 , \16561 , \16562 );
not \U$15880 ( \16564 , \16563 );
nand \U$15881 ( \16565 , \16558 , \16564 );
nand \U$15882 ( \16566 , \16557 , \16563 );
nand \U$15883 ( \16567 , \16482 , \16548 );
xnor \U$15884 ( \16568 , \16544 , \16567 );
buf \U$15885 ( \16569 , \16568 );
not \U$15886 ( \16570 , \16569 );
xor \U$15887 ( \16571 , \16570 , \16563 );
and \U$15888 ( \16572 , \16565 , \16566 , \16571 );
not \U$15889 ( \16573 , \16572 );
not \U$15890 ( \16574 , \16558 );
not \U$15891 ( \16575 , RI9924b38_508);
nor \U$15892 ( \16576 , \16575 , \10823 );
nor \U$15893 ( \16577 , \11586 , \1566 );
nor \U$15894 ( \16578 , \16576 , \16577 );
nor \U$15895 ( \16579 , \11603 , \1552 );
not \U$15896 ( \16580 , RI992abc8_368);
buf \U$15897 ( \16581 , \10880 );
nor \U$15898 ( \16582 , \16580 , \16581 );
nor \U$15899 ( \16583 , \16579 , \16582 );
nand \U$15900 ( \16584 , \16578 , \16583 );
not \U$15901 ( \16585 , \10862 );
not \U$15902 ( \16586 , \1573 );
and \U$15903 ( \16587 , \16585 , \16586 );
and \U$15904 ( \16588 , \11576 , RI992c6f8_348);
nor \U$15905 ( \16589 , \16587 , \16588 );
not \U$15906 ( \16590 , \11032 );
not \U$15907 ( \16591 , \16590 );
not \U$15908 ( \16592 , \1589 );
and \U$15909 ( \16593 , \16591 , \16592 );
not \U$15910 ( \16594 , \10885 );
and \U$15911 ( \16595 , \16594 , RI992ef48_308);
nor \U$15912 ( \16596 , \16593 , \16595 );
nand \U$15913 ( \16597 , \16589 , \16596 );
nor \U$15914 ( \16598 , \16584 , \16597 );
not \U$15915 ( \16599 , RI9931b58_268);
or \U$15916 ( \16600 , \11607 , \16599 );
not \U$15917 ( \16601 , \15797 );
and \U$15918 ( \16602 , \11640 , \16601 );
nor \U$15919 ( \16603 , \16602 , \15810 );
nand \U$15920 ( \16604 , \11648 , \15836 );
and \U$15921 ( \16605 , \16603 , \16604 );
and \U$15922 ( \16606 , \16605 , RI9923878_548);
not \U$15923 ( \16607 , \15817 );
nor \U$15924 ( \16608 , \16607 , \11648 );
or \U$15925 ( \16609 , \16608 , RI9921f28_596);
and \U$15926 ( \16610 , \16609 , RI9922f18_568);
nor \U$15927 ( \16611 , \16606 , \16610 );
nand \U$15928 ( \16612 , \16600 , \16611 );
nor \U$15929 ( \16613 , \10794 , \1546 );
nor \U$15930 ( \16614 , \16612 , \16613 );
and \U$15931 ( \16615 , \11028 , RI9928af8_408);
and \U$15932 ( \16616 , \10931 , RI9928198_428);
nor \U$15933 ( \16617 , \16615 , \16616 );
and \U$15934 ( \16618 , \11030 , RI992f8a8_288);
not \U$15935 ( \16619 , \11568 );
and \U$15936 ( \16620 , \16619 , RI992a268_388);
nor \U$15937 ( \16621 , \16618 , \16620 );
and \U$15938 ( \16622 , \16614 , \16617 , \16621 , \11833 );
nand \U$15939 ( \16623 , \16598 , \16622 );
not \U$15940 ( \16624 , \16623 );
and \U$15941 ( \16625 , \16574 , \16624 );
not \U$15942 ( \16626 , \16574 );
and \U$15943 ( \16627 , \16626 , \16623 );
nor \U$15944 ( \16628 , \16625 , \16627 );
or \U$15945 ( \16629 , \16573 , \16628 );
not \U$15946 ( \16630 , \16571 );
not \U$15947 ( \16631 , \16630 );
or \U$15948 ( \16632 , \16631 , \16626 );
nand \U$15949 ( \16633 , \16629 , \16632 );
buf \U$15951 ( \16634 , \16554 );
not \U$15952 ( \16635 , \16634 );
nand \U$15953 ( \16636 , \16557 , \16635 );
nand \U$15954 ( \16637 , 1'b1 , \16636 );
not \U$15955 ( \16638 , \16637 );
not \U$15956 ( \16639 , \16638 );
not \U$15957 ( \16640 , \16639 );
not \U$15958 ( \16641 , \16640 );
buf \U$15959 ( \16642 , \16635 );
not \U$15960 ( \16643 , \10920 );
and \U$15961 ( \16644 , \16643 , RI9931ae0_269);
nor \U$15962 ( \16645 , \10794 , \1650 );
nor \U$15963 ( \16646 , \16644 , \16645 );
not \U$15964 ( \16647 , \16590 );
not \U$15965 ( \16648 , \1663 );
and \U$15966 ( \16649 , \16647 , \16648 );
and \U$15967 ( \16650 , \11028 , RI9928a80_409);
nor \U$15968 ( \16651 , \16649 , \16650 );
nand \U$15969 ( \16652 , \10931 , RI9928120_429);
nand \U$15970 ( \16653 , \16646 , \16651 , \16652 );
not \U$15971 ( \16654 , \11586 );
and \U$15972 ( \16655 , \16654 , RI9924160_529);
not \U$15973 ( \16656 , \10823 );
and \U$15974 ( \16657 , \16656 , RI9924ac0_509);
nor \U$15975 ( \16658 , \16655 , \16657 );
and \U$15976 ( \16659 , \11576 , RI992b4b0_349);
and \U$15977 ( \16660 , \16594 , RI992eed0_309);
nor \U$15978 ( \16661 , \16659 , \16660 );
nand \U$15979 ( \16662 , \16658 , \16661 );
nor \U$15980 ( \16663 , \16653 , \16662 );
and \U$15981 ( \16664 , \11574 , RI992ab50_369);
and \U$15982 ( \16665 , \10868 , RI9926410_469);
nor \U$15983 ( \16666 , \16664 , \16665 );
and \U$15984 ( \16667 , \11030 , RI992f830_289);
and \U$15985 ( \16668 , \11569 , RI992a1f0_389);
nor \U$15986 ( \16669 , \16667 , \16668 );
nand \U$15987 ( \16670 , \16666 , \16669 );
buf \U$15988 ( \16671 , \10955 );
and \U$15989 ( \16672 , \16671 , RI9925ab0_489);
not \U$15990 ( \16673 , RI9922bd0_569);
not \U$15991 ( \16674 , \16609 );
or \U$15992 ( \16675 , \16673 , \16674 );
not \U$15993 ( \16676 , \16605 );
or \U$15994 ( \16677 , \16676 , \1644 );
nand \U$15995 ( \16678 , \16675 , \16677 );
nor \U$15996 ( \16679 , \16672 , \16678 );
nand \U$15997 ( \16680 , \11752 , \16679 );
nor \U$15998 ( \16681 , \16670 , \16680 );
nand \U$15999 ( \16682 , \16663 , \16681 );
not \U$16000 ( \16683 , \16682 );
and \U$16001 ( \16684 , \16642 , \16683 );
not \U$16002 ( \16685 , \16642 );
not \U$16003 ( \16686 , \16683 );
and \U$16004 ( \16687 , \16685 , \16686 );
nor \U$16005 ( \16688 , \16684 , \16687 );
nand \U$16006 ( \16689 , \16641 , \16688 );
xor \U$16007 ( \16690 , \16633 , \16689 );
not \U$16008 ( \16691 , RI9931a68_270);
nor \U$16009 ( \16692 , \16691 , \11607 );
not \U$16010 ( \16693 , RI9926cf8_450);
nor \U$16011 ( \16694 , \16693 , \10794 );
nor \U$16012 ( \16695 , \16692 , \16694 );
not \U$16013 ( \16696 , RI9928a08_410);
nor \U$16014 ( \16697 , \16696 , \11563 );
not \U$16015 ( \16698 , \11582 );
nor \U$16016 ( \16699 , \16698 , \1687 );
nor \U$16017 ( \16700 , \16697 , \16699 );
nand \U$16018 ( \16701 , \10931 , RI99280a8_430);
nand \U$16019 ( \16702 , \16695 , \16700 , \16701 );
and \U$16020 ( \16703 , \16656 , RI9924a48_510);
not \U$16021 ( \16704 , RI99240e8_530);
nor \U$16022 ( \16705 , \16704 , \11586 );
nor \U$16023 ( \16706 , \16703 , \16705 );
and \U$16024 ( \16707 , \11576 , RI992b438_350);
and \U$16025 ( \16708 , \16594 , RI992ee58_310);
nor \U$16026 ( \16709 , \16707 , \16708 );
nand \U$16027 ( \16710 , \16706 , \16709 );
nor \U$16028 ( \16711 , \16702 , \16710 );
nor \U$16029 ( \16712 , \11573 , \1701 );
not \U$16030 ( \16713 , RI9926398_470);
nor \U$16031 ( \16714 , \16713 , \11603 );
nor \U$16032 ( \16715 , \16712 , \16714 );
and \U$16033 ( \16716 , \16619 , RI992a178_390);
not \U$16034 ( \16717 , RI992f7b8_290);
nor \U$16035 ( \16718 , \16717 , \11599 );
nor \U$16036 ( \16719 , \16716 , \16718 );
nand \U$16037 ( \16720 , \16715 , \16719 );
and \U$16038 ( \16721 , \16671 , RI9925a38_490);
not \U$16039 ( \16722 , RI9923788_550);
not \U$16040 ( \16723 , \16605 );
or \U$16041 ( \16724 , \16722 , \16723 );
nand \U$16042 ( \16725 , \16609 , RI9922b58_570);
nand \U$16043 ( \16726 , \16724 , \16725 );
nor \U$16044 ( \16727 , \16721 , \16726 );
nand \U$16045 ( \16728 , \11941 , \16727 );
nor \U$16046 ( \16729 , \16720 , \16728 );
nand \U$16047 ( \16730 , \16711 , \16729 );
buf \U$16048 ( \16731 , \16730 );
not \U$16049 ( \16732 , \16731 );
and \U$16050 ( \16733 , \16642 , \16732 );
and \U$16051 ( \16734 , \16685 , \16731 );
nor \U$16052 ( \16735 , \16733 , \16734 );
and \U$16053 ( \16736 , \16641 , \16735 );
nand \U$16054 ( \16737 , \16488 , \16539 );
not \U$16055 ( \16738 , \16737 );
not \U$16056 ( \16739 , \16536 );
or \U$16057 ( \16740 , \16738 , \16739 );
or \U$16058 ( \16741 , \16737 , \16536 );
nand \U$16059 ( \16742 , \16740 , \16741 );
nand \U$16060 ( \16743 , \16485 , \16543 );
xnor \U$16061 ( \16744 , \16540 , \16743 );
not \U$16062 ( \16745 , \16744 );
and \U$16063 ( \16746 , \16742 , \16745 );
not \U$16064 ( \16747 , \16742 );
and \U$16065 ( \16748 , \16747 , \16744 );
nor \U$16066 ( \16749 , \16746 , \16748 );
not \U$16067 ( \16750 , \16749 );
not \U$16068 ( \16751 , \16750 );
not \U$16069 ( \16752 , \16751 );
not \U$16070 ( \16753 , \16569 );
nand \U$16071 ( \16754 , \16753 , \16745 );
nand \U$16072 ( \16755 , \16569 , \16744 );
and \U$16073 ( \16756 , \16754 , \16755 , \16749 );
not \U$16074 ( \16757 , \16756 );
not \U$16075 ( \16758 , \16757 );
not \U$16076 ( \16759 , \16758 );
not \U$16077 ( \16760 , \16759 );
or \U$16078 ( \16761 , \16752 , \16760 );
nand \U$16079 ( \16762 , \16761 , \16569 );
xor \U$16080 ( \16763 , \16736 , \16762 );
and \U$16081 ( \16764 , \16574 , \16683 );
buf \U$16082 ( \16765 , \16557 );
buf \U$16083 ( \16766 , \16765 );
not \U$16084 ( \16767 , \16766 );
and \U$16085 ( \16768 , \16767 , \16686 );
nor \U$16086 ( \16769 , \16764 , \16768 );
or \U$16087 ( \16770 , \16573 , \16769 );
or \U$16088 ( \16771 , \16628 , \16631 );
nand \U$16089 ( \16772 , \16770 , \16771 );
and \U$16090 ( \16773 , \16763 , \16772 );
and \U$16091 ( \16774 , \16736 , \16762 );
or \U$16092 ( \16775 , \16773 , \16774 );
xor \U$16093 ( \16776 , \16690 , \16775 );
and \U$16094 ( \16777 , \16569 , \16624 );
and \U$16095 ( \16778 , \16570 , \16623 );
nor \U$16096 ( \16779 , \16777 , \16778 );
or \U$16097 ( \16780 , \16759 , \16779 );
or \U$16098 ( \16781 , \16751 , \16570 );
nand \U$16099 ( \16782 , \16780 , \16781 );
not \U$16100 ( \16783 , \16782 );
not \U$16101 ( \16784 , \10794 );
not \U$16102 ( \16785 , RI9926c80_451);
not \U$16103 ( \16786 , \16785 );
and \U$16104 ( \16787 , \16784 , \16786 );
and \U$16105 ( \16788 , \16643 , RI99319f0_271);
nor \U$16106 ( \16789 , \16787 , \16788 );
not \U$16107 ( \16790 , RI992cef0_331);
nor \U$16108 ( \16791 , \16790 , \16590 );
not \U$16109 ( \16792 , RI9928990_411);
nor \U$16110 ( \16793 , \16792 , \10812 );
nor \U$16111 ( \16794 , \16791 , \16793 );
nand \U$16112 ( \16795 , \10931 , RI9928030_431);
nand \U$16113 ( \16796 , \16789 , \16794 , \16795 );
and \U$16114 ( \16797 , \16656 , RI99249d0_511);
not \U$16115 ( \16798 , RI9924070_531);
nor \U$16116 ( \16799 , \16798 , \11586 );
nor \U$16117 ( \16800 , \16797 , \16799 );
buf \U$16118 ( \16801 , \10873 );
and \U$16119 ( \16802 , \16801 , RI992b3c0_351);
and \U$16120 ( \16803 , \16594 , RI992ede0_311);
nor \U$16121 ( \16804 , \16802 , \16803 );
nand \U$16122 ( \16805 , \16800 , \16804 );
nor \U$16123 ( \16806 , \16796 , \16805 );
and \U$16124 ( \16807 , \10868 , RI9926320_471);
not \U$16125 ( \16808 , RI992aa60_371);
nor \U$16126 ( \16809 , \16808 , \16581 );
nor \U$16127 ( \16810 , \16807 , \16809 );
and \U$16128 ( \16811 , \11030 , RI992f740_291);
and \U$16129 ( \16812 , \11569 , RI992a100_391);
nor \U$16130 ( \16813 , \16811 , \16812 );
nand \U$16131 ( \16814 , \16810 , \16813 );
and \U$16132 ( \16815 , \16671 , RI99259c0_491);
not \U$16133 ( \16816 , RI9923710_551);
not \U$16134 ( \16817 , \16605 );
or \U$16135 ( \16818 , \16816 , \16817 );
nand \U$16136 ( \16819 , \16609 , RI9922ae0_571);
nand \U$16137 ( \16820 , \16818 , \16819 );
nor \U$16138 ( \16821 , \16815 , \16820 );
nand \U$16139 ( \16822 , \12099 , \16821 );
nor \U$16140 ( \16823 , \16814 , \16822 );
nand \U$16141 ( \16824 , \16806 , \16823 );
not \U$16142 ( \16825 , \16824 );
and \U$16143 ( \16826 , \16642 , \16825 );
and \U$16144 ( \16827 , \16685 , \16824 );
nor \U$16145 ( \16828 , \16826 , \16827 );
and \U$16146 ( \16829 , \16641 , \16828 );
xor \U$16147 ( \16830 , \16783 , \16829 );
or \U$16148 ( \16831 , \16767 , \16731 );
or \U$16149 ( \16832 , \16574 , \16732 );
nand \U$16150 ( \16833 , \16831 , \16832 );
not \U$16151 ( \16834 , \16833 );
or \U$16152 ( \16835 , \16573 , \16834 );
or \U$16153 ( \16836 , \16769 , \16631 );
nand \U$16154 ( \16837 , \16835 , \16836 );
and \U$16155 ( \16838 , \16830 , \16837 );
and \U$16156 ( \16839 , \16783 , \16829 );
or \U$16157 ( \16840 , \16838 , \16839 );
xor \U$16158 ( \16841 , \16782 , \16840 );
xor \U$16159 ( \16842 , \16736 , \16762 );
xor \U$16160 ( \16843 , \16842 , \16772 );
and \U$16161 ( \16844 , \16841 , \16843 );
and \U$16162 ( \16845 , \16782 , \16840 );
or \U$16163 ( \16846 , \16844 , \16845 );
xor \U$16164 ( \16847 , \16776 , \16846 );
not \U$16165 ( \16848 , RI9929098_396);
nor \U$16166 ( \16849 , \16848 , \11568 );
nor \U$16167 ( \16850 , \11599 , \2179 );
nor \U$16168 ( \16851 , \16849 , \16850 );
and \U$16169 ( \16852 , \11604 , RI99260c8_476);
nor \U$16170 ( \16853 , \16581 , \2163 );
nor \U$16171 ( \16854 , \16852 , \16853 );
and \U$16172 ( \16855 , \16671 , RI9925768_496);
not \U$16173 ( \16856 , RI99234b8_556);
not \U$16174 ( \16857 , \16605 );
or \U$16175 ( \16858 , \16856 , \16857 );
nand \U$16176 ( \16859 , \16609 , RI9922888_576);
nand \U$16177 ( \16860 , \16858 , \16859 );
nor \U$16178 ( \16861 , \16855 , \16860 );
nand \U$16179 ( \16862 , \16851 , \16854 , \12811 , \16861 );
not \U$16180 ( \16863 , \16862 );
not \U$16181 ( \16864 , RI9931798_276);
nor \U$16182 ( \16865 , \16864 , \11607 );
not \U$16183 ( \16866 , RI9926a28_456);
nor \U$16184 ( \16867 , \16866 , \10794 );
nor \U$16185 ( \16868 , \16865 , \16867 );
not \U$16186 ( \16869 , RI9928738_416);
nor \U$16187 ( \16870 , \16869 , \10812 );
not \U$16188 ( \16871 , RI992cc98_336);
nor \U$16189 ( \16872 , \16871 , \16590 );
nor \U$16190 ( \16873 , \16870 , \16872 );
nand \U$16191 ( \16874 , \10931 , RI9927dd8_436);
nand \U$16192 ( \16875 , \16868 , \16873 , \16874 );
not \U$16193 ( \16876 , RI992b168_356);
nor \U$16194 ( \16877 , \16876 , \10874 );
not \U$16195 ( \16878 , RI992d5f8_316);
nor \U$16196 ( \16879 , \16878 , \10885 );
nor \U$16197 ( \16880 , \16877 , \16879 );
not \U$16198 ( \16881 , \11586 );
not \U$16199 ( \16882 , \2161 );
and \U$16200 ( \16883 , \16881 , \16882 );
and \U$16201 ( \16884 , \16656 , RI9924778_516);
nor \U$16202 ( \16885 , \16883 , \16884 );
nand \U$16203 ( \16886 , \16880 , \16885 );
nor \U$16204 ( \16887 , \16875 , \16886 );
nand \U$16205 ( \16888 , \16863 , \16887 );
not \U$16206 ( \16889 , \16742 );
not \U$16207 ( \16890 , \16889 );
and \U$16208 ( \16891 , \16888 , \16890 );
not \U$16209 ( \16892 , \16888 );
buf \U$16210 ( \16893 , \16742 );
not \U$16211 ( \16894 , \16893 );
and \U$16212 ( \16895 , \16892 , \16894 );
nor \U$16213 ( \16896 , \16891 , \16895 );
not \U$16214 ( \16897 , \16896 );
not \U$16215 ( \16898 , \16529 );
nand \U$16216 ( \16899 , \16898 , \16491 );
not \U$16217 ( \16900 , \16899 );
not \U$16218 ( \16901 , \16493 );
not \U$16219 ( \16902 , \16494 );
not \U$16220 ( \16903 , \16513 );
not \U$16221 ( \16904 , \16512 );
not \U$16222 ( \16905 , \16904 );
or \U$16223 ( \16906 , \16903 , \16905 );
not \U$16224 ( \16907 , \16520 );
nand \U$16225 ( \16908 , \16906 , \16907 );
not \U$16226 ( \16909 , \16908 );
or \U$16227 ( \16910 , \16902 , \16909 );
nand \U$16228 ( \16911 , \16910 , \16524 );
not \U$16229 ( \16912 , \16911 );
or \U$16230 ( \16913 , \16901 , \16912 );
not \U$16231 ( \16914 , \16527 );
nand \U$16232 ( \16915 , \16913 , \16914 );
not \U$16233 ( \16916 , \16915 );
or \U$16234 ( \16917 , \16900 , \16916 );
not \U$16235 ( \16918 , \16915 );
not \U$16236 ( \16919 , \16899 );
nand \U$16237 ( \16920 , \16918 , \16919 );
nand \U$16238 ( \16921 , \16917 , \16920 );
buf \U$16239 ( \16922 , \16921 );
not \U$16240 ( \16923 , \16922 );
nand \U$16241 ( \16924 , \16490 , \16533 );
not \U$16242 ( \16925 , \16924 );
not \U$16243 ( \16926 , \16491 );
not \U$16244 ( \16927 , \16915 );
or \U$16245 ( \16928 , \16926 , \16927 );
nand \U$16246 ( \16929 , \16928 , \16898 );
not \U$16247 ( \16930 , \16929 );
or \U$16248 ( \16931 , \16925 , \16930 );
or \U$16249 ( \16932 , \16929 , \16924 );
nand \U$16250 ( \16933 , \16931 , \16932 );
nand \U$16251 ( \16934 , \16923 , \16933 );
not \U$16252 ( \16935 , \16934 );
not \U$16253 ( \16936 , \16922 );
not \U$16254 ( \16937 , \16742 );
or \U$16255 ( \16938 , \16936 , \16937 );
or \U$16256 ( \16939 , \16933 , \16893 );
nand \U$16257 ( \16940 , \16938 , \16939 );
nor \U$16258 ( \16941 , \16935 , \16940 );
not \U$16259 ( \16942 , \16941 );
or \U$16260 ( \16943 , \16897 , \16942 );
buf \U$16261 ( \16944 , \16922 );
not \U$16262 ( \16945 , \16944 );
not \U$16263 ( \16946 , \16933 );
not \U$16264 ( \16947 , \16946 );
or \U$16265 ( \16948 , \16945 , \16947 );
nand \U$16266 ( \16949 , \16948 , \16934 );
nor \U$16267 ( \16950 , \10812 , \2250 );
not \U$16268 ( \16951 , RI9927e50_435);
nor \U$16269 ( \16952 , \16951 , \10788 );
nor \U$16270 ( \16953 , \16950 , \16952 );
and \U$16271 ( \16954 , \10921 , RI9931810_275);
and \U$16272 ( \16955 , RI9922900_575, \16609 );
and \U$16273 ( \16956 , \16605 , RI9923530_555);
nor \U$16274 ( \16957 , \16954 , \16955 , \16956 );
buf \U$16275 ( \16958 , \10936 );
nand \U$16276 ( \16959 , \16958 , RI9926aa0_455);
nand \U$16277 ( \16960 , \16953 , \16957 , \16959 );
not \U$16278 ( \16961 , \11599 );
not \U$16279 ( \16962 , \2244 );
and \U$16280 ( \16963 , \16961 , \16962 );
and \U$16281 ( \16964 , \16619 , RI9929110_395);
nor \U$16282 ( \16965 , \16963 , \16964 );
nand \U$16283 ( \16966 , \16965 , \12620 );
nor \U$16284 ( \16967 , \16960 , \16966 );
not \U$16285 ( \16968 , RI99247f0_515);
nor \U$16286 ( \16969 , \16968 , \10823 );
nor \U$16287 ( \16970 , \11586 , \2253 );
nor \U$16288 ( \16971 , \16969 , \16970 );
not \U$16289 ( \16972 , \11573 );
not \U$16290 ( \16973 , \2255 );
and \U$16291 ( \16974 , \16972 , \16973 );
and \U$16292 ( \16975 , \11604 , RI9926140_475);
nor \U$16293 ( \16976 , \16974 , \16975 );
nand \U$16294 ( \16977 , \16971 , \16976 );
nor \U$16295 ( \16978 , \10874 , \2237 );
nor \U$16296 ( \16979 , \10862 , \2248 );
nor \U$16297 ( \16980 , \16978 , \16979 );
not \U$16298 ( \16981 , RI992cd10_335);
nor \U$16299 ( \16982 , \16981 , \16698 );
nor \U$16300 ( \16983 , \10885 , \6953 );
nor \U$16301 ( \16984 , \16982 , \16983 );
nand \U$16302 ( \16985 , \16980 , \16984 );
nor \U$16303 ( \16986 , \16977 , \16985 );
nand \U$16304 ( \16987 , \16967 , \16986 );
not \U$16305 ( \16988 , \16987 );
not \U$16306 ( \16989 , \16988 );
or \U$16307 ( \16990 , \16889 , \16989 );
or \U$16308 ( \16991 , \16742 , \16988 );
nand \U$16309 ( \16992 , \16990 , \16991 );
nand \U$16310 ( \16993 , \16949 , \16992 );
nand \U$16311 ( \16994 , \16943 , \16993 );
not \U$16312 ( \16995 , \16922 );
not \U$16313 ( \16996 , \16995 );
not \U$16314 ( \16997 , \11559 );
not \U$16315 ( \16998 , \6783 );
and \U$16316 ( \16999 , \16997 , \16998 );
nor \U$16317 ( \17000 , \10812 , \6787 );
nor \U$16318 ( \17001 , \16999 , \17000 );
and \U$16319 ( \17002 , \16643 , RI9931888_274);
not \U$16320 ( \17003 , RI9922978_574);
not \U$16321 ( \17004 , \16609 );
or \U$16322 ( \17005 , \17003 , \17004 );
or \U$16323 ( \17006 , \16676 , \2036 );
nand \U$16324 ( \17007 , \17005 , \17006 );
nor \U$16325 ( \17008 , \17002 , \17007 );
nand \U$16326 ( \17009 , \16958 , RI9926b18_454);
nand \U$16327 ( \17010 , \17001 , \17008 , \17009 );
not \U$16328 ( \17011 , \11599 );
not \U$16329 ( \17012 , \2043 );
and \U$16330 ( \17013 , \17011 , \17012 );
and \U$16331 ( \17014 , \11569 , RI9929188_394);
nor \U$16332 ( \17015 , \17013 , \17014 );
nand \U$16333 ( \17016 , \17015 , \12457 );
nor \U$16334 ( \17017 , \17010 , \17016 );
nor \U$16335 ( \17018 , \10823 , \6761 );
nor \U$16336 ( \17019 , \11586 , \2064 );
nor \U$16337 ( \17020 , \17018 , \17019 );
not \U$16338 ( \17021 , \16581 );
and \U$16339 ( \17022 , \17021 , RI992a8f8_374);
and \U$16340 ( \17023 , \11604 , RI99261b8_474);
nor \U$16341 ( \17024 , \17022 , \17023 );
nand \U$16342 ( \17025 , \17020 , \17024 );
not \U$16343 ( \17026 , \10862 );
not \U$16344 ( \17027 , \12424 );
and \U$16345 ( \17028 , \17026 , \17027 );
and \U$16346 ( \17029 , \16801 , RI992b258_354);
nor \U$16347 ( \17030 , \17028 , \17029 );
and \U$16348 ( \17031 , \16594 , RI992d6e8_314);
not \U$16349 ( \17032 , RI992cd88_334);
nor \U$16350 ( \17033 , \17032 , \16590 );
nor \U$16351 ( \17034 , \17031 , \17033 );
nand \U$16352 ( \17035 , \17030 , \17034 );
nor \U$16353 ( \17036 , \17025 , \17035 );
and \U$16354 ( \17037 , \17017 , \17036 );
not \U$16355 ( \17038 , \17037 );
not \U$16356 ( \17039 , \17038 );
or \U$16357 ( \17040 , \16996 , \17039 );
nand \U$16358 ( \17041 , \16944 , \17037 );
nand \U$16359 ( \17042 , \17040 , \17041 );
not \U$16360 ( \17043 , \17042 );
not \U$16361 ( \17044 , \16922 );
nand \U$16362 ( \17045 , \16493 , \16914 );
not \U$16363 ( \17046 , \17045 );
not \U$16364 ( \17047 , \16911 );
or \U$16365 ( \17048 , \17046 , \17047 );
or \U$16366 ( \17049 , \16911 , \17045 );
nand \U$16367 ( \17050 , \17048 , \17049 );
not \U$16368 ( \17051 , \17050 );
nand \U$16369 ( \17052 , \17044 , \17051 );
nand \U$16370 ( \17053 , \16922 , \17050 );
nand \U$16371 ( \17054 , \16524 , \16494 );
xnor \U$16372 ( \17055 , \16908 , \17054 );
not \U$16373 ( \17056 , \17055 );
not \U$16374 ( \17057 , \17056 );
not \U$16375 ( \17058 , \17057 );
not \U$16376 ( \17059 , \17051 );
or \U$16377 ( \17060 , \17058 , \17059 );
buf \U$16378 ( \17061 , \17055 );
not \U$16379 ( \17062 , \17061 );
nand \U$16380 ( \17063 , \17050 , \17062 );
nand \U$16381 ( \17064 , \17060 , \17063 );
not \U$16382 ( \17065 , \17064 );
and \U$16383 ( \17066 , \17052 , \17053 , \17065 );
not \U$16384 ( \17067 , \17066 );
or \U$16385 ( \17068 , \17043 , \17067 );
not \U$16386 ( \17069 , \11559 );
not \U$16387 ( \17070 , \12208 );
and \U$16388 ( \17071 , \17069 , \17070 );
nor \U$16389 ( \17072 , \10812 , \12212 );
nor \U$16390 ( \17073 , \17071 , \17072 );
and \U$16391 ( \17074 , \16643 , RI9931900_273);
not \U$16392 ( \17075 , RI99229f0_573);
not \U$16393 ( \17076 , \16609 );
or \U$16394 ( \17077 , \17075 , \17076 );
or \U$16395 ( \17078 , \16676 , \2108 );
nand \U$16396 ( \17079 , \17077 , \17078 );
nor \U$16397 ( \17080 , \17074 , \17079 );
nand \U$16398 ( \17081 , \16958 , RI9926b90_453);
nand \U$16399 ( \17082 , \17073 , \17080 , \17081 );
not \U$16400 ( \17083 , \11599 );
not \U$16401 ( \17084 , \2115 );
and \U$16402 ( \17085 , \17083 , \17084 );
and \U$16403 ( \17086 , \11569 , RI9929200_393);
nor \U$16404 ( \17087 , \17085 , \17086 );
nand \U$16405 ( \17088 , \17087 , \12239 );
nor \U$16406 ( \17089 , \17082 , \17088 );
not \U$16407 ( \17090 , \10823 );
not \U$16408 ( \17091 , \12222 );
and \U$16409 ( \17092 , \17090 , \17091 );
nor \U$16410 ( \17093 , \11586 , \2136 );
nor \U$16411 ( \17094 , \17092 , \17093 );
and \U$16412 ( \17095 , \17021 , RI992a970_373);
and \U$16413 ( \17096 , \11604 , RI9926230_473);
nor \U$16414 ( \17097 , \17095 , \17096 );
nand \U$16415 ( \17098 , \17094 , \17097 );
not \U$16416 ( \17099 , \10862 );
not \U$16417 ( \17100 , \12225 );
and \U$16418 ( \17101 , \17099 , \17100 );
and \U$16419 ( \17102 , \16801 , RI992b2d0_353);
nor \U$16420 ( \17103 , \17101 , \17102 );
and \U$16421 ( \17104 , \16594 , RI992ecf0_313);
not \U$16422 ( \17105 , RI992ce00_333);
nor \U$16423 ( \17106 , \17105 , \16698 );
nor \U$16424 ( \17107 , \17104 , \17106 );
nand \U$16425 ( \17108 , \17103 , \17107 );
nor \U$16426 ( \17109 , \17098 , \17108 );
nand \U$16427 ( \17110 , \17089 , \17109 );
not \U$16428 ( \17111 , \17110 );
not \U$16429 ( \17112 , \17111 );
not \U$16430 ( \17113 , \17112 );
not \U$16431 ( \17114 , \16995 );
or \U$16432 ( \17115 , \17113 , \17114 );
nand \U$16433 ( \17116 , \16922 , \17111 );
nand \U$16434 ( \17117 , \17115 , \17116 );
buf \U$16435 ( \17118 , \17064 );
nand \U$16436 ( \17119 , \17117 , \17118 );
nand \U$16437 ( \17120 , \17068 , \17119 );
or \U$16438 ( \17121 , \16994 , \17120 );
not \U$16439 ( \17122 , \11559 );
not \U$16440 ( \17123 , \2285 );
and \U$16441 ( \17124 , \17122 , \17123 );
nor \U$16442 ( \17125 , \11563 , \7477 );
nor \U$16443 ( \17126 , \17124 , \17125 );
and \U$16444 ( \17127 , \16643 , RI99316a8_278);
not \U$16445 ( \17128 , RI9922798_578);
not \U$16446 ( \17129 , \16609 );
or \U$16447 ( \17130 , \17128 , \17129 );
or \U$16448 ( \17131 , \16676 , \2302 );
nand \U$16449 ( \17132 , \17130 , \17131 );
nor \U$16450 ( \17133 , \17127 , \17132 );
nand \U$16451 ( \17134 , \16958 , RI9926938_458);
nand \U$16452 ( \17135 , \17126 , \17133 , \17134 );
not \U$16453 ( \17136 , \11599 );
not \U$16454 ( \17137 , RI992f3f8_298);
not \U$16455 ( \17138 , \17137 );
and \U$16456 ( \17139 , \17136 , \17138 );
and \U$16457 ( \17140 , \11569 , RI9928fa8_398);
nor \U$16458 ( \17141 , \17139 , \17140 );
nand \U$16459 ( \17142 , \17141 , \13090 );
nor \U$16460 ( \17143 , \17135 , \17142 );
not \U$16461 ( \17144 , \11586 );
not \U$16462 ( \17145 , \2327 );
and \U$16463 ( \17146 , \17144 , \17145 );
and \U$16464 ( \17147 , \16801 , RI992b078_358);
nor \U$16465 ( \17148 , \17146 , \17147 );
and \U$16466 ( \17149 , \11604 , RI9925fd8_478);
nor \U$16467 ( \17150 , \11573 , \2324 );
nor \U$16468 ( \17151 , \17149 , \17150 );
nand \U$16469 ( \17152 , \17148 , \17151 );
not \U$16470 ( \17153 , \16590 );
not \U$16471 ( \17154 , \2308 );
and \U$16472 ( \17155 , \17153 , \17154 );
and \U$16473 ( \17156 , \16594 , RI992d508_318);
nor \U$16474 ( \17157 , \17155 , \17156 );
and \U$16475 ( \17158 , \16671 , RI9925678_498);
and \U$16476 ( \17159 , \16656 , RI9924688_518);
nor \U$16477 ( \17160 , \17158 , \17159 );
nand \U$16478 ( \17161 , \17157 , \17160 );
nor \U$16479 ( \17162 , \17152 , \17161 );
nand \U$16480 ( \17163 , \17143 , \17162 );
buf \U$16481 ( \17164 , \17163 );
not \U$16482 ( \17165 , \17164 );
not \U$16483 ( \17166 , \16569 );
not \U$16484 ( \17167 , \17166 );
or \U$16485 ( \17168 , \17165 , \17167 );
not \U$16486 ( \17169 , \17166 );
not \U$16487 ( \17170 , \17164 );
nand \U$16488 ( \17171 , \17169 , \17170 );
nand \U$16489 ( \17172 , \17168 , \17171 );
not \U$16490 ( \17173 , \17172 );
not \U$16491 ( \17174 , \16758 );
or \U$16492 ( \17175 , \17173 , \17174 );
not \U$16493 ( \17176 , \16570 );
not \U$16494 ( \17177 , \10794 );
not \U$16495 ( \17178 , \2346 );
and \U$16496 ( \17179 , \17177 , \17178 );
and \U$16497 ( \17180 , \16643 , RI9931720_277);
nor \U$16498 ( \17181 , \17179 , \17180 );
nor \U$16499 ( \17182 , \16698 , \2356 );
nor \U$16500 ( \17183 , \10812 , \7268 );
nor \U$16501 ( \17184 , \17182 , \17183 );
nand \U$16502 ( \17185 , \10931 , RI9927d60_437);
nand \U$16503 ( \17186 , \17181 , \17184 , \17185 );
not \U$16504 ( \17187 , \11586 );
not \U$16505 ( \17188 , \2365 );
and \U$16506 ( \17189 , \17187 , \17188 );
and \U$16507 ( \17190 , \16594 , RI992d580_317);
nor \U$16508 ( \17191 , \17189 , \17190 );
and \U$16509 ( \17192 , \11576 , RI992b0f0_357);
and \U$16510 ( \17193 , \16656 , RI9924700_517);
nor \U$16511 ( \17194 , \17192 , \17193 );
nand \U$16512 ( \17195 , \17191 , \17194 );
nor \U$16513 ( \17196 , \17186 , \17195 );
and \U$16514 ( \17197 , \11574 , RI992a790_377);
nor \U$16515 ( \17198 , \11603 , \2349 );
nor \U$16516 ( \17199 , \17197 , \17198 );
and \U$16517 ( \17200 , \11030 , RI992f470_297);
and \U$16518 ( \17201 , \11569 , RI9929020_397);
nor \U$16519 ( \17202 , \17200 , \17201 );
nand \U$16520 ( \17203 , \17199 , \17202 );
and \U$16521 ( \17204 , \16671 , RI99256f0_497);
not \U$16522 ( \17205 , RI9922810_577);
not \U$16523 ( \17206 , \16609 );
or \U$16524 ( \17207 , \17205 , \17206 );
or \U$16525 ( \17208 , \16676 , \2391 );
nand \U$16526 ( \17209 , \17207 , \17208 );
nor \U$16527 ( \17210 , \17204 , \17209 );
nand \U$16528 ( \17211 , \13140 , \17210 );
nor \U$16529 ( \17212 , \17203 , \17211 );
nand \U$16530 ( \17213 , \17196 , \17212 );
buf \U$16531 ( \17214 , \17213 );
not \U$16532 ( \17215 , \17214 );
or \U$16533 ( \17216 , \17176 , \17215 );
not \U$16534 ( \17217 , \17214 );
nand \U$16535 ( \17218 , \16569 , \17217 );
nand \U$16536 ( \17219 , \17216 , \17218 );
nand \U$16537 ( \17220 , \17219 , \16750 );
nand \U$16538 ( \17221 , \17175 , \17220 );
and \U$16539 ( \17222 , \17121 , \17221 );
and \U$16540 ( \17223 , \16994 , \17120 );
nor \U$16541 ( \17224 , \17222 , \17223 );
not \U$16542 ( \17225 , \17224 );
not \U$16543 ( \17226 , \16500 );
nand \U$16544 ( \17227 , \17226 , \16503 );
buf \U$16545 ( \17228 , \16501 );
xor \U$16546 ( \17229 , \17227 , \17228 );
not \U$16547 ( \17230 , \17229 );
not \U$16548 ( \17231 , \17230 );
not \U$16549 ( \17232 , RI994e4d8_13);
not \U$16550 ( \17233 , \16086 );
or \U$16551 ( \17234 , \17232 , \17233 );
not \U$16552 ( \17235 , \17228 );
nand \U$16553 ( \17236 , \17234 , \17235 );
not \U$16554 ( \17237 , \17236 );
not \U$16555 ( \17238 , \17237 );
and \U$16556 ( \17239 , \17231 , \17238 );
not \U$16557 ( \17240 , \17230 );
not \U$16558 ( \17241 , \17240 );
not \U$16559 ( \17242 , \16624 );
or \U$16560 ( \17243 , \17241 , \17242 );
nand \U$16561 ( \17244 , \16623 , \17230 );
nand \U$16562 ( \17245 , \17243 , \17244 );
and \U$16563 ( \17246 , \17240 , \17237 );
and \U$16564 ( \17247 , \17245 , \17246 );
nor \U$16565 ( \17248 , \17239 , \17247 );
not \U$16566 ( \17249 , \17248 );
not \U$16567 ( \17250 , \16511 );
nand \U$16568 ( \17251 , \17250 , \16509 );
not \U$16569 ( \17252 , \17251 );
buf \U$16570 ( \17253 , \16508 );
not \U$16571 ( \17254 , \17253 );
or \U$16572 ( \17255 , \17252 , \17254 );
or \U$16573 ( \17256 , \17253 , \17251 );
nand \U$16574 ( \17257 , \17255 , \17256 );
nand \U$16575 ( \17258 , \16498 , \16507 );
xnor \U$16576 ( \17259 , \16504 , \17258 );
and \U$16577 ( \17260 , \17257 , \17259 );
not \U$16578 ( \17261 , \17257 );
not \U$16579 ( \17262 , \17259 );
and \U$16580 ( \17263 , \17261 , \17262 );
nor \U$16581 ( \17264 , \17260 , \17263 );
and \U$16582 ( \17265 , \17259 , \17229 );
not \U$16583 ( \17266 , \17259 );
and \U$16584 ( \17267 , \17266 , \17230 );
or \U$16585 ( \17268 , \17265 , \17267 );
nand \U$16586 ( \17269 , \17264 , \17268 );
not \U$16587 ( \17270 , \17269 );
not \U$16588 ( \17271 , \17270 );
buf \U$16589 ( \17272 , \17257 );
buf \U$16590 ( \17273 , \17272 );
and \U$16591 ( \17274 , \17273 , \16730 );
not \U$16592 ( \17275 , \17273 );
not \U$16593 ( \17276 , \16730 );
and \U$16594 ( \17277 , \17275 , \17276 );
nor \U$16595 ( \17278 , \17274 , \17277 );
not \U$16596 ( \17279 , \17278 );
or \U$16597 ( \17280 , \17271 , \17279 );
and \U$16598 ( \17281 , \17273 , \16682 );
not \U$16599 ( \17282 , \17273 );
and \U$16600 ( \17283 , \17282 , \16683 );
nor \U$16601 ( \17284 , \17281 , \17283 );
not \U$16602 ( \17285 , \17268 );
nand \U$16603 ( \17286 , \17284 , \17285 );
nand \U$16604 ( \17287 , \17280 , \17286 );
nand \U$16605 ( \17288 , \17249 , \17287 );
not \U$16606 ( \17289 , \17285 );
not \U$16607 ( \17290 , \17273 );
and \U$16608 ( \17291 , \17290 , \16624 );
not \U$16609 ( \17292 , \17290 );
and \U$16610 ( \17293 , \17292 , \16623 );
nor \U$16611 ( \17294 , \17291 , \17293 );
not \U$16612 ( \17295 , \17294 );
or \U$16613 ( \17296 , \17289 , \17295 );
not \U$16614 ( \17297 , \17284 );
or \U$16615 ( \17298 , \17297 , \17269 );
nand \U$16616 ( \17299 , \17296 , \17298 );
xor \U$16617 ( \17300 , \17288 , \17299 );
not \U$16618 ( \17301 , \17300 );
not \U$16619 ( \17302 , \17117 );
buf \U$16620 ( \17303 , \17066 );
not \U$16621 ( \17304 , \17303 );
or \U$16622 ( \17305 , \17302 , \17304 );
not \U$16623 ( \17306 , RI9927fb8_432);
nor \U$16624 ( \17307 , \11559 , \17306 );
not \U$16625 ( \17308 , RI9928918_412);
nor \U$16626 ( \17309 , \17308 , \11563 );
nor \U$16627 ( \17310 , \17307 , \17309 );
and \U$16628 ( \17311 , \16643 , RI9931978_272);
and \U$16629 ( \17312 , RI9923698_552, \16605 );
and \U$16630 ( \17313 , \16609 , RI9922a68_572);
nor \U$16631 ( \17314 , \17311 , \17312 , \17313 );
nand \U$16632 ( \17315 , \16958 , RI9926c08_452);
nand \U$16633 ( \17316 , \17310 , \17314 , \17315 );
not \U$16634 ( \17317 , RI992f6c8_292);
nor \U$16635 ( \17318 , \17317 , \11599 );
not \U$16636 ( \17319 , RI9929278_392);
nor \U$16637 ( \17320 , \17319 , \11568 );
nor \U$16638 ( \17321 , \17318 , \17320 );
nand \U$16639 ( \17322 , \17321 , \12296 );
nor \U$16640 ( \17323 , \17316 , \17322 );
and \U$16641 ( \17324 , \16801 , RI992b348_352);
nor \U$16642 ( \17325 , \11603 , \1884 );
nor \U$16643 ( \17326 , \17324 , \17325 );
and \U$16644 ( \17327 , \11574 , RI992a9e8_372);
not \U$16645 ( \17328 , RI9923ff8_532);
nor \U$16646 ( \17329 , \17328 , \11586 );
nor \U$16647 ( \17330 , \17327 , \17329 );
nand \U$16648 ( \17331 , \17326 , \17330 );
nand \U$16649 ( \17332 , \16656 , RI9924958_512);
nand \U$16650 ( \17333 , \16594 , RI992ed68_312);
nand \U$16651 ( \17334 , \11582 , RI992ce78_332);
nand \U$16652 ( \17335 , \16671 , RI9925948_492);
nand \U$16653 ( \17336 , \17332 , \17333 , \17334 , \17335 );
nor \U$16654 ( \17337 , \17331 , \17336 );
nand \U$16655 ( \17338 , \17323 , \17337 );
not \U$16656 ( \17339 , \17338 );
not \U$16657 ( \17340 , \16995 );
or \U$16658 ( \17341 , \17339 , \17340 );
not \U$16659 ( \17342 , \17338 );
nand \U$16660 ( \17343 , \16944 , \17342 );
nand \U$16661 ( \17344 , \17341 , \17343 );
nand \U$16662 ( \17345 , \17344 , \17118 );
nand \U$16663 ( \17346 , \17305 , \17345 );
not \U$16664 ( \17347 , \17346 );
and \U$16665 ( \17348 , \17301 , \17347 );
and \U$16666 ( \17349 , \17346 , \17300 );
nor \U$16667 ( \17350 , \17348 , \17349 );
not \U$16668 ( \17351 , \17350 );
and \U$16669 ( \17352 , \17225 , \17351 );
not \U$16670 ( \17353 , \17225 );
and \U$16671 ( \17354 , \17353 , \17350 );
nor \U$16672 ( \17355 , \17352 , \17354 );
not \U$16673 ( \17356 , \17230 );
and \U$16674 ( \17357 , \16825 , \17056 );
not \U$16675 ( \17358 , \16825 );
and \U$16676 ( \17359 , \17358 , \17057 );
nor \U$16677 ( \17360 , \17357 , \17359 );
not \U$16678 ( \17361 , \17360 );
not \U$16679 ( \17362 , \16514 );
nand \U$16680 ( \17363 , \17362 , \16907 );
xnor \U$16681 ( \17364 , \16904 , \17363 );
not \U$16682 ( \17365 , \17364 );
and \U$16683 ( \17366 , \17272 , \17365 );
not \U$16684 ( \17367 , \17272 );
and \U$16685 ( \17368 , \17367 , \17364 );
nor \U$16686 ( \17369 , \17366 , \17368 );
nand \U$16687 ( \17370 , \17055 , \17364 );
not \U$16688 ( \17371 , \17055 );
nand \U$16689 ( \17372 , \17371 , \17365 );
and \U$16690 ( \17373 , \17369 , \17370 , \17372 );
not \U$16691 ( \17374 , \17373 );
or \U$16692 ( \17375 , \17361 , \17374 );
and \U$16693 ( \17376 , \17276 , \17056 );
not \U$16694 ( \17377 , \17276 );
and \U$16695 ( \17378 , \17377 , \17057 );
nor \U$16696 ( \17379 , \17376 , \17378 );
buf \U$16697 ( \17380 , \17369 );
not \U$16698 ( \17381 , \17380 );
nand \U$16699 ( \17382 , \17379 , \17381 );
nand \U$16700 ( \17383 , \17375 , \17382 );
not \U$16701 ( \17384 , \17383 );
or \U$16702 ( \17385 , \17356 , \17384 );
not \U$16703 ( \17386 , \17383 );
nand \U$16704 ( \17387 , \17386 , \17240 );
nand \U$16705 ( \17388 , \17385 , \17387 );
not \U$16706 ( \17389 , \17219 );
buf \U$16707 ( \17390 , \16756 );
not \U$16708 ( \17391 , \17390 );
or \U$16709 ( \17392 , \17389 , \17391 );
and \U$16710 ( \17393 , \16888 , \16569 );
not \U$16711 ( \17394 , \16888 );
not \U$16712 ( \17395 , \16569 );
and \U$16713 ( \17396 , \17394 , \17395 );
nor \U$16714 ( \17397 , \17393 , \17396 );
nand \U$16715 ( \17398 , \17397 , \16750 );
nand \U$16716 ( \17399 , \17392 , \17398 );
xor \U$16717 ( \17400 , \17388 , \17399 );
not \U$16718 ( \17401 , \16992 );
buf \U$16719 ( \17402 , \16941 );
not \U$16720 ( \17403 , \17402 );
or \U$16721 ( \17404 , \17401 , \17403 );
buf \U$16722 ( \17405 , \16949 );
buf \U$16723 ( \17406 , \17038 );
and \U$16724 ( \17407 , \17406 , \16893 );
not \U$16725 ( \17408 , \17406 );
and \U$16726 ( \17409 , \17408 , \16894 );
nor \U$16727 ( \17410 , \17407 , \17409 );
nand \U$16728 ( \17411 , \17405 , \17410 );
nand \U$16729 ( \17412 , \17404 , \17411 );
xor \U$16730 ( \17413 , \17400 , \17412 );
xnor \U$16731 ( \17414 , \17355 , \17413 );
not \U$16732 ( \17415 , \17414 );
not \U$16733 ( \17416 , \17110 );
not \U$16734 ( \17417 , \17062 );
or \U$16735 ( \17418 , \17416 , \17417 );
nand \U$16736 ( \17419 , \17061 , \17111 );
nand \U$16737 ( \17420 , \17418 , \17419 );
not \U$16738 ( \17421 , \17420 );
not \U$16739 ( \17422 , \17373 );
or \U$16740 ( \17423 , \17421 , \17422 );
not \U$16741 ( \17424 , \17061 );
and \U$16742 ( \17425 , \17342 , \17424 );
not \U$16743 ( \17426 , \17342 );
and \U$16744 ( \17427 , \17426 , \17061 );
nor \U$16745 ( \17428 , \17425 , \17427 );
nand \U$16746 ( \17429 , \17428 , \17381 );
nand \U$16747 ( \17430 , \17423 , \17429 );
not \U$16748 ( \17431 , \17285 );
not \U$16749 ( \17432 , \17273 );
not \U$16750 ( \17433 , \16825 );
or \U$16751 ( \17434 , \17432 , \17433 );
nand \U$16752 ( \17435 , \16824 , \17290 );
nand \U$16753 ( \17436 , \17434 , \17435 );
not \U$16754 ( \17437 , \17436 );
or \U$16755 ( \17438 , \17431 , \17437 );
xor \U$16756 ( \17439 , \17273 , \17338 );
nand \U$16757 ( \17440 , \17439 , \17270 );
nand \U$16758 ( \17441 , \17438 , \17440 );
not \U$16759 ( \17442 , \17236 );
and \U$16760 ( \17443 , \17240 , \16682 );
not \U$16761 ( \17444 , \17240 );
and \U$16762 ( \17445 , \17444 , \16683 );
nor \U$16763 ( \17446 , \17443 , \17445 );
not \U$16764 ( \17447 , \17446 );
or \U$16765 ( \17448 , \17442 , \17447 );
and \U$16766 ( \17449 , \16730 , \17230 );
not \U$16767 ( \17450 , \16730 );
and \U$16768 ( \17451 , \17450 , \17240 );
or \U$16769 ( \17452 , \17449 , \17451 );
nand \U$16770 ( \17453 , \17452 , \17246 );
nand \U$16771 ( \17454 , \17448 , \17453 );
and \U$16772 ( \17455 , \17441 , \17454 );
xor \U$16773 ( \17456 , \17430 , \17455 );
not \U$16774 ( \17457 , \17270 );
not \U$16775 ( \17458 , \17436 );
or \U$16776 ( \17459 , \17457 , \17458 );
nand \U$16777 ( \17460 , \17278 , \17285 );
nand \U$16778 ( \17461 , \17459 , \17460 );
not \U$16779 ( \17462 , \17246 );
not \U$16780 ( \17463 , \17446 );
or \U$16781 ( \17464 , \17462 , \17463 );
nand \U$16782 ( \17465 , \17245 , \17236 );
nand \U$16783 ( \17466 , \17464 , \17465 );
xor \U$16784 ( \17467 , \17461 , \17466 );
and \U$16785 ( \17468 , \17456 , \17467 );
and \U$16786 ( \17469 , \17430 , \17455 );
or \U$16787 ( \17470 , \17468 , \17469 );
not \U$16788 ( \17471 , RI9931540_281);
nor \U$16789 ( \17472 , \17471 , \10849 );
nor \U$16790 ( \17473 , \10794 , \2563 );
nor \U$16791 ( \17474 , \17472 , \17473 );
not \U$16792 ( \17475 , \11563 );
and \U$16793 ( \17476 , \17475 , RI99284e0_421);
nor \U$16794 ( \17477 , \16698 , \2573 );
nor \U$16795 ( \17478 , \17476 , \17477 );
nand \U$16796 ( \17479 , \10931 , RI9927b80_441);
nand \U$16797 ( \17480 , \17474 , \17478 , \17479 );
and \U$16798 ( \17481 , \16654 , RI9923bc0_541);
nor \U$16799 ( \17482 , \10885 , \2552 );
nor \U$16800 ( \17483 , \17481 , \17482 );
and \U$16801 ( \17484 , \11576 , RI992af10_361);
and \U$16802 ( \17485 , \16656 , RI9924520_521);
nor \U$16803 ( \17486 , \17484 , \17485 );
nand \U$16804 ( \17487 , \17483 , \17486 );
nor \U$16805 ( \17488 , \17480 , \17487 );
and \U$16806 ( \17489 , \11574 , RI992a5b0_381);
and \U$16807 ( \17490 , \11604 , RI9925e70_481);
nor \U$16808 ( \17491 , \17489 , \17490 );
and \U$16809 ( \17492 , \11030 , RI992f290_301);
and \U$16810 ( \17493 , \11569 , RI9928e40_401);
nor \U$16811 ( \17494 , \17492 , \17493 );
nand \U$16812 ( \17495 , \17491 , \17494 );
and \U$16813 ( \17496 , \16671 , RI9925510_501);
not \U$16814 ( \17497 , RI9923260_561);
not \U$16815 ( \17498 , \16605 );
or \U$16816 ( \17499 , \17497 , \17498 );
nand \U$16817 ( \17500 , \16609 , RI9922630_581);
nand \U$16818 ( \17501 , \17499 , \17500 );
nor \U$16819 ( \17502 , \17496 , \17501 );
nand \U$16820 ( \17503 , \13786 , \17502 );
nor \U$16821 ( \17504 , \17495 , \17503 );
nand \U$16822 ( \17505 , \17488 , \17504 );
buf \U$16823 ( \17506 , \17505 );
not \U$16824 ( \17507 , \16635 );
and \U$16825 ( \17508 , \17506 , \17507 );
not \U$16826 ( \17509 , \17506 );
and \U$16827 ( \17510 , \17509 , \16635 );
nor \U$16828 ( \17511 , \17508 , \17510 );
and \U$16829 ( \17512 , \16639 , \17511 );
xor \U$16830 ( \17513 , \17470 , \17512 );
not \U$16831 ( \17514 , \10794 );
not \U$16832 ( \17515 , \2786 );
and \U$16833 ( \17516 , \17514 , \17515 );
and \U$16834 ( \17517 , \16643 , RI99315b8_280);
nor \U$16835 ( \17518 , \17516 , \17517 );
not \U$16836 ( \17519 , \10812 );
not \U$16837 ( \17520 , \2773 );
and \U$16838 ( \17521 , \17519 , \17520 );
nor \U$16839 ( \17522 , \16590 , \2776 );
nor \U$16840 ( \17523 , \17521 , \17522 );
nand \U$16841 ( \17524 , \10931 , RI9927bf8_440);
nand \U$16842 ( \17525 , \17518 , \17523 , \17524 );
nor \U$16843 ( \17526 , \10823 , \7853 );
nor \U$16844 ( \17527 , \10874 , \2764 );
nor \U$16845 ( \17528 , \17526 , \17527 );
not \U$16846 ( \17529 , \11586 );
not \U$16847 ( \17530 , \2790 );
and \U$16848 ( \17531 , \17529 , \17530 );
and \U$16849 ( \17532 , \16594 , RI992d418_320);
nor \U$16850 ( \17533 , \17531 , \17532 );
nand \U$16851 ( \17534 , \17528 , \17533 );
nor \U$16852 ( \17535 , \17525 , \17534 );
not \U$16853 ( \17536 , \11603 );
not \U$16854 ( \17537 , \2783 );
and \U$16855 ( \17538 , \17536 , \17537 );
and \U$16856 ( \17539 , \17021 , RI992a628_380);
nor \U$16857 ( \17540 , \17538 , \17539 );
not \U$16858 ( \17541 , \11599 );
not \U$16859 ( \17542 , \2758 );
and \U$16860 ( \17543 , \17541 , \17542 );
and \U$16861 ( \17544 , \16619 , RI9928eb8_400);
nor \U$16862 ( \17545 , \17543 , \17544 );
nand \U$16863 ( \17546 , \17540 , \17545 );
not \U$16864 ( \17547 , \10862 );
not \U$16865 ( \17548 , \2771 );
and \U$16866 ( \17549 , \17547 , \17548 );
not \U$16867 ( \17550 , RI99232d8_560);
not \U$16868 ( \17551 , \16605 );
or \U$16869 ( \17552 , \17550 , \17551 );
nand \U$16870 ( \17553 , \16609 , RI99226a8_580);
nand \U$16871 ( \17554 , \17552 , \17553 );
nor \U$16872 ( \17555 , \17549 , \17554 );
nand \U$16873 ( \17556 , \13494 , \17555 );
nor \U$16874 ( \17557 , \17546 , \17556 );
nand \U$16875 ( \17558 , \17535 , \17557 );
buf \U$16876 ( \17559 , \17558 );
not \U$16877 ( \17560 , \17559 );
not \U$16878 ( \17561 , \16765 );
not \U$16879 ( \17562 , \17561 );
or \U$16880 ( \17563 , \17560 , \17562 );
not \U$16881 ( \17564 , \17559 );
nand \U$16882 ( \17565 , \16765 , \17564 );
nand \U$16883 ( \17566 , \17563 , \17565 );
not \U$16884 ( \17567 , \17566 );
not \U$16885 ( \17568 , \16572 );
or \U$16886 ( \17569 , \17567 , \17568 );
not \U$16887 ( \17570 , \16571 );
nand \U$16888 ( \17571 , \10931 , RI9927c70_439);
nand \U$16889 ( \17572 , \11028 , RI99285d0_419);
nand \U$16890 ( \17573 , \11582 , RI992cb30_339);
and \U$16891 ( \17574 , \17571 , \17572 , \17573 );
not \U$16892 ( \17575 , \10794 );
not \U$16893 ( \17576 , \13172 );
and \U$16894 ( \17577 , \17575 , \17576 );
and \U$16895 ( \17578 , \16643 , RI9931630_279);
nor \U$16896 ( \17579 , \17577 , \17578 );
not \U$16897 ( \17580 , \10885 );
not \U$16898 ( \17581 , \7634 );
and \U$16899 ( \17582 , \17580 , \17581 );
and \U$16900 ( \17583 , \11576 , RI992b000_359);
nor \U$16901 ( \17584 , \17582 , \17583 );
not \U$16902 ( \17585 , \10823 );
not \U$16903 ( \17586 , \13176 );
and \U$16904 ( \17587 , \17585 , \17586 );
nor \U$16905 ( \17588 , \11586 , \13160 );
nor \U$16906 ( \17589 , \17587 , \17588 );
nand \U$16907 ( \17590 , \17574 , \17579 , \17584 , \17589 );
not \U$16908 ( \17591 , \11599 );
not \U$16909 ( \17592 , \2431 );
and \U$16910 ( \17593 , \17591 , \17592 );
and \U$16911 ( \17594 , \16619 , RI9928f30_399);
nor \U$16912 ( \17595 , \17593 , \17594 );
not \U$16913 ( \17596 , \11603 );
not \U$16914 ( \17597 , \7628 );
and \U$16915 ( \17598 , \17596 , \17597 );
and \U$16916 ( \17599 , \17021 , RI992a6a0_379);
nor \U$16917 ( \17600 , \17598 , \17599 );
not \U$16918 ( \17601 , \10862 );
not \U$16919 ( \17602 , \13179 );
and \U$16920 ( \17603 , \17601 , \17602 );
not \U$16921 ( \17604 , RI9922720_579);
not \U$16922 ( \17605 , \16609 );
or \U$16923 ( \17606 , \17604 , \17605 );
or \U$16924 ( \17607 , \16676 , \2424 );
nand \U$16925 ( \17608 , \17606 , \17607 );
nor \U$16926 ( \17609 , \17603 , \17608 );
nand \U$16927 ( \17610 , \17595 , \17600 , \13191 , \17609 );
nor \U$16928 ( \17611 , \17590 , \17610 );
not \U$16929 ( \17612 , \17611 );
not \U$16930 ( \17613 , \17612 );
not \U$16931 ( \17614 , \16626 );
or \U$16932 ( \17615 , \17613 , \17614 );
not \U$16933 ( \17616 , \17612 );
nand \U$16934 ( \17617 , \16765 , \17616 );
nand \U$16935 ( \17618 , \17615 , \17617 );
nand \U$16936 ( \17619 , \17570 , \17618 );
nand \U$16937 ( \17620 , \17569 , \17619 );
and \U$16938 ( \17621 , \17513 , \17620 );
and \U$16939 ( \17622 , \17470 , \17512 );
or \U$16940 ( \17623 , \17621 , \17622 );
not \U$16941 ( \17624 , \17373 );
not \U$16942 ( \17625 , \17428 );
or \U$16943 ( \17626 , \17624 , \17625 );
nand \U$16944 ( \17627 , \17360 , \17381 );
nand \U$16945 ( \17628 , \17626 , \17627 );
and \U$16946 ( \17629 , \17461 , \17466 );
xor \U$16947 ( \17630 , \17628 , \17629 );
not \U$16948 ( \17631 , \17248 );
not \U$16949 ( \17632 , \17287 );
or \U$16950 ( \17633 , \17631 , \17632 );
or \U$16951 ( \17634 , \17287 , \17248 );
nand \U$16952 ( \17635 , \17633 , \17634 );
and \U$16953 ( \17636 , \17630 , \17635 );
and \U$16954 ( \17637 , \17628 , \17629 );
or \U$16955 ( \17638 , \17636 , \17637 );
not \U$16956 ( \17639 , \16642 );
and \U$16957 ( \17640 , \17559 , \17639 );
not \U$16958 ( \17641 , \17559 );
and \U$16959 ( \17642 , \17641 , \16635 );
nor \U$16960 ( \17643 , \17640 , \17642 );
and \U$16961 ( \17644 , \16637 , \17643 );
xor \U$16962 ( \17645 , \17638 , \17644 );
not \U$16963 ( \17646 , \17618 );
not \U$16964 ( \17647 , \16572 );
or \U$16965 ( \17648 , \17646 , \17647 );
not \U$16966 ( \17649 , \16571 );
not \U$16967 ( \17650 , \17164 );
not \U$16968 ( \17651 , \16626 );
or \U$16969 ( \17652 , \17650 , \17651 );
not \U$16970 ( \17653 , \17561 );
nand \U$16971 ( \17654 , \17653 , \17170 );
nand \U$16972 ( \17655 , \17652 , \17654 );
nand \U$16973 ( \17656 , \17649 , \17655 );
nand \U$16974 ( \17657 , \17648 , \17656 );
xor \U$16975 ( \17658 , \17645 , \17657 );
xor \U$16976 ( \17659 , \17623 , \17658 );
xor \U$16977 ( \17660 , \17628 , \17629 );
xor \U$16978 ( \17661 , \17660 , \17635 );
xor \U$16979 ( \17662 , \17120 , \16994 );
xor \U$16980 ( \17663 , \17662 , \17221 );
xor \U$16981 ( \17664 , \17661 , \17663 );
not \U$16982 ( \17665 , \16989 );
not \U$16983 ( \17666 , \16944 );
not \U$16984 ( \17667 , \17666 );
or \U$16985 ( \17668 , \17665 , \17667 );
nand \U$16986 ( \17669 , \16988 , \16944 );
nand \U$16987 ( \17670 , \17668 , \17669 );
not \U$16988 ( \17671 , \17670 );
not \U$16989 ( \17672 , \17303 );
or \U$16990 ( \17673 , \17671 , \17672 );
nand \U$16991 ( \17674 , \17042 , \17118 );
nand \U$16992 ( \17675 , \17673 , \17674 );
not \U$16993 ( \17676 , \17612 );
not \U$16994 ( \17677 , \16753 );
or \U$16995 ( \17678 , \17676 , \17677 );
nand \U$16996 ( \17679 , \16569 , \17616 );
nand \U$16997 ( \17680 , \17678 , \17679 );
not \U$16998 ( \17681 , \17680 );
not \U$16999 ( \17682 , \17390 );
or \U$17000 ( \17683 , \17681 , \17682 );
nand \U$17001 ( \17684 , \17172 , \16750 );
nand \U$17002 ( \17685 , \17683 , \17684 );
xor \U$17003 ( \17686 , \17675 , \17685 );
not \U$17004 ( \17687 , \16896 );
not \U$17005 ( \17688 , \17405 );
or \U$17006 ( \17689 , \17687 , \17688 );
and \U$17007 ( \17690 , \16890 , \17217 );
and \U$17008 ( \17691 , \16889 , \17214 );
nor \U$17009 ( \17692 , \17690 , \17691 );
not \U$17010 ( \17693 , \17692 );
nand \U$17011 ( \17694 , \17693 , \17402 );
nand \U$17012 ( \17695 , \17689 , \17694 );
and \U$17013 ( \17696 , \17686 , \17695 );
and \U$17014 ( \17697 , \17675 , \17685 );
or \U$17015 ( \17698 , \17696 , \17697 );
and \U$17016 ( \17699 , \17664 , \17698 );
and \U$17017 ( \17700 , \17661 , \17663 );
or \U$17018 ( \17701 , \17699 , \17700 );
xor \U$17019 ( \17702 , \17659 , \17701 );
not \U$17020 ( \17703 , \17702 );
or \U$17021 ( \17704 , \17415 , \17703 );
or \U$17022 ( \17705 , \17414 , \17702 );
nand \U$17023 ( \17706 , \17704 , \17705 );
not \U$17024 ( \17707 , \17373 );
and \U$17025 ( \17708 , \17038 , \17061 );
not \U$17026 ( \17709 , \17038 );
and \U$17027 ( \17710 , \17709 , \17424 );
nor \U$17028 ( \17711 , \17708 , \17710 );
not \U$17029 ( \17712 , \17711 );
or \U$17030 ( \17713 , \17707 , \17712 );
nand \U$17031 ( \17714 , \17420 , \17381 );
nand \U$17032 ( \17715 , \17713 , \17714 );
not \U$17033 ( \17716 , \17285 );
not \U$17034 ( \17717 , \17439 );
or \U$17035 ( \17718 , \17716 , \17717 );
not \U$17036 ( \17719 , \17273 );
not \U$17037 ( \17720 , \17111 );
or \U$17038 ( \17721 , \17719 , \17720 );
nand \U$17039 ( \17722 , \17110 , \17290 );
nand \U$17040 ( \17723 , \17721 , \17722 );
nand \U$17041 ( \17724 , \17723 , \17270 );
nand \U$17042 ( \17725 , \17718 , \17724 );
not \U$17043 ( \17726 , \17246 );
and \U$17044 ( \17727 , \17240 , \16824 );
not \U$17045 ( \17728 , \17240 );
and \U$17046 ( \17729 , \17728 , \16825 );
nor \U$17047 ( \17730 , \17727 , \17729 );
not \U$17048 ( \17731 , \17730 );
or \U$17049 ( \17732 , \17726 , \17731 );
not \U$17050 ( \17733 , \17452 );
or \U$17051 ( \17734 , \17733 , \17237 );
nand \U$17052 ( \17735 , \17732 , \17734 );
and \U$17053 ( \17736 , \17725 , \17735 );
xor \U$17054 ( \17737 , \17715 , \17736 );
xor \U$17055 ( \17738 , \17441 , \17454 );
and \U$17056 ( \17739 , \17737 , \17738 );
and \U$17057 ( \17740 , \17715 , \17736 );
or \U$17058 ( \17741 , \17739 , \17740 );
and \U$17059 ( \17742 , \10931 , RI9927b08_442);
and \U$17060 ( \17743 , \11028 , RI9928468_422);
and \U$17061 ( \17744 , \11032 , RI992c9c8_342);
nor \U$17062 ( \17745 , \17742 , \17743 , \17744 );
not \U$17063 ( \17746 , \10794 );
not \U$17064 ( \17747 , \2508 );
and \U$17065 ( \17748 , \17746 , \17747 );
and \U$17066 ( \17749 , \16643 , RI99314c8_282);
nor \U$17067 ( \17750 , \17748 , \17749 );
not \U$17068 ( \17751 , \16801 );
nor \U$17069 ( \17752 , \17751 , \2512 );
nor \U$17070 ( \17753 , \10823 , \8067 );
nor \U$17071 ( \17754 , \17752 , \17753 );
not \U$17072 ( \17755 , \11586 );
not \U$17073 ( \17756 , RI9923b48_542);
not \U$17074 ( \17757 , \17756 );
and \U$17075 ( \17758 , \17755 , \17757 );
and \U$17076 ( \17759 , \16594 , RI992d328_322);
nor \U$17077 ( \17760 , \17758 , \17759 );
nand \U$17078 ( \17761 , \17745 , \17750 , \17754 , \17760 );
not \U$17079 ( \17762 , \11599 );
not \U$17080 ( \17763 , \2519 );
and \U$17081 ( \17764 , \17762 , \17763 );
and \U$17082 ( \17765 , \11569 , RI9928dc8_402);
nor \U$17083 ( \17766 , \17764 , \17765 );
not \U$17084 ( \17767 , \11603 );
not \U$17085 ( \17768 , \2506 );
and \U$17086 ( \17769 , \17767 , \17768 );
and \U$17087 ( \17770 , \11574 , RI992a538_382);
nor \U$17088 ( \17771 , \17769 , \17770 );
and \U$17089 ( \17772 , \16671 , RI9924e08_502);
not \U$17090 ( \17773 , RI99231e8_562);
not \U$17091 ( \17774 , \16605 );
or \U$17092 ( \17775 , \17773 , \17774 );
nand \U$17093 ( \17776 , \16609 , RI99225b8_582);
nand \U$17094 ( \17777 , \17775 , \17776 );
nor \U$17095 ( \17778 , \17772 , \17777 );
nand \U$17096 ( \17779 , \17766 , \17771 , \13742 , \17778 );
nor \U$17097 ( \17780 , \17761 , \17779 );
not \U$17098 ( \17781 , \17780 );
not \U$17099 ( \17782 , \17781 );
and \U$17100 ( \17783 , \17782 , \16635 );
not \U$17101 ( \17784 , \17782 );
and \U$17102 ( \17785 , \17784 , \17639 );
nor \U$17103 ( \17786 , \17783 , \17785 );
and \U$17104 ( \17787 , \16639 , \17786 );
xor \U$17105 ( \17788 , \17741 , \17787 );
not \U$17106 ( \17789 , \16558 );
not \U$17107 ( \17790 , \17506 );
or \U$17108 ( \17791 , \17789 , \17790 );
not \U$17109 ( \17792 , \17506 );
nand \U$17110 ( \17793 , \16765 , \17792 );
nand \U$17111 ( \17794 , \17791 , \17793 );
not \U$17112 ( \17795 , \17794 );
not \U$17113 ( \17796 , \16572 );
or \U$17114 ( \17797 , \17795 , \17796 );
not \U$17115 ( \17798 , \16571 );
nand \U$17116 ( \17799 , \17798 , \17566 );
nand \U$17117 ( \17800 , \17797 , \17799 );
and \U$17118 ( \17801 , \17788 , \17800 );
and \U$17119 ( \17802 , \17741 , \17787 );
or \U$17120 ( \17803 , \17801 , \17802 );
xor \U$17121 ( \17804 , \17470 , \17512 );
xor \U$17122 ( \17805 , \17804 , \17620 );
xor \U$17123 ( \17806 , \17803 , \17805 );
xor \U$17124 ( \17807 , \17430 , \17455 );
xor \U$17125 ( \17808 , \17807 , \17467 );
not \U$17126 ( \17809 , \17405 );
not \U$17127 ( \17810 , \17809 );
not \U$17128 ( \17811 , \17692 );
and \U$17129 ( \17812 , \17810 , \17811 );
and \U$17130 ( \17813 , \17164 , \16742 );
not \U$17131 ( \17814 , \17164 );
and \U$17132 ( \17815 , \17814 , \16894 );
nor \U$17133 ( \17816 , \17813 , \17815 );
and \U$17134 ( \17817 , \17402 , \17816 );
nor \U$17135 ( \17818 , \17812 , \17817 );
not \U$17136 ( \17819 , \17818 );
not \U$17137 ( \17820 , \17303 );
not \U$17138 ( \17821 , \16888 );
not \U$17139 ( \17822 , \16995 );
or \U$17140 ( \17823 , \17821 , \17822 );
not \U$17141 ( \17824 , \16888 );
nand \U$17142 ( \17825 , \16944 , \17824 );
nand \U$17143 ( \17826 , \17823 , \17825 );
not \U$17144 ( \17827 , \17826 );
or \U$17145 ( \17828 , \17820 , \17827 );
nand \U$17146 ( \17829 , \17670 , \17118 );
nand \U$17147 ( \17830 , \17828 , \17829 );
not \U$17148 ( \17831 , \17830 );
not \U$17149 ( \17832 , \17831 );
or \U$17150 ( \17833 , \17819 , \17832 );
not \U$17151 ( \17834 , \17559 );
not \U$17152 ( \17835 , \16753 );
or \U$17153 ( \17836 , \17834 , \17835 );
nand \U$17154 ( \17837 , \16569 , \17564 );
nand \U$17155 ( \17838 , \17836 , \17837 );
not \U$17156 ( \17839 , \17838 );
not \U$17157 ( \17840 , \16756 );
or \U$17158 ( \17841 , \17839 , \17840 );
nand \U$17159 ( \17842 , \17680 , \16750 );
nand \U$17160 ( \17843 , \17841 , \17842 );
nand \U$17161 ( \17844 , \17833 , \17843 );
not \U$17162 ( \17845 , \17818 );
nand \U$17163 ( \17846 , \17845 , \17830 );
nand \U$17164 ( \17847 , \17844 , \17846 );
xor \U$17165 ( \17848 , \17808 , \17847 );
xor \U$17166 ( \17849 , \17675 , \17685 );
xor \U$17167 ( \17850 , \17849 , \17695 );
and \U$17168 ( \17851 , \17848 , \17850 );
and \U$17169 ( \17852 , \17808 , \17847 );
or \U$17170 ( \17853 , \17851 , \17852 );
and \U$17171 ( \17854 , \17806 , \17853 );
and \U$17172 ( \17855 , \17803 , \17805 );
or \U$17173 ( \17856 , \17854 , \17855 );
not \U$17174 ( \17857 , \17856 );
and \U$17175 ( \17858 , \17706 , \17857 );
not \U$17176 ( \17859 , \17706 );
and \U$17177 ( \17860 , \17859 , \17856 );
nor \U$17178 ( \17861 , \17858 , \17860 );
xor \U$17179 ( \17862 , \17661 , \17663 );
xor \U$17180 ( \17863 , \17862 , \17698 );
not \U$17181 ( \17864 , \17863 );
not \U$17182 ( \17865 , \10794 );
not \U$17183 ( \17866 , \8352 );
and \U$17184 ( \17867 , \17865 , \17866 );
and \U$17185 ( \17868 , \16643 , RI9931450_283);
nor \U$17186 ( \17869 , \17867 , \17868 );
not \U$17187 ( \17870 , \11563 );
not \U$17188 ( \17871 , \8362 );
and \U$17189 ( \17872 , \17870 , \17871 );
nor \U$17190 ( \17873 , \16698 , \8345 );
nor \U$17191 ( \17874 , \17872 , \17873 );
nand \U$17192 ( \17875 , \10931 , RI9927040_443);
nand \U$17193 ( \17876 , \17869 , \17874 , \17875 );
nor \U$17194 ( \17877 , \10823 , \8324 );
nor \U$17195 ( \17878 , \10874 , \2596 );
nor \U$17196 ( \17879 , \17877 , \17878 );
not \U$17197 ( \17880 , \10885 );
not \U$17198 ( \17881 , \8332 );
and \U$17199 ( \17882 , \17880 , \17881 );
and \U$17200 ( \17883 , \16654 , RI9923ad0_543);
nor \U$17201 ( \17884 , \17882 , \17883 );
nand \U$17202 ( \17885 , \17879 , \17884 );
nor \U$17203 ( \17886 , \17876 , \17885 );
not \U$17204 ( \17887 , \11603 );
not \U$17205 ( \17888 , \8368 );
and \U$17206 ( \17889 , \17887 , \17888 );
and \U$17207 ( \17890 , \11574 , RI992a4c0_383);
nor \U$17208 ( \17891 , \17889 , \17890 );
not \U$17209 ( \17892 , \11599 );
not \U$17210 ( \17893 , \2604 );
and \U$17211 ( \17894 , \17892 , \17893 );
and \U$17212 ( \17895 , \11569 , RI9928d50_403);
nor \U$17213 ( \17896 , \17894 , \17895 );
nand \U$17214 ( \17897 , \17891 , \17896 );
and \U$17215 ( \17898 , \16671 , RI9924d90_503);
not \U$17216 ( \17899 , RI9922540_583);
not \U$17217 ( \17900 , \16609 );
or \U$17218 ( \17901 , \17899 , \17900 );
or \U$17219 ( \17902 , \16676 , \2616 );
nand \U$17220 ( \17903 , \17901 , \17902 );
nor \U$17221 ( \17904 , \17898 , \17903 );
nand \U$17222 ( \17905 , \13976 , \17904 );
nor \U$17223 ( \17906 , \17897 , \17905 );
nand \U$17224 ( \17907 , \17886 , \17906 );
not \U$17225 ( \17908 , \17907 );
not \U$17226 ( \17909 , \17908 );
not \U$17227 ( \17910 , \16642 );
and \U$17228 ( \17911 , \17909 , \17910 );
not \U$17229 ( \17912 , \17909 );
and \U$17230 ( \17913 , \17912 , \16635 );
nor \U$17231 ( \17914 , \17911 , \17913 );
and \U$17232 ( \17915 , \16639 , \17914 );
not \U$17233 ( \17916 , \17781 );
not \U$17234 ( \17917 , \17561 );
or \U$17235 ( \17918 , \17916 , \17917 );
nand \U$17236 ( \17919 , \16765 , \17782 );
nand \U$17237 ( \17920 , \17918 , \17919 );
not \U$17238 ( \17921 , \17920 );
and \U$17239 ( \17922 , \16566 , \16565 , \16571 );
not \U$17240 ( \17923 , \17922 );
or \U$17241 ( \17924 , \17921 , \17923 );
nand \U$17242 ( \17925 , \17794 , \16630 );
nand \U$17243 ( \17926 , \17924 , \17925 );
or \U$17244 ( \17927 , \17915 , \17926 );
xor \U$17245 ( \17928 , \17725 , \17735 );
not \U$17246 ( \17929 , \17424 );
not \U$17247 ( \17930 , \16987 );
or \U$17248 ( \17931 , \17929 , \17930 );
nand \U$17249 ( \17932 , \17061 , \16988 );
nand \U$17250 ( \17933 , \17931 , \17932 );
not \U$17251 ( \17934 , \17933 );
not \U$17252 ( \17935 , \17373 );
or \U$17253 ( \17936 , \17934 , \17935 );
nand \U$17254 ( \17937 , \17711 , \17381 );
nand \U$17255 ( \17938 , \17936 , \17937 );
not \U$17256 ( \17939 , \17938 );
not \U$17257 ( \17940 , \17246 );
xor \U$17258 ( \17941 , \17240 , \17338 );
not \U$17259 ( \17942 , \17941 );
or \U$17260 ( \17943 , \17940 , \17942 );
nand \U$17261 ( \17944 , \17730 , \17236 );
nand \U$17262 ( \17945 , \17943 , \17944 );
not \U$17263 ( \17946 , \17270 );
not \U$17264 ( \17947 , \17273 );
not \U$17265 ( \17948 , \17037 );
or \U$17266 ( \17949 , \17947 , \17948 );
nand \U$17267 ( \17950 , \17038 , \17290 );
nand \U$17268 ( \17951 , \17949 , \17950 );
not \U$17269 ( \17952 , \17951 );
or \U$17270 ( \17953 , \17946 , \17952 );
nand \U$17271 ( \17954 , \17723 , \17285 );
nand \U$17272 ( \17955 , \17953 , \17954 );
nand \U$17273 ( \17956 , \17945 , \17955 );
nand \U$17274 ( \17957 , \17939 , \17956 );
and \U$17275 ( \17958 , \17928 , \17957 );
nor \U$17276 ( \17959 , \17939 , \17956 );
nor \U$17277 ( \17960 , \17958 , \17959 );
not \U$17278 ( \17961 , \17960 );
nand \U$17279 ( \17962 , \17927 , \17961 );
nand \U$17280 ( \17963 , \17926 , \17915 );
and \U$17281 ( \17964 , \17962 , \17963 );
not \U$17282 ( \17965 , \17964 );
not \U$17283 ( \17966 , \17965 );
xor \U$17284 ( \17967 , \17741 , \17787 );
xor \U$17285 ( \17968 , \17967 , \17800 );
not \U$17286 ( \17969 , \17968 );
or \U$17287 ( \17970 , \17966 , \17969 );
or \U$17288 ( \17971 , \17965 , \17968 );
not \U$17289 ( \17972 , \17303 );
not \U$17290 ( \17973 , \17214 );
not \U$17291 ( \17974 , \16995 );
or \U$17292 ( \17975 , \17973 , \17974 );
not \U$17293 ( \17976 , \16995 );
nand \U$17294 ( \17977 , \17976 , \17217 );
nand \U$17295 ( \17978 , \17975 , \17977 );
not \U$17296 ( \17979 , \17978 );
or \U$17297 ( \17980 , \17972 , \17979 );
nand \U$17298 ( \17981 , \17826 , \17118 );
nand \U$17299 ( \17982 , \17980 , \17981 );
not \U$17300 ( \17983 , \17982 );
not \U$17301 ( \17984 , \17816 );
not \U$17302 ( \17985 , \17405 );
or \U$17303 ( \17986 , \17984 , \17985 );
or \U$17304 ( \17987 , \16894 , \17612 );
or \U$17305 ( \17988 , \16742 , \17616 );
nand \U$17306 ( \17989 , \17987 , \17988 );
nand \U$17307 ( \17990 , \17402 , \17989 );
nand \U$17308 ( \17991 , \17986 , \17990 );
not \U$17309 ( \17992 , \17991 );
nand \U$17310 ( \17993 , \17983 , \17992 );
not \U$17311 ( \17994 , \17506 );
not \U$17312 ( \17995 , \16753 );
or \U$17313 ( \17996 , \17994 , \17995 );
nand \U$17314 ( \17997 , \16569 , \17792 );
nand \U$17315 ( \17998 , \17996 , \17997 );
not \U$17316 ( \17999 , \17998 );
not \U$17317 ( \18000 , \16756 );
or \U$17318 ( \18001 , \17999 , \18000 );
nand \U$17319 ( \18002 , \17838 , \16750 );
nand \U$17320 ( \18003 , \18001 , \18002 );
and \U$17321 ( \18004 , \17993 , \18003 );
and \U$17322 ( \18005 , \17991 , \17982 );
nor \U$17323 ( \18006 , \18004 , \18005 );
not \U$17324 ( \18007 , \18006 );
xor \U$17325 ( \18008 , \17843 , \17831 );
and \U$17326 ( \18009 , \18008 , \17845 );
not \U$17327 ( \18010 , \18008 );
and \U$17328 ( \18011 , \18010 , \17818 );
nor \U$17329 ( \18012 , \18009 , \18011 );
not \U$17330 ( \18013 , \18012 );
or \U$17331 ( \18014 , \18007 , \18013 );
xor \U$17332 ( \18015 , \17715 , \17736 );
xor \U$17333 ( \18016 , \18015 , \17738 );
nand \U$17334 ( \18017 , \18014 , \18016 );
not \U$17335 ( \18018 , \18006 );
not \U$17336 ( \18019 , \18012 );
nand \U$17337 ( \18020 , \18018 , \18019 );
nand \U$17338 ( \18021 , \18017 , \18020 );
nand \U$17339 ( \18022 , \17971 , \18021 );
nand \U$17340 ( \18023 , \17970 , \18022 );
not \U$17341 ( \18024 , \18023 );
or \U$17342 ( \18025 , \17864 , \18024 );
or \U$17343 ( \18026 , \18023 , \17863 );
xor \U$17344 ( \18027 , \17803 , \17805 );
xor \U$17345 ( \18028 , \18027 , \17853 );
nand \U$17346 ( \18029 , \18026 , \18028 );
nand \U$17347 ( \18030 , \18025 , \18029 );
not \U$17348 ( \18031 , \18030 );
nand \U$17349 ( \18032 , \17861 , \18031 );
xor \U$17350 ( \18033 , \17808 , \17847 );
xor \U$17351 ( \18034 , \18033 , \17850 );
not \U$17352 ( \18035 , \18034 );
not \U$17353 ( \18036 , \17909 );
not \U$17354 ( \18037 , \17561 );
or \U$17355 ( \18038 , \18036 , \18037 );
nand \U$17356 ( \18039 , \16574 , \17908 );
nand \U$17357 ( \18040 , \18038 , \18039 );
not \U$17358 ( \18041 , \18040 );
not \U$17359 ( \18042 , \17922 );
or \U$17360 ( \18043 , \18041 , \18042 );
nand \U$17361 ( \18044 , \17920 , \16630 );
nand \U$17362 ( \18045 , \18043 , \18044 );
not \U$17363 ( \18046 , \18045 );
not \U$17364 ( \18047 , RI9928378_424);
nor \U$17365 ( \18048 , \18047 , \10812 );
nor \U$17366 ( \18049 , \11559 , \3098 );
nor \U$17367 ( \18050 , \18048 , \18049 );
and \U$17368 ( \18051 , \16643 , RI99313d8_284);
not \U$17369 ( \18052 , RI99224c8_584);
not \U$17370 ( \18053 , \16609 );
or \U$17371 ( \18054 , \18052 , \18053 );
nand \U$17372 ( \18055 , \16605 , RI99230f8_564);
nand \U$17373 ( \18056 , \18054 , \18055 );
nor \U$17374 ( \18057 , \18051 , \18056 );
nand \U$17375 ( \18058 , \16958 , RI9926668_464);
nand \U$17376 ( \18059 , \18050 , \18057 , \18058 );
not \U$17377 ( \18060 , \11599 );
not \U$17378 ( \18061 , RI992f128_304);
not \U$17379 ( \18062 , \18061 );
and \U$17380 ( \18063 , \18060 , \18062 );
and \U$17381 ( \18064 , \11569 , RI9928cd8_404);
nor \U$17382 ( \18065 , \18063 , \18064 );
nand \U$17383 ( \18066 , \18065 , \13933 );
nor \U$17384 ( \18067 , \18059 , \18066 );
not \U$17385 ( \18068 , \11603 );
not \U$17386 ( \18069 , \3104 );
and \U$17387 ( \18070 , \18068 , \18069 );
and \U$17388 ( \18071 , \11576 , RI992ada8_364);
nor \U$17389 ( \18072 , \18070 , \18071 );
not \U$17390 ( \18073 , \11586 );
not \U$17391 ( \18074 , \3118 );
and \U$17392 ( \18075 , \18073 , \18074 );
nor \U$17393 ( \18076 , \11573 , \3115 );
nor \U$17394 ( \18077 , \18075 , \18076 );
nand \U$17395 ( \18078 , \18072 , \18077 );
not \U$17396 ( \18079 , \10823 );
not \U$17397 ( \18080 , \8282 );
and \U$17398 ( \18081 , \18079 , \18080 );
nor \U$17399 ( \18082 , \10862 , \8279 );
nor \U$17400 ( \18083 , \18081 , \18082 );
not \U$17401 ( \18084 , \16590 );
not \U$17402 ( \18085 , \3128 );
and \U$17403 ( \18086 , \18084 , \18085 );
and \U$17404 ( \18087 , \16594 , RI992d238_324);
nor \U$17405 ( \18088 , \18086 , \18087 );
nand \U$17406 ( \18089 , \18083 , \18088 );
nor \U$17407 ( \18090 , \18078 , \18089 );
nand \U$17408 ( \18091 , \18067 , \18090 );
not \U$17409 ( \18092 , \18091 );
not \U$17410 ( \18093 , \18092 );
and \U$17411 ( \18094 , \18093 , \17507 );
not \U$17412 ( \18095 , \18093 );
and \U$17413 ( \18096 , \18095 , \16635 );
nor \U$17414 ( \18097 , \18094 , \18096 );
and \U$17415 ( \18098 , \16639 , \18097 );
not \U$17416 ( \18099 , \18098 );
or \U$17417 ( \18100 , \18046 , \18099 );
or \U$17418 ( \18101 , \18045 , \18098 );
not \U$17419 ( \18102 , \16888 );
not \U$17420 ( \18103 , \17424 );
or \U$17421 ( \18104 , \18102 , \18103 );
nand \U$17422 ( \18105 , \17061 , \17824 );
nand \U$17423 ( \18106 , \18104 , \18105 );
not \U$17424 ( \18107 , \18106 );
not \U$17425 ( \18108 , \17373 );
or \U$17426 ( \18109 , \18107 , \18108 );
nand \U$17427 ( \18110 , \17933 , \17381 );
nand \U$17428 ( \18111 , \18109 , \18110 );
not \U$17429 ( \18112 , \17270 );
xor \U$17430 ( \18113 , \17273 , \16987 );
not \U$17431 ( \18114 , \18113 );
or \U$17432 ( \18115 , \18112 , \18114 );
nand \U$17433 ( \18116 , \17951 , \17285 );
nand \U$17434 ( \18117 , \18115 , \18116 );
not \U$17435 ( \18118 , \17236 );
not \U$17436 ( \18119 , \17941 );
or \U$17437 ( \18120 , \18118 , \18119 );
and \U$17438 ( \18121 , \17110 , \17230 );
not \U$17439 ( \18122 , \17110 );
and \U$17440 ( \18123 , \18122 , \17240 );
or \U$17441 ( \18124 , \18121 , \18123 );
nand \U$17442 ( \18125 , \18124 , \17246 );
nand \U$17443 ( \18126 , \18120 , \18125 );
and \U$17444 ( \18127 , \18117 , \18126 );
xor \U$17445 ( \18128 , \18111 , \18127 );
xor \U$17446 ( \18129 , \17955 , \17945 );
and \U$17447 ( \18130 , \18128 , \18129 );
and \U$17448 ( \18131 , \18111 , \18127 );
or \U$17449 ( \18132 , \18130 , \18131 );
nand \U$17450 ( \18133 , \18101 , \18132 );
nand \U$17451 ( \18134 , \18100 , \18133 );
not \U$17452 ( \18135 , \18134 );
not \U$17453 ( \18136 , \17915 );
not \U$17454 ( \18137 , \17960 );
and \U$17455 ( \18138 , \18136 , \18137 );
and \U$17456 ( \18139 , \17915 , \17960 );
nor \U$17457 ( \18140 , \18138 , \18139 );
not \U$17458 ( \18141 , \17926 );
and \U$17459 ( \18142 , \18140 , \18141 );
not \U$17460 ( \18143 , \18140 );
and \U$17461 ( \18144 , \18143 , \17926 );
nor \U$17462 ( \18145 , \18142 , \18144 );
not \U$17463 ( \18146 , \18145 );
or \U$17464 ( \18147 , \18135 , \18146 );
or \U$17465 ( \18148 , \18134 , \18145 );
xor \U$17466 ( \18149 , \17956 , \17938 );
xnor \U$17467 ( \18150 , \18149 , \17928 );
not \U$17468 ( \18151 , \17781 );
not \U$17469 ( \18152 , \17166 );
or \U$17470 ( \18153 , \18151 , \18152 );
nand \U$17471 ( \18154 , \16569 , \17782 );
nand \U$17472 ( \18155 , \18153 , \18154 );
not \U$17473 ( \18156 , \18155 );
not \U$17474 ( \18157 , \16756 );
or \U$17475 ( \18158 , \18156 , \18157 );
nand \U$17476 ( \18159 , \17998 , \16750 );
nand \U$17477 ( \18160 , \18158 , \18159 );
not \U$17478 ( \18161 , \17164 );
not \U$17479 ( \18162 , \17666 );
or \U$17480 ( \18163 , \18161 , \18162 );
nand \U$17481 ( \18164 , \16944 , \17170 );
nand \U$17482 ( \18165 , \18163 , \18164 );
not \U$17483 ( \18166 , \18165 );
not \U$17484 ( \18167 , \17303 );
or \U$17485 ( \18168 , \18166 , \18167 );
nand \U$17486 ( \18169 , \17978 , \17118 );
nand \U$17487 ( \18170 , \18168 , \18169 );
xor \U$17488 ( \18171 , \18160 , \18170 );
not \U$17489 ( \18172 , \17989 );
not \U$17490 ( \18173 , \17405 );
or \U$17491 ( \18174 , \18172 , \18173 );
and \U$17492 ( \18175 , \17559 , \16890 );
not \U$17493 ( \18176 , \17559 );
and \U$17494 ( \18177 , \18176 , \16894 );
nor \U$17495 ( \18178 , \18175 , \18177 );
nand \U$17496 ( \18179 , \17402 , \18178 );
nand \U$17497 ( \18180 , \18174 , \18179 );
and \U$17498 ( \18181 , \18171 , \18180 );
and \U$17499 ( \18182 , \18160 , \18170 );
or \U$17500 ( \18183 , \18181 , \18182 );
xor \U$17501 ( \18184 , \18150 , \18183 );
xor \U$17502 ( \18185 , \17982 , \18003 );
and \U$17503 ( \18186 , \18185 , \17991 );
not \U$17504 ( \18187 , \18185 );
and \U$17505 ( \18188 , \18187 , \17992 );
nor \U$17506 ( \18189 , \18186 , \18188 );
and \U$17507 ( \18190 , \18184 , \18189 );
and \U$17508 ( \18191 , \18150 , \18183 );
or \U$17509 ( \18192 , \18190 , \18191 );
nand \U$17510 ( \18193 , \18148 , \18192 );
nand \U$17511 ( \18194 , \18147 , \18193 );
not \U$17512 ( \18195 , \18194 );
or \U$17513 ( \18196 , \18035 , \18195 );
or \U$17514 ( \18197 , \18034 , \18194 );
xor \U$17515 ( \18198 , \17964 , \17968 );
xnor \U$17516 ( \18199 , \18198 , \18021 );
nand \U$17517 ( \18200 , \18197 , \18199 );
nand \U$17518 ( \18201 , \18196 , \18200 );
not \U$17519 ( \18202 , \18201 );
xor \U$17520 ( \18203 , \17863 , \18023 );
xnor \U$17521 ( \18204 , \18203 , \18028 );
nand \U$17522 ( \18205 , \18202 , \18204 );
and \U$17523 ( \18206 , \18032 , \18205 );
not \U$17524 ( \18207 , \17379 );
not \U$17525 ( \18208 , \17373 );
or \U$17526 ( \18209 , \18207 , \18208 );
and \U$17527 ( \18210 , \17057 , \16682 );
not \U$17528 ( \18211 , \17057 );
and \U$17529 ( \18212 , \18211 , \16683 );
nor \U$17530 ( \18213 , \18210 , \18212 );
nand \U$17531 ( \18214 , \18213 , \17381 );
nand \U$17532 ( \18215 , \18209 , \18214 );
not \U$17533 ( \18216 , \18215 );
not \U$17534 ( \18217 , \17294 );
or \U$17535 ( \18218 , \18217 , \17269 );
or \U$17536 ( \18219 , \17268 , \17290 );
nand \U$17537 ( \18220 , \18218 , \18219 );
xor \U$17538 ( \18221 , \18216 , \18220 );
and \U$17539 ( \18222 , \18221 , \17387 );
and \U$17540 ( \18223 , \18216 , \18220 );
or \U$17541 ( \18224 , \18222 , \18223 );
not \U$17542 ( \18225 , \17397 );
not \U$17543 ( \18226 , \16758 );
or \U$17544 ( \18227 , \18225 , \18226 );
not \U$17545 ( \18228 , \16989 );
not \U$17546 ( \18229 , \17395 );
or \U$17547 ( \18230 , \18228 , \18229 );
not \U$17548 ( \18231 , \16753 );
nand \U$17549 ( \18232 , \18231 , \16988 );
nand \U$17550 ( \18233 , \18230 , \18232 );
nand \U$17551 ( \18234 , \18233 , \16750 );
nand \U$17552 ( \18235 , \18227 , \18234 );
not \U$17553 ( \18236 , \17344 );
not \U$17554 ( \18237 , \17303 );
or \U$17555 ( \18238 , \18236 , \18237 );
not \U$17556 ( \18239 , \16824 );
not \U$17557 ( \18240 , \17666 );
or \U$17558 ( \18241 , \18239 , \18240 );
nand \U$17559 ( \18242 , \16944 , \16825 );
nand \U$17560 ( \18243 , \18241 , \18242 );
nand \U$17561 ( \18244 , \18243 , \17118 );
nand \U$17562 ( \18245 , \18238 , \18244 );
xor \U$17563 ( \18246 , \18235 , \18245 );
not \U$17564 ( \18247 , \17410 );
not \U$17565 ( \18248 , \17402 );
or \U$17566 ( \18249 , \18247 , \18248 );
and \U$17567 ( \18250 , \17112 , \16893 );
not \U$17568 ( \18251 , \17112 );
and \U$17569 ( \18252 , \18251 , \16894 );
nor \U$17570 ( \18253 , \18250 , \18252 );
nand \U$17571 ( \18254 , \17405 , \18253 );
nand \U$17572 ( \18255 , \18249 , \18254 );
and \U$17573 ( \18256 , \18246 , \18255 );
and \U$17574 ( \18257 , \18235 , \18245 );
or \U$17575 ( \18258 , \18256 , \18257 );
xor \U$17576 ( \18259 , \18224 , \18258 );
not \U$17577 ( \18260 , \18233 );
not \U$17578 ( \18261 , \17390 );
or \U$17579 ( \18262 , \18260 , \18261 );
not \U$17580 ( \18263 , \16749 );
not \U$17581 ( \18264 , \17406 );
not \U$17582 ( \18265 , \17166 );
or \U$17583 ( \18266 , \18264 , \18265 );
not \U$17584 ( \18267 , \17406 );
nand \U$17585 ( \18268 , \16569 , \18267 );
nand \U$17586 ( \18269 , \18266 , \18268 );
nand \U$17587 ( \18270 , \18263 , \18269 );
nand \U$17588 ( \18271 , \18262 , \18270 );
not \U$17589 ( \18272 , \18243 );
not \U$17590 ( \18273 , \17303 );
or \U$17591 ( \18274 , \18272 , \18273 );
and \U$17592 ( \18275 , \16732 , \17666 );
not \U$17593 ( \18276 , \16732 );
and \U$17594 ( \18277 , \18276 , \16944 );
nor \U$17595 ( \18278 , \18275 , \18277 );
nand \U$17596 ( \18279 , \18278 , \17118 );
nand \U$17597 ( \18280 , \18274 , \18279 );
xor \U$17598 ( \18281 , \18271 , \18280 );
not \U$17599 ( \18282 , \18253 );
not \U$17600 ( \18283 , \17402 );
or \U$17601 ( \18284 , \18282 , \18283 );
and \U$17602 ( \18285 , \17338 , \16893 );
not \U$17603 ( \18286 , \17338 );
and \U$17604 ( \18287 , \18286 , \16889 );
nor \U$17605 ( \18288 , \18285 , \18287 );
nand \U$17606 ( \18289 , \17405 , \18288 );
nand \U$17607 ( \18290 , \18284 , \18289 );
xor \U$17608 ( \18291 , \18281 , \18290 );
xor \U$17609 ( \18292 , \18259 , \18291 );
not \U$17610 ( \18293 , \17413 );
nand \U$17611 ( \18294 , \17224 , \17350 );
not \U$17612 ( \18295 , \18294 );
or \U$17613 ( \18296 , \18293 , \18295 );
nand \U$17614 ( \18297 , \17225 , \17351 );
nand \U$17615 ( \18298 , \18296 , \18297 );
xor \U$17616 ( \18299 , \17638 , \17644 );
and \U$17617 ( \18300 , \18299 , \17657 );
and \U$17618 ( \18301 , \17638 , \17644 );
or \U$17619 ( \18302 , \18300 , \18301 );
xor \U$17620 ( \18303 , \18298 , \18302 );
nor \U$17621 ( \18304 , \17346 , \17299 );
or \U$17622 ( \18305 , \18304 , \17288 );
nand \U$17623 ( \18306 , \17346 , \17299 );
nand \U$17624 ( \18307 , \18305 , \18306 );
not \U$17625 ( \18308 , \17616 );
not \U$17626 ( \18309 , \16642 );
or \U$17627 ( \18310 , \18308 , \18309 );
nand \U$17628 ( \18311 , \16685 , \17612 );
nand \U$17629 ( \18312 , \18310 , \18311 );
nor \U$17630 ( \18313 , \16640 , \18312 );
xor \U$17631 ( \18314 , \18307 , \18313 );
not \U$17632 ( \18315 , \17655 );
not \U$17633 ( \18316 , \16572 );
or \U$17634 ( \18317 , \18315 , \18316 );
not \U$17635 ( \18318 , \16626 );
not \U$17636 ( \18319 , \17214 );
or \U$17637 ( \18320 , \18318 , \18319 );
nand \U$17638 ( \18321 , \16765 , \17217 );
nand \U$17639 ( \18322 , \18320 , \18321 );
nand \U$17640 ( \18323 , \18322 , \16630 );
nand \U$17641 ( \18324 , \18317 , \18323 );
xor \U$17642 ( \18325 , \18314 , \18324 );
and \U$17643 ( \18326 , \18303 , \18325 );
and \U$17644 ( \18327 , \18298 , \18302 );
or \U$17645 ( \18328 , \18326 , \18327 );
xor \U$17646 ( \18329 , \18292 , \18328 );
xor \U$17647 ( \18330 , \18307 , \18313 );
and \U$17648 ( \18331 , \18330 , \18324 );
and \U$17649 ( \18332 , \18307 , \18313 );
or \U$17650 ( \18333 , \18331 , \18332 );
not \U$17651 ( \18334 , \17268 );
not \U$17652 ( \18335 , \17269 );
or \U$17653 ( \18336 , \18334 , \18335 );
nand \U$17654 ( \18337 , \18336 , \17273 );
xor \U$17655 ( \18338 , \18337 , \18215 );
buf \U$17656 ( \18339 , \17373 );
not \U$17657 ( \18340 , \18339 );
not \U$17658 ( \18341 , \18213 );
or \U$17659 ( \18342 , \18340 , \18341 );
and \U$17660 ( \18343 , \16624 , \17061 );
not \U$17661 ( \18344 , \16624 );
and \U$17662 ( \18345 , \18344 , \17062 );
nor \U$17663 ( \18346 , \18343 , \18345 );
or \U$17664 ( \18347 , \18346 , \17380 );
nand \U$17665 ( \18348 , \18342 , \18347 );
xor \U$17666 ( \18349 , \18338 , \18348 );
not \U$17667 ( \18350 , \18322 );
not \U$17668 ( \18351 , \16572 );
or \U$17669 ( \18352 , \18350 , \18351 );
and \U$17670 ( \18353 , \17824 , \16626 );
not \U$17671 ( \18354 , \17824 );
and \U$17672 ( \18355 , \18354 , \16765 );
nor \U$17673 ( \18356 , \18353 , \18355 );
nand \U$17674 ( \18357 , \18356 , \16630 );
nand \U$17675 ( \18358 , \18352 , \18357 );
xor \U$17676 ( \18359 , \18349 , \18358 );
and \U$17677 ( \18360 , \16642 , \17170 );
and \U$17678 ( \18361 , \17639 , \17164 );
nor \U$17679 ( \18362 , \18360 , \18361 );
and \U$17680 ( \18363 , \16641 , \18362 );
xor \U$17681 ( \18364 , \18359 , \18363 );
xor \U$17682 ( \18365 , \18333 , \18364 );
xor \U$17683 ( \18366 , \18216 , \18220 );
xor \U$17684 ( \18367 , \18366 , \17387 );
xor \U$17685 ( \18368 , \17388 , \17399 );
and \U$17686 ( \18369 , \18368 , \17412 );
and \U$17687 ( \18370 , \17388 , \17399 );
or \U$17688 ( \18371 , \18369 , \18370 );
xor \U$17689 ( \18372 , \18367 , \18371 );
xor \U$17690 ( \18373 , \18235 , \18245 );
xor \U$17691 ( \18374 , \18373 , \18255 );
and \U$17692 ( \18375 , \18372 , \18374 );
and \U$17693 ( \18376 , \18367 , \18371 );
or \U$17694 ( \18377 , \18375 , \18376 );
xor \U$17695 ( \18378 , \18365 , \18377 );
xor \U$17696 ( \18379 , \18329 , \18378 );
xor \U$17697 ( \18380 , \18367 , \18371 );
xor \U$17698 ( \18381 , \18380 , \18374 );
xor \U$17699 ( \18382 , \17623 , \17658 );
and \U$17700 ( \18383 , \18382 , \17701 );
and \U$17701 ( \18384 , \17623 , \17658 );
or \U$17702 ( \18385 , \18383 , \18384 );
xor \U$17703 ( \18386 , \18381 , \18385 );
xor \U$17704 ( \18387 , \18298 , \18302 );
xor \U$17705 ( \18388 , \18387 , \18325 );
and \U$17706 ( \18389 , \18386 , \18388 );
and \U$17707 ( \18390 , \18381 , \18385 );
or \U$17708 ( \18391 , \18389 , \18390 );
nor \U$17709 ( \18392 , \18379 , \18391 );
xor \U$17710 ( \18393 , \18381 , \18385 );
xor \U$17711 ( \18394 , \18393 , \18388 );
not \U$17712 ( \18395 , \17414 );
not \U$17713 ( \18396 , \17857 );
or \U$17714 ( \18397 , \18395 , \18396 );
nand \U$17715 ( \18398 , \18397 , \17702 );
not \U$17716 ( \18399 , \17414 );
nand \U$17717 ( \18400 , \18399 , \17856 );
nand \U$17718 ( \18401 , \18398 , \18400 );
nor \U$17719 ( \18402 , \18394 , \18401 );
nor \U$17720 ( \18403 , \18392 , \18402 );
and \U$17721 ( \18404 , \18206 , \18403 );
not \U$17722 ( \18405 , \18404 );
not \U$17723 ( \18406 , \17612 );
not \U$17724 ( \18407 , \17062 );
or \U$17725 ( \18408 , \18406 , \18407 );
nand \U$17726 ( \18409 , \17061 , \17616 );
nand \U$17727 ( \18410 , \18408 , \18409 );
not \U$17728 ( \18411 , \18410 );
not \U$17729 ( \18412 , \17373 );
or \U$17730 ( \18413 , \18411 , \18412 );
and \U$17731 ( \18414 , \17163 , \17424 );
not \U$17732 ( \18415 , \17163 );
and \U$17733 ( \18416 , \18415 , \17061 );
nor \U$17734 ( \18417 , \18414 , \18416 );
or \U$17735 ( \18418 , \18417 , \17380 );
nand \U$17736 ( \18419 , \18413 , \18418 );
not \U$17737 ( \18420 , \17285 );
and \U$17738 ( \18421 , \17290 , \17824 );
not \U$17739 ( \18422 , \17290 );
and \U$17740 ( \18423 , \18422 , \16888 );
nor \U$17741 ( \18424 , \18421 , \18423 );
not \U$17742 ( \18425 , \18424 );
or \U$17743 ( \18426 , \18420 , \18425 );
xor \U$17744 ( \18427 , \17273 , \17213 );
nand \U$17745 ( \18428 , \18427 , \17270 );
nand \U$17746 ( \18429 , \18426 , \18428 );
xor \U$17747 ( \18430 , \17240 , \16987 );
and \U$17748 ( \18431 , \18430 , \17246 );
not \U$17749 ( \18432 , \17240 );
not \U$17750 ( \18433 , \17037 );
or \U$17751 ( \18434 , \18432 , \18433 );
nand \U$17752 ( \18435 , \17038 , \17230 );
nand \U$17753 ( \18436 , \18434 , \18435 );
and \U$17754 ( \18437 , \18436 , \17236 );
nor \U$17755 ( \18438 , \18431 , \18437 );
xor \U$17756 ( \18439 , \18429 , \18438 );
xor \U$17757 ( \18440 , \18419 , \18439 );
not \U$17758 ( \18441 , \16558 );
nand \U$17759 ( \18442 , \16564 , \16570 );
not \U$17760 ( \18443 , \11599 );
not \U$17761 ( \18444 , \8675 );
and \U$17762 ( \18445 , \18443 , \18444 );
and \U$17763 ( \18446 , \16801 , RI992ac40_367);
nor \U$17764 ( \18447 , \18445 , \18446 );
not \U$17765 ( \18448 , \10794 );
not \U$17766 ( \18449 , \3550 );
and \U$17767 ( \18450 , \18448 , \18449 );
and \U$17768 ( \18451 , \11569 , RI9928b70_407);
nor \U$17769 ( \18452 , \18450 , \18451 );
and \U$17770 ( \18453 , \16671 , RI9924bb0_507);
not \U$17771 ( \18454 , RI9922360_587);
not \U$17772 ( \18455 , \16609 );
or \U$17773 ( \18456 , \18454 , \18455 );
or \U$17774 ( \18457 , \16676 , \8659 );
nand \U$17775 ( \18458 , \18456 , \18457 );
nor \U$17776 ( \18459 , \18453 , \18458 );
nand \U$17777 ( \18460 , \18447 , \18452 , \14267 , \18459 );
not \U$17778 ( \18461 , \18460 );
not \U$17779 ( \18462 , \10849 );
not \U$17780 ( \18463 , \8642 );
and \U$17781 ( \18464 , \18462 , \18463 );
nor \U$17782 ( \18465 , \10885 , \8672 );
nor \U$17783 ( \18466 , \18464 , \18465 );
nor \U$17784 ( \18467 , \11563 , \8655 );
nor \U$17785 ( \18468 , \16590 , \8639 );
nor \U$17786 ( \18469 , \18467 , \18468 );
nand \U$17787 ( \18470 , \16656 , RI9924250_527);
nand \U$17788 ( \18471 , \18466 , \18469 , \18470 );
not \U$17789 ( \18472 , \11586 );
not \U$17790 ( \18473 , \8682 );
and \U$17791 ( \18474 , \18472 , \18473 );
and \U$17792 ( \18475 , \10931 , RI9926e60_447);
nor \U$17793 ( \18476 , \18474 , \18475 );
nor \U$17794 ( \18477 , \11603 , \8662 );
nor \U$17795 ( \18478 , \16581 , \8679 );
nor \U$17796 ( \18479 , \18477 , \18478 );
nand \U$17797 ( \18480 , \18476 , \18479 );
nor \U$17798 ( \18481 , \18471 , \18480 );
nand \U$17799 ( \18482 , \18461 , \18481 );
buf \U$17800 ( \18483 , \18482 );
and \U$17801 ( \18484 , \18442 , \18483 );
and \U$17802 ( \18485 , \16563 , \17169 );
nor \U$17803 ( \18486 , \18484 , \18485 );
nand \U$17804 ( \18487 , \18441 , \18486 );
xnor \U$17805 ( \18488 , \18440 , \18487 );
or \U$17806 ( \18489 , \16894 , \18093 );
or \U$17807 ( \18490 , \16893 , \18092 );
nand \U$17808 ( \18491 , \18489 , \18490 );
not \U$17809 ( \18492 , \18491 );
not \U$17810 ( \18493 , \17402 );
or \U$17811 ( \18494 , \18492 , \18493 );
and \U$17812 ( \18495 , \17909 , \16893 );
not \U$17813 ( \18496 , \17909 );
and \U$17814 ( \18497 , \18496 , \16894 );
nor \U$17815 ( \18498 , \18495 , \18497 );
nand \U$17816 ( \18499 , \17405 , \18498 );
nand \U$17817 ( \18500 , \18494 , \18499 );
not \U$17818 ( \18501 , \16758 );
not \U$17819 ( \18502 , \11559 );
not \U$17820 ( \18503 , \8539 );
and \U$17821 ( \18504 , \18502 , \18503 );
nor \U$17822 ( \18505 , \11563 , \8542 );
nor \U$17823 ( \18506 , \18504 , \18505 );
and \U$17824 ( \18507 , \16643 , RI99312e8_286);
not \U$17825 ( \18508 , RI99223d8_586);
not \U$17826 ( \18509 , \16609 );
or \U$17827 ( \18510 , \18508 , \18509 );
or \U$17828 ( \18511 , \16676 , \3683 );
nand \U$17829 ( \18512 , \18510 , \18511 );
nor \U$17830 ( \18513 , \18507 , \18512 );
nand \U$17831 ( \18514 , \16958 , RI9926578_466);
nand \U$17832 ( \18515 , \18506 , \18513 , \18514 );
and \U$17833 ( \18516 , \11030 , RI992f038_306);
and \U$17834 ( \18517 , \11569 , RI9928be8_406);
nor \U$17835 ( \18518 , \18516 , \18517 );
nand \U$17836 ( \18519 , \18518 , \14160 );
nor \U$17837 ( \18520 , \18515 , \18519 );
not \U$17838 ( \18521 , \11586 );
not \U$17839 ( \18522 , \8535 );
and \U$17840 ( \18523 , \18521 , \18522 );
and \U$17841 ( \18524 , \16801 , RI992acb8_366);
nor \U$17842 ( \18525 , \18523 , \18524 );
and \U$17843 ( \18526 , \11574 , RI992a358_386);
and \U$17844 ( \18527 , \11604 , RI9925c18_486);
nor \U$17845 ( \18528 , \18526 , \18527 );
nand \U$17846 ( \18529 , \18525 , \18528 );
and \U$17847 ( \18530 , \16656 , RI99242c8_526);
nor \U$17848 ( \18531 , \10862 , \14130 );
nor \U$17849 ( \18532 , \18530 , \18531 );
and \U$17850 ( \18533 , \11582 , RI992c7e8_346);
and \U$17851 ( \18534 , \16594 , RI992d148_326);
nor \U$17852 ( \18535 , \18533 , \18534 );
nand \U$17853 ( \18536 , \18532 , \18535 );
nor \U$17854 ( \18537 , \18529 , \18536 );
nand \U$17855 ( \18538 , \18520 , \18537 );
not \U$17856 ( \18539 , \18538 );
not \U$17857 ( \18540 , \18539 );
not \U$17858 ( \18541 , \18540 );
not \U$17859 ( \18542 , \17395 );
or \U$17860 ( \18543 , \18541 , \18542 );
nand \U$17861 ( \18544 , \16569 , \18539 );
nand \U$17862 ( \18545 , \18543 , \18544 );
not \U$17863 ( \18546 , \18545 );
or \U$17864 ( \18547 , \18501 , \18546 );
not \U$17865 ( \18548 , \11603 );
not \U$17866 ( \18549 , \3487 );
and \U$17867 ( \18550 , \18548 , \18549 );
and \U$17868 ( \18551 , \16801 , RI992ad30_365);
nor \U$17869 ( \18552 , \18550 , \18551 );
and \U$17870 ( \18553 , \11574 , RI992a3d0_385);
and \U$17871 ( \18554 , \16654 , RI99239e0_545);
nor \U$17872 ( \18555 , \18553 , \18554 );
nand \U$17873 ( \18556 , \18552 , \18555 );
not \U$17874 ( \18557 , \10823 );
not \U$17875 ( \18558 , \8262 );
and \U$17876 ( \18559 , \18557 , \18558 );
nor \U$17877 ( \18560 , \10862 , \8265 );
nor \U$17878 ( \18561 , \18559 , \18560 );
not \U$17879 ( \18562 , \16590 );
not \U$17880 ( \18563 , \3498 );
and \U$17881 ( \18564 , \18562 , \18563 );
and \U$17882 ( \18565 , \16594 , RI992d1c0_325);
nor \U$17883 ( \18566 , \18564 , \18565 );
nand \U$17884 ( \18567 , \18561 , \18566 );
nor \U$17885 ( \18568 , \18556 , \18567 );
not \U$17886 ( \18569 , \11559 );
not \U$17887 ( \18570 , \8237 );
and \U$17888 ( \18571 , \18569 , \18570 );
nor \U$17889 ( \18572 , \10812 , \8240 );
nor \U$17890 ( \18573 , \18571 , \18572 );
and \U$17891 ( \18574 , \16643 , RI9931360_285);
not \U$17892 ( \18575 , RI9922450_585);
not \U$17893 ( \18576 , \16609 );
or \U$17894 ( \18577 , \18575 , \18576 );
or \U$17895 ( \18578 , \16676 , \3465 );
nand \U$17896 ( \18579 , \18577 , \18578 );
nor \U$17897 ( \18580 , \18574 , \18579 );
nand \U$17898 ( \18581 , \16958 , RI99265f0_465);
nand \U$17899 ( \18582 , \18573 , \18580 , \18581 );
not \U$17900 ( \18583 , \11599 );
not \U$17901 ( \18584 , \3472 );
and \U$17902 ( \18585 , \18583 , \18584 );
and \U$17903 ( \18586 , \16619 , RI9928c60_405);
nor \U$17904 ( \18587 , \18585 , \18586 );
nand \U$17905 ( \18588 , \18587 , \13893 );
nor \U$17906 ( \18589 , \18582 , \18588 );
nand \U$17907 ( \18590 , \18568 , \18589 );
buf \U$17908 ( \18591 , \18590 );
not \U$17909 ( \18592 , \18591 );
not \U$17910 ( \18593 , \17395 );
or \U$17911 ( \18594 , \18592 , \18593 );
not \U$17912 ( \18595 , \18591 );
nand \U$17913 ( \18596 , \16569 , \18595 );
nand \U$17914 ( \18597 , \18594 , \18596 );
nand \U$17915 ( \18598 , \18597 , \16750 );
nand \U$17916 ( \18599 , \18547 , \18598 );
or \U$17917 ( \18600 , \18500 , \18599 );
not \U$17918 ( \18601 , \17236 );
not \U$17919 ( \18602 , \18430 );
or \U$17920 ( \18603 , \18601 , \18602 );
and \U$17921 ( \18604 , \17240 , \16888 );
not \U$17922 ( \18605 , \17240 );
and \U$17923 ( \18606 , \18605 , \17824 );
nor \U$17924 ( \18607 , \18604 , \18606 );
nand \U$17925 ( \18608 , \18607 , \17246 );
nand \U$17926 ( \18609 , \18603 , \18608 );
not \U$17927 ( \18610 , \17285 );
not \U$17928 ( \18611 , \18427 );
or \U$17929 ( \18612 , \18610 , \18611 );
and \U$17930 ( \18613 , \17273 , \17163 );
not \U$17931 ( \18614 , \17273 );
not \U$17932 ( \18615 , \17163 );
and \U$17933 ( \18616 , \18614 , \18615 );
nor \U$17934 ( \18617 , \18613 , \18616 );
nand \U$17935 ( \18618 , \18617 , \17270 );
nand \U$17936 ( \18619 , \18612 , \18618 );
xor \U$17937 ( \18620 , \18609 , \18619 );
not \U$17938 ( \18621 , \17559 );
not \U$17939 ( \18622 , \17062 );
or \U$17940 ( \18623 , \18621 , \18622 );
nand \U$17941 ( \18624 , \17057 , \17564 );
nand \U$17942 ( \18625 , \18623 , \18624 );
not \U$17943 ( \18626 , \18625 );
not \U$17944 ( \18627 , \17373 );
or \U$17945 ( \18628 , \18626 , \18627 );
nand \U$17946 ( \18629 , \18410 , \17381 );
nand \U$17947 ( \18630 , \18628 , \18629 );
xor \U$17948 ( \18631 , \18620 , \18630 );
nand \U$17949 ( \18632 , \18600 , \18631 );
nand \U$17950 ( \18633 , \18500 , \18599 );
and \U$17951 ( \18634 , \18632 , \18633 );
xor \U$17952 ( \18635 , \18488 , \18634 );
xor \U$17953 ( \18636 , \18609 , \18619 );
and \U$17954 ( \18637 , \18636 , \18630 );
and \U$17955 ( \18638 , \18609 , \18619 );
or \U$17956 ( \18639 , \18637 , \18638 );
not \U$17957 ( \18640 , \17303 );
not \U$17958 ( \18641 , \17506 );
not \U$17959 ( \18642 , \17666 );
or \U$17960 ( \18643 , \18641 , \18642 );
nand \U$17961 ( \18644 , \16944 , \17792 );
nand \U$17962 ( \18645 , \18643 , \18644 );
not \U$17963 ( \18646 , \18645 );
or \U$17964 ( \18647 , \18640 , \18646 );
not \U$17965 ( \18648 , \17559 );
not \U$17966 ( \18649 , \16995 );
or \U$17967 ( \18650 , \18648 , \18649 );
nand \U$17968 ( \18651 , \16944 , \17564 );
nand \U$17969 ( \18652 , \18650 , \18651 );
nand \U$17970 ( \18653 , \18652 , \17118 );
nand \U$17971 ( \18654 , \18647 , \18653 );
xor \U$17972 ( \18655 , \18639 , \18654 );
not \U$17973 ( \18656 , \18597 );
not \U$17974 ( \18657 , \16758 );
or \U$17975 ( \18658 , \18656 , \18657 );
and \U$17976 ( \18659 , \18093 , \17169 );
not \U$17977 ( \18660 , \18093 );
and \U$17978 ( \18661 , \18660 , \17395 );
nor \U$17979 ( \18662 , \18659 , \18661 );
nand \U$17980 ( \18663 , \18662 , \16750 );
nand \U$17981 ( \18664 , \18658 , \18663 );
xnor \U$17982 ( \18665 , \18655 , \18664 );
and \U$17983 ( \18666 , \18635 , \18665 );
and \U$17984 ( \18667 , \18488 , \18634 );
or \U$17985 ( \18668 , \18666 , \18667 );
not \U$17986 ( \18669 , \18668 );
not \U$17987 ( \18670 , \18498 );
not \U$17988 ( \18671 , \17402 );
or \U$17989 ( \18672 , \18670 , \18671 );
and \U$17990 ( \18673 , \17781 , \16893 );
not \U$17991 ( \18674 , \17781 );
and \U$17992 ( \18675 , \18674 , \16889 );
nor \U$17993 ( \18676 , \18673 , \18675 );
nand \U$17994 ( \18677 , \17405 , \18676 );
nand \U$17995 ( \18678 , \18672 , \18677 );
not \U$17996 ( \18679 , \18678 );
not \U$17997 ( \18680 , \18679 );
and \U$17998 ( \18681 , \18483 , \16574 );
not \U$17999 ( \18682 , \18483 );
and \U$18000 ( \18683 , \18682 , \16558 );
nor \U$18001 ( \18684 , \18681 , \18683 );
not \U$18002 ( \18685 , \18684 );
not \U$18003 ( \18686 , \17922 );
or \U$18004 ( \18687 , \18685 , \18686 );
and \U$18005 ( \18688 , \18540 , \16574 );
not \U$18006 ( \18689 , \18540 );
and \U$18007 ( \18690 , \18689 , \17561 );
nor \U$18008 ( \18691 , \18688 , \18690 );
nand \U$18009 ( \18692 , \18691 , \16630 );
nand \U$18010 ( \18693 , \18687 , \18692 );
not \U$18011 ( \18694 , \18693 );
not \U$18012 ( \18695 , \18694 );
or \U$18013 ( \18696 , \18680 , \18695 );
or \U$18014 ( \18697 , \16744 , \16893 );
nand \U$18015 ( \18698 , \18697 , \18483 );
nand \U$18016 ( \18699 , \16744 , \16742 );
and \U$18017 ( \18700 , \16569 , \18698 , \18699 );
not \U$18018 ( \18701 , \17246 );
xor \U$18019 ( \18702 , \17240 , \17213 );
not \U$18020 ( \18703 , \18702 );
or \U$18021 ( \18704 , \18701 , \18703 );
nand \U$18022 ( \18705 , \18607 , \17236 );
nand \U$18023 ( \18706 , \18704 , \18705 );
nand \U$18024 ( \18707 , \18700 , \18706 );
nand \U$18025 ( \18708 , \16630 , \18483 );
xor \U$18026 ( \18709 , \18707 , \18708 );
not \U$18027 ( \18710 , \17781 );
not \U$18028 ( \18711 , \17666 );
or \U$18029 ( \18712 , \18710 , \18711 );
not \U$18030 ( \18713 , \16995 );
nand \U$18031 ( \18714 , \18713 , \17782 );
nand \U$18032 ( \18715 , \18712 , \18714 );
and \U$18033 ( \18716 , \18715 , \17303 );
not \U$18034 ( \18717 , \18645 );
not \U$18035 ( \18718 , \17118 );
nor \U$18036 ( \18719 , \18717 , \18718 );
nor \U$18037 ( \18720 , \18716 , \18719 );
and \U$18038 ( \18721 , \18709 , \18720 );
and \U$18039 ( \18722 , \18707 , \18708 );
or \U$18040 ( \18723 , \18721 , \18722 );
not \U$18041 ( \18724 , \18723 );
nand \U$18042 ( \18725 , \18696 , \18724 );
nand \U$18043 ( \18726 , \18693 , \18678 );
nand \U$18044 ( \18727 , \18725 , \18726 );
not \U$18045 ( \18728 , \18727 );
and \U$18046 ( \18729 , \18669 , \18728 );
and \U$18047 ( \18730 , \18668 , \18727 );
nor \U$18048 ( \18731 , \18729 , \18730 );
not \U$18049 ( \18732 , \17246 );
not \U$18050 ( \18733 , \18436 );
or \U$18051 ( \18734 , \18732 , \18733 );
nand \U$18052 ( \18735 , \18124 , \17236 );
nand \U$18053 ( \18736 , \18734 , \18735 );
not \U$18054 ( \18737 , \17270 );
not \U$18055 ( \18738 , \18424 );
or \U$18056 ( \18739 , \18737 , \18738 );
nand \U$18057 ( \18740 , \18113 , \17285 );
nand \U$18058 ( \18741 , \18739 , \18740 );
xor \U$18059 ( \18742 , \18736 , \18741 );
or \U$18060 ( \18743 , \18412 , \18417 );
and \U$18061 ( \18744 , \17213 , \17057 );
not \U$18062 ( \18745 , \17213 );
and \U$18063 ( \18746 , \18745 , \17062 );
nor \U$18064 ( \18747 , \18744 , \18746 );
not \U$18065 ( \18748 , \18747 );
or \U$18066 ( \18749 , \18748 , \17380 );
nand \U$18067 ( \18750 , \18743 , \18749 );
xor \U$18068 ( \18751 , \18742 , \18750 );
not \U$18069 ( \18752 , \18662 );
not \U$18070 ( \18753 , \16758 );
or \U$18071 ( \18754 , \18752 , \18753 );
not \U$18072 ( \18755 , \17909 );
not \U$18073 ( \18756 , \17166 );
or \U$18074 ( \18757 , \18755 , \18756 );
nand \U$18075 ( \18758 , \17169 , \17908 );
nand \U$18076 ( \18759 , \18757 , \18758 );
nand \U$18077 ( \18760 , \18759 , \16750 );
nand \U$18078 ( \18761 , \18754 , \18760 );
xor \U$18079 ( \18762 , \18751 , \18761 );
not \U$18080 ( \18763 , \18676 );
not \U$18081 ( \18764 , \17402 );
or \U$18082 ( \18765 , \18763 , \18764 );
and \U$18083 ( \18766 , \17506 , \16893 );
not \U$18084 ( \18767 , \17506 );
and \U$18085 ( \18768 , \18767 , \16889 );
nor \U$18086 ( \18769 , \18766 , \18768 );
nand \U$18087 ( \18770 , \17405 , \18769 );
nand \U$18088 ( \18771 , \18765 , \18770 );
xor \U$18089 ( \18772 , \18762 , \18771 );
not \U$18090 ( \18773 , \18429 );
nor \U$18091 ( \18774 , \18773 , \18438 );
not \U$18092 ( \18775 , \18652 );
not \U$18093 ( \18776 , \17303 );
or \U$18094 ( \18777 , \18775 , \18776 );
not \U$18095 ( \18778 , \17612 );
not \U$18096 ( \18779 , \17666 );
or \U$18097 ( \18780 , \18778 , \18779 );
nand \U$18098 ( \18781 , \16944 , \17616 );
nand \U$18099 ( \18782 , \18780 , \18781 );
nand \U$18100 ( \18783 , \17118 , \18782 );
nand \U$18101 ( \18784 , \18777 , \18783 );
xor \U$18102 ( \18785 , \18774 , \18784 );
not \U$18103 ( \18786 , \18483 );
nor \U$18104 ( \18787 , \16638 , \18786 );
xor \U$18105 ( \18788 , \18785 , \18787 );
xor \U$18106 ( \18789 , \18772 , \18788 );
not \U$18107 ( \18790 , \18691 );
not \U$18108 ( \18791 , \17922 );
or \U$18109 ( \18792 , \18790 , \18791 );
and \U$18110 ( \18793 , \18591 , \16765 );
not \U$18111 ( \18794 , \18591 );
and \U$18112 ( \18795 , \18794 , \17561 );
nor \U$18113 ( \18796 , \18793 , \18795 );
nand \U$18114 ( \18797 , \18796 , \16630 );
nand \U$18115 ( \18798 , \18792 , \18797 );
not \U$18116 ( \18799 , \18419 );
not \U$18117 ( \18800 , \18799 );
not \U$18118 ( \18801 , \18487 );
or \U$18119 ( \18802 , \18800 , \18801 );
not \U$18120 ( \18803 , \18439 );
nand \U$18121 ( \18804 , \18802 , \18803 );
not \U$18122 ( \18805 , \18487 );
nand \U$18123 ( \18806 , \18805 , \18419 );
nand \U$18124 ( \18807 , \18804 , \18806 );
xor \U$18125 ( \18808 , \18798 , \18807 );
not \U$18126 ( \18809 , \18654 );
not \U$18127 ( \18810 , \18664 );
or \U$18128 ( \18811 , \18809 , \18810 );
or \U$18129 ( \18812 , \18664 , \18654 );
nand \U$18130 ( \18813 , \18812 , \18639 );
nand \U$18131 ( \18814 , \18811 , \18813 );
xor \U$18132 ( \18815 , \18808 , \18814 );
xor \U$18133 ( \18816 , \18789 , \18815 );
xor \U$18134 ( \18817 , \18731 , \18816 );
xor \U$18135 ( \18818 , \18678 , \18693 );
xor \U$18136 ( \18819 , \18818 , \18723 );
xnor \U$18137 ( \18820 , \18700 , \18706 );
and \U$18138 ( \18821 , \17505 , \17424 );
not \U$18139 ( \18822 , \17505 );
and \U$18140 ( \18823 , \18822 , \17057 );
nor \U$18141 ( \18824 , \18821 , \18823 );
not \U$18142 ( \18825 , \18824 );
not \U$18143 ( \18826 , \18825 );
not \U$18144 ( \18827 , \17373 );
or \U$18145 ( \18828 , \18826 , \18827 );
nand \U$18146 ( \18829 , \18625 , \17381 );
nand \U$18147 ( \18830 , \18828 , \18829 );
not \U$18148 ( \18831 , \18830 );
nand \U$18149 ( \18832 , \18820 , \18831 );
not \U$18150 ( \18833 , \17270 );
and \U$18151 ( \18834 , \17273 , \17612 );
not \U$18152 ( \18835 , \17273 );
and \U$18153 ( \18836 , \18835 , \17616 );
nor \U$18154 ( \18837 , \18834 , \18836 );
not \U$18155 ( \18838 , \18837 );
or \U$18156 ( \18839 , \18833 , \18838 );
nand \U$18157 ( \18840 , \18617 , \17285 );
nand \U$18158 ( \18841 , \18839 , \18840 );
and \U$18159 ( \18842 , \18832 , \18841 );
nor \U$18160 ( \18843 , \18820 , \18831 );
nor \U$18161 ( \18844 , \18842 , \18843 );
not \U$18162 ( \18845 , \17303 );
not \U$18163 ( \18846 , \17909 );
not \U$18164 ( \18847 , \17666 );
or \U$18165 ( \18848 , \18846 , \18847 );
nand \U$18166 ( \18849 , \17976 , \17908 );
nand \U$18167 ( \18850 , \18848 , \18849 );
not \U$18168 ( \18851 , \18850 );
or \U$18169 ( \18852 , \18845 , \18851 );
nand \U$18170 ( \18853 , \18715 , \17118 );
nand \U$18171 ( \18854 , \18852 , \18853 );
not \U$18172 ( \18855 , \18483 );
not \U$18173 ( \18856 , \17166 );
or \U$18174 ( \18857 , \18855 , \18856 );
nand \U$18175 ( \18858 , \17169 , \18786 );
nand \U$18176 ( \18859 , \18857 , \18858 );
not \U$18177 ( \18860 , \18859 );
not \U$18178 ( \18861 , \16758 );
or \U$18179 ( \18862 , \18860 , \18861 );
nand \U$18180 ( \18863 , \18545 , \16750 );
nand \U$18181 ( \18864 , \18862 , \18863 );
or \U$18182 ( \18865 , \18854 , \18864 );
not \U$18183 ( \18866 , \17236 );
not \U$18184 ( \18867 , \18702 );
or \U$18185 ( \18868 , \18866 , \18867 );
and \U$18186 ( \18869 , \17240 , \17163 );
not \U$18187 ( \18870 , \17240 );
and \U$18188 ( \18871 , \18870 , \18615 );
nor \U$18189 ( \18872 , \18869 , \18871 );
nand \U$18190 ( \18873 , \18872 , \17246 );
nand \U$18191 ( \18874 , \18868 , \18873 );
not \U$18192 ( \18875 , \17285 );
not \U$18193 ( \18876 , \18837 );
or \U$18194 ( \18877 , \18875 , \18876 );
and \U$18195 ( \18878 , \17559 , \17273 );
not \U$18196 ( \18879 , \17559 );
and \U$18197 ( \18880 , \18879 , \17290 );
nor \U$18198 ( \18881 , \18878 , \18880 );
nand \U$18199 ( \18882 , \18881 , \17270 );
nand \U$18200 ( \18883 , \18877 , \18882 );
xor \U$18201 ( \18884 , \18874 , \18883 );
and \U$18202 ( \18885 , \16750 , \18483 );
and \U$18203 ( \18886 , \18884 , \18885 );
and \U$18204 ( \18887 , \18874 , \18883 );
or \U$18205 ( \18888 , \18886 , \18887 );
nand \U$18206 ( \18889 , \18865 , \18888 );
nand \U$18207 ( \18890 , \18854 , \18864 );
and \U$18208 ( \18891 , \18889 , \18890 );
xor \U$18209 ( \18892 , \18844 , \18891 );
xor \U$18210 ( \18893 , \18707 , \18708 );
xor \U$18211 ( \18894 , \18893 , \18720 );
and \U$18212 ( \18895 , \18892 , \18894 );
and \U$18213 ( \18896 , \18844 , \18891 );
or \U$18214 ( \18897 , \18895 , \18896 );
xor \U$18215 ( \18898 , \18819 , \18897 );
xor \U$18216 ( \18899 , \18488 , \18634 );
xor \U$18217 ( \18900 , \18899 , \18665 );
and \U$18218 ( \18901 , \18898 , \18900 );
and \U$18219 ( \18902 , \18819 , \18897 );
or \U$18220 ( \18903 , \18901 , \18902 );
nand \U$18221 ( \18904 , \18817 , \18903 );
not \U$18222 ( \18905 , \18904 );
and \U$18223 ( \18906 , \18591 , \16890 );
not \U$18224 ( \18907 , \18591 );
and \U$18225 ( \18908 , \18907 , \16894 );
nor \U$18226 ( \18909 , \18906 , \18908 );
not \U$18227 ( \18910 , \18909 );
not \U$18228 ( \18911 , \17402 );
or \U$18229 ( \18912 , \18910 , \18911 );
nand \U$18230 ( \18913 , \17405 , \18491 );
nand \U$18231 ( \18914 , \18912 , \18913 );
xor \U$18232 ( \18915 , \18830 , \18841 );
xnor \U$18233 ( \18916 , \18915 , \18820 );
or \U$18234 ( \18917 , \18914 , \18916 );
and \U$18235 ( \18918 , \17781 , \17061 );
not \U$18236 ( \18919 , \17781 );
and \U$18237 ( \18920 , \18919 , \17056 );
nor \U$18238 ( \18921 , \18918 , \18920 );
not \U$18239 ( \18922 , \18921 );
or \U$18240 ( \18923 , \18340 , \18922 );
or \U$18241 ( \18924 , \18824 , \17380 );
nand \U$18242 ( \18925 , \18923 , \18924 );
not \U$18243 ( \18926 , \17246 );
and \U$18244 ( \18927 , \17240 , \17612 );
not \U$18245 ( \18928 , \17240 );
and \U$18246 ( \18929 , \18928 , \17616 );
nor \U$18247 ( \18930 , \18927 , \18929 );
not \U$18248 ( \18931 , \18930 );
or \U$18249 ( \18932 , \18926 , \18931 );
nand \U$18250 ( \18933 , \18872 , \17236 );
nand \U$18251 ( \18934 , \18932 , \18933 );
not \U$18252 ( \18935 , \17285 );
not \U$18253 ( \18936 , \18881 );
or \U$18254 ( \18937 , \18935 , \18936 );
and \U$18255 ( \18938 , \17273 , \17505 );
not \U$18256 ( \18939 , \17273 );
not \U$18257 ( \18940 , \17505 );
and \U$18258 ( \18941 , \18939 , \18940 );
nor \U$18259 ( \18942 , \18938 , \18941 );
nand \U$18260 ( \18943 , \18942 , \17270 );
nand \U$18261 ( \18944 , \18937 , \18943 );
and \U$18262 ( \18945 , \18934 , \18944 );
xor \U$18263 ( \18946 , \18925 , \18945 );
not \U$18264 ( \18947 , \18093 );
not \U$18265 ( \18948 , \17666 );
or \U$18266 ( \18949 , \18947 , \18948 );
nand \U$18267 ( \18950 , \16944 , \18092 );
nand \U$18268 ( \18951 , \18949 , \18950 );
not \U$18269 ( \18952 , \18951 );
not \U$18270 ( \18953 , \17303 );
or \U$18271 ( \18954 , \18952 , \18953 );
nand \U$18272 ( \18955 , \18850 , \17118 );
nand \U$18273 ( \18956 , \18954 , \18955 );
and \U$18274 ( \18957 , \18946 , \18956 );
and \U$18275 ( \18958 , \18925 , \18945 );
or \U$18276 ( \18959 , \18957 , \18958 );
nand \U$18277 ( \18960 , \18917 , \18959 );
nand \U$18278 ( \18961 , \18914 , \18916 );
and \U$18279 ( \18962 , \18960 , \18961 );
not \U$18280 ( \18963 , \18962 );
xor \U$18281 ( \18964 , \18844 , \18891 );
xor \U$18282 ( \18965 , \18964 , \18894 );
not \U$18283 ( \18966 , \18965 );
or \U$18284 ( \18967 , \18963 , \18966 );
not \U$18285 ( \18968 , \18500 );
not \U$18286 ( \18969 , \18968 );
xor \U$18287 ( \18970 , \18631 , \18599 );
not \U$18288 ( \18971 , \18970 );
or \U$18289 ( \18972 , \18969 , \18971 );
or \U$18290 ( \18973 , \18970 , \18968 );
nand \U$18291 ( \18974 , \18972 , \18973 );
nand \U$18292 ( \18975 , \18967 , \18974 );
not \U$18293 ( \18976 , \18962 );
not \U$18294 ( \18977 , \18965 );
nand \U$18295 ( \18978 , \18976 , \18977 );
nand \U$18296 ( \18979 , \18975 , \18978 );
not \U$18297 ( \18980 , \18979 );
xor \U$18298 ( \18981 , \18819 , \18897 );
xor \U$18299 ( \18982 , \18981 , \18900 );
nand \U$18300 ( \18983 , \18980 , \18982 );
not \U$18301 ( \18984 , \18974 );
not \U$18302 ( \18985 , \18962 );
or \U$18303 ( \18986 , \18984 , \18985 );
or \U$18304 ( \18987 , \18962 , \18974 );
nand \U$18305 ( \18988 , \18986 , \18987 );
xnor \U$18306 ( \18989 , \18988 , \18977 );
xor \U$18307 ( \18990 , \18854 , \18888 );
xor \U$18308 ( \18991 , \18990 , \18864 );
not \U$18309 ( \18992 , \18991 );
not \U$18310 ( \18993 , \18992 );
and \U$18311 ( \18994 , \18540 , \16890 );
not \U$18312 ( \18995 , \18540 );
and \U$18313 ( \18996 , \18995 , \16894 );
nor \U$18314 ( \18997 , \18994 , \18996 );
not \U$18315 ( \18998 , \18997 );
not \U$18316 ( \18999 , \17402 );
or \U$18317 ( \19000 , \18998 , \18999 );
nand \U$18318 ( \19001 , \17405 , \18909 );
nand \U$18319 ( \19002 , \19000 , \19001 );
not \U$18320 ( \19003 , \17909 );
not \U$18321 ( \19004 , \17424 );
or \U$18322 ( \19005 , \19003 , \19004 );
nand \U$18323 ( \19006 , \17057 , \17908 );
nand \U$18324 ( \19007 , \19005 , \19006 );
not \U$18325 ( \19008 , \19007 );
not \U$18326 ( \19009 , \18339 );
or \U$18327 ( \19010 , \19008 , \19009 );
nand \U$18328 ( \19011 , \18921 , \17381 );
nand \U$18329 ( \19012 , \19010 , \19011 );
xor \U$18330 ( \19013 , \18934 , \18944 );
xor \U$18331 ( \19014 , \19012 , \19013 );
not \U$18332 ( \19015 , \16946 );
not \U$18333 ( \19016 , \17666 );
or \U$18334 ( \19017 , \19015 , \19016 );
nand \U$18335 ( \19018 , \19017 , \18483 );
and \U$18336 ( \19019 , \16922 , \16933 );
nor \U$18337 ( \19020 , \19019 , \16889 );
and \U$18338 ( \19021 , \19018 , \19020 );
and \U$18339 ( \19022 , \19014 , \19021 );
and \U$18340 ( \19023 , \19012 , \19013 );
or \U$18341 ( \19024 , \19022 , \19023 );
xor \U$18342 ( \19025 , \19002 , \19024 );
xor \U$18343 ( \19026 , \18874 , \18883 );
xor \U$18344 ( \19027 , \19026 , \18885 );
and \U$18345 ( \19028 , \19025 , \19027 );
and \U$18346 ( \19029 , \19002 , \19024 );
or \U$18347 ( \19030 , \19028 , \19029 );
not \U$18348 ( \19031 , \19030 );
not \U$18349 ( \19032 , \19031 );
or \U$18350 ( \19033 , \18993 , \19032 );
not \U$18351 ( \19034 , \18959 );
not \U$18352 ( \19035 , \19034 );
xor \U$18353 ( \19036 , \18916 , \18914 );
not \U$18354 ( \19037 , \19036 );
or \U$18355 ( \19038 , \19035 , \19037 );
or \U$18356 ( \19039 , \19036 , \19034 );
nand \U$18357 ( \19040 , \19038 , \19039 );
nand \U$18358 ( \19041 , \19033 , \19040 );
nand \U$18359 ( \19042 , \19030 , \18991 );
and \U$18360 ( \19043 , \19041 , \19042 );
nand \U$18361 ( \19044 , \18989 , \19043 );
nand \U$18362 ( \19045 , \18983 , \19044 );
nor \U$18363 ( \19046 , \18905 , \19045 );
not \U$18364 ( \19047 , \18727 );
nand \U$18365 ( \19048 , \19047 , \18668 );
not \U$18366 ( \19049 , \19048 );
not \U$18367 ( \19050 , \18816 );
or \U$18368 ( \19051 , \19049 , \19050 );
not \U$18369 ( \19052 , \18668 );
nand \U$18370 ( \19053 , \19052 , \18727 );
nand \U$18371 ( \19054 , \19051 , \19053 );
not \U$18372 ( \19055 , \19054 );
not \U$18373 ( \19056 , \17373 );
not \U$18374 ( \19057 , \18747 );
or \U$18375 ( \19058 , \19056 , \19057 );
nand \U$18376 ( \19059 , \18106 , \17381 );
nand \U$18377 ( \19060 , \19058 , \19059 );
xor \U$18378 ( \19061 , \18117 , \18126 );
xor \U$18379 ( \19062 , \19060 , \19061 );
xor \U$18381 ( \19063 , \19062 , 1'b0 );
xor \U$18382 ( \19064 , \18736 , \18741 );
and \U$18383 ( \19065 , \19064 , \18750 );
and \U$18384 ( \19066 , \18736 , \18741 );
or \U$18385 ( \19067 , \19065 , \19066 );
not \U$18386 ( \19068 , \18782 );
not \U$18387 ( \19069 , \17303 );
or \U$18388 ( \19070 , \19068 , \19069 );
nand \U$18389 ( \19071 , \18165 , \17118 );
nand \U$18390 ( \19072 , \19070 , \19071 );
xor \U$18391 ( \19073 , \19067 , \19072 );
not \U$18392 ( \19074 , \18759 );
not \U$18393 ( \19075 , \16758 );
or \U$18394 ( \19076 , \19074 , \19075 );
nand \U$18395 ( \19077 , \18155 , \16750 );
nand \U$18396 ( \19078 , \19076 , \19077 );
xor \U$18397 ( \19079 , \19073 , \19078 );
xor \U$18398 ( \19080 , \19063 , \19079 );
xor \U$18399 ( \19081 , \18774 , \18784 );
and \U$18400 ( \19082 , \19081 , \18787 );
and \U$18401 ( \19083 , \18774 , \18784 );
or \U$18402 ( \19084 , \19082 , \19083 );
xor \U$18403 ( \19085 , \19080 , \19084 );
xor \U$18404 ( \19086 , \18772 , \18788 );
and \U$18405 ( \19087 , \19086 , \18815 );
and \U$18406 ( \19088 , \18772 , \18788 );
or \U$18407 ( \19089 , \19087 , \19088 );
xor \U$18408 ( \19090 , \19085 , \19089 );
xor \U$18409 ( \19091 , \18751 , \18761 );
and \U$18410 ( \19092 , \19091 , \18771 );
and \U$18411 ( \19093 , \18751 , \18761 );
or \U$18412 ( \19094 , \19092 , \19093 );
xor \U$18413 ( \19095 , \18798 , \18807 );
and \U$18414 ( \19096 , \19095 , \18814 );
and \U$18415 ( \19097 , \18798 , \18807 );
or \U$18416 ( \19098 , \19096 , \19097 );
xor \U$18417 ( \19099 , \19094 , \19098 );
not \U$18418 ( \19100 , \18769 );
not \U$18419 ( \19101 , \17402 );
or \U$18420 ( \19102 , \19100 , \19101 );
nand \U$18421 ( \19103 , \17405 , \18178 );
nand \U$18422 ( \19104 , \19102 , \19103 );
not \U$18423 ( \19105 , \16638 );
and \U$18424 ( \19106 , \16642 , \18539 );
and \U$18425 ( \19107 , \17910 , \18540 );
nor \U$18426 ( \19108 , \19106 , \19107 );
nand \U$18427 ( \19109 , \19105 , \19108 );
xor \U$18428 ( \19110 , \19104 , \19109 );
not \U$18429 ( \19111 , \18796 );
not \U$18430 ( \19112 , \16572 );
or \U$18431 ( \19113 , \19111 , \19112 );
not \U$18432 ( \19114 , \18093 );
not \U$18433 ( \19115 , \17561 );
or \U$18434 ( \19116 , \19114 , \19115 );
nand \U$18435 ( \19117 , \16574 , \18092 );
nand \U$18436 ( \19118 , \19116 , \19117 );
nand \U$18437 ( \19119 , \19118 , \16630 );
nand \U$18438 ( \19120 , \19113 , \19119 );
xnor \U$18439 ( \19121 , \19110 , \19120 );
xnor \U$18440 ( \19122 , \19099 , \19121 );
not \U$18441 ( \19123 , \19122 );
xnor \U$18442 ( \19124 , \19090 , \19123 );
nand \U$18443 ( \19125 , \19055 , \19124 );
xor \U$18444 ( \19126 , \18925 , \18945 );
xor \U$18445 ( \19127 , \19126 , \18956 );
or \U$18446 ( \19128 , \16889 , \18483 );
or \U$18447 ( \19129 , \18786 , \16890 );
nand \U$18448 ( \19130 , \19128 , \19129 );
not \U$18449 ( \19131 , \19130 );
not \U$18450 ( \19132 , \17402 );
or \U$18451 ( \19133 , \19131 , \19132 );
nand \U$18452 ( \19134 , \17405 , \18997 );
nand \U$18453 ( \19135 , \19133 , \19134 );
not \U$18454 ( \19136 , \18591 );
not \U$18455 ( \19137 , \16995 );
or \U$18456 ( \19138 , \19136 , \19137 );
nand \U$18457 ( \19139 , \16944 , \18595 );
nand \U$18458 ( \19140 , \19138 , \19139 );
not \U$18459 ( \19141 , \19140 );
not \U$18460 ( \19142 , \17303 );
or \U$18461 ( \19143 , \19141 , \19142 );
nand \U$18462 ( \19144 , \18951 , \17118 );
nand \U$18463 ( \19145 , \19143 , \19144 );
xor \U$18464 ( \19146 , \19135 , \19145 );
not \U$18465 ( \19147 , \17236 );
not \U$18466 ( \19148 , \18930 );
or \U$18467 ( \19149 , \19147 , \19148 );
and \U$18468 ( \19150 , \17558 , \17230 );
not \U$18469 ( \19151 , \17558 );
and \U$18470 ( \19152 , \19151 , \17240 );
or \U$18471 ( \19153 , \19150 , \19152 );
nand \U$18472 ( \19154 , \19153 , \17246 );
nand \U$18473 ( \19155 , \19149 , \19154 );
not \U$18474 ( \19156 , \19155 );
not \U$18475 ( \19157 , \17062 );
not \U$18476 ( \19158 , \18093 );
or \U$18477 ( \19159 , \19157 , \19158 );
nand \U$18478 ( \19160 , \18092 , \17057 );
nand \U$18479 ( \19161 , \19159 , \19160 );
not \U$18480 ( \19162 , \19161 );
not \U$18481 ( \19163 , \17373 );
or \U$18482 ( \19164 , \19162 , \19163 );
nand \U$18483 ( \19165 , \19007 , \17381 );
nand \U$18484 ( \19166 , \19164 , \19165 );
not \U$18485 ( \19167 , \19166 );
or \U$18486 ( \19168 , \19156 , \19167 );
or \U$18487 ( \19169 , \19166 , \19155 );
not \U$18488 ( \19170 , \18942 );
not \U$18489 ( \19171 , \19170 );
not \U$18490 ( \19172 , \17268 );
and \U$18491 ( \19173 , \19171 , \19172 );
not \U$18492 ( \19174 , \17273 );
not \U$18493 ( \19175 , \17782 );
or \U$18494 ( \19176 , \19174 , \19175 );
nand \U$18495 ( \19177 , \17781 , \17290 );
nand \U$18496 ( \19178 , \19176 , \19177 );
and \U$18497 ( \19179 , \19178 , \17270 );
nor \U$18498 ( \19180 , \19173 , \19179 );
not \U$18499 ( \19181 , \19180 );
nand \U$18500 ( \19182 , \19169 , \19181 );
nand \U$18501 ( \19183 , \19168 , \19182 );
and \U$18502 ( \19184 , \19146 , \19183 );
and \U$18503 ( \19185 , \19135 , \19145 );
or \U$18504 ( \19186 , \19184 , \19185 );
xor \U$18505 ( \19187 , \19127 , \19186 );
xor \U$18506 ( \19188 , \19002 , \19024 );
xor \U$18507 ( \19189 , \19188 , \19027 );
and \U$18508 ( \19190 , \19187 , \19189 );
and \U$18509 ( \19191 , \19127 , \19186 );
or \U$18510 ( \19192 , \19190 , \19191 );
and \U$18511 ( \19193 , \19030 , \18992 );
not \U$18512 ( \19194 , \19030 );
and \U$18513 ( \19195 , \19194 , \18991 );
nor \U$18514 ( \19196 , \19193 , \19195 );
xnor \U$18515 ( \19197 , \19196 , \19040 );
xor \U$18516 ( \19198 , \19192 , \19197 );
xor \U$18517 ( \19199 , \19012 , \19013 );
xor \U$18518 ( \19200 , \19199 , \19021 );
nand \U$18519 ( \19201 , \17405 , \18483 );
not \U$18520 ( \19202 , \19201 );
not \U$18521 ( \19203 , \17303 );
not \U$18522 ( \19204 , \18540 );
not \U$18523 ( \19205 , \17666 );
or \U$18524 ( \19206 , \19204 , \19205 );
nand \U$18525 ( \19207 , \17976 , \18539 );
nand \U$18526 ( \19208 , \19206 , \19207 );
not \U$18527 ( \19209 , \19208 );
or \U$18528 ( \19210 , \19203 , \19209 );
nand \U$18529 ( \19211 , \19140 , \17118 );
nand \U$18530 ( \19212 , \19210 , \19211 );
nor \U$18531 ( \19213 , \19202 , \19212 );
nand \U$18532 ( \19214 , \17051 , \17062 );
and \U$18533 ( \19215 , \19214 , \18483 );
and \U$18534 ( \19216 , \17057 , \17050 );
nor \U$18535 ( \19217 , \19215 , \19216 );
and \U$18536 ( \19218 , \16922 , \19217 );
not \U$18537 ( \19219 , \17285 );
not \U$18538 ( \19220 , \19178 );
or \U$18539 ( \19221 , \19219 , \19220 );
not \U$18540 ( \19222 , \17273 );
not \U$18541 ( \19223 , \17908 );
or \U$18542 ( \19224 , \19222 , \19223 );
nand \U$18543 ( \19225 , \17907 , \17290 );
nand \U$18544 ( \19226 , \19224 , \19225 );
nand \U$18545 ( \19227 , \19226 , \17270 );
nand \U$18546 ( \19228 , \19221 , \19227 );
nand \U$18547 ( \19229 , \19218 , \19228 );
or \U$18548 ( \19230 , \19213 , \19229 );
not \U$18549 ( \19231 , \19201 );
nand \U$18550 ( \19232 , \19231 , \19212 );
nand \U$18551 ( \19233 , \19230 , \19232 );
xor \U$18552 ( \19234 , \19200 , \19233 );
xor \U$18553 ( \19235 , \19135 , \19145 );
xor \U$18554 ( \19236 , \19235 , \19183 );
and \U$18555 ( \19237 , \19234 , \19236 );
and \U$18556 ( \19238 , \19200 , \19233 );
or \U$18557 ( \19239 , \19237 , \19238 );
xor \U$18558 ( \19240 , \19127 , \19186 );
xor \U$18559 ( \19241 , \19240 , \19189 );
xor \U$18560 ( \19242 , \19239 , \19241 );
xor \U$18561 ( \19243 , \19155 , \19180 );
xor \U$18562 ( \19244 , \19243 , \19166 );
xor \U$18563 ( \19245 , \19218 , \19228 );
not \U$18564 ( \19246 , \17062 );
not \U$18565 ( \19247 , \18591 );
or \U$18566 ( \19248 , \19246 , \19247 );
not \U$18567 ( \19249 , \18590 );
nand \U$18568 ( \19250 , \19249 , \17057 );
nand \U$18569 ( \19251 , \19248 , \19250 );
not \U$18570 ( \19252 , \19251 );
not \U$18571 ( \19253 , \17373 );
or \U$18572 ( \19254 , \19252 , \19253 );
nand \U$18573 ( \19255 , \19161 , \17381 );
nand \U$18574 ( \19256 , \19254 , \19255 );
not \U$18575 ( \19257 , \19256 );
not \U$18576 ( \19258 , \17246 );
and \U$18577 ( \19259 , \17240 , \17505 );
not \U$18578 ( \19260 , \17240 );
and \U$18579 ( \19261 , \19260 , \18940 );
nor \U$18580 ( \19262 , \19259 , \19261 );
not \U$18581 ( \19263 , \19262 );
or \U$18582 ( \19264 , \19258 , \19263 );
nand \U$18583 ( \19265 , \19153 , \17236 );
nand \U$18584 ( \19266 , \19264 , \19265 );
not \U$18585 ( \19267 , \19266 );
nand \U$18586 ( \19268 , \19257 , \19267 );
and \U$18587 ( \19269 , \19245 , \19268 );
nor \U$18588 ( \19270 , \19257 , \19267 );
nor \U$18589 ( \19271 , \19269 , \19270 );
or \U$18590 ( \19272 , \19244 , \19271 );
xor \U$18591 ( \19273 , \19229 , \19201 );
xnor \U$18592 ( \19274 , \19273 , \19212 );
and \U$18593 ( \19275 , \19271 , \19244 );
or \U$18594 ( \19276 , \19274 , \19275 );
nand \U$18595 ( \19277 , \19272 , \19276 );
xor \U$18596 ( \19278 , \19200 , \19233 );
xor \U$18597 ( \19279 , \19278 , \19236 );
xor \U$18598 ( \19280 , \19277 , \19279 );
not \U$18599 ( \19281 , \17285 );
not \U$18600 ( \19282 , \19226 );
or \U$18601 ( \19283 , \19281 , \19282 );
xor \U$18602 ( \19284 , \17273 , \18091 );
nand \U$18603 ( \19285 , \19284 , \17270 );
nand \U$18604 ( \19286 , \19283 , \19285 );
and \U$18605 ( \19287 , \17064 , \18483 );
xor \U$18606 ( \19288 , \19286 , \19287 );
not \U$18607 ( \19289 , \17381 );
not \U$18608 ( \19290 , \19251 );
or \U$18609 ( \19291 , \19289 , \19290 );
not \U$18610 ( \19292 , \17057 );
not \U$18611 ( \19293 , \18539 );
or \U$18612 ( \19294 , \19292 , \19293 );
nand \U$18613 ( \19295 , \18538 , \17056 );
nand \U$18614 ( \19296 , \19294 , \19295 );
nand \U$18615 ( \19297 , \19296 , \17373 );
nand \U$18616 ( \19298 , \19291 , \19297 );
and \U$18617 ( \19299 , \19288 , \19298 );
and \U$18618 ( \19300 , \19286 , \19287 );
or \U$18619 ( \19301 , \19299 , \19300 );
and \U$18620 ( \19302 , \18483 , \17976 );
not \U$18621 ( \19303 , \18483 );
and \U$18622 ( \19304 , \19303 , \17666 );
nor \U$18623 ( \19305 , \19302 , \19304 );
not \U$18624 ( \19306 , \19305 );
not \U$18625 ( \19307 , \17303 );
or \U$18626 ( \19308 , \19306 , \19307 );
nand \U$18627 ( \19309 , \19208 , \17118 );
nand \U$18628 ( \19310 , \19308 , \19309 );
xor \U$18629 ( \19311 , \19301 , \19310 );
not \U$18630 ( \19312 , \19245 );
not \U$18631 ( \19313 , \19267 );
not \U$18632 ( \19314 , \19256 );
and \U$18633 ( \19315 , \19313 , \19314 );
and \U$18634 ( \19316 , \19256 , \19267 );
nor \U$18635 ( \19317 , \19315 , \19316 );
not \U$18636 ( \19318 , \19317 );
or \U$18637 ( \19319 , \19312 , \19318 );
or \U$18638 ( \19320 , \19245 , \19317 );
nand \U$18639 ( \19321 , \19319 , \19320 );
and \U$18640 ( \19322 , \19311 , \19321 );
and \U$18641 ( \19323 , \19301 , \19310 );
or \U$18642 ( \19324 , \19322 , \19323 );
not \U$18643 ( \19325 , \19324 );
not \U$18644 ( \19326 , \19274 );
xor \U$18645 ( \19327 , \19271 , \19244 );
not \U$18646 ( \19328 , \19327 );
and \U$18647 ( \19329 , \19326 , \19328 );
and \U$18648 ( \19330 , \19274 , \19327 );
nor \U$18649 ( \19331 , \19329 , \19330 );
nand \U$18650 ( \19332 , \19325 , \19331 );
not \U$18651 ( \19333 , \19332 );
xor \U$18652 ( \19334 , \19301 , \19310 );
xor \U$18653 ( \19335 , \19334 , \19321 );
not \U$18654 ( \19336 , \17236 );
not \U$18655 ( \19337 , \19262 );
or \U$18656 ( \19338 , \19336 , \19337 );
and \U$18657 ( \19339 , \17240 , \17782 );
not \U$18658 ( \19340 , \17240 );
and \U$18659 ( \19341 , \19340 , \17781 );
nor \U$18660 ( \19342 , \19339 , \19341 );
not \U$18661 ( \19343 , \19342 );
nand \U$18662 ( \19344 , \19343 , \17246 );
nand \U$18663 ( \19345 , \19338 , \19344 );
or \U$18664 ( \19346 , \17364 , \17273 );
nand \U$18665 ( \19347 , \19346 , \18483 );
nand \U$18666 ( \19348 , \17364 , \17273 );
and \U$18667 ( \19349 , \19347 , \17061 , \19348 );
not \U$18668 ( \19350 , \17285 );
not \U$18669 ( \19351 , \19284 );
or \U$18670 ( \19352 , \19350 , \19351 );
and \U$18671 ( \19353 , \17273 , \19249 );
not \U$18672 ( \19354 , \17273 );
and \U$18673 ( \19355 , \19354 , \18590 );
or \U$18674 ( \19356 , \19353 , \19355 );
nand \U$18675 ( \19357 , \19356 , \17270 );
nand \U$18676 ( \19358 , \19352 , \19357 );
and \U$18677 ( \19359 , \19349 , \19358 );
xor \U$18678 ( \19360 , \19345 , \19359 );
xor \U$18679 ( \19361 , \19286 , \19287 );
xor \U$18680 ( \19362 , \19361 , \19298 );
and \U$18681 ( \19363 , \19360 , \19362 );
and \U$18682 ( \19364 , \19345 , \19359 );
or \U$18683 ( \19365 , \19363 , \19364 );
nor \U$18684 ( \19366 , \19335 , \19365 );
nand \U$18685 ( \19367 , \17262 , \17230 );
nand \U$18686 ( \19368 , \18483 , \19367 );
and \U$18687 ( \19369 , \17259 , \17240 );
nor \U$18688 ( \19370 , \19369 , \17290 );
and \U$18689 ( \19371 , \19368 , \19370 );
not \U$18690 ( \19372 , \17236 );
and \U$18691 ( \19373 , \18091 , \17230 );
not \U$18692 ( \19374 , \18091 );
and \U$18693 ( \19375 , \19374 , \17240 );
or \U$18694 ( \19376 , \19373 , \19375 );
not \U$18695 ( \19377 , \19376 );
or \U$18696 ( \19378 , \19372 , \19377 );
and \U$18697 ( \19379 , \18590 , \17230 );
not \U$18698 ( \19380 , \18590 );
and \U$18699 ( \19381 , \19380 , \17240 );
or \U$18700 ( \19382 , \19379 , \19381 );
nand \U$18701 ( \19383 , \19382 , \17246 );
nand \U$18702 ( \19384 , \19378 , \19383 );
and \U$18703 ( \19385 , \19371 , \19384 );
not \U$18704 ( \19386 , \17369 );
nand \U$18705 ( \19387 , \19386 , \18483 );
not \U$18706 ( \19388 , \17246 );
not \U$18707 ( \19389 , \19376 );
or \U$18708 ( \19390 , \19388 , \19389 );
and \U$18709 ( \19391 , \17907 , \17230 );
not \U$18710 ( \19392 , \17907 );
and \U$18711 ( \19393 , \19392 , \17240 );
or \U$18712 ( \19394 , \19391 , \19393 );
nand \U$18713 ( \19395 , \19394 , \17236 );
nand \U$18714 ( \19396 , \19390 , \19395 );
xor \U$18715 ( \19397 , \19387 , \19396 );
not \U$18716 ( \19398 , \17270 );
and \U$18717 ( \19399 , \18538 , \17290 );
not \U$18718 ( \19400 , \18538 );
and \U$18719 ( \19401 , \19400 , \17273 );
or \U$18720 ( \19402 , \19399 , \19401 );
not \U$18721 ( \19403 , \19402 );
or \U$18722 ( \19404 , \19398 , \19403 );
nand \U$18723 ( \19405 , \19356 , \17285 );
nand \U$18724 ( \19406 , \19404 , \19405 );
xnor \U$18725 ( \19407 , \19397 , \19406 );
xor \U$18726 ( \19408 , \19385 , \19407 );
and \U$18727 ( \19409 , \17273 , \18786 );
not \U$18728 ( \19410 , \17273 );
and \U$18729 ( \19411 , \19410 , \18483 );
nor \U$18730 ( \19412 , \19409 , \19411 );
or \U$18731 ( \19413 , \19412 , \17269 );
not \U$18732 ( \19414 , \19402 );
or \U$18733 ( \19415 , \19414 , \17268 );
nand \U$18734 ( \19416 , \19413 , \19415 );
not \U$18735 ( \19417 , \19416 );
xor \U$18736 ( \19418 , \19371 , \19384 );
not \U$18737 ( \19419 , \19418 );
or \U$18738 ( \19420 , \19417 , \19419 );
or \U$18739 ( \19421 , \19418 , \19416 );
not \U$18740 ( \19422 , \17246 );
xor \U$18741 ( \19423 , \17240 , \18538 );
not \U$18742 ( \19424 , \19423 );
or \U$18743 ( \19425 , \19422 , \19424 );
nand \U$18744 ( \19426 , \19382 , \17236 );
nand \U$18745 ( \19427 , \19425 , \19426 );
nor \U$18746 ( \19428 , \18786 , \17268 );
nor \U$18747 ( \19429 , \19427 , \19428 );
not \U$18748 ( \19430 , \17236 );
not \U$18749 ( \19431 , \19423 );
or \U$18750 ( \19432 , \19430 , \19431 );
nand \U$18751 ( \19433 , \18786 , \17246 );
nand \U$18752 ( \19434 , \19432 , \19433 );
nand \U$18753 ( \19435 , \18483 , \17236 );
and \U$18754 ( \19436 , \19435 , \17240 );
nand \U$18755 ( \19437 , \19434 , \19436 );
or \U$18756 ( \19438 , \19429 , \19437 );
nand \U$18757 ( \19439 , \19427 , \19428 );
nand \U$18758 ( \19440 , \19438 , \19439 );
nand \U$18759 ( \19441 , \19421 , \19440 );
nand \U$18760 ( \19442 , \19420 , \19441 );
and \U$18761 ( \19443 , \19408 , \19442 );
and \U$18762 ( \19444 , \19385 , \19407 );
or \U$18763 ( \19445 , \19443 , \19444 );
xor \U$18764 ( \19446 , \19349 , \19358 );
not \U$18765 ( \19447 , \19446 );
not \U$18766 ( \19448 , \17381 );
not \U$18767 ( \19449 , \19296 );
or \U$18768 ( \19450 , \19448 , \19449 );
not \U$18769 ( \19451 , \17056 );
not \U$18770 ( \19452 , \18483 );
or \U$18771 ( \19453 , \19451 , \19452 );
nand \U$18772 ( \19454 , \18786 , \17061 );
nand \U$18773 ( \19455 , \19453 , \19454 );
nand \U$18774 ( \19456 , \17373 , \19455 );
nand \U$18775 ( \19457 , \19450 , \19456 );
not \U$18776 ( \19458 , \19457 );
not \U$18777 ( \19459 , \19342 );
not \U$18778 ( \19460 , \17237 );
and \U$18779 ( \19461 , \19459 , \19460 );
and \U$18780 ( \19462 , \19394 , \17246 );
nor \U$18781 ( \19463 , \19461 , \19462 );
not \U$18782 ( \19464 , \19463 );
and \U$18783 ( \19465 , \19458 , \19464 );
and \U$18784 ( \19466 , \19463 , \19457 );
nor \U$18785 ( \19467 , \19465 , \19466 );
not \U$18786 ( \19468 , \19467 );
and \U$18787 ( \19469 , \19447 , \19468 );
and \U$18788 ( \19470 , \19446 , \19467 );
nor \U$18789 ( \19471 , \19469 , \19470 );
not \U$18790 ( \19472 , \19387 );
or \U$18791 ( \19473 , \19396 , \19472 );
nand \U$18792 ( \19474 , \19473 , \19406 );
nand \U$18793 ( \19475 , \19396 , \19472 );
and \U$18794 ( \19476 , \19474 , \19475 );
nand \U$18795 ( \19477 , \19471 , \19476 );
and \U$18796 ( \19478 , \19445 , \19477 );
nor \U$18797 ( \19479 , \19471 , \19476 );
nor \U$18798 ( \19480 , \19478 , \19479 );
xor \U$18799 ( \19481 , \19345 , \19359 );
xor \U$18800 ( \19482 , \19481 , \19362 );
not \U$18801 ( \19483 , \19457 );
nand \U$18802 ( \19484 , \19483 , \19463 );
not \U$18803 ( \19485 , \19484 );
not \U$18804 ( \19486 , \19446 );
or \U$18805 ( \19487 , \19485 , \19486 );
not \U$18806 ( \19488 , \19463 );
nand \U$18807 ( \19489 , \19488 , \19457 );
nand \U$18808 ( \19490 , \19487 , \19489 );
nor \U$18809 ( \19491 , \19482 , \19490 );
or \U$18810 ( \19492 , \19480 , \19491 );
nand \U$18811 ( \19493 , \19482 , \19490 );
nand \U$18812 ( \19494 , \19492 , \19493 );
not \U$18813 ( \19495 , \19494 );
or \U$18814 ( \19496 , \19366 , \19495 );
nand \U$18815 ( \19497 , \19335 , \19365 );
nand \U$18816 ( \19498 , \19496 , \19497 );
not \U$18817 ( \19499 , \19498 );
or \U$18818 ( \19500 , \19333 , \19499 );
not \U$18819 ( \19501 , \19331 );
nand \U$18820 ( \19502 , \19501 , \19324 );
nand \U$18821 ( \19503 , \19500 , \19502 );
and \U$18822 ( \19504 , \19280 , \19503 );
and \U$18823 ( \19505 , \19277 , \19279 );
or \U$18824 ( \19506 , \19504 , \19505 );
and \U$18825 ( \19507 , \19242 , \19506 );
and \U$18826 ( \19508 , \19239 , \19241 );
or \U$18827 ( \19509 , \19507 , \19508 );
and \U$18828 ( \19510 , \19198 , \19509 );
and \U$18829 ( \19511 , \19192 , \19197 );
or \U$18830 ( \19512 , \19510 , \19511 );
nand \U$18831 ( \19513 , \19046 , \19125 , \19512 );
nor \U$18832 ( \19514 , \18989 , \19043 );
nand \U$18833 ( \19515 , \18983 , \19514 );
not \U$18834 ( \19516 , \18982 );
nand \U$18835 ( \19517 , \19516 , \18979 );
nand \U$18836 ( \19518 , \19515 , \19517 );
nand \U$18837 ( \19519 , \19518 , \18904 );
not \U$18838 ( \19520 , \19519 );
or \U$18839 ( \19521 , \18817 , \18903 );
not \U$18840 ( \19522 , \19521 );
or \U$18841 ( \19523 , \19520 , \19522 );
nand \U$18842 ( \19524 , \19523 , \19125 );
not \U$18843 ( \19525 , \19124 );
nand \U$18844 ( \19526 , \19525 , \19054 );
nand \U$18845 ( \19527 , \19513 , \19524 , \19526 );
xor \U$18846 ( \19528 , \18150 , \18183 );
xor \U$18847 ( \19529 , \19528 , \18189 );
not \U$18848 ( \19530 , \19104 );
nand \U$18849 ( \19531 , \19530 , \19109 );
not \U$18850 ( \19532 , \19531 );
not \U$18851 ( \19533 , \19120 );
or \U$18852 ( \19534 , \19532 , \19533 );
not \U$18853 ( \19535 , \19109 );
nand \U$18854 ( \19536 , \19535 , \19104 );
nand \U$18855 ( \19537 , \19534 , \19536 );
not \U$18856 ( \19538 , \19537 );
and \U$18858 ( \19539 , \19060 , \19061 );
or \U$18859 ( \19540 , 1'b0 , \19539 );
and \U$18860 ( \19541 , \18591 , \17910 );
not \U$18861 ( \19542 , \18591 );
and \U$18862 ( \19543 , \19542 , \16642 );
nor \U$18863 ( \19544 , \19541 , \19543 );
and \U$18864 ( \19545 , \19105 , \19544 );
xor \U$18865 ( \19546 , \19540 , \19545 );
not \U$18866 ( \19547 , \19118 );
not \U$18867 ( \19548 , \17922 );
or \U$18868 ( \19549 , \19547 , \19548 );
nand \U$18869 ( \19550 , \18040 , \16630 );
nand \U$18870 ( \19551 , \19549 , \19550 );
xor \U$18871 ( \19552 , \19546 , \19551 );
not \U$18872 ( \19553 , \19552 );
or \U$18873 ( \19554 , \19538 , \19553 );
or \U$18874 ( \19555 , \19552 , \19537 );
xor \U$18875 ( \19556 , \19063 , \19079 );
and \U$18876 ( \19557 , \19556 , \19084 );
and \U$18877 ( \19558 , \19063 , \19079 );
or \U$18878 ( \19559 , \19557 , \19558 );
nand \U$18879 ( \19560 , \19555 , \19559 );
nand \U$18880 ( \19561 , \19554 , \19560 );
xor \U$18881 ( \19562 , \19529 , \19561 );
not \U$18882 ( \19563 , \19551 );
not \U$18883 ( \19564 , \19545 );
or \U$18884 ( \19565 , \19563 , \19564 );
or \U$18885 ( \19566 , \19545 , \19551 );
nand \U$18886 ( \19567 , \19566 , \19540 );
nand \U$18887 ( \19568 , \19565 , \19567 );
xor \U$18888 ( \19569 , \18132 , \18098 );
xnor \U$18889 ( \19570 , \19569 , \18045 );
xor \U$18890 ( \19571 , \19568 , \19570 );
xor \U$18891 ( \19572 , \18111 , \18127 );
xor \U$18892 ( \19573 , \19572 , \18129 );
xor \U$18893 ( \19574 , \19067 , \19072 );
and \U$18894 ( \19575 , \19574 , \19078 );
and \U$18895 ( \19576 , \19067 , \19072 );
or \U$18896 ( \19577 , \19575 , \19576 );
xor \U$18897 ( \19578 , \19573 , \19577 );
xor \U$18898 ( \19579 , \18160 , \18170 );
xor \U$18899 ( \19580 , \19579 , \18180 );
and \U$18900 ( \19581 , \19578 , \19580 );
and \U$18901 ( \19582 , \19573 , \19577 );
or \U$18902 ( \19583 , \19581 , \19582 );
xnor \U$18903 ( \19584 , \19571 , \19583 );
xor \U$18904 ( \19585 , \19562 , \19584 );
not \U$18905 ( \19586 , \19585 );
xor \U$18906 ( \19587 , \19573 , \19577 );
xor \U$18907 ( \19588 , \19587 , \19580 );
not \U$18908 ( \19589 , \19094 );
not \U$18909 ( \19590 , \19121 );
or \U$18910 ( \19591 , \19589 , \19590 );
or \U$18911 ( \19592 , \19094 , \19121 );
nand \U$18912 ( \19593 , \19592 , \19098 );
nand \U$18913 ( \19594 , \19591 , \19593 );
xor \U$18914 ( \19595 , \19588 , \19594 );
xor \U$18915 ( \19596 , \19537 , \19552 );
xor \U$18916 ( \19597 , \19596 , \19559 );
and \U$18917 ( \19598 , \19595 , \19597 );
and \U$18918 ( \19599 , \19588 , \19594 );
or \U$18919 ( \19600 , \19598 , \19599 );
not \U$18920 ( \19601 , \19600 );
nand \U$18921 ( \19602 , \19586 , \19601 );
xor \U$18922 ( \19603 , \19588 , \19594 );
xor \U$18923 ( \19604 , \19603 , \19597 );
not \U$18924 ( \19605 , \19085 );
not \U$18925 ( \19606 , \19605 );
not \U$18926 ( \19607 , \19122 );
or \U$18927 ( \19608 , \19606 , \19607 );
nand \U$18928 ( \19609 , \19608 , \19089 );
nand \U$18929 ( \19610 , \19123 , \19085 );
nand \U$18930 ( \19611 , \19609 , \19610 );
or \U$18931 ( \19612 , \19604 , \19611 );
nand \U$18932 ( \19613 , \19602 , \19612 );
xor \U$18933 ( \19614 , \18034 , \18194 );
xnor \U$18934 ( \19615 , \19614 , \18199 );
xor \U$18935 ( \19616 , \18016 , \18018 );
xnor \U$18936 ( \19617 , \19616 , \18019 );
not \U$18937 ( \19618 , \19570 );
not \U$18938 ( \19619 , \19568 );
not \U$18939 ( \19620 , \19619 );
or \U$18940 ( \19621 , \19618 , \19620 );
nand \U$18941 ( \19622 , \19621 , \19583 );
not \U$18942 ( \19623 , \19570 );
nand \U$18943 ( \19624 , \19623 , \19568 );
and \U$18944 ( \19625 , \19622 , \19624 );
xor \U$18945 ( \19626 , \19617 , \19625 );
xor \U$18946 ( \19627 , \18134 , \18145 );
xnor \U$18947 ( \19628 , \19627 , \18192 );
and \U$18948 ( \19629 , \19626 , \19628 );
and \U$18949 ( \19630 , \19617 , \19625 );
or \U$18950 ( \19631 , \19629 , \19630 );
nand \U$18951 ( \19632 , \19615 , \19631 );
xor \U$18952 ( \19633 , \19617 , \19625 );
xor \U$18953 ( \19634 , \19633 , \19628 );
not \U$18954 ( \19635 , \19529 );
not \U$18955 ( \19636 , \19584 );
nand \U$18956 ( \19637 , \19635 , \19636 );
and \U$18957 ( \19638 , \19637 , \19561 );
not \U$18958 ( \19639 , \19529 );
nor \U$18959 ( \19640 , \19639 , \19636 );
nor \U$18960 ( \19641 , \19638 , \19640 );
nand \U$18961 ( \19642 , \19634 , \19641 );
nand \U$18962 ( \19643 , \19632 , \19642 );
nor \U$18963 ( \19644 , \19613 , \19643 );
and \U$18964 ( \19645 , \19527 , \19644 );
not \U$18965 ( \19646 , \19645 );
or \U$18966 ( \19647 , \18405 , \19646 );
not \U$18967 ( \19648 , \18201 );
nor \U$18968 ( \19649 , \19648 , \18204 );
and \U$18969 ( \19650 , \18032 , \19649 );
nand \U$18970 ( \19651 , \18379 , \18391 );
not \U$18971 ( \19652 , \19651 );
nor \U$18972 ( \19653 , \19650 , \19652 );
not \U$18973 ( \19654 , \19643 );
nand \U$18974 ( \19655 , \19604 , \19611 );
nand \U$18975 ( \19656 , \19585 , \19600 );
nand \U$18976 ( \19657 , \19655 , \19656 );
and \U$18977 ( \19658 , \19657 , \19602 );
nand \U$18978 ( \19659 , \19654 , \19658 );
nor \U$18979 ( \19660 , \19634 , \19641 );
not \U$18980 ( \19661 , \19660 );
not \U$18981 ( \19662 , \19632 );
or \U$18982 ( \19663 , \19661 , \19662 );
or \U$18983 ( \19664 , \19615 , \19631 );
nand \U$18984 ( \19665 , \19663 , \19664 );
not \U$18985 ( \19666 , \17861 );
nand \U$18986 ( \19667 , \19666 , \18030 );
nand \U$18987 ( \19668 , \18394 , \18401 );
nand \U$18988 ( \19669 , \19667 , \19668 );
nor \U$18989 ( \19670 , \19665 , \19669 );
nand \U$18990 ( \19671 , \19653 , \19659 , \19670 );
nor \U$18991 ( \19672 , \18206 , \19669 );
nand \U$18992 ( \19673 , \19653 , \19672 );
and \U$18993 ( \19674 , \19651 , \18402 );
nor \U$18994 ( \19675 , \19674 , \18392 );
nand \U$18995 ( \19676 , \19671 , \19673 , \19675 );
nand \U$18996 ( \19677 , \19647 , \19676 );
not \U$18997 ( \19678 , \18269 );
not \U$18998 ( \19679 , \17390 );
or \U$18999 ( \19680 , \19678 , \19679 );
and \U$19000 ( \19681 , \17111 , \17169 );
not \U$19001 ( \19682 , \17111 );
and \U$19002 ( \19683 , \19682 , \17166 );
nor \U$19003 ( \19684 , \19681 , \19683 );
not \U$19004 ( \19685 , \19684 );
nand \U$19005 ( \19686 , \19685 , \16750 );
nand \U$19006 ( \19687 , \19680 , \19686 );
not \U$19007 ( \19688 , \18346 );
nand \U$19008 ( \19689 , \19688 , \18339 );
nand \U$19009 ( \19690 , \17061 , \17381 );
and \U$19010 ( \19691 , \19689 , \19690 );
xor \U$19011 ( \19692 , \19687 , \19691 );
not \U$19012 ( \19693 , \18278 );
not \U$19013 ( \19694 , \17303 );
or \U$19014 ( \19695 , \19693 , \19694 );
not \U$19015 ( \19696 , \17666 );
not \U$19016 ( \19697 , \16686 );
or \U$19017 ( \19698 , \19696 , \19697 );
nand \U$19018 ( \19699 , \16944 , \16683 );
nand \U$19019 ( \19700 , \19698 , \19699 );
nand \U$19020 ( \19701 , \19700 , \17118 );
nand \U$19021 ( \19702 , \19695 , \19701 );
xor \U$19022 ( \19703 , \19692 , \19702 );
not \U$19023 ( \19704 , \18356 );
not \U$19024 ( \19705 , \16573 );
not \U$19025 ( \19706 , \19705 );
or \U$19026 ( \19707 , \19704 , \19706 );
and \U$19027 ( \19708 , \16988 , \16574 );
not \U$19028 ( \19709 , \16988 );
and \U$19029 ( \19710 , \19709 , \17561 );
nor \U$19030 ( \19711 , \19708 , \19710 );
not \U$19031 ( \19712 , \19711 );
nand \U$19032 ( \19713 , \19712 , \16630 );
nand \U$19033 ( \19714 , \19707 , \19713 );
xor \U$19034 ( \19715 , \19703 , \19714 );
xor \U$19035 ( \19716 , \18271 , \18280 );
and \U$19036 ( \19717 , \19716 , \18290 );
and \U$19037 ( \19718 , \18271 , \18280 );
or \U$19038 ( \19719 , \19717 , \19718 );
xor \U$19039 ( \19720 , \19715 , \19719 );
xor \U$19040 ( \19721 , \18333 , \18364 );
and \U$19041 ( \19722 , \19721 , \18377 );
and \U$19042 ( \19723 , \18333 , \18364 );
or \U$19043 ( \19724 , \19722 , \19723 );
xor \U$19044 ( \19725 , \19720 , \19724 );
and \U$19045 ( \19726 , \17214 , \17507 );
not \U$19046 ( \19727 , \17214 );
and \U$19047 ( \19728 , \19727 , \16635 );
nor \U$19048 ( \19729 , \19726 , \19728 );
nand \U$19049 ( \19730 , \19105 , \19729 );
xor \U$19050 ( \19731 , \18337 , \18215 );
and \U$19051 ( \19732 , \19731 , \18348 );
and \U$19052 ( \19733 , \18337 , \18215 );
or \U$19053 ( \19734 , \19732 , \19733 );
xor \U$19054 ( \19735 , \19730 , \19734 );
not \U$19055 ( \19736 , \18288 );
not \U$19056 ( \19737 , \17402 );
or \U$19057 ( \19738 , \19736 , \19737 );
and \U$19058 ( \19739 , \16893 , \16825 );
and \U$19059 ( \19740 , \16894 , \16824 );
nor \U$19060 ( \19741 , \19739 , \19740 );
not \U$19061 ( \19742 , \19741 );
nand \U$19062 ( \19743 , \19742 , \17405 );
nand \U$19063 ( \19744 , \19738 , \19743 );
xnor \U$19064 ( \19745 , \19735 , \19744 );
xor \U$19065 ( \19746 , \18349 , \18358 );
and \U$19066 ( \19747 , \19746 , \18363 );
and \U$19067 ( \19748 , \18349 , \18358 );
or \U$19068 ( \19749 , \19747 , \19748 );
xor \U$19069 ( \19750 , \19745 , \19749 );
xor \U$19070 ( \19751 , \18224 , \18258 );
and \U$19071 ( \19752 , \19751 , \18291 );
and \U$19072 ( \19753 , \18224 , \18258 );
or \U$19073 ( \19754 , \19752 , \19753 );
xor \U$19074 ( \19755 , \19750 , \19754 );
xor \U$19075 ( \19756 , \19725 , \19755 );
xor \U$19076 ( \19757 , \18292 , \18328 );
and \U$19077 ( \19758 , \19757 , \18378 );
and \U$19078 ( \19759 , \18292 , \18328 );
or \U$19079 ( \19760 , \19758 , \19759 );
or \U$19080 ( \19761 , \19756 , \19760 );
xor \U$19081 ( \19762 , \19703 , \19714 );
and \U$19082 ( \19763 , \19762 , \19719 );
and \U$19083 ( \19764 , \19703 , \19714 );
or \U$19084 ( \19765 , \19763 , \19764 );
and \U$19085 ( \19766 , \16888 , \17639 );
not \U$19086 ( \19767 , \16888 );
and \U$19087 ( \19768 , \19767 , \16642 );
nor \U$19088 ( \19769 , \19766 , \19768 );
and \U$19089 ( \19770 , \16637 , \19769 );
not \U$19090 ( \19771 , \17402 );
not \U$19091 ( \19772 , \19771 );
not \U$19092 ( \19773 , \19741 );
and \U$19093 ( \19774 , \19772 , \19773 );
and \U$19094 ( \19775 , \16732 , \16894 );
not \U$19095 ( \19776 , \16732 );
and \U$19096 ( \19777 , \19776 , \16893 );
nor \U$19097 ( \19778 , \19775 , \19777 );
and \U$19098 ( \19779 , \17405 , \19778 );
nor \U$19099 ( \19780 , \19774 , \19779 );
xor \U$19100 ( \19781 , \19770 , \19780 );
not \U$19101 ( \19782 , \19700 );
not \U$19102 ( \19783 , \17303 );
or \U$19103 ( \19784 , \19782 , \19783 );
not \U$19104 ( \19785 , \16623 );
not \U$19105 ( \19786 , \17666 );
or \U$19106 ( \19787 , \19785 , \19786 );
nand \U$19107 ( \19788 , \16944 , \16624 );
nand \U$19108 ( \19789 , \19787 , \19788 );
nand \U$19109 ( \19790 , \19789 , \17118 );
nand \U$19110 ( \19791 , \19784 , \19790 );
xnor \U$19111 ( \19792 , \19781 , \19791 );
not \U$19112 ( \19793 , \19792 );
not \U$19113 ( \19794 , \19793 );
not \U$19114 ( \19795 , \19744 );
not \U$19115 ( \19796 , \19795 );
not \U$19116 ( \19797 , \19730 );
or \U$19117 ( \19798 , \19796 , \19797 );
nand \U$19118 ( \19799 , \19798 , \19734 );
not \U$19119 ( \19800 , \19730 );
nand \U$19120 ( \19801 , \19800 , \19744 );
and \U$19121 ( \19802 , \19799 , \19801 );
not \U$19122 ( \19803 , \19802 );
not \U$19123 ( \19804 , \19803 );
or \U$19124 ( \19805 , \19794 , \19804 );
nand \U$19125 ( \19806 , \19792 , \19802 );
nand \U$19126 ( \19807 , \19805 , \19806 );
and \U$19127 ( \19808 , \18340 , \17380 );
nor \U$19128 ( \19809 , \19808 , \17062 );
xor \U$19129 ( \19810 , \19691 , \19809 );
not \U$19130 ( \19811 , \16757 );
not \U$19131 ( \19812 , \19684 );
and \U$19132 ( \19813 , \19811 , \19812 );
and \U$19133 ( \19814 , \17342 , \16569 );
not \U$19134 ( \19815 , \17342 );
and \U$19135 ( \19816 , \19815 , \17166 );
nor \U$19136 ( \19817 , \19814 , \19816 );
nor \U$19137 ( \19818 , \19817 , \16751 );
nor \U$19138 ( \19819 , \19813 , \19818 );
xor \U$19139 ( \19820 , \19810 , \19819 );
or \U$19140 ( \19821 , \19687 , \19691 );
nand \U$19141 ( \19822 , \19821 , \19702 );
nand \U$19142 ( \19823 , \19687 , \19691 );
and \U$19143 ( \19824 , \19822 , \19823 );
xor \U$19144 ( \19825 , \19820 , \19824 );
nor \U$19145 ( \19826 , \16573 , \19711 );
not \U$19146 ( \19827 , \16630 );
and \U$19147 ( \19828 , \18267 , \16765 );
not \U$19148 ( \19829 , \18267 );
and \U$19149 ( \19830 , \19829 , \17561 );
nor \U$19150 ( \19831 , \19828 , \19830 );
nor \U$19151 ( \19832 , \19827 , \19831 );
nor \U$19152 ( \19833 , \19826 , \19832 );
xor \U$19153 ( \19834 , \19825 , \19833 );
not \U$19154 ( \19835 , \19834 );
and \U$19155 ( \19836 , \19807 , \19835 );
not \U$19156 ( \19837 , \19807 );
and \U$19157 ( \19838 , \19837 , \19834 );
nor \U$19158 ( \19839 , \19836 , \19838 );
xor \U$19159 ( \19840 , \19765 , \19839 );
xor \U$19160 ( \19841 , \19745 , \19749 );
and \U$19161 ( \19842 , \19841 , \19754 );
and \U$19162 ( \19843 , \19745 , \19749 );
or \U$19163 ( \19844 , \19842 , \19843 );
xor \U$19164 ( \19845 , \19840 , \19844 );
xor \U$19165 ( \19846 , \19720 , \19724 );
and \U$19166 ( \19847 , \19846 , \19755 );
and \U$19167 ( \19848 , \19720 , \19724 );
or \U$19168 ( \19849 , \19847 , \19848 );
nor \U$19169 ( \19850 , \19845 , \19849 );
not \U$19170 ( \19851 , \19850 );
xor \U$19171 ( \19852 , \19765 , \19839 );
and \U$19172 ( \19853 , \19852 , \19844 );
and \U$19173 ( \19854 , \19765 , \19839 );
or \U$19174 ( \19855 , \19853 , \19854 );
not \U$19175 ( \19856 , \19855 );
or \U$19176 ( \19857 , \16757 , \19817 );
and \U$19177 ( \19858 , \16825 , \17169 );
not \U$19178 ( \19859 , \16825 );
and \U$19179 ( \19860 , \19859 , \17395 );
nor \U$19180 ( \19861 , \19858 , \19860 );
or \U$19181 ( \19862 , \19861 , \16751 );
nand \U$19182 ( \19863 , \19857 , \19862 );
xor \U$19183 ( \19864 , \19691 , \19809 );
and \U$19184 ( \19865 , \19864 , \19819 );
and \U$19185 ( \19866 , \19691 , \19809 );
or \U$19186 ( \19867 , \19865 , \19866 );
xor \U$19187 ( \19868 , \19863 , \19867 );
not \U$19188 ( \19869 , \19831 );
and \U$19189 ( \19870 , \19705 , \19869 );
and \U$19190 ( \19871 , \17112 , \16766 );
not \U$19191 ( \19872 , \17112 );
and \U$19192 ( \19873 , \19872 , \16767 );
nor \U$19193 ( \19874 , \19871 , \19873 );
and \U$19194 ( \19875 , \19874 , \16630 );
nor \U$19195 ( \19876 , \19870 , \19875 );
xor \U$19196 ( \19877 , \19868 , \19876 );
nand \U$19197 ( \19878 , \19802 , \19793 );
nand \U$19198 ( \19879 , \19835 , \19878 );
nand \U$19199 ( \19880 , \19803 , \19792 );
and \U$19200 ( \19881 , \19879 , \19880 );
xor \U$19201 ( \19882 , \19877 , \19881 );
not \U$19202 ( \19883 , \19770 );
nand \U$19203 ( \19884 , \19883 , \19780 );
and \U$19204 ( \19885 , \19884 , \19791 );
nor \U$19205 ( \19886 , \19883 , \19780 );
nor \U$19206 ( \19887 , \19885 , \19886 );
and \U$19207 ( \19888 , \17303 , \19789 );
and \U$19208 ( \19889 , \16944 , \17118 );
nor \U$19209 ( \19890 , \19888 , \19889 );
not \U$19210 ( \19891 , \17809 );
and \U$19211 ( \19892 , \16893 , \16683 );
and \U$19212 ( \19893 , \16889 , \16686 );
nor \U$19213 ( \19894 , \19892 , \19893 );
not \U$19214 ( \19895 , \19894 );
and \U$19215 ( \19896 , \19891 , \19895 );
and \U$19216 ( \19897 , \17402 , \19778 );
nor \U$19217 ( \19898 , \19896 , \19897 );
xor \U$19218 ( \19899 , \19890 , \19898 );
and \U$19219 ( \19900 , \16642 , \16988 );
and \U$19220 ( \19901 , \16685 , \16989 );
nor \U$19221 ( \19902 , \19900 , \19901 );
nand \U$19222 ( \19903 , \16641 , \19902 );
xor \U$19223 ( \19904 , \19899 , \19903 );
xor \U$19224 ( \19905 , \19887 , \19904 );
xor \U$19225 ( \19906 , \19820 , \19824 );
and \U$19226 ( \19907 , \19906 , \19833 );
and \U$19227 ( \19908 , \19820 , \19824 );
or \U$19228 ( \19909 , \19907 , \19908 );
xor \U$19229 ( \19910 , \19905 , \19909 );
xor \U$19230 ( \19911 , \19882 , \19910 );
nand \U$19231 ( \19912 , \19856 , \19911 );
xor \U$19232 ( \19913 , \19877 , \19881 );
and \U$19233 ( \19914 , \19913 , \19910 );
and \U$19234 ( \19915 , \19877 , \19881 );
or \U$19235 ( \19916 , \19914 , \19915 );
not \U$19236 ( \19917 , \19863 );
and \U$19237 ( \19918 , \16642 , \18267 );
and \U$19238 ( \19919 , \17910 , \17406 );
nor \U$19239 ( \19920 , \19918 , \19919 );
nand \U$19240 ( \19921 , \16641 , \19920 );
xor \U$19241 ( \19922 , \19917 , \19921 );
and \U$19242 ( \19923 , \19705 , \19874 );
and \U$19243 ( \19924 , \17338 , \16767 );
not \U$19244 ( \19925 , \17338 );
and \U$19245 ( \19926 , \19925 , \16766 );
nor \U$19246 ( \19927 , \19924 , \19926 );
not \U$19247 ( \19928 , \19927 );
and \U$19248 ( \19929 , \19928 , \16630 );
nor \U$19249 ( \19930 , \19923 , \19929 );
xor \U$19250 ( \19931 , \19922 , \19930 );
xor \U$19251 ( \19932 , \19887 , \19904 );
and \U$19252 ( \19933 , \19932 , \19909 );
and \U$19253 ( \19934 , \19887 , \19904 );
or \U$19254 ( \19935 , \19933 , \19934 );
xor \U$19255 ( \19936 , \19931 , \19935 );
not \U$19256 ( \19937 , \19861 );
not \U$19257 ( \19938 , \19937 );
not \U$19258 ( \19939 , \16758 );
or \U$19259 ( \19940 , \19938 , \19939 );
and \U$19260 ( \19941 , \16731 , \17169 );
not \U$19261 ( \19942 , \16731 );
and \U$19262 ( \19943 , \19942 , \17395 );
nor \U$19263 ( \19944 , \19941 , \19943 );
nand \U$19264 ( \19945 , \19944 , \16750 );
nand \U$19265 ( \19946 , \19940 , \19945 );
not \U$19266 ( \19947 , \19946 );
not \U$19267 ( \19948 , \17303 );
nand \U$19268 ( \19949 , \19948 , \18718 );
and \U$19269 ( \19950 , \19949 , \16944 );
not \U$19270 ( \19951 , \19950 );
or \U$19271 ( \19952 , \19947 , \19951 );
or \U$19272 ( \19953 , \19950 , \19946 );
nand \U$19273 ( \19954 , \19952 , \19953 );
not \U$19274 ( \19955 , \19894 );
not \U$19275 ( \19956 , \19955 );
not \U$19276 ( \19957 , \17402 );
or \U$19277 ( \19958 , \19956 , \19957 );
or \U$19278 ( \19959 , \16889 , \16623 );
or \U$19279 ( \19960 , \16893 , \16624 );
nand \U$19280 ( \19961 , \19959 , \19960 );
nand \U$19281 ( \19962 , \17405 , \19961 );
nand \U$19282 ( \19963 , \19958 , \19962 );
xnor \U$19283 ( \19964 , \19954 , \19963 );
xor \U$19284 ( \19965 , \19890 , \19898 );
and \U$19285 ( \19966 , \19965 , \19903 );
and \U$19286 ( \19967 , \19890 , \19898 );
or \U$19287 ( \19968 , \19966 , \19967 );
xor \U$19288 ( \19969 , \19964 , \19968 );
xor \U$19289 ( \19970 , \19863 , \19867 );
and \U$19290 ( \19971 , \19970 , \19876 );
and \U$19291 ( \19972 , \19863 , \19867 );
or \U$19292 ( \19973 , \19971 , \19972 );
xor \U$19293 ( \19974 , \19969 , \19973 );
xor \U$19294 ( \19975 , \19936 , \19974 );
nand \U$19295 ( \19976 , \19916 , \19975 );
nand \U$19296 ( \19977 , \19761 , \19851 , \19912 , \19976 );
not \U$19297 ( \19978 , \19977 );
nand \U$19298 ( \19979 , \19677 , \19978 );
xor \U$19299 ( \19980 , \16782 , \16840 );
xor \U$19300 ( \19981 , \19980 , \16843 );
not \U$19301 ( \19982 , \19944 );
or \U$19302 ( \19983 , \16759 , \19982 );
and \U$19303 ( \19984 , \16569 , \16683 );
and \U$19304 ( \19985 , \16570 , \16686 );
nor \U$19305 ( \19986 , \19984 , \19985 );
or \U$19306 ( \19987 , \19986 , \16751 );
nand \U$19307 ( \19988 , \19983 , \19987 );
or \U$19308 ( \19989 , \16759 , \19986 );
or \U$19309 ( \19990 , \16779 , \16751 );
nand \U$19310 ( \19991 , \19989 , \19990 );
xor \U$19311 ( \19992 , \19988 , \19991 );
not \U$19312 ( \19993 , \17809 );
not \U$19313 ( \19994 , \19771 );
or \U$19314 ( \19995 , \19993 , \19994 );
nand \U$19315 ( \19996 , \19995 , \16890 );
and \U$19316 ( \19997 , \19992 , \19996 );
and \U$19317 ( \19998 , \19988 , \19991 );
or \U$19318 ( \19999 , \19997 , \19998 );
xor \U$19319 ( \20000 , \16783 , \16829 );
xor \U$19320 ( \20001 , \20000 , \16837 );
xor \U$19321 ( \20002 , \19999 , \20001 );
and \U$19322 ( \20003 , \16642 , \17342 );
and \U$19323 ( \20004 , \16685 , \17338 );
nor \U$19324 ( \20005 , \20003 , \20004 );
and \U$19325 ( \20006 , \16641 , \20005 );
and \U$19326 ( \20007 , \16825 , \16767 );
not \U$19327 ( \20008 , \16825 );
and \U$19328 ( \20009 , \20008 , \16766 );
nor \U$19329 ( \20010 , \20007 , \20009 );
not \U$19330 ( \20011 , \20010 );
not \U$19331 ( \20012 , \19705 );
or \U$19332 ( \20013 , \20011 , \20012 );
nand \U$19333 ( \20014 , \16833 , \16630 );
nand \U$19334 ( \20015 , \20013 , \20014 );
xor \U$19335 ( \20016 , \20006 , \20015 );
not \U$19336 ( \20017 , \19961 );
not \U$19337 ( \20018 , \17402 );
or \U$19338 ( \20019 , \20017 , \20018 );
nand \U$19339 ( \20020 , \17405 , \16890 );
nand \U$19340 ( \20021 , \20019 , \20020 );
not \U$19341 ( \20022 , \20021 );
and \U$19342 ( \20023 , \16642 , \17111 );
and \U$19343 ( \20024 , \17910 , \17112 );
nor \U$19344 ( \20025 , \20023 , \20024 );
nand \U$19345 ( \20026 , \16641 , \20025 );
not \U$19346 ( \20027 , \20026 );
not \U$19347 ( \20028 , \20027 );
or \U$19348 ( \20029 , \20022 , \20028 );
not \U$19349 ( \20030 , \20021 );
not \U$19350 ( \20031 , \20030 );
not \U$19351 ( \20032 , \20026 );
or \U$19352 ( \20033 , \20031 , \20032 );
not \U$19353 ( \20034 , \19988 );
nand \U$19354 ( \20035 , \20033 , \20034 );
nand \U$19355 ( \20036 , \20029 , \20035 );
and \U$19356 ( \20037 , \20016 , \20036 );
and \U$19357 ( \20038 , \20006 , \20015 );
or \U$19358 ( \20039 , \20037 , \20038 );
and \U$19359 ( \20040 , \20002 , \20039 );
and \U$19360 ( \20041 , \19999 , \20001 );
or \U$19361 ( \20042 , \20040 , \20041 );
nor \U$19362 ( \20043 , \19981 , \20042 );
not \U$19363 ( \20044 , \20043 );
xor \U$19364 ( \20045 , \19931 , \19935 );
and \U$19365 ( \20046 , \20045 , \19974 );
and \U$19366 ( \20047 , \19931 , \19935 );
or \U$19367 ( \20048 , \20046 , \20047 );
xor \U$19368 ( \20049 , \19988 , \20021 );
xor \U$19369 ( \20050 , \20049 , \20027 );
xor \U$19370 ( \20051 , \19917 , \19921 );
and \U$19371 ( \20052 , \20051 , \19930 );
and \U$19372 ( \20053 , \19917 , \19921 );
or \U$19373 ( \20054 , \20052 , \20053 );
not \U$19374 ( \20055 , \20054 );
not \U$19375 ( \20056 , \19962 );
not \U$19376 ( \20057 , \17402 );
nor \U$19377 ( \20058 , \20057 , \19894 );
nor \U$19378 ( \20059 , \20056 , \20058 , \19946 );
or \U$19379 ( \20060 , \20059 , \19950 );
nand \U$19380 ( \20061 , \19963 , \19946 );
nand \U$19381 ( \20062 , \20060 , \20061 );
not \U$19382 ( \20063 , \16573 );
not \U$19383 ( \20064 , \19927 );
and \U$19384 ( \20065 , \20063 , \20064 );
and \U$19385 ( \20066 , \20010 , \16630 );
nor \U$19386 ( \20067 , \20065 , \20066 );
xnor \U$19387 ( \20068 , \20062 , \20067 );
not \U$19388 ( \20069 , \20068 );
and \U$19389 ( \20070 , \20055 , \20069 );
and \U$19390 ( \20071 , \20054 , \20068 );
nor \U$19391 ( \20072 , \20070 , \20071 );
xor \U$19392 ( \20073 , \20050 , \20072 );
xor \U$19393 ( \20074 , \19964 , \19968 );
and \U$19394 ( \20075 , \20074 , \19973 );
and \U$19395 ( \20076 , \19964 , \19968 );
or \U$19396 ( \20077 , \20075 , \20076 );
xor \U$19397 ( \20078 , \20073 , \20077 );
nand \U$19398 ( \20079 , \20048 , \20078 );
xor \U$19399 ( \20080 , \19988 , \19991 );
xor \U$19400 ( \20081 , \20080 , \19996 );
xor \U$19401 ( \20082 , \20006 , \20015 );
xor \U$19402 ( \20083 , \20082 , \20036 );
xor \U$19403 ( \20084 , \20081 , \20083 );
not \U$19404 ( \20085 , \20067 );
not \U$19405 ( \20086 , \20054 );
or \U$19406 ( \20087 , \20085 , \20086 );
nand \U$19407 ( \20088 , \20087 , \20062 );
or \U$19408 ( \20089 , \20054 , \20067 );
nand \U$19409 ( \20090 , \20088 , \20089 );
xnor \U$19410 ( \20091 , \20084 , \20090 );
xor \U$19411 ( \20092 , \20050 , \20072 );
and \U$19412 ( \20093 , \20092 , \20077 );
and \U$19413 ( \20094 , \20050 , \20072 );
or \U$19414 ( \20095 , \20093 , \20094 );
nand \U$19415 ( \20096 , \20091 , \20095 );
nand \U$19416 ( \20097 , \20079 , \20096 );
not \U$19417 ( \20098 , \20081 );
not \U$19418 ( \20099 , \20083 );
or \U$19419 ( \20100 , \20098 , \20099 );
or \U$19420 ( \20101 , \20083 , \20081 );
nand \U$19421 ( \20102 , \20101 , \20090 );
nand \U$19422 ( \20103 , \20100 , \20102 );
xor \U$19423 ( \20104 , \19999 , \20001 );
xor \U$19424 ( \20105 , \20104 , \20039 );
nor \U$19425 ( \20106 , \20103 , \20105 );
nor \U$19426 ( \20107 , \20097 , \20106 );
nand \U$19427 ( \20108 , \20044 , \20107 );
or \U$19428 ( \20109 , \19979 , \20108 );
not \U$19429 ( \20110 , \19912 );
nand \U$19430 ( \20111 , \19756 , \19760 );
or \U$19431 ( \20112 , \20111 , \19850 );
nand \U$19432 ( \20113 , \19845 , \19849 );
nand \U$19433 ( \20114 , \20112 , \20113 );
not \U$19434 ( \20115 , \20114 );
or \U$19435 ( \20116 , \20110 , \20115 );
not \U$19436 ( \20117 , \19911 );
nand \U$19437 ( \20118 , \20117 , \19855 );
nand \U$19438 ( \20119 , \20116 , \20118 );
and \U$19439 ( \20120 , \20119 , \19976 );
nor \U$19440 ( \20121 , \19916 , \19975 );
nor \U$19441 ( \20122 , \20120 , \20121 );
not \U$19442 ( \20123 , \20122 );
not \U$19443 ( \20124 , \20108 );
and \U$19444 ( \20125 , \20123 , \20124 );
or \U$19445 ( \20126 , \20048 , \20078 );
not \U$19446 ( \20127 , \20096 );
or \U$19447 ( \20128 , \20126 , \20127 );
or \U$19448 ( \20129 , \20091 , \20095 );
nand \U$19449 ( \20130 , \20128 , \20129 );
not \U$19450 ( \20131 , \20106 );
and \U$19451 ( \20132 , \20130 , \20131 );
and \U$19452 ( \20133 , \20103 , \20105 );
nor \U$19453 ( \20134 , \20132 , \20133 );
or \U$19454 ( \20135 , \20134 , \20043 );
nand \U$19455 ( \20136 , \19981 , \20042 );
nand \U$19456 ( \20137 , \20135 , \20136 );
nor \U$19457 ( \20138 , \20125 , \20137 );
nand \U$19458 ( \20139 , \20109 , \20138 );
and \U$19459 ( \20140 , \16847 , \20139 );
and \U$19460 ( \20141 , \16776 , \16846 );
or \U$19461 ( \20142 , \20140 , \20141 );
xor \U$19462 ( \20143 , \16633 , \16689 );
and \U$19463 ( \20144 , \20143 , \16775 );
and \U$19464 ( \20145 , \16633 , \16689 );
or \U$19465 ( \20146 , \20144 , \20145 );
not \U$19466 ( \20147 , \16689 );
and \U$19467 ( \20148 , \16642 , \16624 );
and \U$19468 ( \20149 , \16685 , \16623 );
nor \U$19469 ( \20150 , \20148 , \20149 , \16640 );
not \U$19470 ( \20151 , \20150 );
and \U$19471 ( \20152 , \16573 , \16631 );
nor \U$19472 ( \20153 , \20152 , \16626 );
not \U$19473 ( \20154 , \20153 );
or \U$19474 ( \20155 , \20151 , \20154 );
or \U$19475 ( \20156 , \20153 , \20150 );
nand \U$19476 ( \20157 , \20155 , \20156 );
not \U$19477 ( \20158 , \20157 );
or \U$19478 ( \20159 , \20147 , \20158 );
or \U$19479 ( \20160 , \20157 , \16689 );
nand \U$19480 ( \20161 , \20159 , \20160 );
xor \U$19481 ( \20162 , \20146 , \20161 );
and \U$19482 ( \20163 , \20142 , \20162 );
not \U$19483 ( \20164 , \20142 );
xnor \U$19484 ( \20165 , \20146 , \20161 );
and \U$19485 ( \20166 , \20164 , \20165 );
nor \U$19486 ( \20167 , \20163 , \20166 );
nand \U$19487 ( \20168 , \16479 , \20167 );
nand \U$19488 ( \20169 , \16478 , \20168 );
buf \U$19489 ( \20170 , \20169 );
xor \U$19490 ( \20171 , \16776 , \16846 );
xor \U$19491 ( \20172 , \20171 , \20139 );
not \U$19492 ( \20173 , \20172 );
and \U$19493 ( \20174 , \16476 , \20173 );
not \U$19494 ( \20175 , \16476 );
nand \U$19495 ( \20176 , \15790 , \12134 );
buf \U$19496 ( \20177 , \15787 );
xor \U$19497 ( \20178 , \20176 , \20177 );
and \U$19498 ( \20179 , \20175 , \20178 );
nor \U$19499 ( \20180 , \20174 , \20179 );
buf \U$19500 ( \20181 , \20180 );
buf \U$19501 ( \20182 , \20122 );
not \U$19502 ( \20183 , \20182 );
not \U$19503 ( \20184 , \19979 );
or \U$19504 ( \20185 , \20183 , \20184 );
nand \U$19505 ( \20186 , \20185 , \20107 );
nand \U$19506 ( \20187 , \20186 , \20134 );
not \U$19507 ( \20188 , \20043 );
nand \U$19508 ( \20189 , \20188 , \20136 );
xor \U$19509 ( \20190 , \20187 , \20189 );
and \U$19510 ( \20191 , \16476 , \20190 );
not \U$19511 ( \20192 , \16476 );
not \U$19512 ( \20193 , \15725 );
and \U$19513 ( \20194 , \13652 , \15731 , \20193 );
buf \U$19514 ( \20195 , \20194 );
and \U$19515 ( \20196 , \14929 , \12901 );
and \U$19516 ( \20197 , \20195 , \20196 );
nand \U$19517 ( \20198 , \13652 , \15743 );
nand \U$19518 ( \20199 , \15741 , \12901 );
nor \U$19519 ( \20200 , \20198 , \20199 );
nor \U$19520 ( \20201 , \20197 , \20200 );
and \U$19521 ( \20202 , \13652 , \12901 );
not \U$19522 ( \20203 , \15221 );
not \U$19523 ( \20204 , \15237 );
and \U$19524 ( \20205 , \20203 , \20204 );
nor \U$19525 ( \20206 , \20205 , \15239 );
and \U$19526 ( \20207 , \20206 , \15731 , \14928 );
buf \U$19527 ( \20208 , \20207 );
and \U$19528 ( \20209 , \20202 , \20208 );
buf \U$19529 ( \20210 , \14780 );
nand \U$19530 ( \20211 , \20210 , \14928 );
not \U$19531 ( \20212 , \20211 );
and \U$19532 ( \20213 , \20202 , \20212 );
nor \U$19533 ( \20214 , \20209 , \20213 );
not \U$19534 ( \20215 , \12901 );
not \U$19535 ( \20216 , \20215 );
and \U$19536 ( \20217 , \20216 , \15766 );
nor \U$19537 ( \20218 , \20217 , \15781 );
nand \U$19538 ( \20219 , \13652 , \15745 );
not \U$19539 ( \20220 , \20219 );
not \U$19540 ( \20221 , \20215 );
and \U$19541 ( \20222 , \20220 , \20221 );
and \U$19542 ( \20223 , \14928 , \14787 );
and \U$19543 ( \20224 , \20202 , \20223 );
nor \U$19544 ( \20225 , \20222 , \20224 );
nand \U$19545 ( \20226 , \20201 , \20214 , \20218 , \20225 );
not \U$19546 ( \20227 , \15783 );
nand \U$19547 ( \20228 , \20227 , \12912 );
xor \U$19548 ( \20229 , \20226 , \20228 );
and \U$19549 ( \20230 , \20192 , \20229 );
nor \U$19550 ( \20231 , \20191 , \20230 );
buf \U$19551 ( \20232 , \20231 );
not \U$19552 ( \20233 , \20097 );
not \U$19553 ( \20234 , \20233 );
not \U$19554 ( \20235 , \19650 );
nand \U$19555 ( \20236 , \20235 , \19667 );
not \U$19556 ( \20237 , \18402 );
nand \U$19557 ( \20238 , \20236 , \20237 );
and \U$19558 ( \20239 , \20238 , \19668 );
buf \U$19559 ( \20240 , \18392 );
nor \U$19560 ( \20241 , \20239 , \20240 );
or \U$19561 ( \20242 , \20241 , \19652 );
nand \U$19562 ( \20243 , \20242 , \19978 );
not \U$19563 ( \20244 , \19645 );
not \U$19564 ( \20245 , \19659 );
nor \U$19565 ( \20246 , \20245 , \19665 );
nand \U$19566 ( \20247 , \20244 , \20246 );
not \U$19567 ( \20248 , \18404 );
nor \U$19568 ( \20249 , \20248 , \19977 );
nand \U$19569 ( \20250 , \20247 , \20249 );
nand \U$19570 ( \20251 , \20243 , \20250 , \20182 );
not \U$19571 ( \20252 , \20251 );
or \U$19572 ( \20253 , \20234 , \20252 );
not \U$19573 ( \20254 , \20130 );
nand \U$19574 ( \20255 , \20253 , \20254 );
nor \U$19575 ( \20256 , \20133 , \20106 );
xor \U$19576 ( \20257 , \20255 , \20256 );
not \U$19577 ( \20258 , \20257 );
not \U$19578 ( \20259 , \16476 );
or \U$19579 ( \20260 , \20258 , \20259 );
nand \U$19580 ( \20261 , \15769 , \15780 );
not \U$19581 ( \20262 , \20261 );
not \U$19582 ( \20263 , \12870 );
not \U$19583 ( \20264 , \20263 );
not \U$19584 ( \20265 , \20211 );
not \U$19585 ( \20266 , \13653 );
and \U$19586 ( \20267 , \20265 , \20266 );
and \U$19587 ( \20268 , \20194 , \14929 );
nor \U$19588 ( \20269 , \20267 , \20268 );
not \U$19589 ( \20270 , \20219 );
nor \U$19590 ( \20271 , \20270 , \15766 );
or \U$19591 ( \20272 , \20207 , \20223 );
not \U$19592 ( \20273 , \13653 );
nand \U$19593 ( \20274 , \20272 , \20273 );
not \U$19594 ( \20275 , \20198 );
nand \U$19595 ( \20276 , \20275 , \15741 );
nand \U$19596 ( \20277 , \20269 , \20271 , \20274 , \20276 );
not \U$19597 ( \20278 , \20277 );
or \U$19598 ( \20279 , \20264 , \20278 );
not \U$19599 ( \20280 , \15777 );
nand \U$19600 ( \20281 , \20279 , \20280 );
not \U$19601 ( \20282 , \20281 );
or \U$19602 ( \20283 , \20262 , \20282 );
or \U$19603 ( \20284 , \20261 , \20281 );
nand \U$19604 ( \20285 , \20283 , \20284 );
nand \U$19605 ( \20286 , \20285 , \16477 );
nand \U$19606 ( \20287 , \20260 , \20286 );
buf \U$19607 ( \20288 , \20287 );
not \U$19608 ( \20289 , \20079 );
buf \U$19609 ( \20290 , \20251 );
not \U$19610 ( \20291 , \20290 );
or \U$19611 ( \20292 , \20289 , \20291 );
nand \U$19612 ( \20293 , \20292 , \20126 );
nand \U$19613 ( \20294 , \20129 , \20096 );
xor \U$19614 ( \20295 , \20293 , \20294 );
and \U$19615 ( \20296 , \16476 , \20295 );
not \U$19616 ( \20297 , \16476 );
not \U$19617 ( \20298 , \12869 );
not \U$19618 ( \20299 , \20277 );
or \U$19619 ( \20300 , \20298 , \20299 );
nand \U$19620 ( \20301 , \20300 , \15773 );
not \U$19621 ( \20302 , \15776 );
nor \U$19622 ( \20303 , \20302 , \15774 );
xnor \U$19623 ( \20304 , \20301 , \20303 );
and \U$19624 ( \20305 , \20297 , \20304 );
nor \U$19625 ( \20306 , \20296 , \20305 );
buf \U$19626 ( \20307 , \20306 );
not \U$19627 ( \20308 , \16477 );
nand \U$19628 ( \20309 , \12869 , \15773 );
not \U$19629 ( \20310 , \20309 );
not \U$19630 ( \20311 , \20277 );
or \U$19631 ( \20312 , \20310 , \20311 );
or \U$19632 ( \20313 , \20277 , \20309 );
nand \U$19633 ( \20314 , \20312 , \20313 );
not \U$19634 ( \20315 , \20314 );
or \U$19635 ( \20316 , \20308 , \20315 );
nand \U$19636 ( \20317 , \20126 , \20079 );
not \U$19637 ( \20318 , \20317 );
not \U$19638 ( \20319 , \20290 );
or \U$19639 ( \20320 , \20318 , \20319 );
or \U$19640 ( \20321 , \20290 , \20317 );
nand \U$19641 ( \20322 , \20320 , \20321 );
nand \U$19642 ( \20323 , \20322 , \16476 );
nand \U$19643 ( \20324 , \20316 , \20323 );
buf \U$19644 ( \20325 , \20324 );
buf \U$19645 ( \20326 , \19761 );
nand \U$19646 ( \20327 , \19677 , \20326 );
not \U$19647 ( \20328 , \20327 );
not \U$19648 ( \20329 , \19850 );
and \U$19649 ( \20330 , \20328 , \20329 );
buf \U$19650 ( \20331 , \20114 );
nor \U$19651 ( \20332 , \20330 , \20331 );
not \U$19652 ( \20333 , \20332 );
and \U$19653 ( \20334 , \20333 , \19912 );
not \U$19654 ( \20335 , \20118 );
nor \U$19655 ( \20336 , \20334 , \20335 );
not \U$19656 ( \20337 , \20121 );
nand \U$19657 ( \20338 , \20337 , \19976 );
and \U$19658 ( \20339 , \20336 , \20338 );
not \U$19659 ( \20340 , \20336 );
not \U$19660 ( \20341 , \20338 );
and \U$19661 ( \20342 , \20340 , \20341 );
or \U$19662 ( \20343 , \20339 , \20342 );
and \U$19663 ( \20344 , \16476 , \20343 );
not \U$19664 ( \20345 , \16476 );
not \U$19665 ( \20346 , \15759 );
not \U$19666 ( \20347 , \20346 );
not \U$19667 ( \20348 , \13617 );
not \U$19668 ( \20349 , \15747 );
or \U$19669 ( \20350 , \20348 , \20349 );
buf \U$19670 ( \20351 , \15758 );
nand \U$19671 ( \20352 , \20350 , \20351 );
not \U$19672 ( \20353 , \20352 );
or \U$19673 ( \20354 , \20347 , \20353 );
nand \U$19674 ( \20355 , \20354 , \15761 );
nand \U$19675 ( \20356 , \15765 , \15752 );
xor \U$19676 ( \20357 , \20355 , \20356 );
and \U$19677 ( \20358 , \20345 , \20357 );
nor \U$19678 ( \20359 , \20344 , \20358 );
buf \U$19679 ( \20360 , \20359 );
nand \U$19680 ( \20361 , \20118 , \19912 );
xnor \U$19681 ( \20362 , \20332 , \20361 );
and \U$19682 ( \20363 , \16476 , \20362 );
not \U$19683 ( \20364 , \16476 );
nand \U$19684 ( \20365 , \15761 , \20346 );
xor \U$19685 ( \20366 , \20352 , \20365 );
and \U$19686 ( \20367 , \20364 , \20366 );
nor \U$19687 ( \20368 , \20363 , \20367 );
buf \U$19688 ( \20369 , \20368 );
nand \U$19689 ( \20370 , \20327 , \20111 );
nand \U$19690 ( \20371 , \20113 , \19851 );
xor \U$19691 ( \20372 , \20370 , \20371 );
and \U$19692 ( \20373 , \16476 , \20372 );
not \U$19693 ( \20374 , \16476 );
not \U$19694 ( \20375 , \13616 );
not \U$19695 ( \20376 , \20375 );
buf \U$19696 ( \20377 , \15747 );
not \U$19697 ( \20378 , \20377 );
or \U$19698 ( \20379 , \20376 , \20378 );
not \U$19699 ( \20380 , \15755 );
nand \U$19700 ( \20381 , \20379 , \20380 );
not \U$19701 ( \20382 , \15754 );
nand \U$19702 ( \20383 , \20382 , \15757 );
xor \U$19703 ( \20384 , \20381 , \20383 );
and \U$19704 ( \20385 , \20374 , \20384 );
nor \U$19705 ( \20386 , \20373 , \20385 );
buf \U$19706 ( \20387 , \20386 );
not \U$19707 ( \20388 , \16475 );
not \U$19708 ( \20389 , \13616 );
nand \U$19709 ( \20390 , \20389 , \20380 );
xnor \U$19710 ( \20391 , \20377 , \20390 );
not \U$19711 ( \20392 , \20391 );
or \U$19712 ( \20393 , \20388 , \20392 );
nand \U$19713 ( \20394 , \20111 , \20326 );
xnor \U$19714 ( \20395 , \19677 , \20394 );
nand \U$19715 ( \20396 , \20395 , \16476 );
nand \U$19716 ( \20397 , \20393 , \20396 );
buf \U$19717 ( \20398 , \20397 );
not \U$19718 ( \20399 , \20237 );
not \U$19719 ( \20400 , \18206 );
not \U$19720 ( \20401 , \20247 );
or \U$19721 ( \20402 , \20400 , \20401 );
not \U$19722 ( \20403 , \20236 );
nand \U$19723 ( \20404 , \20402 , \20403 );
not \U$19724 ( \20405 , \20404 );
or \U$19725 ( \20406 , \20399 , \20405 );
nand \U$19726 ( \20407 , \20406 , \19668 );
nor \U$19727 ( \20408 , \19652 , \20240 );
xnor \U$19728 ( \20409 , \20407 , \20408 );
and \U$19729 ( \20410 , \16476 , \20409 );
not \U$19730 ( \20411 , \16476 );
not \U$19731 ( \20412 , \14912 );
buf \U$19732 ( \20413 , \14887 );
buf \U$19733 ( \20414 , \14919 );
and \U$19734 ( \20415 , \20413 , \20414 );
not \U$19735 ( \20416 , \20415 );
not \U$19736 ( \20417 , \15730 );
nand \U$19737 ( \20418 , \20417 , \15726 );
buf \U$19738 ( \20419 , \14779 );
or \U$19739 ( \20420 , \20418 , \20419 );
not \U$19740 ( \20421 , \14789 );
nand \U$19741 ( \20422 , \20420 , \20421 );
not \U$19742 ( \20423 , \20422 );
or \U$19743 ( \20424 , \20416 , \20423 );
not \U$19744 ( \20425 , \15737 );
nor \U$19745 ( \20426 , \20425 , \15739 );
nand \U$19746 ( \20427 , \20424 , \20426 );
not \U$19747 ( \20428 , \20427 );
or \U$19748 ( \20429 , \20412 , \20428 );
not \U$19749 ( \20430 , \15738 );
nand \U$19750 ( \20431 , \20429 , \20430 );
nand \U$19751 ( \20432 , \15746 , \15742 );
not \U$19752 ( \20433 , \20432 );
and \U$19753 ( \20434 , \20431 , \20433 );
not \U$19754 ( \20435 , \20431 );
and \U$19755 ( \20436 , \20435 , \20432 );
nor \U$19756 ( \20437 , \20434 , \20436 );
not \U$19757 ( \20438 , \20437 );
and \U$19758 ( \20439 , \20411 , \20438 );
nor \U$19759 ( \20440 , \20410 , \20439 );
buf \U$19760 ( \20441 , \20440 );
nand \U$19761 ( \20442 , \19668 , \20237 );
xor \U$19762 ( \20443 , \20404 , \20442 );
and \U$19763 ( \20444 , \16476 , \20443 );
not \U$19764 ( \20445 , \16476 );
nand \U$19765 ( \20446 , \20430 , \14912 );
xor \U$19766 ( \20447 , \20446 , \20427 );
and \U$19767 ( \20448 , \20445 , \20447 );
nor \U$19768 ( \20449 , \20444 , \20448 );
buf \U$19769 ( \20450 , \20449 );
not \U$19770 ( \20451 , \18205 );
not \U$19771 ( \20452 , \20247 );
or \U$19772 ( \20453 , \20451 , \20452 );
not \U$19773 ( \20454 , \19649 );
nand \U$19774 ( \20455 , \20453 , \20454 );
nand \U$19775 ( \20456 , \18032 , \19667 );
xor \U$19776 ( \20457 , \20455 , \20456 );
and \U$19777 ( \20458 , \16476 , \20457 );
not \U$19778 ( \20459 , \16476 );
not \U$19779 ( \20460 , \20414 );
buf \U$19780 ( \20461 , \20422 );
not \U$19781 ( \20462 , \20461 );
or \U$19782 ( \20463 , \20460 , \20462 );
not \U$19783 ( \20464 , \15736 );
nand \U$19784 ( \20465 , \20463 , \20464 );
not \U$19785 ( \20466 , \20413 );
nor \U$19786 ( \20467 , \20466 , \15739 );
and \U$19787 ( \20468 , \20465 , \20467 );
not \U$19788 ( \20469 , \20465 );
not \U$19789 ( \20470 , \20467 );
and \U$19790 ( \20471 , \20469 , \20470 );
nor \U$19791 ( \20472 , \20468 , \20471 );
not \U$19792 ( \20473 , \20472 );
and \U$19793 ( \20474 , \20459 , \20473 );
nor \U$19794 ( \20475 , \20458 , \20474 );
buf \U$19795 ( \20476 , \20475 );
nand \U$19796 ( \20477 , \20454 , \18205 );
xor \U$19797 ( \20478 , \20247 , \20477 );
and \U$19798 ( \20479 , \16476 , \20478 );
not \U$19799 ( \20480 , \16476 );
not \U$19800 ( \20481 , \15736 );
nand \U$19801 ( \20482 , \20481 , \20414 );
xor \U$19802 ( \20483 , \20482 , \20461 );
and \U$19803 ( \20484 , \20480 , \20483 );
nor \U$19804 ( \20485 , \20479 , \20484 );
buf \U$19805 ( \20486 , \20485 );
not \U$19806 ( \20487 , \19642 );
not \U$19807 ( \20488 , \19602 );
and \U$19808 ( \20489 , \19527 , \19612 );
not \U$19809 ( \20490 , \20489 );
or \U$19810 ( \20491 , \20488 , \20490 );
not \U$19811 ( \20492 , \19658 );
nand \U$19812 ( \20493 , \20491 , \20492 );
not \U$19813 ( \20494 , \20493 );
or \U$19814 ( \20495 , \20487 , \20494 );
not \U$19815 ( \20496 , \19660 );
nand \U$19816 ( \20497 , \20495 , \20496 );
nand \U$19817 ( \20498 , \19664 , \19632 );
xor \U$19818 ( \20499 , \20497 , \20498 );
and \U$19819 ( \20500 , \16476 , \20499 );
not \U$19820 ( \20501 , \16476 );
buf \U$19821 ( \20502 , \14689 );
not \U$19822 ( \20503 , \20502 );
buf \U$19823 ( \20504 , \14449 );
nand \U$19824 ( \20505 , \20504 , \14569 );
nand \U$19825 ( \20506 , \20418 , \20505 );
not \U$19826 ( \20507 , \20506 );
or \U$19827 ( \20508 , \20503 , \20507 );
not \U$19828 ( \20509 , \14782 );
nand \U$19829 ( \20510 , \20508 , \20509 );
nand \U$19830 ( \20511 , \14786 , \14778 );
xor \U$19831 ( \20512 , \20510 , \20511 );
and \U$19832 ( \20513 , \20501 , \20512 );
nor \U$19833 ( \20514 , \20500 , \20513 );
buf \U$19834 ( \20515 , \20514 );
and \U$19835 ( \20516 , \20496 , \19642 );
xnor \U$19836 ( \20517 , \20516 , \20493 );
and \U$19837 ( \20518 , \16476 , \20517 );
not \U$19838 ( \20519 , \16476 );
nand \U$19839 ( \20520 , \20509 , \20502 );
xor \U$19840 ( \20521 , \20506 , \20520 );
and \U$19841 ( \20522 , \20519 , \20521 );
nor \U$19842 ( \20523 , \20518 , \20522 );
buf \U$19843 ( \20524 , \20523 );
not \U$19844 ( \20525 , \20489 );
nand \U$19845 ( \20526 , \20525 , \19655 );
nand \U$19846 ( \20527 , \19602 , \19656 );
xor \U$19847 ( \20528 , \20526 , \20527 );
and \U$19848 ( \20529 , \16476 , \20528 );
not \U$19849 ( \20530 , \16476 );
not \U$19850 ( \20531 , \15729 );
not \U$19851 ( \20532 , \15726 );
or \U$19852 ( \20533 , \20531 , \20532 );
nand \U$19853 ( \20534 , \20533 , \14568 );
nand \U$19854 ( \20535 , \20504 , \14450 );
xor \U$19855 ( \20536 , \20534 , \20535 );
and \U$19856 ( \20537 , \20530 , \20536 );
nor \U$19857 ( \20538 , \20529 , \20537 );
buf \U$19858 ( \20539 , \20538 );
not \U$19859 ( \20540 , \16475 );
nand \U$19860 ( \20541 , \14568 , \15729 );
not \U$19861 ( \20542 , \20541 );
not \U$19862 ( \20543 , \15726 );
or \U$19863 ( \20544 , \20542 , \20543 );
or \U$19864 ( \20545 , \20541 , \15726 );
nand \U$19865 ( \20546 , \20544 , \20545 );
not \U$19866 ( \20547 , \20546 );
or \U$19867 ( \20548 , \20540 , \20547 );
nand \U$19868 ( \20549 , \19655 , \19612 );
not \U$19869 ( \20550 , \20549 );
buf \U$19870 ( \20551 , \19527 );
not \U$19871 ( \20552 , \20551 );
or \U$19872 ( \20553 , \20550 , \20552 );
or \U$19873 ( \20554 , \20551 , \20549 );
nand \U$19874 ( \20555 , \20553 , \20554 );
nand \U$19875 ( \20556 , \20555 , \16476 );
nand \U$19876 ( \20557 , \20548 , \20556 );
buf \U$19877 ( \20558 , \20557 );
not \U$19878 ( \20559 , \19045 );
not \U$19879 ( \20560 , \20559 );
not \U$19880 ( \20561 , \19512 );
or \U$19881 ( \20562 , \20560 , \20561 );
not \U$19882 ( \20563 , \19518 );
nand \U$19883 ( \20564 , \20562 , \20563 );
not \U$19884 ( \20565 , \18905 );
and \U$19885 ( \20566 , \20564 , \20565 );
not \U$19886 ( \20567 , \19521 );
nor \U$19887 ( \20568 , \20566 , \20567 );
nand \U$19888 ( \20569 , \19125 , \19526 );
xor \U$19889 ( \20570 , \20568 , \20569 );
not \U$19890 ( \20571 , \20570 );
nor \U$19891 ( \20572 , \20571 , \16475 );
not \U$19892 ( \20573 , \20572 );
nand \U$19893 ( \20574 , \15236 , \15240 );
not \U$19894 ( \20575 , \20574 );
buf \U$19895 ( \20576 , \15062 );
not \U$19896 ( \20577 , \20576 );
not \U$19897 ( \20578 , \15724 );
not \U$19898 ( \20579 , \15720 );
or \U$19899 ( \20580 , \20578 , \20579 );
nand \U$19900 ( \20581 , \20580 , \15220 );
not \U$19901 ( \20582 , \20581 );
or \U$19902 ( \20583 , \20577 , \20582 );
buf \U$19903 ( \20584 , \15223 );
nand \U$19904 ( \20585 , \20583 , \20584 );
not \U$19905 ( \20586 , \20585 );
or \U$19906 ( \20587 , \20575 , \20586 );
or \U$19907 ( \20588 , \20585 , \20574 );
nand \U$19908 ( \20589 , \20587 , \20588 );
nand \U$19909 ( \20590 , \20589 , \16475 );
nand \U$19910 ( \20591 , \20573 , \20590 );
buf \U$19911 ( \20592 , \20591 );
nand \U$19912 ( \20593 , \20565 , \19521 );
xnor \U$19913 ( \20594 , \20564 , \20593 );
and \U$19914 ( \20595 , \16476 , \20594 );
not \U$19915 ( \20596 , \16476 );
nand \U$19916 ( \20597 , \20576 , \20584 );
not \U$19917 ( \20598 , \20597 );
not \U$19918 ( \20599 , \20581 );
or \U$19919 ( \20600 , \20598 , \20599 );
or \U$19920 ( \20601 , \20597 , \20581 );
nand \U$19921 ( \20602 , \20600 , \20601 );
and \U$19922 ( \20603 , \20596 , \20602 );
or \U$19923 ( \20604 , \20595 , \20603 );
buf \U$19924 ( \20605 , \20604 );
and \U$19925 ( \20606 , \19512 , \19044 );
nor \U$19926 ( \20607 , \20606 , \19514 );
nand \U$19927 ( \20608 , \19517 , \18983 );
and \U$19928 ( \20609 , \20607 , \20608 );
not \U$19929 ( \20610 , \20607 );
not \U$19930 ( \20611 , \20608 );
and \U$19931 ( \20612 , \20610 , \20611 );
nor \U$19932 ( \20613 , \20609 , \20612 );
not \U$19933 ( \20614 , \20613 );
nor \U$19934 ( \20615 , \20614 , \16475 );
not \U$19935 ( \20616 , \20615 );
nand \U$19936 ( \20617 , \15154 , \15219 );
not \U$19937 ( \20618 , \20617 );
not \U$19938 ( \20619 , \15723 );
not \U$19939 ( \20620 , \15720 );
or \U$19940 ( \20621 , \20619 , \20620 );
buf \U$19941 ( \20622 , \15216 );
nand \U$19942 ( \20623 , \20621 , \20622 );
not \U$19943 ( \20624 , \20623 );
or \U$19944 ( \20625 , \20618 , \20624 );
or \U$19945 ( \20626 , \20623 , \20617 );
nand \U$19946 ( \20627 , \20625 , \20626 );
nand \U$19947 ( \20628 , \20627 , \16475 );
nand \U$19948 ( \20629 , \20616 , \20628 );
buf \U$19949 ( \20630 , \20629 );
not \U$19950 ( \20631 , \19514 );
nand \U$19951 ( \20632 , \20631 , \19044 );
xnor \U$19952 ( \20633 , \19512 , \20632 );
and \U$19953 ( \20634 , \16476 , \20633 );
not \U$19954 ( \20635 , \16476 );
nand \U$19955 ( \20636 , \20622 , \15723 );
not \U$19956 ( \20637 , \20636 );
and \U$19957 ( \20638 , \15720 , \20637 );
not \U$19958 ( \20639 , \15720 );
and \U$19959 ( \20640 , \20639 , \20636 );
nor \U$19960 ( \20641 , \20638 , \20640 );
and \U$19961 ( \20642 , \20635 , \20641 );
or \U$19962 ( \20643 , \20634 , \20642 );
buf \U$19963 ( \20644 , \20643 );
not \U$19964 ( \20645 , \16475 );
nand \U$19965 ( \20646 , \15306 , \15719 );
not \U$19966 ( \20647 , \20646 );
or \U$19967 ( \20648 , \15705 , \15714 );
not \U$19968 ( \20649 , \20648 );
not \U$19969 ( \20650 , \15703 );
or \U$19970 ( \20651 , \20649 , \20650 );
not \U$19971 ( \20652 , \15717 );
nand \U$19972 ( \20653 , \20651 , \20652 );
not \U$19973 ( \20654 , \20653 );
or \U$19974 ( \20655 , \20647 , \20654 );
or \U$19975 ( \20656 , \20653 , \20646 );
nand \U$19976 ( \20657 , \20655 , \20656 );
not \U$19977 ( \20658 , \20657 );
or \U$19978 ( \20659 , \20645 , \20658 );
xor \U$19979 ( \20660 , \19192 , \19197 );
xor \U$19980 ( \20661 , \20660 , \19509 );
nand \U$19981 ( \20662 , \20661 , \16476 );
nand \U$19982 ( \20663 , \20659 , \20662 );
buf \U$19983 ( \20664 , \20663 );
not \U$19984 ( \20665 , \16475 );
nand \U$19985 ( \20666 , \20652 , \15715 );
xnor \U$19986 ( \20667 , \15703 , \20666 );
not \U$19987 ( \20668 , \20667 );
or \U$19988 ( \20669 , \20665 , \20668 );
xor \U$19989 ( \20670 , \19239 , \19241 );
xor \U$19990 ( \20671 , \20670 , \19506 );
nand \U$19991 ( \20672 , \20671 , \16476 );
nand \U$19992 ( \20673 , \20669 , \20672 );
buf \U$19993 ( \20674 , \20673 );
xor \U$19994 ( \20675 , \19277 , \19279 );
xor \U$19995 ( \20676 , \20675 , \19503 );
and \U$19996 ( \20677 , \16476 , \20676 );
not \U$19997 ( \20678 , \16476 );
xor \U$19998 ( \20679 , \15390 , \15423 );
xor \U$19999 ( \20680 , \20679 , \15700 );
and \U$20000 ( \20681 , \20678 , \20680 );
or \U$20001 ( \20682 , \20677 , \20681 );
buf \U$20002 ( \20683 , \20682 );
not \U$20003 ( \20684 , \16475 );
nand \U$20004 ( \20685 , \15699 , \15489 );
not \U$20005 ( \20686 , \20685 );
buf \U$20006 ( \20687 , \15695 );
not \U$20007 ( \20688 , \20687 );
or \U$20008 ( \20689 , \20686 , \20688 );
or \U$20009 ( \20690 , \20687 , \20685 );
nand \U$20010 ( \20691 , \20689 , \20690 );
not \U$20011 ( \20692 , \20691 );
or \U$20012 ( \20693 , \20684 , \20692 );
nand \U$20013 ( \20694 , \19332 , \19502 );
buf \U$20014 ( \20695 , \19498 );
xnor \U$20015 ( \20696 , \20694 , \20695 );
nand \U$20016 ( \20697 , \20696 , \16476 );
nand \U$20017 ( \20698 , \20693 , \20697 );
buf \U$20018 ( \20699 , \20698 );
and \U$20019 ( \20700 , \15694 , \15690 );
buf \U$20020 ( \20701 , \15674 );
xor \U$20021 ( \20702 , \20700 , \20701 );
and \U$20022 ( \20703 , \16475 , \20702 );
not \U$20023 ( \20704 , \16475 );
not \U$20024 ( \20705 , \19366 );
nand \U$20025 ( \20706 , \20705 , \19497 );
and \U$20026 ( \20707 , \20706 , \19495 );
not \U$20027 ( \20708 , \20706 );
and \U$20028 ( \20709 , \20708 , \19494 );
nor \U$20029 ( \20710 , \20707 , \20709 );
and \U$20030 ( \20711 , \20704 , \20710 );
or \U$20031 ( \20712 , \20703 , \20711 );
buf \U$20032 ( \20713 , \20712 );
endmodule

