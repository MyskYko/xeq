//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RI994e3e8_15,RI994e370_16,RI994e2f8_17,RI994e280_18,RI994e208_19,RI994e190_20,RI994e118_21,RI994e0a0_22,RI994e028_23,
        RI994dfb0_24,RI994df38_25,RI995e450_236,RI9921730_613,RI99217a8_612,RI9921820_611,RI9921898_610,RI9921910_609,RI9921988_608,RI9921a00_607,
        RI9921a78_606,RI9921af0_605,RI9921b68_604,RI9921be0_603,RI9921c58_602,RI9921cd0_601,RI9967078_223,RI9967690_210,RI890fba0_197,RI8918b88_184,
        RI89253b0_171,RI8930dc8_158,RI8939db0_145,RI89465d8_132,RI89ec640_119,RI9776f80_106,RI9808480_93,RI9808a98_80,RI9819730_67,RI98abc38_54,
        RI98bc8d0_41,RI994ddd0_28,RI995e3d8_237,RI99669e8_224,RI9967618_211,RI890fb28_198,RI8918b10_185,RI8925338_172,RI8930d50_159,RI8939d38_146,
        RI8946560_133,RI89ec5c8_120,RI9776f08_107,RI9808408_94,RI9808a20_81,RI98196b8_68,RI98abbc0_55,RI98bc858_42,RI994dd58_29,RI9959fe0_238,
        RI995e978_225,RI99675a0_212,RI890fab0_199,RI8918a98_186,RI89252c0_173,RI8930cd8_160,RI8939cc0_147,RI89464e8_134,RI89ec550_121,RI9776e90_108,
        RI9808390_95,RI98089a8_82,RI9819640_69,RI98abb48_56,RI98bc7e0_43,RI994dce0_30,RI9959f68_239,RI995e900_226,RI9967528_213,RI890fa38_200,
        RI8918a20_187,RI8925248_174,RI8930c60_161,RI8939c48_148,RI8946470_135,RI89ec4d8_122,RI9776e18_109,RI9808318_96,RI9808930_83,RI98195c8_70,
        RI98abad0_57,RI98bc768_44,RI994dc68_31,RI9959860_240,RI995e888_227,RI99674b0_214,RI890f9c0_201,RI89189a8_188,RI89251d0_175,RI8930be8_162,
        RI8939bd0_149,RI89463f8_136,RI89ec460_123,RI9776da0_110,RI98082a0_97,RI98088b8_84,RI9819550_71,RI98aba58_58,RI98bc6f0_45,RI994dbf0_32,
        RI994d998_241,RI995e810_228,RI9967438_215,RI890f948_202,RI8918930_189,RI8925158_176,RI8930b70_163,RI8939b58_150,RI8946380_137,RI89ec3e8_124,
        RI9776d28_111,RI9808228_98,RI9808840_85,RI98194d8_72,RI98ab9e0_59,RI98abff8_46,RI98bcc90_33,RI994d920_242,RI995e798_229,RI99673c0_216,
        RI890f8d0_203,RI89188b8_190,RI89250e0_177,RI8930af8_164,RI8939ae0_151,RI8946308_138,RI89ec370_125,RI89ec988_112,RI97772c8_99,RI98087c8_86,
        RI9819460_73,RI98ab968_60,RI98abf80_47,RI98bcc18_34,RI994d8a8_243,RI995e720_230,RI9967348_217,RI890f858_204,RI8918840_191,RI8925068_178,
        RI8930a80_165,RI8939a68_152,RI8946290_139,RI89ec2f8_126,RI89ec910_113,RI9777250_100,RI9808750_87,RI98193e8_74,RI98ab8f0_61,RI98abf08_48,
        RI98bcba0_35,RI994d830_244,RI995e6a8_231,RI99672d0_218,RI890f7e0_205,RI89187c8_192,RI8924ff0_179,RI8930a08_166,RI89399f0_153,RI8946218_140,
        RI89ec280_127,RI89ec898_114,RI97771d8_101,RI98086d8_88,RI9819370_75,RI98ab878_62,RI98abe90_49,RI98bcb28_36,RI994d7b8_245,RI995e630_232,
        RI9967258_219,RI890f768_206,RI8918750_193,RI8924f78_180,RI8930990_167,RI8939978_154,RI89461a0_141,RI89ec208_128,RI89ec820_115,RI9777160_102,
        RI9808660_89,RI98192f8_76,RI98ab800_63,RI98abe18_50,RI98bcab0_37,RI994d740_246,RI995e5b8_233,RI99671e0_220,RI890f6f0_207,RI89186d8_194,
        RI8924f00_181,RI8930918_168,RI8939900_155,RI8946128_142,RI89ec190_129,RI89ec7a8_116,RI97770e8_103,RI98085e8_90,RI9819280_77,RI98ab788_64,
        RI98abda0_51,RI98bca38_38,RI994dec0_26,RI994d6c8_247,RI995e540_234,RI9967168_221,RI890f678_208,RI8918660_195,RI8924e88_182,RI89308a0_169,
        RI8939888_156,RI89460b0_143,RI89ec118_130,RI89ec730_117,RI9777070_104,RI9808570_91,RI9819208_78,RI98ab710_65,RI98abd28_52,RI98bc9c0_39,
        RI9922bd0_569,RI9923800_549,RI9924160_529,RI9924ac0_509,RI9925ab0_489,RI9926410_469,RI9926d70_449,RI9928120_429,RI9928a80_409,RI992a1f0_389,
        RI992ab50_369,RI992b4b0_349,RI992cfe0_329,RI992eed0_309,RI992f830_289,RI9931ae0_269,RI994d5d8_249,RI994e460_14,RI995e4c8_235,RI99670f0_222,
        RI890f600_209,RI89185e8_196,RI8924e10_183,RI8930828_170,RI8939810_157,RI8946038_144,RI89ec0a0_131,RI89ec6b8_118,RI9776ff8_105,RI98084f8_92,
        RI9808b10_79,RI98197a8_66,RI98abcb0_53,RI98bc948_40,RI994de48_27,RI9922f18_568,RI9923878_548,RI99241d8_528,RI9924b38_508,RI9925b28_488,
        RI9926488_468,RI9926de8_448,RI9928198_428,RI9928af8_408,RI992a268_388,RI992abc8_368,RI992c6f8_348,RI992d058_328,RI992ef48_308,RI992f8a8_288,
        RI9931b58_268,RI994d650_248,RI9922b58_570,RI9923788_550,RI99240e8_530,RI9924a48_510,RI9925a38_490,RI9926398_470,RI9926cf8_450,RI99280a8_430,
        RI9928a08_410,RI992a178_390,RI992aad8_370,RI992b438_350,RI992cf68_330,RI992ee58_310,RI992f7b8_290,RI9931a68_270,RI994d560_250,RI9922a68_572,
        RI9923698_552,RI9923ff8_532,RI9924958_512,RI9925948_492,RI99262a8_472,RI9926c08_452,RI9927fb8_432,RI9928918_412,RI9929278_392,RI992a9e8_372,
        RI992b348_352,RI992ce78_332,RI992ed68_312,RI992f6c8_292,RI9931978_272,RI994d470_252,RI9922ae0_571,RI9923710_551,RI9924070_531,RI99249d0_511,
        RI99259c0_491,RI9926320_471,RI9926c80_451,RI9928030_431,RI9928990_411,RI992a100_391,RI992aa60_371,RI992b3c0_351,RI992cef0_331,RI992ede0_311,
        RI992f740_291,RI99319f0_271,RI994d4e8_251,RI99229f0_573,RI9923620_553,RI9923f80_533,RI99248e0_513,RI99258d0_493,RI9926230_473,RI9926b90_453,
        RI9927f40_433,RI99288a0_413,RI9929200_393,RI992a970_373,RI992b2d0_353,RI992ce00_333,RI992ecf0_313,RI992f650_293,RI9931900_273,RI994d3f8_253,
        RI9922900_575,RI9923530_555,RI9923e90_535,RI99247f0_515,RI99257e0_495,RI9926140_475,RI9926aa0_455,RI9927e50_435,RI99287b0_415,RI9929110_395,
        RI992a880_375,RI992b1e0_355,RI992cd10_335,RI992d670_315,RI992f560_295,RI9931810_275,RI9935f50_255,RI9922978_574,RI99235a8_554,RI9923f08_534,
        RI9924868_514,RI9925858_494,RI99261b8_474,RI9926b18_454,RI9927ec8_434,RI9928828_414,RI9929188_394,RI992a8f8_374,RI992b258_354,RI992cd88_334,
        RI992d6e8_314,RI992f5d8_294,RI9931888_274,RI9935fc8_254,RI9922810_577,RI9923440_557,RI9923da0_537,RI9924700_517,RI99256f0_497,RI9926050_477,
        RI99269b0_457,RI9927d60_437,RI99286c0_417,RI9929020_397,RI992a790_377,RI992b0f0_357,RI992cc20_337,RI992d580_317,RI992f470_297,RI9931720_277,
        RI9933d90_257,RI9922888_576,RI99234b8_556,RI9923e18_536,RI9924778_516,RI9925768_496,RI99260c8_476,RI9926a28_456,RI9927dd8_436,RI9928738_416,
        RI9929098_396,RI992a808_376,RI992b168_356,RI992cc98_336,RI992d5f8_316,RI992f4e8_296,RI9931798_276,RI9935ed8_256,RI9922720_579,RI9923350_559,
        RI9923cb0_539,RI9924610_519,RI9925600_499,RI9925f60_479,RI99268c0_459,RI9927c70_439,RI99285d0_419,RI9928f30_399,RI992a6a0_379,RI992b000_359,
        RI992cb30_339,RI992d490_319,RI992f380_299,RI9931630_279,RI9933ca0_259,RI9922798_578,RI99233c8_558,RI9923d28_538,RI9924688_518,RI9925678_498,
        RI9925fd8_478,RI9926938_458,RI9927ce8_438,RI9928648_418,RI9928fa8_398,RI992a718_378,RI992b078_358,RI992cba8_338,RI992d508_318,RI992f3f8_298,
        RI99316a8_278,RI9933d18_258,RI9922630_581,RI9923260_561,RI9923bc0_541,RI9924520_521,RI9925510_501,RI9925e70_481,RI99267d0_461,RI9927b80_441,
        RI99284e0_421,RI9928e40_401,RI992a5b0_381,RI992af10_361,RI992ca40_341,RI992d3a0_321,RI992f290_301,RI9931540_281,RI9933bb0_261,RI99226a8_580,
        RI99232d8_560,RI9923c38_540,RI9924598_520,RI9925588_500,RI9925ee8_480,RI9926848_460,RI9927bf8_440,RI9928558_420,RI9928eb8_400,RI992a628_380,
        RI992af88_360,RI992cab8_340,RI992d418_320,RI992f308_300,RI99315b8_280,RI9933c28_260,RI9922540_583,RI9923170_563,RI9923ad0_543,RI9924430_523,
        RI9924d90_503,RI9925d80_483,RI99266e0_463,RI9927040_443,RI99283f0_423,RI9928d50_403,RI992a4c0_383,RI992ae20_363,RI992c950_343,RI992d2b0_323,
        RI992f1a0_303,RI9931450_283,RI9933ac0_263,RI99225b8_582,RI99231e8_562,RI9923b48_542,RI99244a8_522,RI9924e08_502,RI9925df8_482,RI9926758_462,
        RI9927b08_442,RI9928468_422,RI9928dc8_402,RI992a538_382,RI992ae98_362,RI992c9c8_342,RI992d328_322,RI992f218_302,RI99314c8_282,RI9933b38_262,
        RI9922450_585,RI9923080_565,RI99239e0_545,RI9924340_525,RI9924ca0_505,RI9925c90_485,RI99265f0_465,RI9926f50_445,RI9928300_425,RI9928c60_405,
        RI992a3d0_385,RI992ad30_365,RI992c860_345,RI992d1c0_325,RI992f0b0_305,RI9931360_285,RI99339d0_265,RI99224c8_584,RI99230f8_564,RI9923a58_544,
        RI99243b8_524,RI9924d18_504,RI9925d08_484,RI9926668_464,RI9926fc8_444,RI9928378_424,RI9928cd8_404,RI992a448_384,RI992ada8_364,RI992c8d8_344,
        RI992d238_324,RI992f128_304,RI99313d8_284,RI9933a48_264,RI99223d8_586,RI9923008_566,RI9923968_546,RI99242c8_526,RI9924c28_506,RI9925c18_486,
        RI9926578_466,RI9926ed8_446,RI9928288_426,RI9928be8_406,RI992a358_386,RI992acb8_366,RI992c7e8_346,RI992d148_326,RI992f038_306,RI99312e8_286,
        RI9933958_266,RI9922360_587,RI9922f90_567,RI99238f0_547,RI9924250_527,RI9924bb0_507,RI9925ba0_487,RI9926500_467,RI9926e60_447,RI9928210_427,
        RI9928b70_407,RI992a2e0_387,RI992ac40_367,RI992c770_347,RI992d0d0_327,RI992efc0_307,RI992f920_287,RI99338e0_267,RI99216b8_614,RI995f080_2,
        RI995f008_3,RI995ef90_4,RI995ef18_5,RI995eea0_6,RI995ee28_7,RI995edb0_8,RI995ed38_9,RI995ecc0_10,RI995ec48_11,RI995ebd0_12,
        RI9921d48_600,RI9921dc0_599,RI9921e38_598,RI9921eb0_597,RI9921f28_596,RI9921fa0_595,RI9922018_594,RI9922090_593,RI9922108_592,RI9922180_591,
        RI99221f8_590,RI9922270_589,RI99222e8_588,RI994e4d8_13,RI995f0f8_1,R_289_8400778,R_28a_8401e70,R_28b_8401f18,R_28c_8401fc0,R_28d_8402068,
        R_28e_8402110,R_28f_84021b8,R_290_8402260,R_291_8402308,R_292_84023b0,R_293_8402458,R_294_8402500,R_295_84025a8,R_296_8402650,R_297_84026f8,
        R_298_84027a0,R_299_8402848,R_29a_84028f0,R_29b_8402998,R_29c_8402a40,R_29d_8402ae8,R_29e_8402b90,R_29f_8402c38,R_2a0_8402ce0,R_2a1_8402d88,
        R_2a2_8402e30,R_2a3_8402ed8,R_267_8403418,R_268_8400820,R_269_84008c8,R_26a_8400970,R_26b_8400a18,R_26c_8400ac0,R_26d_8400b68,R_26e_8400c10,
        R_26f_8400cb8,R_270_8400d60,R_271_8400e08,R_272_8400eb0,R_273_8400f58,R_274_8401000,R_275_84010a8,R_276_8401150,R_277_84011f8,R_278_84012a0,
        R_279_8401348,R_27a_84013f0,R_27b_8401498,R_27c_8401540,R_27d_84015e8,R_27e_8401690,R_27f_8401738,R_280_84017e0,R_281_8401888);
input RI994e3e8_15,RI994e370_16,RI994e2f8_17,RI994e280_18,RI994e208_19,RI994e190_20,RI994e118_21,RI994e0a0_22,RI994e028_23,
        RI994dfb0_24,RI994df38_25,RI995e450_236,RI9921730_613,RI99217a8_612,RI9921820_611,RI9921898_610,RI9921910_609,RI9921988_608,RI9921a00_607,
        RI9921a78_606,RI9921af0_605,RI9921b68_604,RI9921be0_603,RI9921c58_602,RI9921cd0_601,RI9967078_223,RI9967690_210,RI890fba0_197,RI8918b88_184,
        RI89253b0_171,RI8930dc8_158,RI8939db0_145,RI89465d8_132,RI89ec640_119,RI9776f80_106,RI9808480_93,RI9808a98_80,RI9819730_67,RI98abc38_54,
        RI98bc8d0_41,RI994ddd0_28,RI995e3d8_237,RI99669e8_224,RI9967618_211,RI890fb28_198,RI8918b10_185,RI8925338_172,RI8930d50_159,RI8939d38_146,
        RI8946560_133,RI89ec5c8_120,RI9776f08_107,RI9808408_94,RI9808a20_81,RI98196b8_68,RI98abbc0_55,RI98bc858_42,RI994dd58_29,RI9959fe0_238,
        RI995e978_225,RI99675a0_212,RI890fab0_199,RI8918a98_186,RI89252c0_173,RI8930cd8_160,RI8939cc0_147,RI89464e8_134,RI89ec550_121,RI9776e90_108,
        RI9808390_95,RI98089a8_82,RI9819640_69,RI98abb48_56,RI98bc7e0_43,RI994dce0_30,RI9959f68_239,RI995e900_226,RI9967528_213,RI890fa38_200,
        RI8918a20_187,RI8925248_174,RI8930c60_161,RI8939c48_148,RI8946470_135,RI89ec4d8_122,RI9776e18_109,RI9808318_96,RI9808930_83,RI98195c8_70,
        RI98abad0_57,RI98bc768_44,RI994dc68_31,RI9959860_240,RI995e888_227,RI99674b0_214,RI890f9c0_201,RI89189a8_188,RI89251d0_175,RI8930be8_162,
        RI8939bd0_149,RI89463f8_136,RI89ec460_123,RI9776da0_110,RI98082a0_97,RI98088b8_84,RI9819550_71,RI98aba58_58,RI98bc6f0_45,RI994dbf0_32,
        RI994d998_241,RI995e810_228,RI9967438_215,RI890f948_202,RI8918930_189,RI8925158_176,RI8930b70_163,RI8939b58_150,RI8946380_137,RI89ec3e8_124,
        RI9776d28_111,RI9808228_98,RI9808840_85,RI98194d8_72,RI98ab9e0_59,RI98abff8_46,RI98bcc90_33,RI994d920_242,RI995e798_229,RI99673c0_216,
        RI890f8d0_203,RI89188b8_190,RI89250e0_177,RI8930af8_164,RI8939ae0_151,RI8946308_138,RI89ec370_125,RI89ec988_112,RI97772c8_99,RI98087c8_86,
        RI9819460_73,RI98ab968_60,RI98abf80_47,RI98bcc18_34,RI994d8a8_243,RI995e720_230,RI9967348_217,RI890f858_204,RI8918840_191,RI8925068_178,
        RI8930a80_165,RI8939a68_152,RI8946290_139,RI89ec2f8_126,RI89ec910_113,RI9777250_100,RI9808750_87,RI98193e8_74,RI98ab8f0_61,RI98abf08_48,
        RI98bcba0_35,RI994d830_244,RI995e6a8_231,RI99672d0_218,RI890f7e0_205,RI89187c8_192,RI8924ff0_179,RI8930a08_166,RI89399f0_153,RI8946218_140,
        RI89ec280_127,RI89ec898_114,RI97771d8_101,RI98086d8_88,RI9819370_75,RI98ab878_62,RI98abe90_49,RI98bcb28_36,RI994d7b8_245,RI995e630_232,
        RI9967258_219,RI890f768_206,RI8918750_193,RI8924f78_180,RI8930990_167,RI8939978_154,RI89461a0_141,RI89ec208_128,RI89ec820_115,RI9777160_102,
        RI9808660_89,RI98192f8_76,RI98ab800_63,RI98abe18_50,RI98bcab0_37,RI994d740_246,RI995e5b8_233,RI99671e0_220,RI890f6f0_207,RI89186d8_194,
        RI8924f00_181,RI8930918_168,RI8939900_155,RI8946128_142,RI89ec190_129,RI89ec7a8_116,RI97770e8_103,RI98085e8_90,RI9819280_77,RI98ab788_64,
        RI98abda0_51,RI98bca38_38,RI994dec0_26,RI994d6c8_247,RI995e540_234,RI9967168_221,RI890f678_208,RI8918660_195,RI8924e88_182,RI89308a0_169,
        RI8939888_156,RI89460b0_143,RI89ec118_130,RI89ec730_117,RI9777070_104,RI9808570_91,RI9819208_78,RI98ab710_65,RI98abd28_52,RI98bc9c0_39,
        RI9922bd0_569,RI9923800_549,RI9924160_529,RI9924ac0_509,RI9925ab0_489,RI9926410_469,RI9926d70_449,RI9928120_429,RI9928a80_409,RI992a1f0_389,
        RI992ab50_369,RI992b4b0_349,RI992cfe0_329,RI992eed0_309,RI992f830_289,RI9931ae0_269,RI994d5d8_249,RI994e460_14,RI995e4c8_235,RI99670f0_222,
        RI890f600_209,RI89185e8_196,RI8924e10_183,RI8930828_170,RI8939810_157,RI8946038_144,RI89ec0a0_131,RI89ec6b8_118,RI9776ff8_105,RI98084f8_92,
        RI9808b10_79,RI98197a8_66,RI98abcb0_53,RI98bc948_40,RI994de48_27,RI9922f18_568,RI9923878_548,RI99241d8_528,RI9924b38_508,RI9925b28_488,
        RI9926488_468,RI9926de8_448,RI9928198_428,RI9928af8_408,RI992a268_388,RI992abc8_368,RI992c6f8_348,RI992d058_328,RI992ef48_308,RI992f8a8_288,
        RI9931b58_268,RI994d650_248,RI9922b58_570,RI9923788_550,RI99240e8_530,RI9924a48_510,RI9925a38_490,RI9926398_470,RI9926cf8_450,RI99280a8_430,
        RI9928a08_410,RI992a178_390,RI992aad8_370,RI992b438_350,RI992cf68_330,RI992ee58_310,RI992f7b8_290,RI9931a68_270,RI994d560_250,RI9922a68_572,
        RI9923698_552,RI9923ff8_532,RI9924958_512,RI9925948_492,RI99262a8_472,RI9926c08_452,RI9927fb8_432,RI9928918_412,RI9929278_392,RI992a9e8_372,
        RI992b348_352,RI992ce78_332,RI992ed68_312,RI992f6c8_292,RI9931978_272,RI994d470_252,RI9922ae0_571,RI9923710_551,RI9924070_531,RI99249d0_511,
        RI99259c0_491,RI9926320_471,RI9926c80_451,RI9928030_431,RI9928990_411,RI992a100_391,RI992aa60_371,RI992b3c0_351,RI992cef0_331,RI992ede0_311,
        RI992f740_291,RI99319f0_271,RI994d4e8_251,RI99229f0_573,RI9923620_553,RI9923f80_533,RI99248e0_513,RI99258d0_493,RI9926230_473,RI9926b90_453,
        RI9927f40_433,RI99288a0_413,RI9929200_393,RI992a970_373,RI992b2d0_353,RI992ce00_333,RI992ecf0_313,RI992f650_293,RI9931900_273,RI994d3f8_253,
        RI9922900_575,RI9923530_555,RI9923e90_535,RI99247f0_515,RI99257e0_495,RI9926140_475,RI9926aa0_455,RI9927e50_435,RI99287b0_415,RI9929110_395,
        RI992a880_375,RI992b1e0_355,RI992cd10_335,RI992d670_315,RI992f560_295,RI9931810_275,RI9935f50_255,RI9922978_574,RI99235a8_554,RI9923f08_534,
        RI9924868_514,RI9925858_494,RI99261b8_474,RI9926b18_454,RI9927ec8_434,RI9928828_414,RI9929188_394,RI992a8f8_374,RI992b258_354,RI992cd88_334,
        RI992d6e8_314,RI992f5d8_294,RI9931888_274,RI9935fc8_254,RI9922810_577,RI9923440_557,RI9923da0_537,RI9924700_517,RI99256f0_497,RI9926050_477,
        RI99269b0_457,RI9927d60_437,RI99286c0_417,RI9929020_397,RI992a790_377,RI992b0f0_357,RI992cc20_337,RI992d580_317,RI992f470_297,RI9931720_277,
        RI9933d90_257,RI9922888_576,RI99234b8_556,RI9923e18_536,RI9924778_516,RI9925768_496,RI99260c8_476,RI9926a28_456,RI9927dd8_436,RI9928738_416,
        RI9929098_396,RI992a808_376,RI992b168_356,RI992cc98_336,RI992d5f8_316,RI992f4e8_296,RI9931798_276,RI9935ed8_256,RI9922720_579,RI9923350_559,
        RI9923cb0_539,RI9924610_519,RI9925600_499,RI9925f60_479,RI99268c0_459,RI9927c70_439,RI99285d0_419,RI9928f30_399,RI992a6a0_379,RI992b000_359,
        RI992cb30_339,RI992d490_319,RI992f380_299,RI9931630_279,RI9933ca0_259,RI9922798_578,RI99233c8_558,RI9923d28_538,RI9924688_518,RI9925678_498,
        RI9925fd8_478,RI9926938_458,RI9927ce8_438,RI9928648_418,RI9928fa8_398,RI992a718_378,RI992b078_358,RI992cba8_338,RI992d508_318,RI992f3f8_298,
        RI99316a8_278,RI9933d18_258,RI9922630_581,RI9923260_561,RI9923bc0_541,RI9924520_521,RI9925510_501,RI9925e70_481,RI99267d0_461,RI9927b80_441,
        RI99284e0_421,RI9928e40_401,RI992a5b0_381,RI992af10_361,RI992ca40_341,RI992d3a0_321,RI992f290_301,RI9931540_281,RI9933bb0_261,RI99226a8_580,
        RI99232d8_560,RI9923c38_540,RI9924598_520,RI9925588_500,RI9925ee8_480,RI9926848_460,RI9927bf8_440,RI9928558_420,RI9928eb8_400,RI992a628_380,
        RI992af88_360,RI992cab8_340,RI992d418_320,RI992f308_300,RI99315b8_280,RI9933c28_260,RI9922540_583,RI9923170_563,RI9923ad0_543,RI9924430_523,
        RI9924d90_503,RI9925d80_483,RI99266e0_463,RI9927040_443,RI99283f0_423,RI9928d50_403,RI992a4c0_383,RI992ae20_363,RI992c950_343,RI992d2b0_323,
        RI992f1a0_303,RI9931450_283,RI9933ac0_263,RI99225b8_582,RI99231e8_562,RI9923b48_542,RI99244a8_522,RI9924e08_502,RI9925df8_482,RI9926758_462,
        RI9927b08_442,RI9928468_422,RI9928dc8_402,RI992a538_382,RI992ae98_362,RI992c9c8_342,RI992d328_322,RI992f218_302,RI99314c8_282,RI9933b38_262,
        RI9922450_585,RI9923080_565,RI99239e0_545,RI9924340_525,RI9924ca0_505,RI9925c90_485,RI99265f0_465,RI9926f50_445,RI9928300_425,RI9928c60_405,
        RI992a3d0_385,RI992ad30_365,RI992c860_345,RI992d1c0_325,RI992f0b0_305,RI9931360_285,RI99339d0_265,RI99224c8_584,RI99230f8_564,RI9923a58_544,
        RI99243b8_524,RI9924d18_504,RI9925d08_484,RI9926668_464,RI9926fc8_444,RI9928378_424,RI9928cd8_404,RI992a448_384,RI992ada8_364,RI992c8d8_344,
        RI992d238_324,RI992f128_304,RI99313d8_284,RI9933a48_264,RI99223d8_586,RI9923008_566,RI9923968_546,RI99242c8_526,RI9924c28_506,RI9925c18_486,
        RI9926578_466,RI9926ed8_446,RI9928288_426,RI9928be8_406,RI992a358_386,RI992acb8_366,RI992c7e8_346,RI992d148_326,RI992f038_306,RI99312e8_286,
        RI9933958_266,RI9922360_587,RI9922f90_567,RI99238f0_547,RI9924250_527,RI9924bb0_507,RI9925ba0_487,RI9926500_467,RI9926e60_447,RI9928210_427,
        RI9928b70_407,RI992a2e0_387,RI992ac40_367,RI992c770_347,RI992d0d0_327,RI992efc0_307,RI992f920_287,RI99338e0_267,RI99216b8_614,RI995f080_2,
        RI995f008_3,RI995ef90_4,RI995ef18_5,RI995eea0_6,RI995ee28_7,RI995edb0_8,RI995ed38_9,RI995ecc0_10,RI995ec48_11,RI995ebd0_12,
        RI9921d48_600,RI9921dc0_599,RI9921e38_598,RI9921eb0_597,RI9921f28_596,RI9921fa0_595,RI9922018_594,RI9922090_593,RI9922108_592,RI9922180_591,
        RI99221f8_590,RI9922270_589,RI99222e8_588,RI994e4d8_13,RI995f0f8_1;
output R_289_8400778,R_28a_8401e70,R_28b_8401f18,R_28c_8401fc0,R_28d_8402068,R_28e_8402110,R_28f_84021b8,R_290_8402260,R_291_8402308,
        R_292_84023b0,R_293_8402458,R_294_8402500,R_295_84025a8,R_296_8402650,R_297_84026f8,R_298_84027a0,R_299_8402848,R_29a_84028f0,R_29b_8402998,
        R_29c_8402a40,R_29d_8402ae8,R_29e_8402b90,R_29f_8402c38,R_2a0_8402ce0,R_2a1_8402d88,R_2a2_8402e30,R_2a3_8402ed8,R_267_8403418,R_268_8400820,
        R_269_84008c8,R_26a_8400970,R_26b_8400a18,R_26c_8400ac0,R_26d_8400b68,R_26e_8400c10,R_26f_8400cb8,R_270_8400d60,R_271_8400e08,R_272_8400eb0,
        R_273_8400f58,R_274_8401000,R_275_84010a8,R_276_8401150,R_277_84011f8,R_278_84012a0,R_279_8401348,R_27a_84013f0,R_27b_8401498,R_27c_8401540,
        R_27d_84015e8,R_27e_8401690,R_27f_8401738,R_280_84017e0,R_281_8401888;

wire \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 ,
         \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 ,
         \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 ,
         \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 ,
         \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 ,
         \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 ,
         \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 ,
         \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 ,
         \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 ,
         \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 ,
         \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 ,
         \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 ,
         \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 ,
         \1368 , \1369 , \1370 , \1371 , \1372 , \1373_N$1 , \1374_N$2 , \1375_N$3 , \1376_N$4 , \1377_N$5 ,
         \1378_N$6 , \1379_N$7 , \1380_N$8 , \1381_N$9 , \1382_N$10 , \1383_N$11 , \1384_N$12 , \1385_N$13 , \1386_N$14 , \1387_N$15 ,
         \1388_N$16 , \1389_N$17 , \1390_N$18 , \1391_N$20 , \1392_N$21 , \1393_N$22 , \1394_N$23 , \1395_N$24 , \1396_N$25 , \1397_N$26 ,
         \1398_N$27 , \1399_N$28 , \1400_N$29 , \1401_N$30 , \1402_N$31 , \1403_N$32 , \1404_N$33 , \1405_N$34 , \1406_N$35 , \1407_N$36 ,
         \1408_N$37 , \1409_N$38 , \1410_N$39 , \1411_N$40 , \1412_N$41 , \1413_N$42 , \1414_N$43 , \1415_N$45 , \1416_N$46 , \1417_N$47 ,
         \1418_N$48 , \1419_N$49 , \1420_N$50 , \1421_N$51 , \1422_N$52 , \1423_N$53 , \1424_N$54 , \1425_N$55 , \1426_N$56 , \1427_N$57 ,
         \1428_N$58 , \1429_N$59 , \1430_N$60 , \1431_N$61 , \1432_N$62 , \1433_N$63 , \1434_N$64 , \1435_N$65 , \1436_N$66 , \1437_N$67 ,
         \1438_N$68 , \1439_N$69 , \1440_N$70 , \1441_N$71 , \1442_N$72 , \1443_N$73 , \1444_N$74 , \1445_N$75 , \1446_N$76 , \1447_N$77 ,
         \1448_N$78 , \1449_N$79 , \1450_N$80 , \1451_N$81 , \1452_N$82 , \1453_N$83 , \1454_N$85 , \1455_N$86 , \1456_N$87 , \1457_N$88 ,
         \1458_N$90 , \1459_N$91 , \1460_N$92 , \1461_N$93 , \1462_N$94 , \1463_N$95 , \1464_N$96 , \1465_N$98 , \1466_N$99 , \1467_N$100 ,
         \1468_N$101 , \1469_N$102 , \1470_N$103 , \1471_N$104 , \1472_N$105 , \1473_N$106 , \1474_N$107 , \1475_N$108 , \1476_N$109 , \1477_N$110 ,
         \1478_N$111 , \1479_N$112 , \1480_N$113 , \1481_N$114 , \1482_N$115 , \1483_N$116 , \1484_N$117 , \1485_N$118 , \1486_N$119 , \1487_N$120 ,
         \1488_N$121 , \1489_N$122 , \1490_N$123 , \1491_N$124 , \1492_N$125 , \1493_N$126 , \1494_N$127 , \1495_N$128 , \1496_N$129 , \1497_N$130 ,
         \1498_N$131 , \1499_N$132 , \1500_N$133 , \1501_N$134 , \1502_N$135 , \1503_N$137 , \1504_N$138 , \1505_N$139 , \1506_N$140 , \1507_N$141 ,
         \1508_N$142 , \1509_N$143 , \1510_N$144 , \1511_N$145 , \1512_N$146 , \1513_N$147 , \1514_N$148 , \1515_N$149 , \1516_N$150 , \1517_N$151 ,
         \1518_N$152 , \1519_N$153 , \1520_N$154 , \1521_N$155 , \1522_N$156 , \1523_N$157 , \1524_N$158 , \1525_N$159 , \1526_N$160 , \1527_N$161 ,
         \1528_N$162 , \1529_N$163 , \1530_N$164 , \1531_N$165 , \1532_N$166 , \1533_N$167 , \1534_N$168 , \1535_N$169 , \1536_N$171 , \1537_N$172 ,
         \1538_N$173 , \1539_N$174 , \1540_N$175 , \1541_N$176 , \1542_N$177 , \1543_N$178 , \1544_N$179 , \1545_N$180 , \1546_N$181 , \1547_N$182 ,
         \1548_N$183 , \1549_N$184 , \1550_N$185 , \1551_N$186 , \1552_N$187 , \1553_N$188 , \1554_N$189 , \1555_N$190 , \1556_N$191 , \1557_N$192 ,
         \1558_N$193 , \1559_N$194 , \1560_N$195 , \1561_N$196 , \1562_N$197 , \1563_N$198 , \1564_N$199 , \1565_N$200 , \1566_N$201 , \1567_N$203 ,
         \1568_N$204 , \1569_N$205 , \1570_N$206 , \1571_N$207 , \1572_N$208 , \1573_N$209 , \1574_N$210 , \1575_N$211 , \1576_N$212 , \1577_N$213 ,
         \1578_N$214 , \1579_N$215 , \1580_N$216 , \1581_N$217 , \1582_N$218 , \1583_N$219 , \1584_N$220 , \1585_N$221 , \1586_N$222 , \1587_N$223 ,
         \1588_N$224 , \1589_N$225 , \1590_N$226 , \1591_N$228 , \1592_N$229 , \1593_N$230 , \1594_N$231 , \1595_N$232 , \1596_N$233 , \1597_N$234 ,
         \1598_N$235 , \1599_N$236 , \1600_N$237 , \1601_N$238 , \1602_N$239 , \1603_N$240 , \1604_N$241 , \1605_N$242 , \1606_N$243 , \1607_N$244 ,
         \1608_N$245 , \1609_N$246 , \1610_N$247 , \1611_N$248 , \1612_N$249 , \1613_N$250 , \1614_N$251 , \1615_N$252 , \1616_N$253 , \1617_N$254 ,
         \1618_N$255 , \1619_N$256 , \1620_N$257 , \1621_N$258 , \1622_N$259 , \1623_N$260 , \1624_N$261 , \1625_N$262 , \1626_N$263 , \1627_N$264 ,
         \1628_N$265 , \1629_N$266 , \1630_N$268 , \1631_N$269 , \1632_N$270 , \1633_N$271 , \1634_N$273 , \1635_N$274 , \1636_N$275 , \1637_N$276 ,
         \1638_N$277 , \1639_N$278 , \1640_N$279 , \1641_N$281 , \1642_N$282 , \1643_N$283 , \1644_N$284 , \1645_N$285 , \1646_N$286 , \1647_N$287 ,
         \1648_N$288 , \1649_N$289 , \1650_N$290 , \1651_N$291 , \1652_N$292 , \1653_N$293 , \1654_N$294 , \1655_N$295 , \1656_N$296 , \1657_N$297 ,
         \1658_N$298 , \1659_N$299 , \1660_N$300 , \1661_N$301 , \1662_N$302 , \1663_N$303 , \1664_N$304 , \1665_N$305 , \1666_N$306 , \1667_N$307 ,
         \1668_N$308 , \1669_N$309 , \1670_N$310 , \1671_N$311 , \1672_N$312 , \1673_N$313 , \1674_N$314 , \1675_N$315 , \1676_N$316 , \1677_N$317 ,
         \1678_N$318 , \1679_N$320 , \1680_N$321 , \1681_N$322 , \1682_N$323 , \1683_N$324 , \1684_N$325 , \1685_N$326 , \1686_N$327 , \1687_N$328 ,
         \1688_N$329 , \1689_N$330 , \1690_N$331 , \1691_N$332 , \1692_N$333 , \1693_N$334 , \1694_N$335 , \1695_N$336 , \1696_N$337 , \1697_N$338 ,
         \1698_N$339 , \1699_N$340 , \1700_N$341 , \1701_N$342 , \1702_N$343 , \1703_N$344 , \1704_N$345 , \1705_N$346 , \1706_N$347 , \1707_N$348 ,
         \1708_N$349 , \1709_N$350 , \1710_N$351 , \1711_N$352 , \1712_N$354 , \1713_N$355 , \1714_N$356 , \1715_N$357 , \1716_N$358 , \1717_N$359 ,
         \1718_N$360 , \1719_N$361 , \1720_N$362 , \1721_N$363 , \1722_N$364 , \1723_N$365 , \1724_N$366 , \1725_N$367 , \1726_N$368 , \1727_N$369 ,
         \1728_N$370 , \1729_N$371 , \1730_N$372 , \1731_N$373 , \1732_N$374 , \1733_N$375 , \1734_N$376 , \1735_N$377 , \1736_N$378 , \1737_N$379 ,
         \1738_N$380 , \1739_N$381 , \1740_N$382 , \1741_N$383 , \1742_N$384 , \1743_N$386 , \1744_N$387 , \1745_N$388 , \1746_N$389 , \1747_N$390 ,
         \1748_N$391 , \1749_N$392 , \1750_N$393 , \1751_N$394 , \1752_N$395 , \1753_N$396 , \1754_N$397 , \1755_N$398 , \1756_N$399 , \1757_N$400 ,
         \1758_N$401 , \1759_N$402 , \1760_N$403 , \1761_N$404 , \1762_N$405 , \1763_N$406 , \1764_N$407 , \1765_N$408 , \1766_N$409 , \1767_N$411 ,
         \1768_N$412 , \1769_N$413 , \1770_N$414 , \1771_N$415 , \1772_N$416 , \1773_N$417 , \1774_N$418 , \1775_N$419 , \1776_N$420 , \1777_N$421 ,
         \1778_N$422 , \1779_N$423 , \1780_N$424 , \1781_N$425 , \1782_N$426 , \1783_N$427 , \1784_N$428 , \1785_N$429 , \1786_N$430 , \1787_N$431 ,
         \1788_N$432 , \1789_N$433 , \1790_N$434 , \1791_N$435 , \1792_N$436 , \1793_N$437 , \1794_N$438 , \1795_N$439 , \1796_N$440 , \1797_N$441 ,
         \1798_N$442 , \1799_N$443 , \1800_N$444 , \1801_N$445 , \1802_N$446 , \1803_N$447 , \1804_N$448 , \1805_N$449 , \1806_N$451 , \1807_N$452 ,
         \1808_N$453 , \1809_N$454 , \1810_N$456 , \1811_N$457 , \1812_N$458 , \1813_N$459 , \1814_N$460 , \1815_N$461 , \1816_N$462 , \1817_N$464 ,
         \1818_N$465 , \1819_N$466 , \1820_N$467 , \1821_N$468 , \1822_N$469 , \1823_N$470 , \1824_N$471 , \1825_N$472 , \1826_N$473 , \1827_N$474 ,
         \1828_N$475 , \1829_N$476 , \1830_N$477 , \1831_N$478 , \1832_N$479 , \1833_N$480 , \1834_N$481 , \1835_N$482 , \1836_N$483 , \1837_N$484 ,
         \1838_N$485 , \1839_N$486 , \1840_N$487 , \1841_N$488 , \1842_N$489 , \1843_N$490 , \1844_N$491 , \1845_N$492 , \1846_N$493 , \1847_N$494 ,
         \1848_N$495 , \1849_N$496 , \1850_N$497 , \1851_N$498 , \1852_N$499 , \1853_N$500 , \1854_N$501 , \1855_N$503 , \1856_N$504 , \1857_N$505 ,
         \1858_N$506 , \1859_N$507 , \1860_N$508 , \1861_N$509 , \1862_N$510 , \1863_N$511 , \1864_N$512 , \1865_N$513 , \1866_N$514 , \1867_N$515 ,
         \1868_N$516 , \1869_N$517 , \1870_N$518 , \1871_N$519 , \1872_N$520 , \1873_N$521 , \1874_N$522 , \1875_N$523 , \1876_N$524 , \1877_N$525 ,
         \1878_N$526 , \1879_N$527 , \1880_N$528 , \1881_N$529 , \1882_N$530 , \1883_N$531 , \1884_N$532 , \1885_N$533 , \1886_N$534 , \1887_N$535 ,
         \1888_N$537 , \1889_N$538 , \1890_N$539 , \1891_N$540 , \1892_N$541 , \1893_N$542 , \1894_N$543 , \1895_N$544 , \1896_N$545 , \1897_N$546 ,
         \1898_N$547 , \1899_N$548 , \1900_N$549 , \1901_N$550 , \1902_N$551 , \1903_N$552 , \1904_N$553 , \1905_N$554 , \1906_N$555 , \1907_N$556 ,
         \1908_N$557 , \1909_N$558 , \1910_N$559 , \1911_N$560 , \1912_N$561 , \1913_N$562 , \1914_N$563 , \1915_N$564 , \1916_N$565 , \1917_N$566 ,
         \1918_N$567 , \1919_N$569 , \1920_N$570 , \1921_N$571 , \1922_N$572 , \1923_N$573 , \1924_N$574 , \1925_N$575 , \1926_N$576 , \1927_N$577 ,
         \1928_N$578 , \1929_N$579 , \1930_N$580 , \1931_N$581 , \1932_N$582 , \1933_N$583 , \1934_N$584 , \1935_N$585 , \1936_N$586 , \1937_N$587 ,
         \1938_N$588 , \1939_N$589 , \1940_N$590 , \1941_N$591 , \1942_N$592 , \1943_N$594 , \1944_N$595 , \1945_N$596 , \1946_N$597 , \1947_N$598 ,
         \1948_N$599 , \1949_N$600 , \1950_N$601 , \1951_N$602 , \1952_N$603 , \1953_N$604 , \1954_N$605 , \1955_N$606 , \1956_N$607 , \1957_N$608 ,
         \1958_N$609 , \1959_N$610 , \1960_N$611 , \1961_N$612 , \1962_N$613 , \1963_N$614 , \1964_N$615 , \1965_N$616 , \1966_N$617 , \1967_N$618 ,
         \1968_N$619 , \1969_N$620 , \1970_N$621 , \1971_N$622 , \1972_N$623 , \1973_N$624 , \1974_N$625 , \1975_N$626 , \1976_N$627 , \1977_N$628 ,
         \1978_N$629 , \1979_N$630 , \1980_N$631 , \1981_N$632 , \1982_N$634 , \1983_N$635 , \1984_N$636 , \1985_N$637 , \1986_N$639 , \1987_N$640 ,
         \1988_N$641 , \1989_N$642 , \1990_N$643 , \1991_N$644 , \1992_N$645 , \1993_N$647 , \1994_N$648 , \1995_N$649 , \1996_N$650 , \1997_N$651 ,
         \1998_N$652 , \1999_N$653 , \2000_N$654 , \2001_N$655 , \2002_N$656 , \2003_N$657 , \2004_N$658 , \2005_N$659 , \2006_N$660 , \2007_N$661 ,
         \2008_N$662 , \2009_N$663 , \2010_N$664 , \2011_N$665 , \2012_N$666 , \2013_N$667 , \2014_N$668 , \2015_N$669 , \2016_N$670 , \2017_N$671 ,
         \2018_N$672 , \2019_N$673 , \2020_N$674 , \2021_N$675 , \2022_N$676 , \2023_N$677 , \2024_N$678 , \2025_N$679 , \2026_N$680 , \2027_N$681 ,
         \2028_N$682 , \2029_N$683 , \2030_N$684 , \2031_N$686 , \2032_N$687 , \2033_N$688 , \2034_N$689 , \2035_N$690 , \2036_N$691 , \2037_N$692 ,
         \2038_N$693 , \2039_N$694 , \2040_N$695 , \2041_N$696 , \2042_N$697 , \2043_N$698 , \2044_N$699 , \2045_N$700 , \2046_N$701 , \2047_N$702 ,
         \2048_N$703 , \2049_N$704 , \2050_N$705 , \2051_N$706 , \2052_N$707 , \2053_N$708 , \2054_N$709 , \2055_N$710 , \2056_N$711 , \2057_N$712 ,
         \2058_N$713 , \2059_N$714 , \2060_N$715 , \2061_N$716 , \2062_N$717 , \2063_N$718 , \2064_N$720 , \2065_N$721 , \2066_N$722 , \2067_N$723 ,
         \2068_N$724 , \2069_N$725 , \2070_N$726 , \2071_N$727 , \2072_N$728 , \2073_N$729 , \2074_N$730 , \2075_N$731 , \2076_N$732 , \2077_ZERO ,
         \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 ,
         \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 ,
         \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106_N$19 , \2107_N$44 ,
         \2108_N$84 , \2109_N$89 , \2110_N$97 , \2111_N$136 , \2112_N$170 , \2113_N$202 , \2114_N$227 , \2115_N$267 , \2116_N$272 , \2117_N$280 ,
         \2118_N$319 , \2119_N$353 , \2120_N$385 , \2121_N$410 , \2122_N$450 , \2123_N$455 , \2124_N$463 , \2125_N$502 , \2126_N$536 , \2127_N$568 ,
         \2128_N$593 , \2129_N$633 , \2130_N$638 , \2131_N$646 , \2132_N$685 , \2133_N$719 , \2134_ONE , \2135 , \2136 , \2137 ,
         \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 ,
         \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 ,
         \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 ,
         \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 ,
         \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 ,
         \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 ,
         \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 ,
         \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215_nG2199 , \2216 , \2217 ,
         \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 ,
         \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 ,
         \2238 , \2239 , \2240_nG2175 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 ,
         \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 ,
         \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265_nG1fee , \2266 , \2267 ,
         \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 ,
         \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 ,
         \2288 , \2289 , \2290_nG1fca , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 ,
         \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 ,
         \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315_nG1e55 , \2316 , \2317 ,
         \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 ,
         \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 ,
         \2338 , \2339 , \2340_nG1e31 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 ,
         \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 ,
         \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365_nG1cf3 , \2366 , \2367 ,
         \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 ,
         \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 ,
         \2388 , \2389 , \2390_nG1ccf , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 ,
         \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 ,
         \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415_nG1bc2 , \2416 , \2417 ,
         \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 ,
         \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 ,
         \2438 , \2439 , \2440_nG1bdb , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 ,
         \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 ,
         \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465_nG1aa5 , \2466 , \2467 ,
         \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 ,
         \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 ,
         \2488 , \2489_nG1a89 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 ,
         \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 ,
         \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 ,
         \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524_nG21a2 , \2525 , \2526 , \2527 ,
         \2528_nG217e , \2529 , \2530 , \2531 , \2532_nG1ff7 , \2533 , \2534 , \2535 , \2536 , \2537 ,
         \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 ,
         \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 ,
         \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 ,
         \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 ,
         \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 ,
         \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 ,
         \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 ,
         \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 ,
         \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 ,
         \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 ,
         \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 ,
         \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 ,
         \2658_nG2899 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 ,
         \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 ,
         \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686_nG2361 , \2687 ,
         \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 ,
         \2698_nG2376 , \2699 , \2700 , \2701 , \2702_nG236a , \2703 , \2704 , \2705 , \2706 , \2707 ,
         \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 ,
         \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727_nG298d ,
         \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 ,
         \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 ,
         \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754_nG27d7 , \2755 , \2756 , \2757 ,
         \2758_nG2572 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 ,
         \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 ,
         \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 ,
         \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 ,
         \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 ,
         \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 ,
         \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825_nG1fd3 , \2826 , \2827 ,
         \2828 , \2829 , \2830_nG1e5e , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 ,
         \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 ,
         \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 ,
         \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865_nG263c , \2866 , \2867 ,
         \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 ,
         \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886_nG2716 , \2887 ,
         \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 ,
         \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 ,
         \2908 , \2909_nG2551 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 ,
         \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 ,
         \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 ,
         \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 ,
         \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 ,
         \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 ,
         \2968 , \2969 , \2970 , \2971 , \2972_nG1aac , \2973 , \2974 , \2975_nG1a8c , \2976 , \2977 ,
         \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 ,
         \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 ,
         \2998 , \2999 , \3000 , \3001 , \3002_nG239e , \3003 , \3004 , \3005 , \3006_nG1be7 , \3007 ,
         \3008 , \3009 , \3010_nG1beb , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 ,
         \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 ,
         \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035_nG2472 , \3036 , \3037 ,
         \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 ,
         \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 ,
         \3058 , \3059 , \3060 , \3061 , \3062_nG21d1 , \3063 , \3064 , \3065 , \3066_nG1cfc , \3067 ,
         \3068 , \3069 , \3070_nG1cd8 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 ,
         \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 ,
         \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095_nG22a8 , \3096 , \3097 ,
         \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 ,
         \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 ,
         \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124_nG2012 , \3125 , \3126 , \3127 ,
         \3128_nG1e3a , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 ,
         \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 ,
         \3148 , \3149 , \3150 , \3151 , \3152 , \3153_nG20db , \3154 , \3155 , \3156 , \3157 ,
         \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 ,
         \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 ,
         \3178 , \3179_nG1e79 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 ,
         \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 ,
         \3198 , \3199 , \3200_nG1f2c , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 ,
         \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 ,
         \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224_nG1d15 , \3225 , \3226 , \3227 ,
         \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 ,
         \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245_nG1dbc , \3246 , \3247 ,
         \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 ,
         \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 ,
         \3268 , \3269 , \3270 , \3271 , \3272_nG1ba5 , \3273 , \3274 , \3275 , \3276 , \3277 ,
         \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 ,
         \3288 , \3289 , \3290 , \3291 , \3292 , \3293_nG1c76 , \3294 , \3295 , \3296 , \3297 ,
         \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 ,
         \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316_nG1b63 , \3317 ,
         \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 ,
         \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 ,
         \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 ,
         \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 ,
         \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 ,
         \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 ,
         \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 ,
         \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 ,
         \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 ,
         \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 ,
         \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 ,
         \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 ,
         \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 ,
         \3448 , \3449_nG1a4f , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 ,
         \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 ,
         \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 ,
         \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 ,
         \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 ,
         \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 ,
         \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 ,
         \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 ,
         \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 ,
         \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 ,
         \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 ,
         \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 ,
         \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 ,
         \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 ,
         \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 ,
         \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 ,
         \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 ,
         \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 ,
         \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 ,
         \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 ,
         \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 ,
         \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 ,
         \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 ,
         \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 ,
         \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 ,
         \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 ,
         \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 ,
         \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 ,
         \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 ,
         \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 ,
         \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 ,
         \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 ,
         \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 ,
         \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 ,
         \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 ,
         \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 ,
         \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 ,
         \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 ,
         \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 ,
         \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 ,
         \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 ,
         \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 ,
         \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 ,
         \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 ,
         \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 ,
         \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 ,
         \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 ,
         \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 ,
         \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 ,
         \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 ,
         \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 ,
         \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 ,
         \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 ,
         \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 ,
         \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 ,
         \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 ,
         \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 ,
         \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 ,
         \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 ,
         \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 ,
         \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 ,
         \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 ,
         \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 ,
         \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 ,
         \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 ,
         \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 ,
         \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 ,
         \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 ,
         \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 ,
         \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 ,
         \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 ,
         \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 ,
         \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 ,
         \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 ,
         \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 ,
         \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 ,
         \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 ,
         \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 ,
         \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 ,
         \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 ,
         \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 ,
         \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 ,
         \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 ,
         \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 ,
         \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 ,
         \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 ,
         \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 ,
         \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 ,
         \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 ,
         \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 ,
         \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 ,
         \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 ,
         \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 ,
         \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 ,
         \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 ,
         \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 ,
         \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 ,
         \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 ,
         \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 ,
         \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 ,
         \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 ,
         \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 ,
         \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 ,
         \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 ,
         \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 ,
         \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 ,
         \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 ,
         \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 ,
         \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 ,
         \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 ,
         \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 ,
         \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 ,
         \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 ,
         \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 ,
         \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 ,
         \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 ,
         \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 ,
         \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 ,
         \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 ,
         \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 ,
         \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 ,
         \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 ,
         \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 ,
         \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 ,
         \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 ,
         \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 ,
         \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 ,
         \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 ,
         \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 ,
         \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 ,
         \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 ,
         \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 ,
         \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 ,
         \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 ,
         \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 ,
         \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 ,
         \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 ,
         \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 ,
         \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 ,
         \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 ,
         \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 ,
         \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 ,
         \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 ,
         \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 ,
         \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 ,
         \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 ,
         \4908 , \4909 , \4910 , \4911 , \4912_nG3284 , \4913 , \4914 , \4915 , \4916 , \4917 ,
         \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 ,
         \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 ,
         \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 ,
         \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 ,
         \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 ,
         \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 ,
         \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 ,
         \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 ,
         \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 ,
         \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 ,
         \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 ,
         \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 ,
         \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 ,
         \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 ,
         \5058 , \5059 , \5060 , \5061_nG2232 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 ,
         \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 ,
         \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086_nG220e , \5087 ,
         \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 ,
         \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 ,
         \5108 , \5109 , \5110 , \5111_nG207b , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 ,
         \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 ,
         \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136_nG2057 , \5137 ,
         \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 ,
         \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 ,
         \5158 , \5159 , \5160 , \5161_nG1ed8 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 ,
         \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 ,
         \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186_nG1eb4 , \5187 ,
         \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 ,
         \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 ,
         \5208 , \5209 , \5210 , \5211_nG1d69 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 ,
         \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 ,
         \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236_nG1d45 , \5237 ,
         \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 ,
         \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 ,
         \5258 , \5259 , \5260 , \5261_nG1c2a , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 ,
         \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 ,
         \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286_nG1c43 , \5287 ,
         \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 ,
         \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 ,
         \5308 , \5309 , \5310 , \5311_nG1b40 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 ,
         \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 ,
         \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335_nG1b24 , \5336 , \5337 ,
         \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 ,
         \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 ,
         \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 ,
         \5368 , \5369 , \5370_nG223b , \5371 , \5372 , \5373 , \5374_nG2217 , \5375 , \5376 , \5377 ,
         \5378_nG2084 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 ,
         \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 ,
         \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 ,
         \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 ,
         \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 ,
         \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 ,
         \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 ,
         \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 ,
         \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 ,
         \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 ,
         \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 ,
         \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 ,
         \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504_nG290c , \5505 , \5506 , \5507 ,
         \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 ,
         \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 ,
         \5528 , \5529 , \5530 , \5531 , \5532_nG23ed , \5533 , \5534 , \5535 , \5536 , \5537 ,
         \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544_nG2402 , \5545 , \5546 , \5547 ,
         \5548_nG23f6 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 ,
         \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 ,
         \5568 , \5569 , \5570 , \5571 , \5572 , \5573_nG2a01 , \5574 , \5575 , \5576 , \5577 ,
         \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 ,
         \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 ,
         \5598 , \5599 , \5600_nG2843 , \5601 , \5602 , \5603 , \5604_nG25dc , \5605 , \5606 , \5607 ,
         \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 ,
         \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 ,
         \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 ,
         \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 ,
         \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 ,
         \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 ,
         \5668 , \5669 , \5670 , \5671_nG2060 , \5672 , \5673 , \5674 , \5675 , \5676_nG1ee1 , \5677 ,
         \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 ,
         \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 ,
         \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 ,
         \5708 , \5709 , \5710 , \5711_nG26a4 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 ,
         \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 ,
         \5728 , \5729 , \5730 , \5731 , \5732_nG2782 , \5733 , \5734 , \5735 , \5736 , \5737 ,
         \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 ,
         \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755_nG25bb , \5756 , \5757 ,
         \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 ,
         \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 ,
         \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 ,
         \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 ,
         \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 ,
         \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 ,
         \5818_nG1b47 , \5819 , \5820 , \5821_nG1b27 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 ,
         \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 ,
         \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 ,
         \5848_nG242a , \5849 , \5850 , \5851 , \5852_nG1c4f , \5853 , \5854 , \5855 , \5856_nG1c53 , \5857 ,
         \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 ,
         \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 ,
         \5878 , \5879 , \5880 , \5881_nG24d7 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 ,
         \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 ,
         \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 ,
         \5908_nG226a , \5909 , \5910 , \5911 , \5912_nG1d72 , \5913 , \5914 , \5915 , \5916_nG1d4e , \5917 ,
         \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 ,
         \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 ,
         \5938 , \5939 , \5940 , \5941_nG2302 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 ,
         \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 ,
         \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 ,
         \5968 , \5969 , \5970_nG209f , \5971 , \5972 , \5973 , \5974_nG1ebd , \5975 , \5976 , \5977 ,
         \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 ,
         \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 ,
         \5998 , \5999_nG2129 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 ,
         \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 ,
         \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025_nG1efc , \6026 , \6027 ,
         \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 ,
         \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046_nG1f70 , \6047 ,
         \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 ,
         \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 ,
         \6068 , \6069 , \6070_nG1d8b , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 ,
         \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 ,
         \6088 , \6089 , \6090 , \6091_nG1df2 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 ,
         \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 ,
         \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 ,
         \6118_nG1c0d , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 ,
         \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 ,
         \6138 , \6139_nG1ca0 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 ,
         \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 ,
         \6158 , \6159 , \6160 , \6161 , \6162_nG1b85 , \6163 , \6164 , \6165 , \6166 , \6167 ,
         \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 ,
         \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 ,
         \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 ,
         \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 ,
         \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 ,
         \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 ,
         \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 ,
         \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 ,
         \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 ,
         \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 ,
         \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 ,
         \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 ,
         \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295_nG1aea , \6296 , \6297 ,
         \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 ,
         \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 ,
         \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 ,
         \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 ,
         \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 ,
         \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 ,
         \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 ,
         \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 ,
         \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 ,
         \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 ,
         \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 ,
         \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 ,
         \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 ,
         \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 ,
         \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 ,
         \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 ,
         \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 ,
         \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 ,
         \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 ,
         \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 ,
         \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 ,
         \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 ,
         \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 ,
         \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 ,
         \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 ,
         \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 ,
         \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 ,
         \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 ,
         \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 ,
         \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 ,
         \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 ,
         \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 ,
         \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 ,
         \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 ,
         \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 ,
         \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 ,
         \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 ,
         \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 ,
         \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 ,
         \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 ,
         \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 ,
         \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 ,
         \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 ,
         \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 ,
         \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 ,
         \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 ,
         \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 ,
         \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 ,
         \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 ,
         \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 ,
         \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 ,
         \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 ,
         \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 ,
         \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 ,
         \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 ,
         \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 ,
         \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 ,
         \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 ,
         \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 ,
         \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 ,
         \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 ,
         \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 ,
         \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 ,
         \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 ,
         \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 ,
         \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 ,
         \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 ,
         \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 ,
         \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 ,
         \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 ,
         \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 ,
         \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 ,
         \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 ,
         \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 ,
         \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 ,
         \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 ,
         \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 ,
         \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 ,
         \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 ,
         \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 ,
         \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 ,
         \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 ,
         \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 ,
         \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 ,
         \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 ,
         \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 ,
         \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 ,
         \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 ,
         \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 ,
         \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 ,
         \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 ,
         \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 ,
         \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 ,
         \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 ,
         \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 ,
         \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 ,
         \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 ,
         \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 ,
         \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 ,
         \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 ,
         \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 ,
         \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 ,
         \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 ,
         \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 ,
         \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 ,
         \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 ,
         \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 ,
         \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 ,
         \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 ,
         \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 ,
         \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 ,
         \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 ,
         \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 ,
         \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 ,
         \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 ,
         \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 ,
         \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 ,
         \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 ,
         \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 ,
         \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 ,
         \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 ,
         \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 ,
         \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 ,
         \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 ,
         \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 ,
         \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 ,
         \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 ,
         \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 ,
         \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 ,
         \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 ,
         \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
         \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 ,
         \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 ,
         \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 ,
         \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 ,
         \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 ,
         \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 ,
         \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 ,
         \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 ,
         \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 ,
         \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 ,
         \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 ,
         \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 ,
         \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 ,
         \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 ,
         \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 ,
         \7758_nG32b2 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 ,
         \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 ,
         \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 ,
         \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 ,
         \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 ,
         \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 ,
         \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 ,
         \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 ,
         \7838 , \7839 , \7840_nG1080 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 ,
         \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 ,
         \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 , \7865_nG1099 , \7866 , \7867 ,
         \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 ,
         \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 ,
         \7888 , \7889 , \7890_nG10b2 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 ,
         \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 ,
         \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915_nG10cb , \7916 , \7917 ,
         \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 ,
         \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 ,
         \7938 , \7939 , \7940_nG10e4 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 ,
         \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 ,
         \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965_nG10fd , \7966 , \7967 ,
         \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 ,
         \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 ,
         \7988 , \7989 , \7990_nG1116 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 ,
         \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 ,
         \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015_nG112f , \8016 , \8017 ,
         \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 ,
         \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 ,
         \8038 , \8039 , \8040_nG1148 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 ,
         \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 ,
         \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065_nG1161 , \8066 , \8067 ,
         \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 ,
         \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 ,
         \8088 , \8089 , \8090_nG117a , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 ,
         \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 ,
         \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 , \8115_nG1193 , \8116 , \8117 ,
         \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 ,
         \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 ,
         \8138 , \8139_nG11ad , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 ,
         \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 ,
         \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 ,
         \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 ,
         \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 ,
         \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 ,
         \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 ,
         \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 ,
         \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 ,
         \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 ,
         \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 ,
         \8248 , \8249_nG1220 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 ,
         \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 ,
         \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 ,
         \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 ,
         \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 ,
         \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304_nG1257 , \8305 , \8306 , \8307 ,
         \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 ,
         \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325_nG126c , \8326 , \8327 ,
         \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 ,
         \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346_nG1281 , \8347 ,
         \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 ,
         \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367_nG1296 ,
         \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 ,
         \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 ,
         \8388_nG12ab , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 ,
         \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 ,
         \8408 , \8409_nG12c0 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 ,
         \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 ,
         \8428 , \8429 , \8430_nG12d5 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 ,
         \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 ,
         \8448 , \8449 , \8450 , \8451_nG12ea , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 ,
         \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 ,
         \8468 , \8469 , \8470 , \8471 , \8472_nG12ff , \8473 , \8474 , \8475 , \8476 , \8477 ,
         \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 ,
         \8488 , \8489 , \8490 , \8491 , \8492 , \8493_nG1314 , \8494 , \8495 , \8496 , \8497 ,
         \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 ,
         \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514_nG1329 , \8515 , \8516 , \8517 ,
         \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 ,
         \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535_nG133e , \8536 , \8537 ,
         \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 ,
         \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556_nG1353 , \8557 ,
         \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 ,
         \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577_nG1368 ,
         \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 ,
         \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 ,
         \8598_nG137d , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 ,
         \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 ,
         \8618 , \8619_nG1392 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 ,
         \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 ,
         \8638 , \8639 , \8640_nG13a7 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 ,
         \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 ,
         \8658 , \8659 , \8660 , \8661_nG13bc , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 ,
         \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 ,
         \8678 , \8679 , \8680 , \8681 , \8682_nG13d1 , \8683 , \8684 , \8685 , \8686 , \8687 ,
         \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 ,
         \8698 , \8699 , \8700 , \8701 , \8702 , \8703_nG13e6 , \8704 , \8705 , \8706 , \8707 ,
         \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 ,
         \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724_nG13fb , \8725 , \8726 , \8727 ,
         \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 ,
         \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745_nG1410 , \8746 , \8747 ,
         \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 ,
         \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766_nG1425 , \8767 ,
         \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 ,
         \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787_nG143a ,
         \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 ,
         \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 ,
         \8808_nG144f , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 ,
         \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 ,
         \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 ,
         \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 ,
         \8848 , \8849_nG32b3 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 ,
         \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 ,
         \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 ,
         \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 ,
         \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 ,
         \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 ,
         \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 ,
         \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 ,
         \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 ,
         \8938 , \8939 , \8940 , \8941 , \8942_nG3221 , \8943 , \8944 , \8945 , \8946 , \8947 ,
         \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 ,
         \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 ,
         \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 ,
         \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 ,
         \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 ,
         \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 ,
         \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 ,
         \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 ,
         \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034_nG3255 , \9035_nG3256 , \9036 , \9037 ,
         \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 ,
         \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 ,
         \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 ,
         \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 ,
         \9078 , \9079 , \9080 , \9081_nG31b2 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 ,
         \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 ,
         \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 ,
         \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 ,
         \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126_nG31ec , \9127_nG31ed ,
         \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 ,
         \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 ,
         \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 ,
         \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 ,
         \9168 , \9169 , \9170 , \9171 , \9172_nG3135 , \9173 , \9174 , \9175 , \9176 , \9177 ,
         \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 ,
         \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 ,
         \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 ,
         \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216_nG3177 , \9217_nG3178 ,
         \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 ,
         \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 ,
         \9238 , \9239 , \9240_nG30ac , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 ,
         \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 ,
         \9258 , \9259 , \9260 , \9261 , \9262_nG30f2 , \9263_nG30f3 , \9264 , \9265 , \9266 , \9267 ,
         \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 ,
         \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286_nG301d , \9287 ,
         \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 ,
         \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 ,
         \9308_nG3065 , \9309_nG3066 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 ,
         \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 ,
         \9328 , \9329 , \9330 , \9331_nG2f88 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 ,
         \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 ,
         \9348 , \9349 , \9350 , \9351 , \9352_nG2fd4 , \9353_nG2fd5 , \9354 , \9355 , \9356 , \9357 ,
         \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 ,
         \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375_nG2eeb , \9376 , \9377 ,
         \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 ,
         \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396_nG2f3b , \9397_nG2f3c ,
         \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 ,
         \9408 , \9409_nG2e49 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 ,
         \9418 , \9419 , \9420_nG2e9a , \9421_nG2e9b , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 ,
         \9428 , \9429 , \9430 , \9431 , \9432 , \9433_nG2d9e , \9434 , \9435 , \9436 , \9437 ,
         \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444_nG2df7 , \9445_nG2df8 , \9446 , \9447 ,
         \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457_nG2ce8 ,
         \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 ,
         \9468_nG2d44 , \9469_nG2d45 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 ,
         \9478 , \9479 , \9480 , \9481_nG2c2b , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 ,
         \9488 , \9489 , \9490 , \9491 , \9492_nG2c8b , \9493_nG2c8c , \9494 , \9495 , \9496 , \9497 ,
         \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504_nG2b6b , \9505 , \9506 , \9507 ,
         \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514_nG2bca , \9515_nG2bcb , \9516 , \9517 ,
         \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526_nG2aac , \9527 ,
         \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536_nG2b0b , \9537_nG2b0c ,
         \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 ,
         \9548_nG29d8 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 ,
         \9558_nG2a4c , \9559_nG2a4d , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 ,
         \9568 , \9569 , \9570_nG28f0 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 ,
         \9578 , \9579 , \9580_nG2963 , \9581_nG2964 , \9582 , \9583 , \9584 , \9585 , \9586_nG2810 , \9587 ,
         \9588 , \9589 , \9590_nG287c , \9591_nG287d , \9592 , \9593 , \9594 , \9595 , \9596_nG2737 , \9597 ,
         \9598 , \9599 , \9600_nG27a3 , \9601_nG27a4 , \9602 , \9603 , \9604 , \9605 , \9606_nG2662 , \9607 ,
         \9608 , \9609 , \9610_nG26ca , \9611_nG26cb , \9612 , \9613 , \9614 , \9615 , \9616_nG258f , \9617 ,
         \9618 , \9619 , \9620_nG25f9 , \9621_nG25fa , \9622 , \9623 , \9624 , \9625 , \9626_nG24bf , \9627 ,
         \9628 , \9629 , \9630_nG2524 , \9631_nG2525 , \9632 , \9633 , \9634 , \9635 , \9636_nG23cd , \9637 ,
         \9638 , \9639 , \9640_nG2459 , \9641_nG245a , \9642 , \9643 , \9644 , \9645 , \9646_nG22e6 , \9647 ,
         \9648 , \9649 , \9650_nG2340 , \9651_nG2341 , \9652 , \9653 , \9654 , \9655 , \9656_nG21f2 , \9657 ,
         \9658 , \9659 , \9660_nG228b , \9661_nG228c , \9662 , \9663 , \9664 , \9665 , \9666_nG210a , \9667 ,
         \9668 , \9669 , \9670_nG2158 , \9671_nG2159 , \9672 , \9673 , \9674 , \9675 , \9676_nG202e , \9677 ,
         \9678 , \9679 , \9680_nG20bb , \9681_nG20bc , \9682 , \9683 , \9684 , \9685 , \9686_nG1f5c , \9687 ,
         \9688 , \9689 , \9690_nG1fa0 , \9691_nG1fa1 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 ,
         \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 ,
         \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 ,
         \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 ,
         \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 ,
         \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 ,
         \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 ,
         \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 ,
         \9768 , \9769 , \9770 , \9771 , \9772 , \9773_nG3a87 , \9774 , \9775 , \9776 , \9777 ,
         \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 ,
         \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 ,
         \9798_nG3a63 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 ,
         \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 ,
         \9818 , \9819 , \9820 , \9821 , \9822 , \9823_nG38dc , \9824 , \9825 , \9826 , \9827 ,
         \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 ,
         \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 ,
         \9848_nG38b8 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 ,
         \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 ,
         \9868 , \9869 , \9870 , \9871 , \9872 , \9873_nG3743 , \9874 , \9875 , \9876 , \9877 ,
         \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 ,
         \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 ,
         \9898_nG371f , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 ,
         \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 ,
         \9918 , \9919 , \9920 , \9921 , \9922 , \9923_nG35e1 , \9924 , \9925 , \9926 , \9927 ,
         \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 ,
         \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 ,
         \9948_nG35bd , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 ,
         \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 ,
         \9968 , \9969 , \9970 , \9971 , \9972 , \9973_nG34b0 , \9974 , \9975 , \9976 , \9977 ,
         \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 ,
         \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 ,
         \9998_nG34c9 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 ,
         \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 ,
         \10018 , \10019 , \10020 , \10021 , \10022 , \10023_nG3393 , \10024 , \10025 , \10026 , \10027 ,
         \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 ,
         \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047_nG3377 ,
         \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 ,
         \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 ,
         \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 ,
         \10078 , \10079 , \10080 , \10081 , \10082_nG3a90 , \10083 , \10084 , \10085 , \10086_nG3a6c , \10087 ,
         \10088 , \10089 , \10090_nG38e5 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 ,
         \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 ,
         \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 ,
         \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 ,
         \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 ,
         \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 ,
         \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 ,
         \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 ,
         \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 ,
         \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 ,
         \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 ,
         \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 ,
         \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216_nG4187 , \10217 ,
         \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 ,
         \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 ,
         \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244_nG3c4f , \10245 , \10246 , \10247 ,
         \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256_nG3c64 , \10257 ,
         \10258 , \10259 , \10260_nG3c58 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 ,
         \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 ,
         \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285_nG427b , \10286 , \10287 ,
         \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 ,
         \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 ,
         \10308 , \10309 , \10310 , \10311 , \10312_nG40c5 , \10313 , \10314 , \10315 , \10316_nG3e60 , \10317 ,
         \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 ,
         \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 ,
         \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 ,
         \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 ,
         \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 ,
         \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 ,
         \10378 , \10379 , \10380 , \10381 , \10382 , \10383_nG38c1 , \10384 , \10385 , \10386 , \10387 ,
         \10388_nG374c , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 ,
         \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 ,
         \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 ,
         \10418 , \10419 , \10420 , \10421 , \10422 , \10423_nG3f2a , \10424 , \10425 , \10426 , \10427 ,
         \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 ,
         \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444_nG4004 , \10445 , \10446 , \10447 ,
         \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 ,
         \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467_nG3e3f ,
         \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 ,
         \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 ,
         \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 ,
         \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 ,
         \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 ,
         \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 ,
         \10528 , \10529 , \10530_nG339a , \10531 , \10532 , \10533_nG337a , \10534 , \10535 , \10536 , \10537 ,
         \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 ,
         \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 ,
         \10558 , \10559 , \10560_nG3c8c , \10561 , \10562 , \10563 , \10564_nG34d5 , \10565 , \10566 , \10567 ,
         \10568_nG34d9 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 ,
         \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 ,
         \10588 , \10589 , \10590 , \10591 , \10592 , \10593_nG3d60 , \10594 , \10595 , \10596 , \10597 ,
         \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 ,
         \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 ,
         \10618 , \10619 , \10620_nG3abf , \10621 , \10622 , \10623 , \10624_nG35ea , \10625 , \10626 , \10627 ,
         \10628_nG35c6 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 ,
         \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 ,
         \10648 , \10649 , \10650 , \10651 , \10652 , \10653_nG3b96 , \10654 , \10655 , \10656 , \10657 ,
         \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 ,
         \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 ,
         \10678 , \10679 , \10680 , \10681 , \10682_nG3900 , \10683 , \10684 , \10685 , \10686_nG3728 , \10687 ,
         \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 ,
         \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 ,
         \10708 , \10709 , \10710 , \10711_nG39c9 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 ,
         \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 ,
         \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737_nG3767 ,
         \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 ,
         \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 ,
         \10758_nG381a , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 ,
         \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 ,
         \10778 , \10779 , \10780 , \10781 , \10782_nG3603 , \10783 , \10784 , \10785 , \10786 , \10787 ,
         \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 ,
         \10798 , \10799 , \10800 , \10801 , \10802 , \10803_nG36aa , \10804 , \10805 , \10806 , \10807 ,
         \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 ,
         \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 ,
         \10828 , \10829 , \10830_nG3493 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 ,
         \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 ,
         \10848 , \10849 , \10850 , \10851_nG3564 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 ,
         \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 ,
         \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874_nG3451 , \10875 , \10876 , \10877 ,
         \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 ,
         \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 ,
         \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 ,
         \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 ,
         \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 ,
         \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 ,
         \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 ,
         \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 ,
         \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 ,
         \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 ,
         \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 ,
         \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 ,
         \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007_nG333d ,
         \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 ,
         \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 ,
         \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 ,
         \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 ,
         \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 ,
         \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 ,
         \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 ,
         \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 ,
         \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 ,
         \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 ,
         \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 ,
         \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 ,
         \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 ,
         \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 ,
         \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 ,
         \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 ,
         \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 ,
         \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 ,
         \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 ,
         \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 ,
         \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 ,
         \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 ,
         \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 ,
         \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 ,
         \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 ,
         \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 ,
         \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 ,
         \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 ,
         \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 ,
         \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 ,
         \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 ,
         \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 ,
         \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 ,
         \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 ,
         \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 ,
         \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 ,
         \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 ,
         \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 ,
         \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 ,
         \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 ,
         \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 ,
         \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 ,
         \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 ,
         \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 ,
         \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 ,
         \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 ,
         \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 ,
         \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 ,
         \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 ,
         \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 ,
         \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 ,
         \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 ,
         \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 ,
         \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 ,
         \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 ,
         \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 ,
         \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 ,
         \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 ,
         \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 ,
         \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 ,
         \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 ,
         \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 ,
         \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 ,
         \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 ,
         \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 ,
         \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 ,
         \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 ,
         \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 ,
         \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 ,
         \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 ,
         \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 ,
         \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 ,
         \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 ,
         \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 ,
         \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 ,
         \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 ,
         \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 ,
         \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 ,
         \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 ,
         \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 ,
         \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 ,
         \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 ,
         \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 ,
         \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 ,
         \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 ,
         \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 ,
         \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 ,
         \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 ,
         \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 ,
         \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 ,
         \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 ,
         \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 ,
         \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 ,
         \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 ,
         \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 ,
         \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 ,
         \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 ,
         \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 ,
         \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 ,
         \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 ,
         \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 ,
         \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 ,
         \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 ,
         \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 ,
         \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 ,
         \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 ,
         \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 ,
         \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 ,
         \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 ,
         \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 ,
         \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 ,
         \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 ,
         \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 ,
         \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 ,
         \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 ,
         \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 ,
         \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 ,
         \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 ,
         \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 ,
         \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 ,
         \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 ,
         \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 ,
         \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 ,
         \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 ,
         \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 ,
         \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 ,
         \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 ,
         \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 ,
         \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 ,
         \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 ,
         \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 ,
         \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 ,
         \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 ,
         \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 ,
         \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 ,
         \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 ,
         \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 ,
         \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 ,
         \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 ,
         \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 ,
         \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 ,
         \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 ,
         \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 ,
         \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 ,
         \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 ,
         \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 ,
         \12468 , \12469 , \12470_nG4b72 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 ,
         \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 ,
         \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 ,
         \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 ,
         \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 ,
         \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 ,
         \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 ,
         \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 ,
         \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 ,
         \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 ,
         \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 ,
         \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 ,
         \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 ,
         \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 ,
         \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 ,
         \12618 , \12619_nG3b20 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 ,
         \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 ,
         \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644_nG3afc , \12645 , \12646 , \12647 ,
         \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 ,
         \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 ,
         \12668 , \12669_nG3969 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 ,
         \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 ,
         \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694_nG3945 , \12695 , \12696 , \12697 ,
         \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 ,
         \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 ,
         \12718 , \12719_nG37c6 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 ,
         \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 ,
         \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744_nG37a2 , \12745 , \12746 , \12747 ,
         \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 ,
         \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 ,
         \12768 , \12769_nG3657 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 ,
         \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 ,
         \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794_nG3633 , \12795 , \12796 , \12797 ,
         \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 ,
         \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 ,
         \12818 , \12819_nG3518 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 ,
         \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 ,
         \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844_nG3531 , \12845 , \12846 , \12847 ,
         \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 ,
         \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 ,
         \12868 , \12869_nG342e , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 ,
         \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 ,
         \12888 , \12889 , \12890 , \12891 , \12892 , \12893_nG3412 , \12894 , \12895 , \12896 , \12897 ,
         \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 ,
         \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 ,
         \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 ,
         \12928_nG3b29 , \12929 , \12930 , \12931 , \12932_nG3b05 , \12933 , \12934 , \12935 , \12936_nG3972 , \12937 ,
         \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 ,
         \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 ,
         \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 ,
         \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 ,
         \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 ,
         \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 ,
         \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 ,
         \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 ,
         \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 ,
         \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 ,
         \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 ,
         \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 ,
         \13058 , \13059 , \13060 , \13061 , \13062_nG41fa , \13063 , \13064 , \13065 , \13066 , \13067 ,
         \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 ,
         \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 ,
         \13088 , \13089 , \13090_nG3cdb , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 ,
         \13098 , \13099 , \13100 , \13101 , \13102_nG3cf0 , \13103 , \13104 , \13105 , \13106_nG3ce4 , \13107 ,
         \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 ,
         \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 ,
         \13128 , \13129 , \13130 , \13131_nG42ef , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 ,
         \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 ,
         \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 ,
         \13158_nG4131 , \13159 , \13160 , \13161 , \13162_nG3eca , \13163 , \13164 , \13165 , \13166 , \13167 ,
         \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 ,
         \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 ,
         \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 ,
         \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 ,
         \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 ,
         \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 ,
         \13228 , \13229_nG394e , \13230 , \13231 , \13232 , \13233 , \13234_nG37cf , \13235 , \13236 , \13237 ,
         \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 ,
         \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 ,
         \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 ,
         \13268 , \13269_nG3f92 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 ,
         \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 ,
         \13288 , \13289 , \13290_nG4070 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 ,
         \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 ,
         \13308 , \13309 , \13310 , \13311 , \13312 , \13313_nG3ea9 , \13314 , \13315 , \13316 , \13317 ,
         \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 ,
         \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 ,
         \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 ,
         \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 ,
         \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 ,
         \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376_nG3435 , \13377 ,
         \13378 , \13379_nG3415 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 ,
         \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 ,
         \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406_nG3d18 , \13407 ,
         \13408 , \13409 , \13410_nG353d , \13411 , \13412 , \13413 , \13414_nG3541 , \13415 , \13416 , \13417 ,
         \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 ,
         \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 ,
         \13438 , \13439_nG3dc5 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 ,
         \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 ,
         \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466_nG3b58 , \13467 ,
         \13468 , \13469 , \13470_nG3660 , \13471 , \13472 , \13473 , \13474_nG363c , \13475 , \13476 , \13477 ,
         \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 ,
         \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 ,
         \13498 , \13499_nG3bf0 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 ,
         \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 ,
         \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 ,
         \13528_nG398d , \13529 , \13530 , \13531 , \13532_nG37ab , \13533 , \13534 , \13535 , \13536 , \13537 ,
         \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 ,
         \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557_nG3a17 ,
         \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 ,
         \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 ,
         \13578 , \13579 , \13580 , \13581 , \13582 , \13583_nG37ea , \13584 , \13585 , \13586 , \13587 ,
         \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 ,
         \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604_nG385e , \13605 , \13606 , \13607 ,
         \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 ,
         \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 ,
         \13628_nG3679 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 ,
         \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 ,
         \13648 , \13649_nG36e0 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 ,
         \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 ,
         \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676_nG34fb , \13677 ,
         \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 ,
         \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697_nG358e ,
         \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 ,
         \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 ,
         \13718 , \13719 , \13720_nG3473 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 ,
         \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 ,
         \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 ,
         \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 ,
         \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 ,
         \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 ,
         \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 ,
         \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 ,
         \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 ,
         \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 ,
         \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 ,
         \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 ,
         \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 ,
         \13848 , \13849 , \13850 , \13851 , \13852 , \13853_nG33d8 , \13854 , \13855 , \13856 , \13857 ,
         \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 ,
         \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 ,
         \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 ,
         \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 ,
         \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 ,
         \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 ,
         \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 ,
         \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 ,
         \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 ,
         \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 ,
         \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 ,
         \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 ,
         \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 ,
         \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 ,
         \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 ,
         \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 ,
         \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 ,
         \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 ,
         \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 ,
         \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 ,
         \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 ,
         \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 ,
         \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 ,
         \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 ,
         \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 ,
         \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 ,
         \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 ,
         \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 ,
         \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 ,
         \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 ,
         \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 ,
         \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 ,
         \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 ,
         \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 ,
         \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 ,
         \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 ,
         \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 ,
         \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 ,
         \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 ,
         \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 ,
         \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 ,
         \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 ,
         \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 ,
         \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 ,
         \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 ,
         \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 ,
         \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 ,
         \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 ,
         \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 ,
         \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 ,
         \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 ,
         \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 ,
         \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 ,
         \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 ,
         \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 ,
         \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 ,
         \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 ,
         \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 ,
         \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 ,
         \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 ,
         \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 ,
         \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 ,
         \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 ,
         \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 ,
         \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 ,
         \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 ,
         \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 ,
         \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 ,
         \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 ,
         \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 ,
         \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 ,
         \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 ,
         \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 ,
         \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 ,
         \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 ,
         \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 ,
         \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 ,
         \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 ,
         \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 ,
         \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 ,
         \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 ,
         \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 ,
         \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 ,
         \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 ,
         \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 ,
         \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 ,
         \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 ,
         \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 ,
         \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 ,
         \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 ,
         \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 ,
         \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 ,
         \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 ,
         \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 ,
         \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 ,
         \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 ,
         \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 ,
         \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 ,
         \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 ,
         \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 ,
         \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 ,
         \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 ,
         \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 ,
         \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 ,
         \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 ,
         \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 ,
         \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 ,
         \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 ,
         \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 ,
         \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 ,
         \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 ,
         \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 ,
         \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 ,
         \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 ,
         \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 ,
         \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 ,
         \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 ,
         \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 ,
         \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 ,
         \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 ,
         \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 ,
         \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 ,
         \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 ,
         \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 ,
         \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 ,
         \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 ,
         \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 ,
         \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 ,
         \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 ,
         \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 ,
         \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 ,
         \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 ,
         \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 ,
         \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 ,
         \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 ,
         \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 ,
         \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 ,
         \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 ,
         \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 ,
         \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 ,
         \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 ,
         \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 ,
         \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 ,
         \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 ,
         \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 ,
         \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316_nG4ba0 , \15317 ,
         \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 ,
         \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 ,
         \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 ,
         \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 ,
         \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 ,
         \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 ,
         \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 ,
         \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 ,
         \15398_nG1512 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 ,
         \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 ,
         \15418 , \15419 , \15420 , \15421 , \15422 , \15423_nG152b , \15424 , \15425 , \15426 , \15427 ,
         \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 ,
         \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 ,
         \15448_nG1544 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 ,
         \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 ,
         \15468 , \15469 , \15470 , \15471 , \15472 , \15473_nG155d , \15474 , \15475 , \15476 , \15477 ,
         \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 ,
         \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 ,
         \15498_nG1576 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 ,
         \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 ,
         \15518 , \15519 , \15520 , \15521 , \15522 , \15523_nG158f , \15524 , \15525 , \15526 , \15527 ,
         \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 ,
         \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 ,
         \15548_nG15a8 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 ,
         \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 ,
         \15568 , \15569 , \15570 , \15571 , \15572 , \15573_nG15c1 , \15574 , \15575 , \15576 , \15577 ,
         \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 ,
         \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 ,
         \15598_nG15da , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 ,
         \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 ,
         \15618 , \15619 , \15620 , \15621 , \15622 , \15623_nG15f3 , \15624 , \15625 , \15626 , \15627 ,
         \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 ,
         \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 ,
         \15648_nG160c , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 ,
         \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 ,
         \15668 , \15669 , \15670 , \15671 , \15672 , \15673_nG1625 , \15674 , \15675 , \15676 , \15677 ,
         \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 ,
         \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697_nG163f ,
         \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 ,
         \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 ,
         \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 ,
         \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 ,
         \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 ,
         \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 ,
         \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 ,
         \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 ,
         \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 ,
         \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 ,
         \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807_nG16b2 ,
         \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 ,
         \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 ,
         \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 ,
         \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 ,
         \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 ,
         \15858 , \15859 , \15860 , \15861 , \15862_nG16e9 , \15863 , \15864 , \15865 , \15866 , \15867 ,
         \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 ,
         \15878 , \15879 , \15880 , \15881 , \15882 , \15883_nG16fe , \15884 , \15885 , \15886 , \15887 ,
         \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 ,
         \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904_nG1713 , \15905 , \15906 , \15907 ,
         \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 ,
         \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925_nG1728 , \15926 , \15927 ,
         \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 ,
         \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946_nG173d , \15947 ,
         \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 ,
         \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967_nG1752 ,
         \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 ,
         \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 ,
         \15988_nG1767 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 ,
         \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 ,
         \16008 , \16009_nG177c , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 ,
         \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 ,
         \16028 , \16029 , \16030_nG1791 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 ,
         \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 ,
         \16048 , \16049 , \16050 , \16051_nG17a6 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 ,
         \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 ,
         \16068 , \16069 , \16070 , \16071 , \16072_nG17bb , \16073 , \16074 , \16075 , \16076 , \16077 ,
         \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 ,
         \16088 , \16089 , \16090 , \16091 , \16092 , \16093_nG17d0 , \16094 , \16095 , \16096 , \16097 ,
         \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 ,
         \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114_nG17e5 , \16115 , \16116 , \16117 ,
         \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 ,
         \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135_nG17fa , \16136 , \16137 ,
         \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 ,
         \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156_nG180f , \16157 ,
         \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 ,
         \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177_nG1824 ,
         \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 ,
         \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 ,
         \16198_nG1839 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 ,
         \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 ,
         \16218 , \16219_nG184e , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 ,
         \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 ,
         \16238 , \16239 , \16240_nG1863 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 ,
         \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 ,
         \16258 , \16259 , \16260 , \16261_nG1878 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 ,
         \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 ,
         \16278 , \16279 , \16280 , \16281 , \16282_nG188d , \16283 , \16284 , \16285 , \16286 , \16287 ,
         \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 ,
         \16298 , \16299 , \16300 , \16301 , \16302 , \16303_nG18a2 , \16304 , \16305 , \16306 , \16307 ,
         \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 ,
         \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324_nG18b7 , \16325 , \16326 , \16327 ,
         \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 ,
         \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345_nG18cc , \16346 , \16347 ,
         \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 ,
         \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366_nG18e1 , \16367 ,
         \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 ,
         \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 ,
         \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 ,
         \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407_nG4ba1 ,
         \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 ,
         \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 ,
         \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 ,
         \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 ,
         \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 ,
         \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 ,
         \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 ,
         \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 ,
         \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 ,
         \16498 , \16499 , \16500_nG4b0f , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 ,
         \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 ,
         \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 ,
         \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 ,
         \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 ,
         \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 ,
         \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 ,
         \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 ,
         \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 ,
         \16588 , \16589 , \16590 , \16591 , \16592_nG4b43 , \16593_nG4b44 , \16594 , \16595 , \16596 , \16597 ,
         \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 ,
         \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 ,
         \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 ,
         \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 ,
         \16638 , \16639_nG4aa0 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 ,
         \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 ,
         \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 ,
         \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 ,
         \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684_nG4ada , \16685_nG4adb , \16686 , \16687 ,
         \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 ,
         \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 ,
         \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 ,
         \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 ,
         \16728 , \16729 , \16730_nG4a23 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 ,
         \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 ,
         \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 ,
         \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 ,
         \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774_nG4a65 , \16775_nG4a66 , \16776 , \16777 ,
         \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 ,
         \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 ,
         \16798_nG499a , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 ,
         \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 ,
         \16818 , \16819 , \16820_nG49e0 , \16821_nG49e1 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 ,
         \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 ,
         \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844_nG490b , \16845 , \16846 , \16847 ,
         \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 ,
         \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866_nG4953 , \16867_nG4954 ,
         \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 ,
         \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 ,
         \16888 , \16889_nG4876 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 ,
         \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 ,
         \16908 , \16909 , \16910_nG48c2 , \16911_nG48c3 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 ,
         \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 ,
         \16928 , \16929 , \16930 , \16931 , \16932 , \16933_nG47d9 , \16934 , \16935 , \16936 , \16937 ,
         \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 ,
         \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954_nG4829 , \16955_nG482a , \16956 , \16957 ,
         \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967_nG4737 ,
         \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 ,
         \16978_nG4788 , \16979_nG4789 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 ,
         \16988 , \16989 , \16990 , \16991_nG468c , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 ,
         \16998 , \16999 , \17000 , \17001 , \17002_nG46e5 , \17003_nG46e6 , \17004 , \17005 , \17006 , \17007 ,
         \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 , \17015_nG45d6 , \17016 , \17017 ,
         \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026_nG4632 , \17027_nG4633 ,
         \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 ,
         \17038 , \17039_nG4519 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 ,
         \17048 , \17049 , \17050_nG4579 , \17051_nG457a , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 ,
         \17058 , \17059 , \17060 , \17061 , \17062_nG4459 , \17063 , \17064 , \17065 , \17066 , \17067 ,
         \17068 , \17069 , \17070 , \17071 , \17072_nG44b8 , \17073_nG44b9 , \17074 , \17075 , \17076 , \17077 ,
         \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084_nG439a , \17085 , \17086 , \17087 ,
         \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094_nG43f9 , \17095_nG43fa , \17096 , \17097 ,
         \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106_nG42c6 , \17107 ,
         \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116_nG433a , \17117_nG433b ,
         \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 ,
         \17128_nG41de , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 ,
         \17138_nG4251 , \17139_nG4252 , \17140 , \17141 , \17142 , \17143 , \17144_nG40fe , \17145 , \17146 , \17147 ,
         \17148_nG416a , \17149_nG416b , \17150 , \17151 , \17152 , \17153 , \17154_nG4025 , \17155 , \17156 , \17157 ,
         \17158_nG4091 , \17159_nG4092 , \17160 , \17161 , \17162 , \17163 , \17164_nG3f50 , \17165 , \17166 , \17167 ,
         \17168_nG3fb8 , \17169_nG3fb9 , \17170 , \17171 , \17172 , \17173 , \17174_nG3e7d , \17175 , \17176 , \17177 ,
         \17178_nG3ee7 , \17179_nG3ee8 , \17180 , \17181 , \17182 , \17183 , \17184_nG3dad , \17185 , \17186 , \17187 ,
         \17188_nG3e12 , \17189_nG3e13 , \17190 , \17191 , \17192 , \17193 , \17194_nG3cbb , \17195 , \17196 , \17197 ,
         \17198_nG3d47 , \17199_nG3d48 , \17200 , \17201 , \17202 , \17203 , \17204_nG3bd4 , \17205 , \17206 , \17207 ,
         \17208_nG3c2e , \17209_nG3c2f , \17210 , \17211 , \17212 , \17213 , \17214_nG3ae0 , \17215 , \17216 , \17217 ,
         \17218_nG3b79 , \17219_nG3b7a , \17220 , \17221 , \17222 , \17223 , \17224_nG39f8 , \17225 , \17226 , \17227 ,
         \17228_nG3a46 , \17229_nG3a47 , \17230 , \17231 , \17232 , \17233 , \17234_nG391c , \17235 , \17236 , \17237 ,
         \17238_nG39a9 , \17239_nG39aa , \17240 , \17241 , \17242 , \17243 , \17244_nG384a , \17245 , \17246 , \17247 ,
         \17248_nG388e , \17249_nG388f , \17250 ;
buf \U$labaj1799 ( R_289_8400778, \8850 );
buf \U$labaj1800 ( R_28a_8401e70, \9036 );
buf \U$labaj1801 ( R_28b_8401f18, \9128 );
buf \U$labaj1802 ( R_28c_8401fc0, \9218 );
buf \U$labaj1803 ( R_28d_8402068, \9264 );
buf \U$labaj1804 ( R_28e_8402110, \9310 );
buf \U$labaj1805 ( R_28f_84021b8, \9354 );
buf \U$labaj1806 ( R_290_8402260, \9398 );
buf \U$labaj1807 ( R_291_8402308, \9422 );
buf \U$labaj1808 ( R_292_84023b0, \9446 );
buf \U$labaj1809 ( R_293_8402458, \9470 );
buf \U$labaj1810 ( R_294_8402500, \9494 );
buf \U$labaj1811 ( R_295_84025a8, \9516 );
buf \U$labaj1812 ( R_296_8402650, \9538 );
buf \U$labaj1813 ( R_297_84026f8, \9560 );
buf \U$labaj1814 ( R_298_84027a0, \9582 );
buf \U$labaj1815 ( R_299_8402848, \9592 );
buf \U$labaj1816 ( R_29a_84028f0, \9602 );
buf \U$labaj1817 ( R_29b_8402998, \9612 );
buf \U$labaj1818 ( R_29c_8402a40, \9622 );
buf \U$labaj1819 ( R_29d_8402ae8, \9632 );
buf \U$labaj1820 ( R_29e_8402b90, \9642 );
buf \U$labaj1821 ( R_29f_8402c38, \9652 );
buf \U$labaj1822 ( R_2a0_8402ce0, \9662 );
buf \U$labaj1823 ( R_2a1_8402d88, \9672 );
buf \U$labaj1824 ( R_2a2_8402e30, \9682 );
buf \U$labaj1825 ( R_2a3_8402ed8, \9692 );
buf \U$labaj1826 ( R_267_8403418, \16408 );
buf \U$labaj1827 ( R_268_8400820, \16594 );
buf \U$labaj1828 ( R_269_84008c8, \16686 );
buf \U$labaj1829 ( R_26a_8400970, \16776 );
buf \U$labaj1830 ( R_26b_8400a18, \16822 );
buf \U$labaj1831 ( R_26c_8400ac0, \16868 );
buf \U$labaj1832 ( R_26d_8400b68, \16912 );
buf \U$labaj1833 ( R_26e_8400c10, \16956 );
buf \U$labaj1834 ( R_26f_8400cb8, \16980 );
buf \U$labaj1835 ( R_270_8400d60, \17004 );
buf \U$labaj1836 ( R_271_8400e08, \17028 );
buf \U$labaj1837 ( R_272_8400eb0, \17052 );
buf \U$labaj1838 ( R_273_8400f58, \17074 );
buf \U$labaj1839 ( R_274_8401000, \17096 );
buf \U$labaj1840 ( R_275_84010a8, \17118 );
buf \U$labaj1841 ( R_276_8401150, \17140 );
buf \U$labaj1842 ( R_277_84011f8, \17150 );
buf \U$labaj1843 ( R_278_84012a0, \17160 );
buf \U$labaj1844 ( R_279_8401348, \17170 );
buf \U$labaj1845 ( R_27a_84013f0, \17180 );
buf \U$labaj1846 ( R_27b_8401498, \17190 );
buf \U$labaj1847 ( R_27c_8401540, \17200 );
buf \U$labaj1848 ( R_27d_84015e8, \17210 );
buf \U$labaj1849 ( R_27e_8401690, \17220 );
buf \U$labaj1850 ( R_27f_8401738, \17230 );
buf \U$labaj1851 ( R_280_84017e0, \17240 );
buf \U$labaj1852 ( R_281_8401888, \17250 );
buf \U$5 ( \2135 , RI994e3e8_15);
buf \U$6 ( \2136 , RI994e370_16);
buf \U$7 ( \2137 , RI994e2f8_17);
buf \U$8 ( \2138 , RI994e280_18);
buf \U$9 ( \2139 , RI994e208_19);
buf \U$10 ( \2140 , RI994e190_20);
buf \U$11 ( \2141 , RI994e118_21);
buf \U$12 ( \2142 , RI994e0a0_22);
buf \U$13 ( \2143 , RI994e028_23);
buf \U$14 ( \2144 , RI994dfb0_24);
buf \U$15 ( \2145 , RI994df38_25);
and \U$16 ( \2146 , \2144 , \2145 );
and \U$17 ( \2147 , \2143 , \2146 );
and \U$18 ( \2148 , \2142 , \2147 );
and \U$19 ( \2149 , \2141 , \2148 );
and \U$20 ( \2150 , \2140 , \2149 );
and \U$21 ( \2151 , \2139 , \2150 );
and \U$22 ( \2152 , \2138 , \2151 );
and \U$23 ( \2153 , \2137 , \2152 );
and \U$24 ( \2154 , \2136 , \2153 );
xor \U$25 ( \2155 , \2135 , \2154 );
buf \U$26 ( \2156 , \2155 );
buf \U$27 ( \2157 , \2156 );
not \U$28 ( \2158 , RI9921910_609);
nor \U$29 ( \2159 , RI9921730_613, RI99217a8_612, RI9921820_611, RI9921898_610, \2158 , RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$30 ( \2160 , RI995e450_236, \2159 );
not \U$31 ( \2161 , RI9921730_613);
not \U$32 ( \2162 , RI99217a8_612);
not \U$33 ( \2163 , RI9921820_611);
not \U$34 ( \2164 , RI9921898_610);
nor \U$35 ( \2165 , \2161 , \2162 , \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$36 ( \2166 , RI9967078_223, \2165 );
nor \U$37 ( \2167 , RI9921730_613, \2162 , \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$38 ( \2168 , RI9967690_210, \2167 );
nor \U$39 ( \2169 , \2161 , RI99217a8_612, \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$40 ( \2170 , RI890fba0_197, \2169 );
nor \U$41 ( \2171 , RI9921730_613, RI99217a8_612, \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$42 ( \2172 , RI8918b88_184, \2171 );
nor \U$43 ( \2173 , \2161 , \2162 , RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$44 ( \2174 , RI89253b0_171, \2173 );
nor \U$45 ( \2175 , RI9921730_613, \2162 , RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$46 ( \2176 , RI8930dc8_158, \2175 );
nor \U$47 ( \2177 , \2161 , RI99217a8_612, RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$48 ( \2178 , RI8939db0_145, \2177 );
nor \U$49 ( \2179 , RI9921730_613, RI99217a8_612, RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$50 ( \2180 , RI89465d8_132, \2179 );
nor \U$51 ( \2181 , \2161 , \2162 , \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$52 ( \2182 , RI89ec640_119, \2181 );
nor \U$53 ( \2183 , RI9921730_613, \2162 , \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$54 ( \2184 , RI9776f80_106, \2183 );
nor \U$55 ( \2185 , \2161 , RI99217a8_612, \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$56 ( \2186 , RI9808480_93, \2185 );
nor \U$57 ( \2187 , RI9921730_613, RI99217a8_612, \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$58 ( \2188 , RI9808a98_80, \2187 );
nor \U$59 ( \2189 , \2161 , \2162 , RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$60 ( \2190 , RI9819730_67, \2189 );
nor \U$61 ( \2191 , RI9921730_613, \2162 , RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$62 ( \2192 , RI98abc38_54, \2191 );
nor \U$63 ( \2193 , \2161 , RI99217a8_612, RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$64 ( \2194 , RI98bc8d0_41, \2193 );
nor \U$65 ( \2195 , RI9921730_613, RI99217a8_612, RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$66 ( \2196 , RI994ddd0_28, \2195 );
or \U$67 ( \2197 , \2160 , \2166 , \2168 , \2170 , \2172 , \2174 , \2176 , \2178 , \2180 , \2182 , \2184 , \2186 , \2188 , \2190 , \2192 , \2194 , \2196 );
buf \U$68 ( \2198 , RI9921988_608);
buf \U$69 ( \2199 , RI9921a00_607);
buf \U$70 ( \2200 , RI9921a78_606);
buf \U$71 ( \2201 , RI9921af0_605);
buf \U$72 ( \2202 , RI9921b68_604);
buf \U$73 ( \2203 , RI9921be0_603);
buf \U$74 ( \2204 , RI9921c58_602);
buf \U$75 ( \2205 , RI9921cd0_601);
buf \U$76 ( \2206 , RI9921910_609);
buf \U$77 ( \2207 , RI9921730_613);
buf \U$78 ( \2208 , RI99217a8_612);
buf \U$79 ( \2209 , RI9921820_611);
buf \U$80 ( \2210 , RI9921898_610);
or \U$81 ( \2211 , \2207 , \2208 , \2209 , \2210 );
and \U$82 ( \2212 , \2206 , \2211 );
or \U$83 ( \2213 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2212 );
buf \U$84 ( \2214 , \2213 );
_DC g2199 ( \2215_nG2199 , \2197 , \2214 );
buf \U$85 ( \2216 , \2215_nG2199 );
not \U$86 ( \2217 , \2216 );
xor \U$87 ( \2218 , \2157 , \2217 );
xor \U$88 ( \2219 , \2136 , \2153 );
buf \U$89 ( \2220 , \2219 );
buf \U$90 ( \2221 , \2220 );
and \U$91 ( \2222 , RI995e3d8_237, \2159 );
and \U$92 ( \2223 , RI99669e8_224, \2165 );
and \U$93 ( \2224 , RI9967618_211, \2167 );
and \U$94 ( \2225 , RI890fb28_198, \2169 );
and \U$95 ( \2226 , RI8918b10_185, \2171 );
and \U$96 ( \2227 , RI8925338_172, \2173 );
and \U$97 ( \2228 , RI8930d50_159, \2175 );
and \U$98 ( \2229 , RI8939d38_146, \2177 );
and \U$99 ( \2230 , RI8946560_133, \2179 );
and \U$100 ( \2231 , RI89ec5c8_120, \2181 );
and \U$101 ( \2232 , RI9776f08_107, \2183 );
and \U$102 ( \2233 , RI9808408_94, \2185 );
and \U$103 ( \2234 , RI9808a20_81, \2187 );
and \U$104 ( \2235 , RI98196b8_68, \2189 );
and \U$105 ( \2236 , RI98abbc0_55, \2191 );
and \U$106 ( \2237 , RI98bc858_42, \2193 );
and \U$107 ( \2238 , RI994dd58_29, \2195 );
or \U$108 ( \2239 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 );
_DC g2175 ( \2240_nG2175 , \2239 , \2214 );
buf \U$109 ( \2241 , \2240_nG2175 );
not \U$110 ( \2242 , \2241 );
and \U$111 ( \2243 , \2221 , \2242 );
xor \U$112 ( \2244 , \2137 , \2152 );
buf \U$113 ( \2245 , \2244 );
buf \U$114 ( \2246 , \2245 );
and \U$115 ( \2247 , RI9959fe0_238, \2159 );
and \U$116 ( \2248 , RI995e978_225, \2165 );
and \U$117 ( \2249 , RI99675a0_212, \2167 );
and \U$118 ( \2250 , RI890fab0_199, \2169 );
and \U$119 ( \2251 , RI8918a98_186, \2171 );
and \U$120 ( \2252 , RI89252c0_173, \2173 );
and \U$121 ( \2253 , RI8930cd8_160, \2175 );
and \U$122 ( \2254 , RI8939cc0_147, \2177 );
and \U$123 ( \2255 , RI89464e8_134, \2179 );
and \U$124 ( \2256 , RI89ec550_121, \2181 );
and \U$125 ( \2257 , RI9776e90_108, \2183 );
and \U$126 ( \2258 , RI9808390_95, \2185 );
and \U$127 ( \2259 , RI98089a8_82, \2187 );
and \U$128 ( \2260 , RI9819640_69, \2189 );
and \U$129 ( \2261 , RI98abb48_56, \2191 );
and \U$130 ( \2262 , RI98bc7e0_43, \2193 );
and \U$131 ( \2263 , RI994dce0_30, \2195 );
or \U$132 ( \2264 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 );
_DC g1fee ( \2265_nG1fee , \2264 , \2214 );
buf \U$133 ( \2266 , \2265_nG1fee );
not \U$134 ( \2267 , \2266 );
and \U$135 ( \2268 , \2246 , \2267 );
xor \U$136 ( \2269 , \2138 , \2151 );
buf \U$137 ( \2270 , \2269 );
buf \U$138 ( \2271 , \2270 );
and \U$139 ( \2272 , RI9959f68_239, \2159 );
and \U$140 ( \2273 , RI995e900_226, \2165 );
and \U$141 ( \2274 , RI9967528_213, \2167 );
and \U$142 ( \2275 , RI890fa38_200, \2169 );
and \U$143 ( \2276 , RI8918a20_187, \2171 );
and \U$144 ( \2277 , RI8925248_174, \2173 );
and \U$145 ( \2278 , RI8930c60_161, \2175 );
and \U$146 ( \2279 , RI8939c48_148, \2177 );
and \U$147 ( \2280 , RI8946470_135, \2179 );
and \U$148 ( \2281 , RI89ec4d8_122, \2181 );
and \U$149 ( \2282 , RI9776e18_109, \2183 );
and \U$150 ( \2283 , RI9808318_96, \2185 );
and \U$151 ( \2284 , RI9808930_83, \2187 );
and \U$152 ( \2285 , RI98195c8_70, \2189 );
and \U$153 ( \2286 , RI98abad0_57, \2191 );
and \U$154 ( \2287 , RI98bc768_44, \2193 );
and \U$155 ( \2288 , RI994dc68_31, \2195 );
or \U$156 ( \2289 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 );
_DC g1fca ( \2290_nG1fca , \2289 , \2214 );
buf \U$157 ( \2291 , \2290_nG1fca );
not \U$158 ( \2292 , \2291 );
and \U$159 ( \2293 , \2271 , \2292 );
xor \U$160 ( \2294 , \2139 , \2150 );
buf \U$161 ( \2295 , \2294 );
buf \U$162 ( \2296 , \2295 );
and \U$163 ( \2297 , RI9959860_240, \2159 );
and \U$164 ( \2298 , RI995e888_227, \2165 );
and \U$165 ( \2299 , RI99674b0_214, \2167 );
and \U$166 ( \2300 , RI890f9c0_201, \2169 );
and \U$167 ( \2301 , RI89189a8_188, \2171 );
and \U$168 ( \2302 , RI89251d0_175, \2173 );
and \U$169 ( \2303 , RI8930be8_162, \2175 );
and \U$170 ( \2304 , RI8939bd0_149, \2177 );
and \U$171 ( \2305 , RI89463f8_136, \2179 );
and \U$172 ( \2306 , RI89ec460_123, \2181 );
and \U$173 ( \2307 , RI9776da0_110, \2183 );
and \U$174 ( \2308 , RI98082a0_97, \2185 );
and \U$175 ( \2309 , RI98088b8_84, \2187 );
and \U$176 ( \2310 , RI9819550_71, \2189 );
and \U$177 ( \2311 , RI98aba58_58, \2191 );
and \U$178 ( \2312 , RI98bc6f0_45, \2193 );
and \U$179 ( \2313 , RI994dbf0_32, \2195 );
or \U$180 ( \2314 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 );
_DC g1e55 ( \2315_nG1e55 , \2314 , \2214 );
buf \U$181 ( \2316 , \2315_nG1e55 );
not \U$182 ( \2317 , \2316 );
and \U$183 ( \2318 , \2296 , \2317 );
xor \U$184 ( \2319 , \2140 , \2149 );
buf \U$185 ( \2320 , \2319 );
buf \U$186 ( \2321 , \2320 );
and \U$187 ( \2322 , RI994d998_241, \2159 );
and \U$188 ( \2323 , RI995e810_228, \2165 );
and \U$189 ( \2324 , RI9967438_215, \2167 );
and \U$190 ( \2325 , RI890f948_202, \2169 );
and \U$191 ( \2326 , RI8918930_189, \2171 );
and \U$192 ( \2327 , RI8925158_176, \2173 );
and \U$193 ( \2328 , RI8930b70_163, \2175 );
and \U$194 ( \2329 , RI8939b58_150, \2177 );
and \U$195 ( \2330 , RI8946380_137, \2179 );
and \U$196 ( \2331 , RI89ec3e8_124, \2181 );
and \U$197 ( \2332 , RI9776d28_111, \2183 );
and \U$198 ( \2333 , RI9808228_98, \2185 );
and \U$199 ( \2334 , RI9808840_85, \2187 );
and \U$200 ( \2335 , RI98194d8_72, \2189 );
and \U$201 ( \2336 , RI98ab9e0_59, \2191 );
and \U$202 ( \2337 , RI98abff8_46, \2193 );
and \U$203 ( \2338 , RI98bcc90_33, \2195 );
or \U$204 ( \2339 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 );
_DC g1e31 ( \2340_nG1e31 , \2339 , \2214 );
buf \U$205 ( \2341 , \2340_nG1e31 );
not \U$206 ( \2342 , \2341 );
and \U$207 ( \2343 , \2321 , \2342 );
xor \U$208 ( \2344 , \2141 , \2148 );
buf \U$209 ( \2345 , \2344 );
buf \U$210 ( \2346 , \2345 );
and \U$211 ( \2347 , RI994d920_242, \2159 );
and \U$212 ( \2348 , RI995e798_229, \2165 );
and \U$213 ( \2349 , RI99673c0_216, \2167 );
and \U$214 ( \2350 , RI890f8d0_203, \2169 );
and \U$215 ( \2351 , RI89188b8_190, \2171 );
and \U$216 ( \2352 , RI89250e0_177, \2173 );
and \U$217 ( \2353 , RI8930af8_164, \2175 );
and \U$218 ( \2354 , RI8939ae0_151, \2177 );
and \U$219 ( \2355 , RI8946308_138, \2179 );
and \U$220 ( \2356 , RI89ec370_125, \2181 );
and \U$221 ( \2357 , RI89ec988_112, \2183 );
and \U$222 ( \2358 , RI97772c8_99, \2185 );
and \U$223 ( \2359 , RI98087c8_86, \2187 );
and \U$224 ( \2360 , RI9819460_73, \2189 );
and \U$225 ( \2361 , RI98ab968_60, \2191 );
and \U$226 ( \2362 , RI98abf80_47, \2193 );
and \U$227 ( \2363 , RI98bcc18_34, \2195 );
or \U$228 ( \2364 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 );
_DC g1cf3 ( \2365_nG1cf3 , \2364 , \2214 );
buf \U$229 ( \2366 , \2365_nG1cf3 );
not \U$230 ( \2367 , \2366 );
and \U$231 ( \2368 , \2346 , \2367 );
xor \U$232 ( \2369 , \2142 , \2147 );
buf \U$233 ( \2370 , \2369 );
buf \U$234 ( \2371 , \2370 );
and \U$235 ( \2372 , RI994d8a8_243, \2159 );
and \U$236 ( \2373 , RI995e720_230, \2165 );
and \U$237 ( \2374 , RI9967348_217, \2167 );
and \U$238 ( \2375 , RI890f858_204, \2169 );
and \U$239 ( \2376 , RI8918840_191, \2171 );
and \U$240 ( \2377 , RI8925068_178, \2173 );
and \U$241 ( \2378 , RI8930a80_165, \2175 );
and \U$242 ( \2379 , RI8939a68_152, \2177 );
and \U$243 ( \2380 , RI8946290_139, \2179 );
and \U$244 ( \2381 , RI89ec2f8_126, \2181 );
and \U$245 ( \2382 , RI89ec910_113, \2183 );
and \U$246 ( \2383 , RI9777250_100, \2185 );
and \U$247 ( \2384 , RI9808750_87, \2187 );
and \U$248 ( \2385 , RI98193e8_74, \2189 );
and \U$249 ( \2386 , RI98ab8f0_61, \2191 );
and \U$250 ( \2387 , RI98abf08_48, \2193 );
and \U$251 ( \2388 , RI98bcba0_35, \2195 );
or \U$252 ( \2389 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 );
_DC g1ccf ( \2390_nG1ccf , \2389 , \2214 );
buf \U$253 ( \2391 , \2390_nG1ccf );
not \U$254 ( \2392 , \2391 );
and \U$255 ( \2393 , \2371 , \2392 );
xor \U$256 ( \2394 , \2143 , \2146 );
buf \U$257 ( \2395 , \2394 );
buf \U$258 ( \2396 , \2395 );
and \U$259 ( \2397 , RI994d830_244, \2159 );
and \U$260 ( \2398 , RI995e6a8_231, \2165 );
and \U$261 ( \2399 , RI99672d0_218, \2167 );
and \U$262 ( \2400 , RI890f7e0_205, \2169 );
and \U$263 ( \2401 , RI89187c8_192, \2171 );
and \U$264 ( \2402 , RI8924ff0_179, \2173 );
and \U$265 ( \2403 , RI8930a08_166, \2175 );
and \U$266 ( \2404 , RI89399f0_153, \2177 );
and \U$267 ( \2405 , RI8946218_140, \2179 );
and \U$268 ( \2406 , RI89ec280_127, \2181 );
and \U$269 ( \2407 , RI89ec898_114, \2183 );
and \U$270 ( \2408 , RI97771d8_101, \2185 );
and \U$271 ( \2409 , RI98086d8_88, \2187 );
and \U$272 ( \2410 , RI9819370_75, \2189 );
and \U$273 ( \2411 , RI98ab878_62, \2191 );
and \U$274 ( \2412 , RI98abe90_49, \2193 );
and \U$275 ( \2413 , RI98bcb28_36, \2195 );
or \U$276 ( \2414 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 );
_DC g1bc2 ( \2415_nG1bc2 , \2414 , \2214 );
buf \U$277 ( \2416 , \2415_nG1bc2 );
not \U$278 ( \2417 , \2416 );
and \U$279 ( \2418 , \2396 , \2417 );
xor \U$280 ( \2419 , \2144 , \2145 );
buf \U$281 ( \2420 , \2419 );
buf \U$282 ( \2421 , \2420 );
and \U$283 ( \2422 , RI994d7b8_245, \2159 );
and \U$284 ( \2423 , RI995e630_232, \2165 );
and \U$285 ( \2424 , RI9967258_219, \2167 );
and \U$286 ( \2425 , RI890f768_206, \2169 );
and \U$287 ( \2426 , RI8918750_193, \2171 );
and \U$288 ( \2427 , RI8924f78_180, \2173 );
and \U$289 ( \2428 , RI8930990_167, \2175 );
and \U$290 ( \2429 , RI8939978_154, \2177 );
and \U$291 ( \2430 , RI89461a0_141, \2179 );
and \U$292 ( \2431 , RI89ec208_128, \2181 );
and \U$293 ( \2432 , RI89ec820_115, \2183 );
and \U$294 ( \2433 , RI9777160_102, \2185 );
and \U$295 ( \2434 , RI9808660_89, \2187 );
and \U$296 ( \2435 , RI98192f8_76, \2189 );
and \U$297 ( \2436 , RI98ab800_63, \2191 );
and \U$298 ( \2437 , RI98abe18_50, \2193 );
and \U$299 ( \2438 , RI98bcab0_37, \2195 );
or \U$300 ( \2439 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 );
_DC g1bdb ( \2440_nG1bdb , \2439 , \2214 );
buf \U$301 ( \2441 , \2440_nG1bdb );
not \U$302 ( \2442 , \2441 );
and \U$303 ( \2443 , \2421 , \2442 );
not \U$304 ( \2444 , \2145 );
buf \U$305 ( \2445 , \2444 );
buf \U$306 ( \2446 , \2445 );
and \U$307 ( \2447 , RI994d740_246, \2159 );
and \U$308 ( \2448 , RI995e5b8_233, \2165 );
and \U$309 ( \2449 , RI99671e0_220, \2167 );
and \U$310 ( \2450 , RI890f6f0_207, \2169 );
and \U$311 ( \2451 , RI89186d8_194, \2171 );
and \U$312 ( \2452 , RI8924f00_181, \2173 );
and \U$313 ( \2453 , RI8930918_168, \2175 );
and \U$314 ( \2454 , RI8939900_155, \2177 );
and \U$315 ( \2455 , RI8946128_142, \2179 );
and \U$316 ( \2456 , RI89ec190_129, \2181 );
and \U$317 ( \2457 , RI89ec7a8_116, \2183 );
and \U$318 ( \2458 , RI97770e8_103, \2185 );
and \U$319 ( \2459 , RI98085e8_90, \2187 );
and \U$320 ( \2460 , RI9819280_77, \2189 );
and \U$321 ( \2461 , RI98ab788_64, \2191 );
and \U$322 ( \2462 , RI98abda0_51, \2193 );
and \U$323 ( \2463 , RI98bca38_38, \2195 );
or \U$324 ( \2464 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 );
_DC g1aa5 ( \2465_nG1aa5 , \2464 , \2214 );
buf \U$325 ( \2466 , \2465_nG1aa5 );
not \U$326 ( \2467 , \2466 );
and \U$327 ( \2468 , \2446 , \2467 );
buf \U$328 ( \2469 , RI994dec0_26);
buf \U$331 ( \2470 , \2469 );
and \U$332 ( \2471 , RI994d6c8_247, \2159 );
and \U$333 ( \2472 , RI995e540_234, \2165 );
and \U$334 ( \2473 , RI9967168_221, \2167 );
and \U$335 ( \2474 , RI890f678_208, \2169 );
and \U$336 ( \2475 , RI8918660_195, \2171 );
and \U$337 ( \2476 , RI8924e88_182, \2173 );
and \U$338 ( \2477 , RI89308a0_169, \2175 );
and \U$339 ( \2478 , RI8939888_156, \2177 );
and \U$340 ( \2479 , RI89460b0_143, \2179 );
and \U$341 ( \2480 , RI89ec118_130, \2181 );
and \U$342 ( \2481 , RI89ec730_117, \2183 );
and \U$343 ( \2482 , RI9777070_104, \2185 );
and \U$344 ( \2483 , RI9808570_91, \2187 );
and \U$345 ( \2484 , RI9819208_78, \2189 );
and \U$346 ( \2485 , RI98ab710_65, \2191 );
and \U$347 ( \2486 , RI98abd28_52, \2193 );
and \U$348 ( \2487 , RI98bc9c0_39, \2195 );
or \U$349 ( \2488 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 );
_DC g1a89 ( \2489_nG1a89 , \2488 , \2214 );
buf \U$350 ( \2490 , \2489_nG1a89 );
not \U$351 ( \2491 , \2490 );
or \U$352 ( \2492 , \2470 , \2491 );
and \U$353 ( \2493 , \2467 , \2492 );
and \U$354 ( \2494 , \2446 , \2492 );
or \U$355 ( \2495 , \2468 , \2493 , \2494 );
and \U$356 ( \2496 , \2442 , \2495 );
and \U$357 ( \2497 , \2421 , \2495 );
or \U$358 ( \2498 , \2443 , \2496 , \2497 );
and \U$359 ( \2499 , \2417 , \2498 );
and \U$360 ( \2500 , \2396 , \2498 );
or \U$361 ( \2501 , \2418 , \2499 , \2500 );
and \U$362 ( \2502 , \2392 , \2501 );
and \U$363 ( \2503 , \2371 , \2501 );
or \U$364 ( \2504 , \2393 , \2502 , \2503 );
and \U$365 ( \2505 , \2367 , \2504 );
and \U$366 ( \2506 , \2346 , \2504 );
or \U$367 ( \2507 , \2368 , \2505 , \2506 );
and \U$368 ( \2508 , \2342 , \2507 );
and \U$369 ( \2509 , \2321 , \2507 );
or \U$370 ( \2510 , \2343 , \2508 , \2509 );
and \U$371 ( \2511 , \2317 , \2510 );
and \U$372 ( \2512 , \2296 , \2510 );
or \U$373 ( \2513 , \2318 , \2511 , \2512 );
and \U$374 ( \2514 , \2292 , \2513 );
and \U$375 ( \2515 , \2271 , \2513 );
or \U$376 ( \2516 , \2293 , \2514 , \2515 );
and \U$377 ( \2517 , \2267 , \2516 );
and \U$378 ( \2518 , \2246 , \2516 );
or \U$379 ( \2519 , \2268 , \2517 , \2518 );
and \U$380 ( \2520 , \2242 , \2519 );
and \U$381 ( \2521 , \2221 , \2519 );
or \U$382 ( \2522 , \2243 , \2520 , \2521 );
xor \U$383 ( \2523 , \2218 , \2522 );
buf g21a2_GF_PartitionCandidate( \2524_nG21a2 , \2523 );
buf \U$384 ( \2525 , \2524_nG21a2 );
xor \U$385 ( \2526 , \2221 , \2242 );
xor \U$386 ( \2527 , \2526 , \2519 );
buf g217e_GF_PartitionCandidate( \2528_nG217e , \2527 );
buf \U$387 ( \2529 , \2528_nG217e );
xor \U$388 ( \2530 , \2246 , \2267 );
xor \U$389 ( \2531 , \2530 , \2516 );
buf g1ff7_GF_PartitionCandidate( \2532_nG1ff7 , \2531 );
buf \U$390 ( \2533 , \2532_nG1ff7 );
and \U$391 ( \2534 , \2529 , \2533 );
not \U$392 ( \2535 , \2534 );
and \U$393 ( \2536 , \2525 , \2535 );
not \U$394 ( \2537 , \2536 );
buf \U$395 ( \2538 , RI9921730_613);
buf \U$396 ( \2539 , RI9921988_608);
buf \U$397 ( \2540 , RI9921a00_607);
buf \U$398 ( \2541 , RI9921a78_606);
buf \U$399 ( \2542 , RI9921af0_605);
buf \U$400 ( \2543 , RI9921b68_604);
buf \U$401 ( \2544 , RI9921be0_603);
buf \U$402 ( \2545 , RI9921c58_602);
buf \U$403 ( \2546 , RI9921cd0_601);
buf \U$404 ( \2547 , RI9921910_609);
nor \U$405 ( \2548 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 );
buf \U$406 ( \2549 , \2548 );
buf \U$407 ( \2550 , \2549 );
xor \U$408 ( \2551 , \2538 , \2550 );
buf \U$409 ( \2552 , \2551 );
buf \U$410 ( \2553 , RI99217a8_612);
and \U$411 ( \2554 , \2538 , \2550 );
xor \U$412 ( \2555 , \2553 , \2554 );
buf \U$413 ( \2556 , \2555 );
buf \U$414 ( \2557 , RI9921820_611);
and \U$415 ( \2558 , \2553 , \2554 );
xor \U$416 ( \2559 , \2557 , \2558 );
buf \U$417 ( \2560 , \2559 );
buf \U$418 ( \2561 , RI9921898_610);
and \U$419 ( \2562 , \2557 , \2558 );
xor \U$420 ( \2563 , \2561 , \2562 );
buf \U$421 ( \2564 , \2563 );
buf \U$422 ( \2565 , RI9921910_609);
and \U$423 ( \2566 , \2561 , \2562 );
xor \U$424 ( \2567 , \2565 , \2566 );
buf \U$425 ( \2568 , \2567 );
not \U$426 ( \2569 , \2568 );
buf \U$427 ( \2570 , RI9921988_608);
and \U$428 ( \2571 , \2565 , \2566 );
xor \U$429 ( \2572 , \2570 , \2571 );
buf \U$430 ( \2573 , \2572 );
buf \U$431 ( \2574 , RI9921a00_607);
and \U$432 ( \2575 , \2570 , \2571 );
xor \U$433 ( \2576 , \2574 , \2575 );
buf \U$434 ( \2577 , \2576 );
buf \U$435 ( \2578 , RI9921a78_606);
and \U$436 ( \2579 , \2574 , \2575 );
xor \U$437 ( \2580 , \2578 , \2579 );
buf \U$438 ( \2581 , \2580 );
buf \U$439 ( \2582 , RI9921af0_605);
and \U$440 ( \2583 , \2578 , \2579 );
xor \U$441 ( \2584 , \2582 , \2583 );
buf \U$442 ( \2585 , \2584 );
buf \U$443 ( \2586 , RI9921b68_604);
and \U$444 ( \2587 , \2582 , \2583 );
xor \U$445 ( \2588 , \2586 , \2587 );
buf \U$446 ( \2589 , \2588 );
buf \U$447 ( \2590 , RI9921be0_603);
and \U$448 ( \2591 , \2586 , \2587 );
xor \U$449 ( \2592 , \2590 , \2591 );
buf \U$450 ( \2593 , \2592 );
buf \U$451 ( \2594 , RI9921c58_602);
and \U$452 ( \2595 , \2590 , \2591 );
xor \U$453 ( \2596 , \2594 , \2595 );
buf \U$454 ( \2597 , \2596 );
buf \U$455 ( \2598 , RI9921cd0_601);
and \U$456 ( \2599 , \2594 , \2595 );
xor \U$457 ( \2600 , \2598 , \2599 );
buf \U$458 ( \2601 , \2600 );
nor \U$459 ( \2602 , \2552 , \2556 , \2560 , \2564 , \2569 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$460 ( \2603 , RI9922bd0_569, \2602 );
not \U$461 ( \2604 , \2552 );
not \U$462 ( \2605 , \2556 );
not \U$463 ( \2606 , \2560 );
not \U$464 ( \2607 , \2564 );
nor \U$465 ( \2608 , \2604 , \2605 , \2606 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$466 ( \2609 , RI9923800_549, \2608 );
nor \U$467 ( \2610 , \2552 , \2605 , \2606 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$468 ( \2611 , RI9924160_529, \2610 );
nor \U$469 ( \2612 , \2604 , \2556 , \2606 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$470 ( \2613 , RI9924ac0_509, \2612 );
nor \U$471 ( \2614 , \2552 , \2556 , \2606 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$472 ( \2615 , RI9925ab0_489, \2614 );
nor \U$473 ( \2616 , \2604 , \2605 , \2560 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$474 ( \2617 , RI9926410_469, \2616 );
nor \U$475 ( \2618 , \2552 , \2605 , \2560 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$476 ( \2619 , RI9926d70_449, \2618 );
nor \U$477 ( \2620 , \2604 , \2556 , \2560 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$478 ( \2621 , RI9928120_429, \2620 );
nor \U$479 ( \2622 , \2552 , \2556 , \2560 , \2607 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$480 ( \2623 , RI9928a80_409, \2622 );
nor \U$481 ( \2624 , \2604 , \2605 , \2606 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$482 ( \2625 , RI992a1f0_389, \2624 );
nor \U$483 ( \2626 , \2552 , \2605 , \2606 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$484 ( \2627 , RI992ab50_369, \2626 );
nor \U$485 ( \2628 , \2604 , \2556 , \2606 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$486 ( \2629 , RI992b4b0_349, \2628 );
nor \U$487 ( \2630 , \2552 , \2556 , \2606 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$488 ( \2631 , RI992cfe0_329, \2630 );
nor \U$489 ( \2632 , \2604 , \2605 , \2560 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$490 ( \2633 , RI992eed0_309, \2632 );
nor \U$491 ( \2634 , \2552 , \2605 , \2560 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$492 ( \2635 , RI992f830_289, \2634 );
nor \U$493 ( \2636 , \2604 , \2556 , \2560 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$494 ( \2637 , RI9931ae0_269, \2636 );
nor \U$495 ( \2638 , \2552 , \2556 , \2560 , \2564 , \2568 , \2573 , \2577 , \2581 , \2585 , \2589 , \2593 , \2597 , \2601 );
and \U$496 ( \2639 , RI994d5d8_249, \2638 );
or \U$497 ( \2640 , \2603 , \2609 , \2611 , \2613 , \2615 , \2617 , \2619 , \2621 , \2623 , \2625 , \2627 , \2629 , \2631 , \2633 , \2635 , \2637 , \2639 );
buf \U$498 ( \2641 , \2573 );
buf \U$499 ( \2642 , \2577 );
buf \U$500 ( \2643 , \2581 );
buf \U$501 ( \2644 , \2585 );
buf \U$502 ( \2645 , \2589 );
buf \U$503 ( \2646 , \2593 );
buf \U$504 ( \2647 , \2597 );
buf \U$505 ( \2648 , \2601 );
buf \U$506 ( \2649 , \2568 );
buf \U$507 ( \2650 , \2552 );
buf \U$508 ( \2651 , \2556 );
buf \U$509 ( \2652 , \2560 );
buf \U$510 ( \2653 , \2564 );
or \U$511 ( \2654 , \2650 , \2651 , \2652 , \2653 );
and \U$512 ( \2655 , \2649 , \2654 );
or \U$513 ( \2656 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2655 );
buf \U$514 ( \2657 , \2656 );
_DC g2899 ( \2658_nG2899 , \2640 , \2657 );
buf \U$515 ( \2659 , \2658_nG2899 );
buf \U$516 ( \2660 , RI994e460_14);
and \U$517 ( \2661 , \2135 , \2154 );
and \U$518 ( \2662 , \2660 , \2661 );
buf \U$519 ( \2663 , \2662 );
buf \U$520 ( \2664 , \2663 );
xor \U$521 ( \2665 , \2660 , \2661 );
buf \U$522 ( \2666 , \2665 );
buf \U$523 ( \2667 , \2666 );
and \U$524 ( \2668 , RI995e4c8_235, \2159 );
and \U$525 ( \2669 , RI99670f0_222, \2165 );
and \U$526 ( \2670 , RI890f600_209, \2167 );
and \U$527 ( \2671 , RI89185e8_196, \2169 );
and \U$528 ( \2672 , RI8924e10_183, \2171 );
and \U$529 ( \2673 , RI8930828_170, \2173 );
and \U$530 ( \2674 , RI8939810_157, \2175 );
and \U$531 ( \2675 , RI8946038_144, \2177 );
and \U$532 ( \2676 , RI89ec0a0_131, \2179 );
and \U$533 ( \2677 , RI89ec6b8_118, \2181 );
and \U$534 ( \2678 , RI9776ff8_105, \2183 );
and \U$535 ( \2679 , RI98084f8_92, \2185 );
and \U$536 ( \2680 , RI9808b10_79, \2187 );
and \U$537 ( \2681 , RI98197a8_66, \2189 );
and \U$538 ( \2682 , RI98abcb0_53, \2191 );
and \U$539 ( \2683 , RI98bc948_40, \2193 );
and \U$540 ( \2684 , RI994de48_27, \2195 );
or \U$541 ( \2685 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 );
_DC g2361 ( \2686_nG2361 , \2685 , \2214 );
buf \U$542 ( \2687 , \2686_nG2361 );
not \U$543 ( \2688 , \2687 );
and \U$544 ( \2689 , \2667 , \2688 );
and \U$545 ( \2690 , \2157 , \2217 );
and \U$546 ( \2691 , \2217 , \2522 );
and \U$547 ( \2692 , \2157 , \2522 );
or \U$548 ( \2693 , \2690 , \2691 , \2692 );
and \U$549 ( \2694 , \2688 , \2693 );
and \U$550 ( \2695 , \2667 , \2693 );
or \U$551 ( \2696 , \2689 , \2694 , \2695 );
xnor \U$552 ( \2697 , \2664 , \2696 );
buf g2376_GF_PartitionCandidate( \2698_nG2376 , \2697 );
buf \U$553 ( \2699 , \2698_nG2376 );
xor \U$554 ( \2700 , \2667 , \2688 );
xor \U$555 ( \2701 , \2700 , \2693 );
buf g236a_GF_PartitionCandidate( \2702_nG236a , \2701 );
buf \U$556 ( \2703 , \2702_nG236a );
xor \U$557 ( \2704 , \2699 , \2703 );
xor \U$558 ( \2705 , \2703 , \2525 );
not \U$559 ( \2706 , \2705 );
and \U$560 ( \2707 , \2704 , \2706 );
and \U$561 ( \2708 , \2659 , \2707 );
and \U$562 ( \2709 , RI9922f18_568, \2602 );
and \U$563 ( \2710 , RI9923878_548, \2608 );
and \U$564 ( \2711 , RI99241d8_528, \2610 );
and \U$565 ( \2712 , RI9924b38_508, \2612 );
and \U$566 ( \2713 , RI9925b28_488, \2614 );
and \U$567 ( \2714 , RI9926488_468, \2616 );
and \U$568 ( \2715 , RI9926de8_448, \2618 );
and \U$569 ( \2716 , RI9928198_428, \2620 );
and \U$570 ( \2717 , RI9928af8_408, \2622 );
and \U$571 ( \2718 , RI992a268_388, \2624 );
and \U$572 ( \2719 , RI992abc8_368, \2626 );
and \U$573 ( \2720 , RI992c6f8_348, \2628 );
and \U$574 ( \2721 , RI992d058_328, \2630 );
and \U$575 ( \2722 , RI992ef48_308, \2632 );
and \U$576 ( \2723 , RI992f8a8_288, \2634 );
and \U$577 ( \2724 , RI9931b58_268, \2636 );
and \U$578 ( \2725 , RI994d650_248, \2638 );
or \U$579 ( \2726 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 );
_DC g298d ( \2727_nG298d , \2726 , \2657 );
buf \U$580 ( \2728 , \2727_nG298d );
and \U$581 ( \2729 , \2728 , \2705 );
nor \U$582 ( \2730 , \2708 , \2729 );
and \U$583 ( \2731 , \2703 , \2525 );
not \U$584 ( \2732 , \2731 );
and \U$585 ( \2733 , \2699 , \2732 );
xnor \U$586 ( \2734 , \2730 , \2733 );
xor \U$587 ( \2735 , \2537 , \2734 );
and \U$589 ( \2736 , RI9922b58_570, \2602 );
and \U$590 ( \2737 , RI9923788_550, \2608 );
and \U$591 ( \2738 , RI99240e8_530, \2610 );
and \U$592 ( \2739 , RI9924a48_510, \2612 );
and \U$593 ( \2740 , RI9925a38_490, \2614 );
and \U$594 ( \2741 , RI9926398_470, \2616 );
and \U$595 ( \2742 , RI9926cf8_450, \2618 );
and \U$596 ( \2743 , RI99280a8_430, \2620 );
and \U$597 ( \2744 , RI9928a08_410, \2622 );
and \U$598 ( \2745 , RI992a178_390, \2624 );
and \U$599 ( \2746 , RI992aad8_370, \2626 );
and \U$600 ( \2747 , RI992b438_350, \2628 );
and \U$601 ( \2748 , RI992cf68_330, \2630 );
and \U$602 ( \2749 , RI992ee58_310, \2632 );
and \U$603 ( \2750 , RI992f7b8_290, \2634 );
and \U$604 ( \2751 , RI9931a68_270, \2636 );
and \U$605 ( \2752 , RI994d560_250, \2638 );
or \U$606 ( \2753 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 );
_DC g27d7 ( \2754_nG27d7 , \2753 , \2657 );
buf \U$607 ( \2755 , \2754_nG27d7 );
or \U$608 ( \2756 , \2664 , \2696 );
not \U$609 ( \2757 , \2756 );
buf g2572_GF_PartitionCandidate( \2758_nG2572 , \2757 );
buf \U$610 ( \2759 , \2758_nG2572 );
xor \U$611 ( \2760 , \2759 , \2699 );
and \U$612 ( \2761 , \2755 , \2760 );
nor \U$613 ( \2762 , 1'b0 , \2761 );
xnor \U$615 ( \2763 , \2762 , 1'b0 );
xor \U$616 ( \2764 , \2735 , \2763 );
xor \U$617 ( \2765 , 1'b0 , \2764 );
xor \U$619 ( \2766 , \2525 , \2529 );
xor \U$620 ( \2767 , \2529 , \2533 );
not \U$621 ( \2768 , \2767 );
and \U$622 ( \2769 , \2766 , \2768 );
and \U$623 ( \2770 , \2728 , \2769 );
not \U$624 ( \2771 , \2770 );
xnor \U$625 ( \2772 , \2771 , \2536 );
and \U$626 ( \2773 , \2755 , \2707 );
and \U$627 ( \2774 , \2659 , \2705 );
nor \U$628 ( \2775 , \2773 , \2774 );
xnor \U$629 ( \2776 , \2775 , \2733 );
and \U$630 ( \2777 , \2772 , \2776 );
or \U$632 ( \2778 , 1'b0 , \2777 , 1'b0 );
xor \U$634 ( \2779 , \2778 , 1'b0 );
xor \U$636 ( \2780 , \2779 , 1'b0 );
and \U$637 ( \2781 , \2765 , \2780 );
or \U$638 ( \2782 , 1'b0 , 1'b0 , \2781 );
and \U$641 ( \2783 , \2728 , \2707 );
not \U$642 ( \2784 , \2783 );
xnor \U$643 ( \2785 , \2784 , \2733 );
xor \U$644 ( \2786 , 1'b0 , \2785 );
and \U$646 ( \2787 , \2659 , \2760 );
nor \U$647 ( \2788 , 1'b0 , \2787 );
xnor \U$648 ( \2789 , \2788 , 1'b0 );
xor \U$649 ( \2790 , \2786 , \2789 );
xor \U$650 ( \2791 , 1'b0 , \2790 );
xor \U$652 ( \2792 , \2791 , 1'b1 );
and \U$653 ( \2793 , \2537 , \2734 );
and \U$654 ( \2794 , \2734 , \2763 );
and \U$655 ( \2795 , \2537 , \2763 );
or \U$656 ( \2796 , \2793 , \2794 , \2795 );
xor \U$658 ( \2797 , \2796 , 1'b0 );
xor \U$660 ( \2798 , \2797 , 1'b0 );
xor \U$661 ( \2799 , \2792 , \2798 );
and \U$662 ( \2800 , \2782 , \2799 );
or \U$664 ( \2801 , 1'b0 , \2800 , 1'b0 );
xor \U$666 ( \2802 , \2801 , 1'b0 );
and \U$668 ( \2803 , \2791 , 1'b1 );
and \U$669 ( \2804 , 1'b1 , \2798 );
and \U$670 ( \2805 , \2791 , \2798 );
or \U$671 ( \2806 , \2803 , \2804 , \2805 );
xor \U$672 ( \2807 , 1'b0 , \2806 );
not \U$674 ( \2808 , \2733 );
and \U$676 ( \2809 , \2728 , \2760 );
nor \U$677 ( \2810 , 1'b0 , \2809 );
xnor \U$678 ( \2811 , \2810 , 1'b0 );
xor \U$679 ( \2812 , \2808 , \2811 );
xor \U$681 ( \2813 , \2812 , 1'b0 );
xor \U$682 ( \2814 , 1'b0 , \2813 );
xor \U$684 ( \2815 , \2814 , 1'b0 );
and \U$686 ( \2816 , \2785 , \2789 );
or \U$688 ( \2817 , 1'b0 , \2816 , 1'b0 );
xor \U$690 ( \2818 , \2817 , 1'b0 );
xor \U$692 ( \2819 , \2818 , 1'b0 );
xor \U$693 ( \2820 , \2815 , \2819 );
xor \U$694 ( \2821 , \2807 , \2820 );
xor \U$695 ( \2822 , \2802 , \2821 );
xor \U$701 ( \2823 , \2271 , \2292 );
xor \U$702 ( \2824 , \2823 , \2513 );
buf g1fd3_GF_PartitionCandidate( \2825_nG1fd3 , \2824 );
buf \U$703 ( \2826 , \2825_nG1fd3 );
xor \U$704 ( \2827 , \2533 , \2826 );
xor \U$705 ( \2828 , \2296 , \2317 );
xor \U$706 ( \2829 , \2828 , \2510 );
buf g1e5e_GF_PartitionCandidate( \2830_nG1e5e , \2829 );
buf \U$707 ( \2831 , \2830_nG1e5e );
xor \U$708 ( \2832 , \2826 , \2831 );
not \U$709 ( \2833 , \2832 );
and \U$710 ( \2834 , \2827 , \2833 );
and \U$711 ( \2835 , \2728 , \2834 );
not \U$712 ( \2836 , \2835 );
and \U$713 ( \2837 , \2826 , \2831 );
not \U$714 ( \2838 , \2837 );
and \U$715 ( \2839 , \2533 , \2838 );
xnor \U$716 ( \2840 , \2836 , \2839 );
and \U$717 ( \2841 , \2755 , \2769 );
and \U$718 ( \2842 , \2659 , \2767 );
nor \U$719 ( \2843 , \2841 , \2842 );
xnor \U$720 ( \2844 , \2843 , \2536 );
and \U$721 ( \2845 , \2840 , \2844 );
or \U$723 ( \2846 , 1'b0 , \2845 , 1'b0 );
and \U$724 ( \2847 , RI9922a68_572, \2602 );
and \U$725 ( \2848 , RI9923698_552, \2608 );
and \U$726 ( \2849 , RI9923ff8_532, \2610 );
and \U$727 ( \2850 , RI9924958_512, \2612 );
and \U$728 ( \2851 , RI9925948_492, \2614 );
and \U$729 ( \2852 , RI99262a8_472, \2616 );
and \U$730 ( \2853 , RI9926c08_452, \2618 );
and \U$731 ( \2854 , RI9927fb8_432, \2620 );
and \U$732 ( \2855 , RI9928918_412, \2622 );
and \U$733 ( \2856 , RI9929278_392, \2624 );
and \U$734 ( \2857 , RI992a9e8_372, \2626 );
and \U$735 ( \2858 , RI992b348_352, \2628 );
and \U$736 ( \2859 , RI992ce78_332, \2630 );
and \U$737 ( \2860 , RI992ed68_312, \2632 );
and \U$738 ( \2861 , RI992f6c8_292, \2634 );
and \U$739 ( \2862 , RI9931978_272, \2636 );
and \U$740 ( \2863 , RI994d470_252, \2638 );
or \U$741 ( \2864 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 );
_DC g263c ( \2865_nG263c , \2864 , \2657 );
buf \U$742 ( \2866 , \2865_nG263c );
and \U$743 ( \2867 , \2866 , \2707 );
and \U$744 ( \2868 , RI9922ae0_571, \2602 );
and \U$745 ( \2869 , RI9923710_551, \2608 );
and \U$746 ( \2870 , RI9924070_531, \2610 );
and \U$747 ( \2871 , RI99249d0_511, \2612 );
and \U$748 ( \2872 , RI99259c0_491, \2614 );
and \U$749 ( \2873 , RI9926320_471, \2616 );
and \U$750 ( \2874 , RI9926c80_451, \2618 );
and \U$751 ( \2875 , RI9928030_431, \2620 );
and \U$752 ( \2876 , RI9928990_411, \2622 );
and \U$753 ( \2877 , RI992a100_391, \2624 );
and \U$754 ( \2878 , RI992aa60_371, \2626 );
and \U$755 ( \2879 , RI992b3c0_351, \2628 );
and \U$756 ( \2880 , RI992cef0_331, \2630 );
and \U$757 ( \2881 , RI992ede0_311, \2632 );
and \U$758 ( \2882 , RI992f740_291, \2634 );
and \U$759 ( \2883 , RI99319f0_271, \2636 );
and \U$760 ( \2884 , RI994d4e8_251, \2638 );
or \U$761 ( \2885 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 );
_DC g2716 ( \2886_nG2716 , \2885 , \2657 );
buf \U$762 ( \2887 , \2886_nG2716 );
and \U$763 ( \2888 , \2887 , \2705 );
nor \U$764 ( \2889 , \2867 , \2888 );
xnor \U$765 ( \2890 , \2889 , \2733 );
and \U$767 ( \2891 , RI99229f0_573, \2602 );
and \U$768 ( \2892 , RI9923620_553, \2608 );
and \U$769 ( \2893 , RI9923f80_533, \2610 );
and \U$770 ( \2894 , RI99248e0_513, \2612 );
and \U$771 ( \2895 , RI99258d0_493, \2614 );
and \U$772 ( \2896 , RI9926230_473, \2616 );
and \U$773 ( \2897 , RI9926b90_453, \2618 );
and \U$774 ( \2898 , RI9927f40_433, \2620 );
and \U$775 ( \2899 , RI99288a0_413, \2622 );
and \U$776 ( \2900 , RI9929200_393, \2624 );
and \U$777 ( \2901 , RI992a970_373, \2626 );
and \U$778 ( \2902 , RI992b2d0_353, \2628 );
and \U$779 ( \2903 , RI992ce00_333, \2630 );
and \U$780 ( \2904 , RI992ecf0_313, \2632 );
and \U$781 ( \2905 , RI992f650_293, \2634 );
and \U$782 ( \2906 , RI9931900_273, \2636 );
and \U$783 ( \2907 , RI994d3f8_253, \2638 );
or \U$784 ( \2908 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 );
_DC g2551 ( \2909_nG2551 , \2908 , \2657 );
buf \U$785 ( \2910 , \2909_nG2551 );
and \U$786 ( \2911 , \2910 , \2760 );
nor \U$787 ( \2912 , 1'b0 , \2911 );
xnor \U$788 ( \2913 , \2912 , 1'b0 );
and \U$789 ( \2914 , \2890 , \2913 );
or \U$792 ( \2915 , \2914 , 1'b0 , 1'b0 );
and \U$793 ( \2916 , \2846 , \2915 );
or \U$796 ( \2917 , \2916 , 1'b0 , 1'b0 );
and \U$799 ( \2918 , \2866 , \2760 );
nor \U$800 ( \2919 , 1'b0 , \2918 );
xnor \U$801 ( \2920 , \2919 , 1'b0 );
xor \U$803 ( \2921 , \2920 , 1'b0 );
xor \U$805 ( \2922 , \2921 , 1'b0 );
not \U$806 ( \2923 , \2839 );
and \U$807 ( \2924 , \2659 , \2769 );
and \U$808 ( \2925 , \2728 , \2767 );
nor \U$809 ( \2926 , \2924 , \2925 );
xnor \U$810 ( \2927 , \2926 , \2536 );
xor \U$811 ( \2928 , \2923 , \2927 );
and \U$812 ( \2929 , \2887 , \2707 );
and \U$813 ( \2930 , \2755 , \2705 );
nor \U$814 ( \2931 , \2929 , \2930 );
xnor \U$815 ( \2932 , \2931 , \2733 );
xor \U$816 ( \2933 , \2928 , \2932 );
and \U$817 ( \2934 , \2922 , \2933 );
or \U$819 ( \2935 , 1'b0 , \2934 , 1'b0 );
and \U$820 ( \2936 , \2917 , \2935 );
or \U$821 ( \2937 , 1'b0 , 1'b0 , \2936 );
and \U$823 ( \2938 , \2887 , \2760 );
nor \U$824 ( \2939 , 1'b0 , \2938 );
xnor \U$825 ( \2940 , \2939 , 1'b0 );
xor \U$827 ( \2941 , \2940 , 1'b0 );
xor \U$829 ( \2942 , \2941 , 1'b0 );
xor \U$831 ( \2943 , 1'b0 , \2772 );
xor \U$832 ( \2944 , \2943 , \2776 );
xor \U$833 ( \2945 , \2942 , \2944 );
and \U$835 ( \2946 , \2945 , 1'b1 );
and \U$836 ( \2947 , \2923 , \2927 );
and \U$837 ( \2948 , \2927 , \2932 );
and \U$838 ( \2949 , \2923 , \2932 );
or \U$839 ( \2950 , \2947 , \2948 , \2949 );
xor \U$841 ( \2951 , \2950 , 1'b0 );
xor \U$843 ( \2952 , \2951 , 1'b0 );
and \U$844 ( \2953 , 1'b1 , \2952 );
and \U$845 ( \2954 , \2945 , \2952 );
or \U$846 ( \2955 , \2946 , \2953 , \2954 );
and \U$847 ( \2956 , \2937 , \2955 );
xor \U$849 ( \2957 , \2765 , 1'b0 );
xor \U$850 ( \2958 , \2957 , \2780 );
and \U$851 ( \2959 , \2955 , \2958 );
and \U$852 ( \2960 , \2937 , \2958 );
or \U$853 ( \2961 , \2956 , \2959 , \2960 );
xor \U$855 ( \2962 , 1'b0 , \2782 );
xor \U$856 ( \2963 , \2962 , \2799 );
and \U$857 ( \2964 , \2961 , \2963 );
or \U$858 ( \2965 , 1'b0 , 1'b0 , \2964 );
nand \U$859 ( \2966 , \2822 , \2965 );
nor \U$860 ( \2967 , \2822 , \2965 );
not \U$861 ( \2968 , \2967 );
nand \U$862 ( \2969 , \2966 , \2968 );
xor \U$863 ( \2970 , \2446 , \2467 );
xor \U$864 ( \2971 , \2970 , \2492 );
buf g1aac_GF_PartitionCandidate( \2972_nG1aac , \2971 );
buf \U$865 ( \2973 , \2972_nG1aac );
xor \U$866 ( \2974 , \2470 , \2490 );
buf g1a8c_GF_PartitionCandidate( \2975_nG1a8c , \2974 );
buf \U$867 ( \2976 , \2975_nG1a8c );
xor \U$868 ( \2977 , \2973 , \2976 );
not \U$869 ( \2978 , \2976 );
and \U$870 ( \2979 , \2977 , \2978 );
and \U$871 ( \2980 , \2910 , \2979 );
and \U$872 ( \2981 , \2866 , \2976 );
nor \U$873 ( \2982 , \2980 , \2981 );
xnor \U$874 ( \2983 , \2982 , \2973 );
and \U$875 ( \2984 , RI9922900_575, \2602 );
and \U$876 ( \2985 , RI9923530_555, \2608 );
and \U$877 ( \2986 , RI9923e90_535, \2610 );
and \U$878 ( \2987 , RI99247f0_515, \2612 );
and \U$879 ( \2988 , RI99257e0_495, \2614 );
and \U$880 ( \2989 , RI9926140_475, \2616 );
and \U$881 ( \2990 , RI9926aa0_455, \2618 );
and \U$882 ( \2991 , RI9927e50_435, \2620 );
and \U$883 ( \2992 , RI99287b0_415, \2622 );
and \U$884 ( \2993 , RI9929110_395, \2624 );
and \U$885 ( \2994 , RI992a880_375, \2626 );
and \U$886 ( \2995 , RI992b1e0_355, \2628 );
and \U$887 ( \2996 , RI992cd10_335, \2630 );
and \U$888 ( \2997 , RI992d670_315, \2632 );
and \U$889 ( \2998 , RI992f560_295, \2634 );
and \U$890 ( \2999 , RI9931810_275, \2636 );
and \U$891 ( \3000 , RI9935f50_255, \2638 );
or \U$892 ( \3001 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 );
_DC g239e ( \3002_nG239e , \3001 , \2657 );
buf \U$893 ( \3003 , \3002_nG239e );
xor \U$894 ( \3004 , \2396 , \2417 );
xor \U$895 ( \3005 , \3004 , \2498 );
buf g1be7_GF_PartitionCandidate( \3006_nG1be7 , \3005 );
buf \U$896 ( \3007 , \3006_nG1be7 );
xor \U$897 ( \3008 , \2421 , \2442 );
xor \U$898 ( \3009 , \3008 , \2495 );
buf g1beb_GF_PartitionCandidate( \3010_nG1beb , \3009 );
buf \U$899 ( \3011 , \3010_nG1beb );
xor \U$900 ( \3012 , \3007 , \3011 );
xor \U$901 ( \3013 , \3011 , \2973 );
not \U$902 ( \3014 , \3013 );
and \U$903 ( \3015 , \3012 , \3014 );
and \U$904 ( \3016 , \3003 , \3015 );
and \U$905 ( \3017 , RI9922978_574, \2602 );
and \U$906 ( \3018 , RI99235a8_554, \2608 );
and \U$907 ( \3019 , RI9923f08_534, \2610 );
and \U$908 ( \3020 , RI9924868_514, \2612 );
and \U$909 ( \3021 , RI9925858_494, \2614 );
and \U$910 ( \3022 , RI99261b8_474, \2616 );
and \U$911 ( \3023 , RI9926b18_454, \2618 );
and \U$912 ( \3024 , RI9927ec8_434, \2620 );
and \U$913 ( \3025 , RI9928828_414, \2622 );
and \U$914 ( \3026 , RI9929188_394, \2624 );
and \U$915 ( \3027 , RI992a8f8_374, \2626 );
and \U$916 ( \3028 , RI992b258_354, \2628 );
and \U$917 ( \3029 , RI992cd88_334, \2630 );
and \U$918 ( \3030 , RI992d6e8_314, \2632 );
and \U$919 ( \3031 , RI992f5d8_294, \2634 );
and \U$920 ( \3032 , RI9931888_274, \2636 );
and \U$921 ( \3033 , RI9935fc8_254, \2638 );
or \U$922 ( \3034 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 );
_DC g2472 ( \3035_nG2472 , \3034 , \2657 );
buf \U$923 ( \3036 , \3035_nG2472 );
and \U$924 ( \3037 , \3036 , \3013 );
nor \U$925 ( \3038 , \3016 , \3037 );
and \U$926 ( \3039 , \3011 , \2973 );
not \U$927 ( \3040 , \3039 );
and \U$928 ( \3041 , \3007 , \3040 );
xnor \U$929 ( \3042 , \3038 , \3041 );
and \U$930 ( \3043 , \2983 , \3042 );
and \U$931 ( \3044 , RI9922810_577, \2602 );
and \U$932 ( \3045 , RI9923440_557, \2608 );
and \U$933 ( \3046 , RI9923da0_537, \2610 );
and \U$934 ( \3047 , RI9924700_517, \2612 );
and \U$935 ( \3048 , RI99256f0_497, \2614 );
and \U$936 ( \3049 , RI9926050_477, \2616 );
and \U$937 ( \3050 , RI99269b0_457, \2618 );
and \U$938 ( \3051 , RI9927d60_437, \2620 );
and \U$939 ( \3052 , RI99286c0_417, \2622 );
and \U$940 ( \3053 , RI9929020_397, \2624 );
and \U$941 ( \3054 , RI992a790_377, \2626 );
and \U$942 ( \3055 , RI992b0f0_357, \2628 );
and \U$943 ( \3056 , RI992cc20_337, \2630 );
and \U$944 ( \3057 , RI992d580_317, \2632 );
and \U$945 ( \3058 , RI992f470_297, \2634 );
and \U$946 ( \3059 , RI9931720_277, \2636 );
and \U$947 ( \3060 , RI9933d90_257, \2638 );
or \U$948 ( \3061 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 );
_DC g21d1 ( \3062_nG21d1 , \3061 , \2657 );
buf \U$949 ( \3063 , \3062_nG21d1 );
xor \U$950 ( \3064 , \2346 , \2367 );
xor \U$951 ( \3065 , \3064 , \2504 );
buf g1cfc_GF_PartitionCandidate( \3066_nG1cfc , \3065 );
buf \U$952 ( \3067 , \3066_nG1cfc );
xor \U$953 ( \3068 , \2371 , \2392 );
xor \U$954 ( \3069 , \3068 , \2501 );
buf g1cd8_GF_PartitionCandidate( \3070_nG1cd8 , \3069 );
buf \U$955 ( \3071 , \3070_nG1cd8 );
xor \U$956 ( \3072 , \3067 , \3071 );
xor \U$957 ( \3073 , \3071 , \3007 );
not \U$958 ( \3074 , \3073 );
and \U$959 ( \3075 , \3072 , \3074 );
and \U$960 ( \3076 , \3063 , \3075 );
and \U$961 ( \3077 , RI9922888_576, \2602 );
and \U$962 ( \3078 , RI99234b8_556, \2608 );
and \U$963 ( \3079 , RI9923e18_536, \2610 );
and \U$964 ( \3080 , RI9924778_516, \2612 );
and \U$965 ( \3081 , RI9925768_496, \2614 );
and \U$966 ( \3082 , RI99260c8_476, \2616 );
and \U$967 ( \3083 , RI9926a28_456, \2618 );
and \U$968 ( \3084 , RI9927dd8_436, \2620 );
and \U$969 ( \3085 , RI9928738_416, \2622 );
and \U$970 ( \3086 , RI9929098_396, \2624 );
and \U$971 ( \3087 , RI992a808_376, \2626 );
and \U$972 ( \3088 , RI992b168_356, \2628 );
and \U$973 ( \3089 , RI992cc98_336, \2630 );
and \U$974 ( \3090 , RI992d5f8_316, \2632 );
and \U$975 ( \3091 , RI992f4e8_296, \2634 );
and \U$976 ( \3092 , RI9931798_276, \2636 );
and \U$977 ( \3093 , RI9935ed8_256, \2638 );
or \U$978 ( \3094 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 );
_DC g22a8 ( \3095_nG22a8 , \3094 , \2657 );
buf \U$979 ( \3096 , \3095_nG22a8 );
and \U$980 ( \3097 , \3096 , \3073 );
nor \U$981 ( \3098 , \3076 , \3097 );
and \U$982 ( \3099 , \3071 , \3007 );
not \U$983 ( \3100 , \3099 );
and \U$984 ( \3101 , \3067 , \3100 );
xnor \U$985 ( \3102 , \3098 , \3101 );
and \U$986 ( \3103 , \3042 , \3102 );
and \U$987 ( \3104 , \2983 , \3102 );
or \U$988 ( \3105 , \3043 , \3103 , \3104 );
and \U$989 ( \3106 , RI9922720_579, \2602 );
and \U$990 ( \3107 , RI9923350_559, \2608 );
and \U$991 ( \3108 , RI9923cb0_539, \2610 );
and \U$992 ( \3109 , RI9924610_519, \2612 );
and \U$993 ( \3110 , RI9925600_499, \2614 );
and \U$994 ( \3111 , RI9925f60_479, \2616 );
and \U$995 ( \3112 , RI99268c0_459, \2618 );
and \U$996 ( \3113 , RI9927c70_439, \2620 );
and \U$997 ( \3114 , RI99285d0_419, \2622 );
and \U$998 ( \3115 , RI9928f30_399, \2624 );
and \U$999 ( \3116 , RI992a6a0_379, \2626 );
and \U$1000 ( \3117 , RI992b000_359, \2628 );
and \U$1001 ( \3118 , RI992cb30_339, \2630 );
and \U$1002 ( \3119 , RI992d490_319, \2632 );
and \U$1003 ( \3120 , RI992f380_299, \2634 );
and \U$1004 ( \3121 , RI9931630_279, \2636 );
and \U$1005 ( \3122 , RI9933ca0_259, \2638 );
or \U$1006 ( \3123 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 );
_DC g2012 ( \3124_nG2012 , \3123 , \2657 );
buf \U$1007 ( \3125 , \3124_nG2012 );
xor \U$1008 ( \3126 , \2321 , \2342 );
xor \U$1009 ( \3127 , \3126 , \2507 );
buf g1e3a_GF_PartitionCandidate( \3128_nG1e3a , \3127 );
buf \U$1010 ( \3129 , \3128_nG1e3a );
xor \U$1011 ( \3130 , \2831 , \3129 );
xor \U$1012 ( \3131 , \3129 , \3067 );
not \U$1013 ( \3132 , \3131 );
and \U$1014 ( \3133 , \3130 , \3132 );
and \U$1015 ( \3134 , \3125 , \3133 );
and \U$1016 ( \3135 , RI9922798_578, \2602 );
and \U$1017 ( \3136 , RI99233c8_558, \2608 );
and \U$1018 ( \3137 , RI9923d28_538, \2610 );
and \U$1019 ( \3138 , RI9924688_518, \2612 );
and \U$1020 ( \3139 , RI9925678_498, \2614 );
and \U$1021 ( \3140 , RI9925fd8_478, \2616 );
and \U$1022 ( \3141 , RI9926938_458, \2618 );
and \U$1023 ( \3142 , RI9927ce8_438, \2620 );
and \U$1024 ( \3143 , RI9928648_418, \2622 );
and \U$1025 ( \3144 , RI9928fa8_398, \2624 );
and \U$1026 ( \3145 , RI992a718_378, \2626 );
and \U$1027 ( \3146 , RI992b078_358, \2628 );
and \U$1028 ( \3147 , RI992cba8_338, \2630 );
and \U$1029 ( \3148 , RI992d508_318, \2632 );
and \U$1030 ( \3149 , RI992f3f8_298, \2634 );
and \U$1031 ( \3150 , RI99316a8_278, \2636 );
and \U$1032 ( \3151 , RI9933d18_258, \2638 );
or \U$1033 ( \3152 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 );
_DC g20db ( \3153_nG20db , \3152 , \2657 );
buf \U$1034 ( \3154 , \3153_nG20db );
and \U$1035 ( \3155 , \3154 , \3131 );
nor \U$1036 ( \3156 , \3134 , \3155 );
and \U$1037 ( \3157 , \3129 , \3067 );
not \U$1038 ( \3158 , \3157 );
and \U$1039 ( \3159 , \2831 , \3158 );
xnor \U$1040 ( \3160 , \3156 , \3159 );
and \U$1041 ( \3161 , RI9922630_581, \2602 );
and \U$1042 ( \3162 , RI9923260_561, \2608 );
and \U$1043 ( \3163 , RI9923bc0_541, \2610 );
and \U$1044 ( \3164 , RI9924520_521, \2612 );
and \U$1045 ( \3165 , RI9925510_501, \2614 );
and \U$1046 ( \3166 , RI9925e70_481, \2616 );
and \U$1047 ( \3167 , RI99267d0_461, \2618 );
and \U$1048 ( \3168 , RI9927b80_441, \2620 );
and \U$1049 ( \3169 , RI99284e0_421, \2622 );
and \U$1050 ( \3170 , RI9928e40_401, \2624 );
and \U$1051 ( \3171 , RI992a5b0_381, \2626 );
and \U$1052 ( \3172 , RI992af10_361, \2628 );
and \U$1053 ( \3173 , RI992ca40_341, \2630 );
and \U$1054 ( \3174 , RI992d3a0_321, \2632 );
and \U$1055 ( \3175 , RI992f290_301, \2634 );
and \U$1056 ( \3176 , RI9931540_281, \2636 );
and \U$1057 ( \3177 , RI9933bb0_261, \2638 );
or \U$1058 ( \3178 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 );
_DC g1e79 ( \3179_nG1e79 , \3178 , \2657 );
buf \U$1059 ( \3180 , \3179_nG1e79 );
and \U$1060 ( \3181 , \3180 , \2834 );
and \U$1061 ( \3182 , RI99226a8_580, \2602 );
and \U$1062 ( \3183 , RI99232d8_560, \2608 );
and \U$1063 ( \3184 , RI9923c38_540, \2610 );
and \U$1064 ( \3185 , RI9924598_520, \2612 );
and \U$1065 ( \3186 , RI9925588_500, \2614 );
and \U$1066 ( \3187 , RI9925ee8_480, \2616 );
and \U$1067 ( \3188 , RI9926848_460, \2618 );
and \U$1068 ( \3189 , RI9927bf8_440, \2620 );
and \U$1069 ( \3190 , RI9928558_420, \2622 );
and \U$1070 ( \3191 , RI9928eb8_400, \2624 );
and \U$1071 ( \3192 , RI992a628_380, \2626 );
and \U$1072 ( \3193 , RI992af88_360, \2628 );
and \U$1073 ( \3194 , RI992cab8_340, \2630 );
and \U$1074 ( \3195 , RI992d418_320, \2632 );
and \U$1075 ( \3196 , RI992f308_300, \2634 );
and \U$1076 ( \3197 , RI99315b8_280, \2636 );
and \U$1077 ( \3198 , RI9933c28_260, \2638 );
or \U$1078 ( \3199 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 );
_DC g1f2c ( \3200_nG1f2c , \3199 , \2657 );
buf \U$1079 ( \3201 , \3200_nG1f2c );
and \U$1080 ( \3202 , \3201 , \2832 );
nor \U$1081 ( \3203 , \3181 , \3202 );
xnor \U$1082 ( \3204 , \3203 , \2839 );
and \U$1083 ( \3205 , \3160 , \3204 );
and \U$1084 ( \3206 , RI9922540_583, \2602 );
and \U$1085 ( \3207 , RI9923170_563, \2608 );
and \U$1086 ( \3208 , RI9923ad0_543, \2610 );
and \U$1087 ( \3209 , RI9924430_523, \2612 );
and \U$1088 ( \3210 , RI9924d90_503, \2614 );
and \U$1089 ( \3211 , RI9925d80_483, \2616 );
and \U$1090 ( \3212 , RI99266e0_463, \2618 );
and \U$1091 ( \3213 , RI9927040_443, \2620 );
and \U$1092 ( \3214 , RI99283f0_423, \2622 );
and \U$1093 ( \3215 , RI9928d50_403, \2624 );
and \U$1094 ( \3216 , RI992a4c0_383, \2626 );
and \U$1095 ( \3217 , RI992ae20_363, \2628 );
and \U$1096 ( \3218 , RI992c950_343, \2630 );
and \U$1097 ( \3219 , RI992d2b0_323, \2632 );
and \U$1098 ( \3220 , RI992f1a0_303, \2634 );
and \U$1099 ( \3221 , RI9931450_283, \2636 );
and \U$1100 ( \3222 , RI9933ac0_263, \2638 );
or \U$1101 ( \3223 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 );
_DC g1d15 ( \3224_nG1d15 , \3223 , \2657 );
buf \U$1102 ( \3225 , \3224_nG1d15 );
and \U$1103 ( \3226 , \3225 , \2769 );
and \U$1104 ( \3227 , RI99225b8_582, \2602 );
and \U$1105 ( \3228 , RI99231e8_562, \2608 );
and \U$1106 ( \3229 , RI9923b48_542, \2610 );
and \U$1107 ( \3230 , RI99244a8_522, \2612 );
and \U$1108 ( \3231 , RI9924e08_502, \2614 );
and \U$1109 ( \3232 , RI9925df8_482, \2616 );
and \U$1110 ( \3233 , RI9926758_462, \2618 );
and \U$1111 ( \3234 , RI9927b08_442, \2620 );
and \U$1112 ( \3235 , RI9928468_422, \2622 );
and \U$1113 ( \3236 , RI9928dc8_402, \2624 );
and \U$1114 ( \3237 , RI992a538_382, \2626 );
and \U$1115 ( \3238 , RI992ae98_362, \2628 );
and \U$1116 ( \3239 , RI992c9c8_342, \2630 );
and \U$1117 ( \3240 , RI992d328_322, \2632 );
and \U$1118 ( \3241 , RI992f218_302, \2634 );
and \U$1119 ( \3242 , RI99314c8_282, \2636 );
and \U$1120 ( \3243 , RI9933b38_262, \2638 );
or \U$1121 ( \3244 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 );
_DC g1dbc ( \3245_nG1dbc , \3244 , \2657 );
buf \U$1122 ( \3246 , \3245_nG1dbc );
and \U$1123 ( \3247 , \3246 , \2767 );
nor \U$1124 ( \3248 , \3226 , \3247 );
xnor \U$1125 ( \3249 , \3248 , \2536 );
and \U$1126 ( \3250 , \3204 , \3249 );
and \U$1127 ( \3251 , \3160 , \3249 );
or \U$1128 ( \3252 , \3205 , \3250 , \3251 );
and \U$1129 ( \3253 , \3105 , \3252 );
and \U$1130 ( \3254 , RI9922450_585, \2602 );
and \U$1131 ( \3255 , RI9923080_565, \2608 );
and \U$1132 ( \3256 , RI99239e0_545, \2610 );
and \U$1133 ( \3257 , RI9924340_525, \2612 );
and \U$1134 ( \3258 , RI9924ca0_505, \2614 );
and \U$1135 ( \3259 , RI9925c90_485, \2616 );
and \U$1136 ( \3260 , RI99265f0_465, \2618 );
and \U$1137 ( \3261 , RI9926f50_445, \2620 );
and \U$1138 ( \3262 , RI9928300_425, \2622 );
and \U$1139 ( \3263 , RI9928c60_405, \2624 );
and \U$1140 ( \3264 , RI992a3d0_385, \2626 );
and \U$1141 ( \3265 , RI992ad30_365, \2628 );
and \U$1142 ( \3266 , RI992c860_345, \2630 );
and \U$1143 ( \3267 , RI992d1c0_325, \2632 );
and \U$1144 ( \3268 , RI992f0b0_305, \2634 );
and \U$1145 ( \3269 , RI9931360_285, \2636 );
and \U$1146 ( \3270 , RI99339d0_265, \2638 );
or \U$1147 ( \3271 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 );
_DC g1ba5 ( \3272_nG1ba5 , \3271 , \2657 );
buf \U$1148 ( \3273 , \3272_nG1ba5 );
and \U$1149 ( \3274 , \3273 , \2707 );
and \U$1150 ( \3275 , RI99224c8_584, \2602 );
and \U$1151 ( \3276 , RI99230f8_564, \2608 );
and \U$1152 ( \3277 , RI9923a58_544, \2610 );
and \U$1153 ( \3278 , RI99243b8_524, \2612 );
and \U$1154 ( \3279 , RI9924d18_504, \2614 );
and \U$1155 ( \3280 , RI9925d08_484, \2616 );
and \U$1156 ( \3281 , RI9926668_464, \2618 );
and \U$1157 ( \3282 , RI9926fc8_444, \2620 );
and \U$1158 ( \3283 , RI9928378_424, \2622 );
and \U$1159 ( \3284 , RI9928cd8_404, \2624 );
and \U$1160 ( \3285 , RI992a448_384, \2626 );
and \U$1161 ( \3286 , RI992ada8_364, \2628 );
and \U$1162 ( \3287 , RI992c8d8_344, \2630 );
and \U$1163 ( \3288 , RI992d238_324, \2632 );
and \U$1164 ( \3289 , RI992f128_304, \2634 );
and \U$1165 ( \3290 , RI99313d8_284, \2636 );
and \U$1166 ( \3291 , RI9933a48_264, \2638 );
or \U$1167 ( \3292 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 );
_DC g1c76 ( \3293_nG1c76 , \3292 , \2657 );
buf \U$1168 ( \3294 , \3293_nG1c76 );
and \U$1169 ( \3295 , \3294 , \2705 );
nor \U$1170 ( \3296 , \3274 , \3295 );
xnor \U$1171 ( \3297 , \3296 , \2733 );
and \U$1173 ( \3298 , RI99223d8_586, \2602 );
and \U$1174 ( \3299 , RI9923008_566, \2608 );
and \U$1175 ( \3300 , RI9923968_546, \2610 );
and \U$1176 ( \3301 , RI99242c8_526, \2612 );
and \U$1177 ( \3302 , RI9924c28_506, \2614 );
and \U$1178 ( \3303 , RI9925c18_486, \2616 );
and \U$1179 ( \3304 , RI9926578_466, \2618 );
and \U$1180 ( \3305 , RI9926ed8_446, \2620 );
and \U$1181 ( \3306 , RI9928288_426, \2622 );
and \U$1182 ( \3307 , RI9928be8_406, \2624 );
and \U$1183 ( \3308 , RI992a358_386, \2626 );
and \U$1184 ( \3309 , RI992acb8_366, \2628 );
and \U$1185 ( \3310 , RI992c7e8_346, \2630 );
and \U$1186 ( \3311 , RI992d148_326, \2632 );
and \U$1187 ( \3312 , RI992f038_306, \2634 );
and \U$1188 ( \3313 , RI99312e8_286, \2636 );
and \U$1189 ( \3314 , RI9933958_266, \2638 );
or \U$1190 ( \3315 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 );
_DC g1b63 ( \3316_nG1b63 , \3315 , \2657 );
buf \U$1191 ( \3317 , \3316_nG1b63 );
and \U$1192 ( \3318 , \3317 , \2760 );
nor \U$1193 ( \3319 , 1'b0 , \3318 );
xnor \U$1194 ( \3320 , \3319 , 1'b0 );
and \U$1195 ( \3321 , \3297 , \3320 );
and \U$1196 ( \3322 , \3252 , \3321 );
and \U$1197 ( \3323 , \3105 , \3321 );
or \U$1198 ( \3324 , \3253 , \3322 , \3323 );
and \U$1200 ( \3325 , \3246 , \2769 );
and \U$1201 ( \3326 , \3180 , \2767 );
nor \U$1202 ( \3327 , \3325 , \3326 );
xnor \U$1203 ( \3328 , \3327 , \2536 );
and \U$1204 ( \3329 , \3294 , \2707 );
and \U$1205 ( \3330 , \3225 , \2705 );
nor \U$1206 ( \3331 , \3329 , \3330 );
xnor \U$1207 ( \3332 , \3331 , \2733 );
xor \U$1208 ( \3333 , \3328 , \3332 );
and \U$1210 ( \3334 , \3273 , \2760 );
nor \U$1211 ( \3335 , 1'b0 , \3334 );
xnor \U$1212 ( \3336 , \3335 , 1'b0 );
xor \U$1213 ( \3337 , \3333 , \3336 );
and \U$1214 ( \3338 , \3096 , \3075 );
and \U$1215 ( \3339 , \3003 , \3073 );
nor \U$1216 ( \3340 , \3338 , \3339 );
xnor \U$1217 ( \3341 , \3340 , \3101 );
and \U$1218 ( \3342 , \3154 , \3133 );
and \U$1219 ( \3343 , \3063 , \3131 );
nor \U$1220 ( \3344 , \3342 , \3343 );
xnor \U$1221 ( \3345 , \3344 , \3159 );
xor \U$1222 ( \3346 , \3341 , \3345 );
and \U$1223 ( \3347 , \3201 , \2834 );
and \U$1224 ( \3348 , \3125 , \2832 );
nor \U$1225 ( \3349 , \3347 , \3348 );
xnor \U$1226 ( \3350 , \3349 , \2839 );
xor \U$1227 ( \3351 , \3346 , \3350 );
and \U$1228 ( \3352 , \3337 , \3351 );
or \U$1230 ( \3353 , 1'b0 , \3352 , 1'b0 );
xor \U$1231 ( \3354 , \3324 , \3353 );
and \U$1232 ( \3355 , \3225 , \2707 );
and \U$1233 ( \3356 , \3246 , \2705 );
nor \U$1234 ( \3357 , \3355 , \3356 );
xnor \U$1235 ( \3358 , \3357 , \2733 );
and \U$1237 ( \3359 , \3294 , \2760 );
nor \U$1238 ( \3360 , 1'b0 , \3359 );
xnor \U$1239 ( \3361 , \3360 , 1'b0 );
xor \U$1240 ( \3362 , \3358 , \3361 );
xor \U$1242 ( \3363 , \3362 , 1'b0 );
and \U$1243 ( \3364 , \3063 , \3133 );
and \U$1244 ( \3365 , \3096 , \3131 );
nor \U$1245 ( \3366 , \3364 , \3365 );
xnor \U$1246 ( \3367 , \3366 , \3159 );
and \U$1247 ( \3368 , \3125 , \2834 );
and \U$1248 ( \3369 , \3154 , \2832 );
nor \U$1249 ( \3370 , \3368 , \3369 );
xnor \U$1250 ( \3371 , \3370 , \2839 );
xor \U$1251 ( \3372 , \3367 , \3371 );
and \U$1252 ( \3373 , \3180 , \2769 );
and \U$1253 ( \3374 , \3201 , \2767 );
nor \U$1254 ( \3375 , \3373 , \3374 );
xnor \U$1255 ( \3376 , \3375 , \2536 );
xor \U$1256 ( \3377 , \3372 , \3376 );
xor \U$1257 ( \3378 , \3363 , \3377 );
and \U$1258 ( \3379 , \2887 , \2979 );
and \U$1259 ( \3380 , \2755 , \2976 );
nor \U$1260 ( \3381 , \3379 , \3380 );
xnor \U$1261 ( \3382 , \3381 , \2973 );
and \U$1262 ( \3383 , \2910 , \3015 );
and \U$1263 ( \3384 , \2866 , \3013 );
nor \U$1264 ( \3385 , \3383 , \3384 );
xnor \U$1265 ( \3386 , \3385 , \3041 );
xor \U$1266 ( \3387 , \3382 , \3386 );
and \U$1267 ( \3388 , \3003 , \3075 );
and \U$1268 ( \3389 , \3036 , \3073 );
nor \U$1269 ( \3390 , \3388 , \3389 );
xnor \U$1270 ( \3391 , \3390 , \3101 );
xor \U$1271 ( \3392 , \3387 , \3391 );
xor \U$1272 ( \3393 , \3378 , \3392 );
xor \U$1273 ( \3394 , \3354 , \3393 );
and \U$1275 ( \3395 , \3036 , \2979 );
and \U$1276 ( \3396 , \2910 , \2976 );
nor \U$1277 ( \3397 , \3395 , \3396 );
xnor \U$1278 ( \3398 , \3397 , \2973 );
and \U$1279 ( \3399 , \3096 , \3015 );
and \U$1280 ( \3400 , \3003 , \3013 );
nor \U$1281 ( \3401 , \3399 , \3400 );
xnor \U$1282 ( \3402 , \3401 , \3041 );
and \U$1283 ( \3403 , \3398 , \3402 );
or \U$1285 ( \3404 , 1'b0 , \3403 , 1'b0 );
and \U$1286 ( \3405 , \3154 , \3075 );
and \U$1287 ( \3406 , \3063 , \3073 );
nor \U$1288 ( \3407 , \3405 , \3406 );
xnor \U$1289 ( \3408 , \3407 , \3101 );
and \U$1290 ( \3409 , \3201 , \3133 );
and \U$1291 ( \3410 , \3125 , \3131 );
nor \U$1292 ( \3411 , \3409 , \3410 );
xnor \U$1293 ( \3412 , \3411 , \3159 );
and \U$1294 ( \3413 , \3408 , \3412 );
and \U$1295 ( \3414 , \3246 , \2834 );
and \U$1296 ( \3415 , \3180 , \2832 );
nor \U$1297 ( \3416 , \3414 , \3415 );
xnor \U$1298 ( \3417 , \3416 , \2839 );
and \U$1299 ( \3418 , \3412 , \3417 );
and \U$1300 ( \3419 , \3408 , \3417 );
or \U$1301 ( \3420 , \3413 , \3418 , \3419 );
and \U$1302 ( \3421 , \3404 , \3420 );
and \U$1303 ( \3422 , \3294 , \2769 );
and \U$1304 ( \3423 , \3225 , \2767 );
nor \U$1305 ( \3424 , \3422 , \3423 );
xnor \U$1306 ( \3425 , \3424 , \2536 );
and \U$1307 ( \3426 , \3317 , \2707 );
and \U$1308 ( \3427 , \3273 , \2705 );
nor \U$1309 ( \3428 , \3426 , \3427 );
xnor \U$1310 ( \3429 , \3428 , \2733 );
and \U$1311 ( \3430 , \3425 , \3429 );
and \U$1312 ( \3431 , RI9922360_587, \2602 );
and \U$1313 ( \3432 , RI9922f90_567, \2608 );
and \U$1314 ( \3433 , RI99238f0_547, \2610 );
and \U$1315 ( \3434 , RI9924250_527, \2612 );
and \U$1316 ( \3435 , RI9924bb0_507, \2614 );
and \U$1317 ( \3436 , RI9925ba0_487, \2616 );
and \U$1318 ( \3437 , RI9926500_467, \2618 );
and \U$1319 ( \3438 , RI9926e60_447, \2620 );
and \U$1320 ( \3439 , RI9928210_427, \2622 );
and \U$1321 ( \3440 , RI9928b70_407, \2624 );
and \U$1322 ( \3441 , RI992a2e0_387, \2626 );
and \U$1323 ( \3442 , RI992ac40_367, \2628 );
and \U$1324 ( \3443 , RI992c770_347, \2630 );
and \U$1325 ( \3444 , RI992d0d0_327, \2632 );
and \U$1326 ( \3445 , RI992efc0_307, \2634 );
and \U$1327 ( \3446 , RI992f920_287, \2636 );
and \U$1328 ( \3447 , RI99338e0_267, \2638 );
or \U$1329 ( \3448 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 );
_DC g1a4f ( \3449_nG1a4f , \3448 , \2657 );
buf \U$1330 ( \3450 , \3449_nG1a4f );
nand \U$1331 ( \3451 , \3450 , \2760 );
xnor \U$1332 ( \3452 , \3451 , 1'b0 );
and \U$1333 ( \3453 , \3429 , \3452 );
and \U$1334 ( \3454 , \3425 , \3452 );
or \U$1335 ( \3455 , \3430 , \3453 , \3454 );
and \U$1336 ( \3456 , \3420 , \3455 );
and \U$1337 ( \3457 , \3404 , \3455 );
or \U$1338 ( \3458 , \3421 , \3456 , \3457 );
xor \U$1339 ( \3459 , \3297 , \3320 );
xor \U$1340 ( \3460 , \3160 , \3204 );
xor \U$1341 ( \3461 , \3460 , \3249 );
and \U$1342 ( \3462 , \3459 , \3461 );
xor \U$1343 ( \3463 , \2983 , \3042 );
xor \U$1344 ( \3464 , \3463 , \3102 );
and \U$1345 ( \3465 , \3461 , \3464 );
and \U$1346 ( \3466 , \3459 , \3464 );
or \U$1347 ( \3467 , \3462 , \3465 , \3466 );
and \U$1348 ( \3468 , \3458 , \3467 );
and \U$1350 ( \3469 , \2866 , \2979 );
and \U$1351 ( \3470 , \2887 , \2976 );
nor \U$1352 ( \3471 , \3469 , \3470 );
xnor \U$1353 ( \3472 , \3471 , \2973 );
xor \U$1354 ( \3473 , 1'b0 , \3472 );
and \U$1355 ( \3474 , \3036 , \3015 );
and \U$1356 ( \3475 , \2910 , \3013 );
nor \U$1357 ( \3476 , \3474 , \3475 );
xnor \U$1358 ( \3477 , \3476 , \3041 );
xor \U$1359 ( \3478 , \3473 , \3477 );
and \U$1360 ( \3479 , \3467 , \3478 );
and \U$1361 ( \3480 , \3458 , \3478 );
or \U$1362 ( \3481 , \3468 , \3479 , \3480 );
xor \U$1364 ( \3482 , 1'b0 , \3337 );
xor \U$1365 ( \3483 , \3482 , \3351 );
xor \U$1366 ( \3484 , \3105 , \3252 );
xor \U$1367 ( \3485 , \3484 , \3321 );
and \U$1368 ( \3486 , \3483 , \3485 );
xor \U$1369 ( \3487 , \3481 , \3486 );
and \U$1371 ( \3488 , \3472 , \3477 );
or \U$1373 ( \3489 , 1'b0 , \3488 , 1'b0 );
and \U$1374 ( \3490 , \3341 , \3345 );
and \U$1375 ( \3491 , \3345 , \3350 );
and \U$1376 ( \3492 , \3341 , \3350 );
or \U$1377 ( \3493 , \3490 , \3491 , \3492 );
xor \U$1378 ( \3494 , \3489 , \3493 );
and \U$1379 ( \3495 , \3328 , \3332 );
and \U$1380 ( \3496 , \3332 , \3336 );
and \U$1381 ( \3497 , \3328 , \3336 );
or \U$1382 ( \3498 , \3495 , \3496 , \3497 );
xor \U$1383 ( \3499 , \3494 , \3498 );
xor \U$1384 ( \3500 , \3487 , \3499 );
xor \U$1385 ( \3501 , \3394 , \3500 );
and \U$1386 ( \3502 , \3003 , \2979 );
and \U$1387 ( \3503 , \3036 , \2976 );
nor \U$1388 ( \3504 , \3502 , \3503 );
xnor \U$1389 ( \3505 , \3504 , \2973 );
and \U$1390 ( \3506 , \3063 , \3015 );
and \U$1391 ( \3507 , \3096 , \3013 );
nor \U$1392 ( \3508 , \3506 , \3507 );
xnor \U$1393 ( \3509 , \3508 , \3041 );
and \U$1394 ( \3510 , \3505 , \3509 );
and \U$1395 ( \3511 , \3125 , \3075 );
and \U$1396 ( \3512 , \3154 , \3073 );
nor \U$1397 ( \3513 , \3511 , \3512 );
xnor \U$1398 ( \3514 , \3513 , \3101 );
and \U$1399 ( \3515 , \3509 , \3514 );
and \U$1400 ( \3516 , \3505 , \3514 );
or \U$1401 ( \3517 , \3510 , \3515 , \3516 );
and \U$1402 ( \3518 , \3180 , \3133 );
and \U$1403 ( \3519 , \3201 , \3131 );
nor \U$1404 ( \3520 , \3518 , \3519 );
xnor \U$1405 ( \3521 , \3520 , \3159 );
and \U$1406 ( \3522 , \3225 , \2834 );
and \U$1407 ( \3523 , \3246 , \2832 );
nor \U$1408 ( \3524 , \3522 , \3523 );
xnor \U$1409 ( \3525 , \3524 , \2839 );
and \U$1410 ( \3526 , \3521 , \3525 );
and \U$1411 ( \3527 , \3273 , \2769 );
and \U$1412 ( \3528 , \3294 , \2767 );
nor \U$1413 ( \3529 , \3527 , \3528 );
xnor \U$1414 ( \3530 , \3529 , \2536 );
and \U$1415 ( \3531 , \3525 , \3530 );
and \U$1416 ( \3532 , \3521 , \3530 );
or \U$1417 ( \3533 , \3526 , \3531 , \3532 );
and \U$1418 ( \3534 , \3517 , \3533 );
xor \U$1419 ( \3535 , \3425 , \3429 );
xor \U$1420 ( \3536 , \3535 , \3452 );
and \U$1421 ( \3537 , \3533 , \3536 );
and \U$1422 ( \3538 , \3517 , \3536 );
or \U$1423 ( \3539 , \3534 , \3537 , \3538 );
xor \U$1424 ( \3540 , \3408 , \3412 );
xor \U$1425 ( \3541 , \3540 , \3417 );
xor \U$1426 ( \3542 , 1'b0 , \3398 );
xor \U$1427 ( \3543 , \3542 , \3402 );
and \U$1428 ( \3544 , \3541 , \3543 );
and \U$1429 ( \3545 , \3539 , \3544 );
xor \U$1430 ( \3546 , \3459 , \3461 );
xor \U$1431 ( \3547 , \3546 , \3464 );
and \U$1432 ( \3548 , \3544 , \3547 );
and \U$1433 ( \3549 , \3539 , \3547 );
or \U$1434 ( \3550 , \3545 , \3548 , \3549 );
xor \U$1435 ( \3551 , \3483 , \3485 );
and \U$1436 ( \3552 , \3550 , \3551 );
xor \U$1437 ( \3553 , \3458 , \3467 );
xor \U$1438 ( \3554 , \3553 , \3478 );
and \U$1439 ( \3555 , \3551 , \3554 );
and \U$1440 ( \3556 , \3550 , \3554 );
or \U$1441 ( \3557 , \3552 , \3555 , \3556 );
nor \U$1442 ( \3558 , \3501 , \3557 );
and \U$1443 ( \3559 , \3481 , \3486 );
and \U$1444 ( \3560 , \3486 , \3499 );
and \U$1445 ( \3561 , \3481 , \3499 );
or \U$1446 ( \3562 , \3559 , \3560 , \3561 );
and \U$1447 ( \3563 , \3324 , \3353 );
and \U$1448 ( \3564 , \3353 , \3393 );
and \U$1449 ( \3565 , \3324 , \3393 );
or \U$1450 ( \3566 , \3563 , \3564 , \3565 );
and \U$1452 ( \3567 , \2755 , \2979 );
and \U$1453 ( \3568 , \2659 , \2976 );
nor \U$1454 ( \3569 , \3567 , \3568 );
xnor \U$1455 ( \3570 , \3569 , \2973 );
xor \U$1456 ( \3571 , 1'b0 , \3570 );
and \U$1457 ( \3572 , \2866 , \3015 );
and \U$1458 ( \3573 , \2887 , \3013 );
nor \U$1459 ( \3574 , \3572 , \3573 );
xnor \U$1460 ( \3575 , \3574 , \3041 );
xor \U$1461 ( \3576 , \3571 , \3575 );
and \U$1463 ( \3577 , \3201 , \2769 );
and \U$1464 ( \3578 , \3125 , \2767 );
nor \U$1465 ( \3579 , \3577 , \3578 );
xnor \U$1466 ( \3580 , \3579 , \2536 );
and \U$1467 ( \3581 , \3246 , \2707 );
and \U$1468 ( \3582 , \3180 , \2705 );
nor \U$1469 ( \3583 , \3581 , \3582 );
xnor \U$1470 ( \3584 , \3583 , \2733 );
xor \U$1471 ( \3585 , \3580 , \3584 );
and \U$1473 ( \3586 , \3225 , \2760 );
nor \U$1474 ( \3587 , 1'b0 , \3586 );
xnor \U$1475 ( \3588 , \3587 , 1'b0 );
xor \U$1476 ( \3589 , \3585 , \3588 );
xor \U$1477 ( \3590 , 1'b0 , \3589 );
xor \U$1478 ( \3591 , \3576 , \3590 );
and \U$1479 ( \3592 , \3382 , \3386 );
and \U$1480 ( \3593 , \3386 , \3391 );
and \U$1481 ( \3594 , \3382 , \3391 );
or \U$1482 ( \3595 , \3592 , \3593 , \3594 );
and \U$1483 ( \3596 , \3367 , \3371 );
and \U$1484 ( \3597 , \3371 , \3376 );
and \U$1485 ( \3598 , \3367 , \3376 );
or \U$1486 ( \3599 , \3596 , \3597 , \3598 );
xor \U$1487 ( \3600 , \3595 , \3599 );
and \U$1488 ( \3601 , \3358 , \3361 );
or \U$1491 ( \3602 , \3601 , 1'b0 , 1'b0 );
xor \U$1492 ( \3603 , \3600 , \3602 );
xor \U$1493 ( \3604 , \3591 , \3603 );
xor \U$1494 ( \3605 , \3566 , \3604 );
and \U$1495 ( \3606 , \3489 , \3493 );
and \U$1496 ( \3607 , \3493 , \3498 );
and \U$1497 ( \3608 , \3489 , \3498 );
or \U$1498 ( \3609 , \3606 , \3607 , \3608 );
and \U$1499 ( \3610 , \3363 , \3377 );
and \U$1500 ( \3611 , \3377 , \3392 );
and \U$1501 ( \3612 , \3363 , \3392 );
or \U$1502 ( \3613 , \3610 , \3611 , \3612 );
xor \U$1503 ( \3614 , \3609 , \3613 );
and \U$1504 ( \3615 , \3036 , \3075 );
and \U$1505 ( \3616 , \2910 , \3073 );
nor \U$1506 ( \3617 , \3615 , \3616 );
xnor \U$1507 ( \3618 , \3617 , \3101 );
and \U$1508 ( \3619 , \3096 , \3133 );
and \U$1509 ( \3620 , \3003 , \3131 );
nor \U$1510 ( \3621 , \3619 , \3620 );
xnor \U$1511 ( \3622 , \3621 , \3159 );
xor \U$1512 ( \3623 , \3618 , \3622 );
and \U$1513 ( \3624 , \3154 , \2834 );
and \U$1514 ( \3625 , \3063 , \2832 );
nor \U$1515 ( \3626 , \3624 , \3625 );
xnor \U$1516 ( \3627 , \3626 , \2839 );
xor \U$1517 ( \3628 , \3623 , \3627 );
xor \U$1518 ( \3629 , \3614 , \3628 );
xor \U$1519 ( \3630 , \3605 , \3629 );
xor \U$1520 ( \3631 , \3562 , \3630 );
and \U$1521 ( \3632 , \3394 , \3500 );
nor \U$1522 ( \3633 , \3631 , \3632 );
nor \U$1523 ( \3634 , \3558 , \3633 );
and \U$1524 ( \3635 , \3566 , \3604 );
and \U$1525 ( \3636 , \3604 , \3629 );
and \U$1526 ( \3637 , \3566 , \3629 );
or \U$1527 ( \3638 , \3635 , \3636 , \3637 );
and \U$1529 ( \3639 , \3570 , \3575 );
or \U$1531 ( \3640 , 1'b0 , \3639 , 1'b0 );
and \U$1532 ( \3641 , \3618 , \3622 );
and \U$1533 ( \3642 , \3622 , \3627 );
and \U$1534 ( \3643 , \3618 , \3627 );
or \U$1535 ( \3644 , \3641 , \3642 , \3643 );
xor \U$1536 ( \3645 , \3640 , \3644 );
and \U$1537 ( \3646 , \3580 , \3584 );
and \U$1538 ( \3647 , \3584 , \3588 );
and \U$1539 ( \3648 , \3580 , \3588 );
or \U$1540 ( \3649 , \3646 , \3647 , \3648 );
xor \U$1541 ( \3650 , \3645 , \3649 );
and \U$1542 ( \3651 , \3595 , \3599 );
and \U$1543 ( \3652 , \3599 , \3602 );
and \U$1544 ( \3653 , \3595 , \3602 );
or \U$1545 ( \3654 , \3651 , \3652 , \3653 );
xor \U$1547 ( \3655 , \3654 , 1'b0 );
and \U$1548 ( \3656 , \2659 , \2979 );
and \U$1549 ( \3657 , \2728 , \2976 );
nor \U$1550 ( \3658 , \3656 , \3657 );
xnor \U$1551 ( \3659 , \3658 , \2973 );
and \U$1552 ( \3660 , \2887 , \3015 );
and \U$1553 ( \3661 , \2755 , \3013 );
nor \U$1554 ( \3662 , \3660 , \3661 );
xnor \U$1555 ( \3663 , \3662 , \3041 );
xor \U$1556 ( \3664 , \3659 , \3663 );
and \U$1557 ( \3665 , \2910 , \3075 );
and \U$1558 ( \3666 , \2866 , \3073 );
nor \U$1559 ( \3667 , \3665 , \3666 );
xnor \U$1560 ( \3668 , \3667 , \3101 );
xor \U$1561 ( \3669 , \3664 , \3668 );
xor \U$1562 ( \3670 , \3655 , \3669 );
xor \U$1563 ( \3671 , \3650 , \3670 );
xor \U$1564 ( \3672 , \3638 , \3671 );
and \U$1565 ( \3673 , \3609 , \3613 );
and \U$1566 ( \3674 , \3613 , \3628 );
and \U$1567 ( \3675 , \3609 , \3628 );
or \U$1568 ( \3676 , \3673 , \3674 , \3675 );
and \U$1569 ( \3677 , \3576 , \3590 );
and \U$1570 ( \3678 , \3590 , \3603 );
and \U$1571 ( \3679 , \3576 , \3603 );
or \U$1572 ( \3680 , \3677 , \3678 , \3679 );
xor \U$1573 ( \3681 , \3676 , \3680 );
and \U$1575 ( \3682 , \3180 , \2707 );
and \U$1576 ( \3683 , \3201 , \2705 );
nor \U$1577 ( \3684 , \3682 , \3683 );
xnor \U$1578 ( \3685 , \3684 , \2733 );
and \U$1580 ( \3686 , \3246 , \2760 );
nor \U$1581 ( \3687 , 1'b0 , \3686 );
xnor \U$1582 ( \3688 , \3687 , 1'b0 );
xor \U$1583 ( \3689 , \3685 , \3688 );
xor \U$1585 ( \3690 , \3689 , 1'b0 );
xor \U$1586 ( \3691 , 1'b0 , \3690 );
and \U$1587 ( \3692 , \3003 , \3133 );
and \U$1588 ( \3693 , \3036 , \3131 );
nor \U$1589 ( \3694 , \3692 , \3693 );
xnor \U$1590 ( \3695 , \3694 , \3159 );
and \U$1591 ( \3696 , \3063 , \2834 );
and \U$1592 ( \3697 , \3096 , \2832 );
nor \U$1593 ( \3698 , \3696 , \3697 );
xnor \U$1594 ( \3699 , \3698 , \2839 );
xor \U$1595 ( \3700 , \3695 , \3699 );
and \U$1596 ( \3701 , \3125 , \2769 );
and \U$1597 ( \3702 , \3154 , \2767 );
nor \U$1598 ( \3703 , \3701 , \3702 );
xnor \U$1599 ( \3704 , \3703 , \2536 );
xor \U$1600 ( \3705 , \3700 , \3704 );
xor \U$1601 ( \3706 , \3691 , \3705 );
xor \U$1602 ( \3707 , \3681 , \3706 );
xor \U$1603 ( \3708 , \3672 , \3707 );
and \U$1604 ( \3709 , \3562 , \3630 );
nor \U$1605 ( \3710 , \3708 , \3709 );
and \U$1606 ( \3711 , \3676 , \3680 );
and \U$1607 ( \3712 , \3680 , \3706 );
and \U$1608 ( \3713 , \3676 , \3706 );
or \U$1609 ( \3714 , \3711 , \3712 , \3713 );
and \U$1610 ( \3715 , \3650 , \3670 );
xor \U$1611 ( \3716 , \3714 , \3715 );
and \U$1614 ( \3717 , \3654 , \3669 );
or \U$1615 ( \3718 , 1'b0 , 1'b0 , \3717 );
and \U$1617 ( \3719 , \3154 , \2769 );
and \U$1618 ( \3720 , \3063 , \2767 );
nor \U$1619 ( \3721 , \3719 , \3720 );
xnor \U$1620 ( \3722 , \3721 , \2536 );
and \U$1621 ( \3723 , \3201 , \2707 );
and \U$1622 ( \3724 , \3125 , \2705 );
nor \U$1623 ( \3725 , \3723 , \3724 );
xnor \U$1624 ( \3726 , \3725 , \2733 );
xor \U$1625 ( \3727 , \3722 , \3726 );
and \U$1627 ( \3728 , \3180 , \2760 );
nor \U$1628 ( \3729 , 1'b0 , \3728 );
xnor \U$1629 ( \3730 , \3729 , 1'b0 );
xor \U$1630 ( \3731 , \3727 , \3730 );
xor \U$1631 ( \3732 , 1'b0 , \3731 );
and \U$1632 ( \3733 , \2866 , \3075 );
and \U$1633 ( \3734 , \2887 , \3073 );
nor \U$1634 ( \3735 , \3733 , \3734 );
xnor \U$1635 ( \3736 , \3735 , \3101 );
and \U$1636 ( \3737 , \3036 , \3133 );
and \U$1637 ( \3738 , \2910 , \3131 );
nor \U$1638 ( \3739 , \3737 , \3738 );
xnor \U$1639 ( \3740 , \3739 , \3159 );
xor \U$1640 ( \3741 , \3736 , \3740 );
and \U$1641 ( \3742 , \3096 , \2834 );
and \U$1642 ( \3743 , \3003 , \2832 );
nor \U$1643 ( \3744 , \3742 , \3743 );
xnor \U$1644 ( \3745 , \3744 , \2839 );
xor \U$1645 ( \3746 , \3741 , \3745 );
xor \U$1646 ( \3747 , \3732 , \3746 );
and \U$1647 ( \3748 , \3659 , \3663 );
and \U$1648 ( \3749 , \3663 , \3668 );
and \U$1649 ( \3750 , \3659 , \3668 );
or \U$1650 ( \3751 , \3748 , \3749 , \3750 );
and \U$1651 ( \3752 , \3695 , \3699 );
and \U$1652 ( \3753 , \3699 , \3704 );
and \U$1653 ( \3754 , \3695 , \3704 );
or \U$1654 ( \3755 , \3752 , \3753 , \3754 );
xor \U$1655 ( \3756 , \3751 , \3755 );
and \U$1656 ( \3757 , \3685 , \3688 );
or \U$1659 ( \3758 , \3757 , 1'b0 , 1'b0 );
xor \U$1660 ( \3759 , \3756 , \3758 );
xor \U$1661 ( \3760 , \3747 , \3759 );
xor \U$1662 ( \3761 , \3718 , \3760 );
and \U$1663 ( \3762 , \3640 , \3644 );
and \U$1664 ( \3763 , \3644 , \3649 );
and \U$1665 ( \3764 , \3640 , \3649 );
or \U$1666 ( \3765 , \3762 , \3763 , \3764 );
and \U$1668 ( \3766 , \3690 , \3705 );
or \U$1670 ( \3767 , 1'b0 , \3766 , 1'b0 );
xor \U$1671 ( \3768 , \3765 , \3767 );
and \U$1673 ( \3769 , \2728 , \2979 );
not \U$1674 ( \3770 , \3769 );
xnor \U$1675 ( \3771 , \3770 , \2973 );
xor \U$1676 ( \3772 , 1'b0 , \3771 );
and \U$1677 ( \3773 , \2755 , \3015 );
and \U$1678 ( \3774 , \2659 , \3013 );
nor \U$1679 ( \3775 , \3773 , \3774 );
xnor \U$1680 ( \3776 , \3775 , \3041 );
xor \U$1681 ( \3777 , \3772 , \3776 );
xor \U$1682 ( \3778 , \3768 , \3777 );
xor \U$1683 ( \3779 , \3761 , \3778 );
xor \U$1684 ( \3780 , \3716 , \3779 );
and \U$1685 ( \3781 , \3638 , \3671 );
and \U$1686 ( \3782 , \3671 , \3707 );
and \U$1687 ( \3783 , \3638 , \3707 );
or \U$1688 ( \3784 , \3781 , \3782 , \3783 );
nor \U$1689 ( \3785 , \3780 , \3784 );
nor \U$1690 ( \3786 , \3710 , \3785 );
nand \U$1691 ( \3787 , \3634 , \3786 );
and \U$1692 ( \3788 , \3718 , \3760 );
and \U$1693 ( \3789 , \3760 , \3778 );
and \U$1694 ( \3790 , \3718 , \3778 );
or \U$1695 ( \3791 , \3788 , \3789 , \3790 );
and \U$1696 ( \3792 , \3751 , \3755 );
and \U$1697 ( \3793 , \3755 , \3758 );
and \U$1698 ( \3794 , \3751 , \3758 );
or \U$1699 ( \3795 , \3792 , \3793 , \3794 );
and \U$1701 ( \3796 , \3731 , \3746 );
or \U$1703 ( \3797 , 1'b0 , \3796 , 1'b0 );
xor \U$1704 ( \3798 , \3795 , \3797 );
and \U$1705 ( \3799 , \2910 , \3133 );
and \U$1706 ( \3800 , \2866 , \3131 );
nor \U$1707 ( \3801 , \3799 , \3800 );
xnor \U$1708 ( \3802 , \3801 , \3159 );
and \U$1709 ( \3803 , \3003 , \2834 );
and \U$1710 ( \3804 , \3036 , \2832 );
nor \U$1711 ( \3805 , \3803 , \3804 );
xnor \U$1712 ( \3806 , \3805 , \2839 );
xor \U$1713 ( \3807 , \3802 , \3806 );
and \U$1714 ( \3808 , \3063 , \2769 );
and \U$1715 ( \3809 , \3096 , \2767 );
nor \U$1716 ( \3810 , \3808 , \3809 );
xnor \U$1717 ( \3811 , \3810 , \2536 );
xor \U$1718 ( \3812 , \3807 , \3811 );
xor \U$1719 ( \3813 , \3798 , \3812 );
xor \U$1720 ( \3814 , \3791 , \3813 );
and \U$1721 ( \3815 , \3765 , \3767 );
and \U$1722 ( \3816 , \3767 , \3777 );
and \U$1723 ( \3817 , \3765 , \3777 );
or \U$1724 ( \3818 , \3815 , \3816 , \3817 );
and \U$1725 ( \3819 , \3747 , \3759 );
xor \U$1726 ( \3820 , \3818 , \3819 );
not \U$1727 ( \3821 , \2973 );
and \U$1728 ( \3822 , \2659 , \3015 );
and \U$1729 ( \3823 , \2728 , \3013 );
nor \U$1730 ( \3824 , \3822 , \3823 );
xnor \U$1731 ( \3825 , \3824 , \3041 );
xor \U$1732 ( \3826 , \3821 , \3825 );
and \U$1733 ( \3827 , \2887 , \3075 );
and \U$1734 ( \3828 , \2755 , \3073 );
nor \U$1735 ( \3829 , \3827 , \3828 );
xnor \U$1736 ( \3830 , \3829 , \3101 );
xor \U$1737 ( \3831 , \3826 , \3830 );
and \U$1739 ( \3832 , \3125 , \2707 );
and \U$1740 ( \3833 , \3154 , \2705 );
nor \U$1741 ( \3834 , \3832 , \3833 );
xnor \U$1742 ( \3835 , \3834 , \2733 );
and \U$1744 ( \3836 , \3201 , \2760 );
nor \U$1745 ( \3837 , 1'b0 , \3836 );
xnor \U$1746 ( \3838 , \3837 , 1'b0 );
xor \U$1747 ( \3839 , \3835 , \3838 );
xor \U$1749 ( \3840 , \3839 , 1'b0 );
xor \U$1750 ( \3841 , 1'b1 , \3840 );
xor \U$1751 ( \3842 , \3831 , \3841 );
and \U$1753 ( \3843 , \3771 , \3776 );
or \U$1755 ( \3844 , 1'b0 , \3843 , 1'b0 );
and \U$1756 ( \3845 , \3736 , \3740 );
and \U$1757 ( \3846 , \3740 , \3745 );
and \U$1758 ( \3847 , \3736 , \3745 );
or \U$1759 ( \3848 , \3845 , \3846 , \3847 );
xor \U$1760 ( \3849 , \3844 , \3848 );
and \U$1761 ( \3850 , \3722 , \3726 );
and \U$1762 ( \3851 , \3726 , \3730 );
and \U$1763 ( \3852 , \3722 , \3730 );
or \U$1764 ( \3853 , \3850 , \3851 , \3852 );
xor \U$1765 ( \3854 , \3849 , \3853 );
xor \U$1766 ( \3855 , \3842 , \3854 );
xor \U$1767 ( \3856 , \3820 , \3855 );
xor \U$1768 ( \3857 , \3814 , \3856 );
and \U$1769 ( \3858 , \3714 , \3715 );
and \U$1770 ( \3859 , \3715 , \3779 );
and \U$1771 ( \3860 , \3714 , \3779 );
or \U$1772 ( \3861 , \3858 , \3859 , \3860 );
nor \U$1773 ( \3862 , \3857 , \3861 );
and \U$1774 ( \3863 , \3818 , \3819 );
and \U$1775 ( \3864 , \3819 , \3855 );
and \U$1776 ( \3865 , \3818 , \3855 );
or \U$1777 ( \3866 , \3863 , \3864 , \3865 );
and \U$1778 ( \3867 , \3821 , \3825 );
and \U$1779 ( \3868 , \3825 , \3830 );
and \U$1780 ( \3869 , \3821 , \3830 );
or \U$1781 ( \3870 , \3867 , \3868 , \3869 );
and \U$1782 ( \3871 , \3802 , \3806 );
and \U$1783 ( \3872 , \3806 , \3811 );
and \U$1784 ( \3873 , \3802 , \3811 );
or \U$1785 ( \3874 , \3871 , \3872 , \3873 );
xor \U$1786 ( \3875 , \3870 , \3874 );
and \U$1787 ( \3876 , \3835 , \3838 );
or \U$1790 ( \3877 , \3876 , 1'b0 , 1'b0 );
xor \U$1791 ( \3878 , \3875 , \3877 );
and \U$1792 ( \3879 , \3844 , \3848 );
and \U$1793 ( \3880 , \3848 , \3853 );
and \U$1794 ( \3881 , \3844 , \3853 );
or \U$1795 ( \3882 , \3879 , \3880 , \3881 );
and \U$1798 ( \3883 , 1'b1 , \3840 );
or \U$1800 ( \3884 , 1'b0 , \3883 , 1'b0 );
xor \U$1801 ( \3885 , \3882 , \3884 );
and \U$1802 ( \3886 , \3154 , \2707 );
and \U$1803 ( \3887 , \3063 , \2705 );
nor \U$1804 ( \3888 , \3886 , \3887 );
xnor \U$1805 ( \3889 , \3888 , \2733 );
and \U$1807 ( \3890 , \3125 , \2760 );
nor \U$1808 ( \3891 , 1'b0 , \3890 );
xnor \U$1809 ( \3892 , \3891 , 1'b0 );
xor \U$1810 ( \3893 , \3889 , \3892 );
xor \U$1812 ( \3894 , \3893 , 1'b0 );
and \U$1813 ( \3895 , \2866 , \3133 );
and \U$1814 ( \3896 , \2887 , \3131 );
nor \U$1815 ( \3897 , \3895 , \3896 );
xnor \U$1816 ( \3898 , \3897 , \3159 );
and \U$1817 ( \3899 , \3036 , \2834 );
and \U$1818 ( \3900 , \2910 , \2832 );
nor \U$1819 ( \3901 , \3899 , \3900 );
xnor \U$1820 ( \3902 , \3901 , \2839 );
xor \U$1821 ( \3903 , \3898 , \3902 );
and \U$1822 ( \3904 , \3096 , \2769 );
and \U$1823 ( \3905 , \3003 , \2767 );
nor \U$1824 ( \3906 , \3904 , \3905 );
xnor \U$1825 ( \3907 , \3906 , \2536 );
xor \U$1826 ( \3908 , \3903 , \3907 );
xor \U$1827 ( \3909 , \3894 , \3908 );
and \U$1829 ( \3910 , \2728 , \3015 );
not \U$1830 ( \3911 , \3910 );
xnor \U$1831 ( \3912 , \3911 , \3041 );
xor \U$1832 ( \3913 , 1'b0 , \3912 );
and \U$1833 ( \3914 , \2755 , \3075 );
and \U$1834 ( \3915 , \2659 , \3073 );
nor \U$1835 ( \3916 , \3914 , \3915 );
xnor \U$1836 ( \3917 , \3916 , \3101 );
xor \U$1837 ( \3918 , \3913 , \3917 );
xor \U$1838 ( \3919 , \3909 , \3918 );
xor \U$1839 ( \3920 , \3885 , \3919 );
xor \U$1840 ( \3921 , \3878 , \3920 );
xor \U$1841 ( \3922 , \3866 , \3921 );
and \U$1842 ( \3923 , \3795 , \3797 );
and \U$1843 ( \3924 , \3797 , \3812 );
and \U$1844 ( \3925 , \3795 , \3812 );
or \U$1845 ( \3926 , \3923 , \3924 , \3925 );
and \U$1846 ( \3927 , \3831 , \3841 );
and \U$1847 ( \3928 , \3841 , \3854 );
and \U$1848 ( \3929 , \3831 , \3854 );
or \U$1849 ( \3930 , \3927 , \3928 , \3929 );
xor \U$1850 ( \3931 , \3926 , \3930 );
xor \U$1852 ( \3932 , \3931 , 1'b1 );
xor \U$1853 ( \3933 , \3922 , \3932 );
and \U$1854 ( \3934 , \3791 , \3813 );
and \U$1855 ( \3935 , \3813 , \3856 );
and \U$1856 ( \3936 , \3791 , \3856 );
or \U$1857 ( \3937 , \3934 , \3935 , \3936 );
nor \U$1858 ( \3938 , \3933 , \3937 );
nor \U$1859 ( \3939 , \3862 , \3938 );
and \U$1860 ( \3940 , \3926 , \3930 );
and \U$1861 ( \3941 , \3930 , 1'b1 );
and \U$1862 ( \3942 , \3926 , 1'b1 );
or \U$1863 ( \3943 , \3940 , \3941 , \3942 );
and \U$1864 ( \3944 , \3878 , \3920 );
xor \U$1865 ( \3945 , \3943 , \3944 );
and \U$1866 ( \3946 , \3882 , \3884 );
and \U$1867 ( \3947 , \3884 , \3919 );
and \U$1868 ( \3948 , \3882 , \3919 );
or \U$1869 ( \3949 , \3946 , \3947 , \3948 );
and \U$1871 ( \3950 , \3154 , \2760 );
nor \U$1872 ( \3951 , 1'b0 , \3950 );
xnor \U$1873 ( \3952 , \3951 , 1'b0 );
xor \U$1875 ( \3953 , \3952 , 1'b0 );
xor \U$1877 ( \3954 , \3953 , 1'b0 );
and \U$1878 ( \3955 , \2910 , \2834 );
and \U$1879 ( \3956 , \2866 , \2832 );
nor \U$1880 ( \3957 , \3955 , \3956 );
xnor \U$1881 ( \3958 , \3957 , \2839 );
and \U$1882 ( \3959 , \3003 , \2769 );
and \U$1883 ( \3960 , \3036 , \2767 );
nor \U$1884 ( \3961 , \3959 , \3960 );
xnor \U$1885 ( \3962 , \3961 , \2536 );
xor \U$1886 ( \3963 , \3958 , \3962 );
and \U$1887 ( \3964 , \3063 , \2707 );
and \U$1888 ( \3965 , \3096 , \2705 );
nor \U$1889 ( \3966 , \3964 , \3965 );
xnor \U$1890 ( \3967 , \3966 , \2733 );
xor \U$1891 ( \3968 , \3963 , \3967 );
xor \U$1892 ( \3969 , \3954 , \3968 );
not \U$1893 ( \3970 , \3041 );
and \U$1894 ( \3971 , \2659 , \3075 );
and \U$1895 ( \3972 , \2728 , \3073 );
nor \U$1896 ( \3973 , \3971 , \3972 );
xnor \U$1897 ( \3974 , \3973 , \3101 );
xor \U$1898 ( \3975 , \3970 , \3974 );
and \U$1899 ( \3976 , \2887 , \3133 );
and \U$1900 ( \3977 , \2755 , \3131 );
nor \U$1901 ( \3978 , \3976 , \3977 );
xnor \U$1902 ( \3979 , \3978 , \3159 );
xor \U$1903 ( \3980 , \3975 , \3979 );
xor \U$1904 ( \3981 , \3969 , \3980 );
xor \U$1906 ( \3982 , \3981 , 1'b0 );
and \U$1908 ( \3983 , \3912 , \3917 );
or \U$1910 ( \3984 , 1'b0 , \3983 , 1'b0 );
and \U$1911 ( \3985 , \3898 , \3902 );
and \U$1912 ( \3986 , \3902 , \3907 );
and \U$1913 ( \3987 , \3898 , \3907 );
or \U$1914 ( \3988 , \3985 , \3986 , \3987 );
xor \U$1915 ( \3989 , \3984 , \3988 );
and \U$1916 ( \3990 , \3889 , \3892 );
or \U$1919 ( \3991 , \3990 , 1'b0 , 1'b0 );
xor \U$1920 ( \3992 , \3989 , \3991 );
xor \U$1921 ( \3993 , \3982 , \3992 );
xor \U$1922 ( \3994 , \3949 , \3993 );
and \U$1923 ( \3995 , \3870 , \3874 );
and \U$1924 ( \3996 , \3874 , \3877 );
and \U$1925 ( \3997 , \3870 , \3877 );
or \U$1926 ( \3998 , \3995 , \3996 , \3997 );
xor \U$1928 ( \3999 , \3998 , 1'b0 );
and \U$1929 ( \4000 , \3894 , \3908 );
and \U$1930 ( \4001 , \3908 , \3918 );
and \U$1931 ( \4002 , \3894 , \3918 );
or \U$1932 ( \4003 , \4000 , \4001 , \4002 );
xor \U$1933 ( \4004 , \3999 , \4003 );
xor \U$1934 ( \4005 , \3994 , \4004 );
xor \U$1935 ( \4006 , \3945 , \4005 );
and \U$1936 ( \4007 , \3866 , \3921 );
and \U$1937 ( \4008 , \3921 , \3932 );
and \U$1938 ( \4009 , \3866 , \3932 );
or \U$1939 ( \4010 , \4007 , \4008 , \4009 );
nor \U$1940 ( \4011 , \4006 , \4010 );
and \U$1941 ( \4012 , \3949 , \3993 );
and \U$1942 ( \4013 , \3993 , \4004 );
and \U$1943 ( \4014 , \3949 , \4004 );
or \U$1944 ( \4015 , \4012 , \4013 , \4014 );
and \U$1945 ( \4016 , \3984 , \3988 );
and \U$1946 ( \4017 , \3988 , \3991 );
and \U$1947 ( \4018 , \3984 , \3991 );
or \U$1948 ( \4019 , \4016 , \4017 , \4018 );
xor \U$1950 ( \4020 , \4019 , 1'b0 );
and \U$1951 ( \4021 , \3954 , \3968 );
and \U$1952 ( \4022 , \3968 , \3980 );
and \U$1953 ( \4023 , \3954 , \3980 );
or \U$1954 ( \4024 , \4021 , \4022 , \4023 );
xor \U$1955 ( \4025 , \4020 , \4024 );
xor \U$1956 ( \4026 , \4015 , \4025 );
and \U$1959 ( \4027 , \3998 , \4003 );
or \U$1960 ( \4028 , 1'b0 , 1'b0 , \4027 );
and \U$1963 ( \4029 , \3981 , \3992 );
or \U$1964 ( \4030 , 1'b0 , 1'b0 , \4029 );
xor \U$1965 ( \4031 , \4028 , \4030 );
and \U$1966 ( \4032 , \2866 , \2834 );
and \U$1967 ( \4033 , \2887 , \2832 );
nor \U$1968 ( \4034 , \4032 , \4033 );
xnor \U$1969 ( \4035 , \4034 , \2839 );
and \U$1970 ( \4036 , \3036 , \2769 );
and \U$1971 ( \4037 , \2910 , \2767 );
nor \U$1972 ( \4038 , \4036 , \4037 );
xnor \U$1973 ( \4039 , \4038 , \2536 );
xor \U$1974 ( \4040 , \4035 , \4039 );
and \U$1975 ( \4041 , \3096 , \2707 );
and \U$1976 ( \4042 , \3003 , \2705 );
nor \U$1977 ( \4043 , \4041 , \4042 );
xnor \U$1978 ( \4044 , \4043 , \2733 );
xor \U$1979 ( \4045 , \4040 , \4044 );
and \U$1981 ( \4046 , \2728 , \3075 );
not \U$1982 ( \4047 , \4046 );
xnor \U$1983 ( \4048 , \4047 , \3101 );
xor \U$1984 ( \4049 , 1'b0 , \4048 );
and \U$1985 ( \4050 , \2755 , \3133 );
and \U$1986 ( \4051 , \2659 , \3131 );
nor \U$1987 ( \4052 , \4050 , \4051 );
xnor \U$1988 ( \4053 , \4052 , \3159 );
xor \U$1989 ( \4054 , \4049 , \4053 );
xor \U$1990 ( \4055 , \4045 , \4054 );
and \U$1993 ( \4056 , \3063 , \2760 );
nor \U$1994 ( \4057 , 1'b0 , \4056 );
xnor \U$1995 ( \4058 , \4057 , 1'b0 );
xor \U$1997 ( \4059 , \4058 , 1'b0 );
xor \U$1999 ( \4060 , \4059 , 1'b0 );
xnor \U$2000 ( \4061 , 1'b0 , \4060 );
xor \U$2001 ( \4062 , \4055 , \4061 );
and \U$2002 ( \4063 , \3970 , \3974 );
and \U$2003 ( \4064 , \3974 , \3979 );
and \U$2004 ( \4065 , \3970 , \3979 );
or \U$2005 ( \4066 , \4063 , \4064 , \4065 );
and \U$2006 ( \4067 , \3958 , \3962 );
and \U$2007 ( \4068 , \3962 , \3967 );
and \U$2008 ( \4069 , \3958 , \3967 );
or \U$2009 ( \4070 , \4067 , \4068 , \4069 );
xor \U$2010 ( \4071 , \4066 , \4070 );
xor \U$2012 ( \4072 , \4071 , 1'b0 );
xor \U$2013 ( \4073 , \4062 , \4072 );
xor \U$2014 ( \4074 , \4031 , \4073 );
xor \U$2015 ( \4075 , \4026 , \4074 );
and \U$2016 ( \4076 , \3943 , \3944 );
and \U$2017 ( \4077 , \3944 , \4005 );
and \U$2018 ( \4078 , \3943 , \4005 );
or \U$2019 ( \4079 , \4076 , \4077 , \4078 );
nor \U$2020 ( \4080 , \4075 , \4079 );
nor \U$2021 ( \4081 , \4011 , \4080 );
nand \U$2022 ( \4082 , \3939 , \4081 );
nor \U$2023 ( \4083 , \3787 , \4082 );
and \U$2024 ( \4084 , \4028 , \4030 );
and \U$2025 ( \4085 , \4030 , \4073 );
and \U$2026 ( \4086 , \4028 , \4073 );
or \U$2027 ( \4087 , \4084 , \4085 , \4086 );
and \U$2028 ( \4088 , \4066 , \4070 );
or \U$2031 ( \4089 , \4088 , 1'b0 , 1'b0 );
or \U$2032 ( \4090 , 1'b0 , \4060 );
xor \U$2033 ( \4091 , \4089 , \4090 );
and \U$2034 ( \4092 , \4045 , \4054 );
xor \U$2035 ( \4093 , \4091 , \4092 );
xor \U$2036 ( \4094 , \4087 , \4093 );
and \U$2039 ( \4095 , \4019 , \4024 );
or \U$2040 ( \4096 , 1'b0 , 1'b0 , \4095 );
and \U$2041 ( \4097 , \4055 , \4061 );
and \U$2042 ( \4098 , \4061 , \4072 );
and \U$2043 ( \4099 , \4055 , \4072 );
or \U$2044 ( \4100 , \4097 , \4098 , \4099 );
xor \U$2045 ( \4101 , \4096 , \4100 );
and \U$2047 ( \4102 , \2910 , \2769 );
and \U$2048 ( \4103 , \2866 , \2767 );
nor \U$2049 ( \4104 , \4102 , \4103 );
xnor \U$2050 ( \4105 , \4104 , \2536 );
and \U$2051 ( \4106 , \3003 , \2707 );
and \U$2052 ( \4107 , \3036 , \2705 );
nor \U$2053 ( \4108 , \4106 , \4107 );
xnor \U$2054 ( \4109 , \4108 , \2733 );
xor \U$2055 ( \4110 , \4105 , \4109 );
and \U$2057 ( \4111 , \3096 , \2760 );
nor \U$2058 ( \4112 , 1'b0 , \4111 );
xnor \U$2059 ( \4113 , \4112 , 1'b0 );
xor \U$2060 ( \4114 , \4110 , \4113 );
xor \U$2061 ( \4115 , 1'b0 , \4114 );
not \U$2062 ( \4116 , \3101 );
and \U$2063 ( \4117 , \2659 , \3133 );
and \U$2064 ( \4118 , \2728 , \3131 );
nor \U$2065 ( \4119 , \4117 , \4118 );
xnor \U$2066 ( \4120 , \4119 , \3159 );
xor \U$2067 ( \4121 , \4116 , \4120 );
and \U$2068 ( \4122 , \2887 , \2834 );
and \U$2069 ( \4123 , \2755 , \2832 );
nor \U$2070 ( \4124 , \4122 , \4123 );
xnor \U$2071 ( \4125 , \4124 , \2839 );
xor \U$2072 ( \4126 , \4121 , \4125 );
xor \U$2073 ( \4127 , \4115 , \4126 );
xor \U$2075 ( \4128 , \4127 , 1'b0 );
and \U$2077 ( \4129 , \4048 , \4053 );
or \U$2079 ( \4130 , 1'b0 , \4129 , 1'b0 );
and \U$2080 ( \4131 , \4035 , \4039 );
and \U$2081 ( \4132 , \4039 , \4044 );
and \U$2082 ( \4133 , \4035 , \4044 );
or \U$2083 ( \4134 , \4131 , \4132 , \4133 );
xor \U$2084 ( \4135 , \4130 , \4134 );
xor \U$2086 ( \4136 , \4135 , 1'b0 );
xor \U$2087 ( \4137 , \4128 , \4136 );
xor \U$2088 ( \4138 , \4101 , \4137 );
xor \U$2089 ( \4139 , \4094 , \4138 );
and \U$2090 ( \4140 , \4015 , \4025 );
and \U$2091 ( \4141 , \4025 , \4074 );
and \U$2092 ( \4142 , \4015 , \4074 );
or \U$2093 ( \4143 , \4140 , \4141 , \4142 );
nor \U$2094 ( \4144 , \4139 , \4143 );
and \U$2095 ( \4145 , \4096 , \4100 );
and \U$2096 ( \4146 , \4100 , \4137 );
and \U$2097 ( \4147 , \4096 , \4137 );
or \U$2098 ( \4148 , \4145 , \4146 , \4147 );
and \U$2099 ( \4149 , \4130 , \4134 );
or \U$2102 ( \4150 , \4149 , 1'b0 , 1'b0 );
xor \U$2104 ( \4151 , \4150 , 1'b0 );
and \U$2106 ( \4152 , \4114 , \4126 );
or \U$2108 ( \4153 , 1'b0 , \4152 , 1'b0 );
xor \U$2109 ( \4154 , \4151 , \4153 );
xor \U$2110 ( \4155 , \4148 , \4154 );
and \U$2111 ( \4156 , \4089 , \4090 );
and \U$2112 ( \4157 , \4090 , \4092 );
and \U$2113 ( \4158 , \4089 , \4092 );
or \U$2114 ( \4159 , \4156 , \4157 , \4158 );
and \U$2117 ( \4160 , \4127 , \4136 );
or \U$2118 ( \4161 , 1'b0 , 1'b0 , \4160 );
xor \U$2119 ( \4162 , \4159 , \4161 );
and \U$2120 ( \4163 , \2866 , \2769 );
and \U$2121 ( \4164 , \2887 , \2767 );
nor \U$2122 ( \4165 , \4163 , \4164 );
xnor \U$2123 ( \4166 , \4165 , \2536 );
and \U$2124 ( \4167 , \3036 , \2707 );
and \U$2125 ( \4168 , \2910 , \2705 );
nor \U$2126 ( \4169 , \4167 , \4168 );
xnor \U$2127 ( \4170 , \4169 , \2733 );
xor \U$2128 ( \4171 , \4166 , \4170 );
and \U$2130 ( \4172 , \3003 , \2760 );
nor \U$2131 ( \4173 , 1'b0 , \4172 );
xnor \U$2132 ( \4174 , \4173 , 1'b0 );
xor \U$2133 ( \4175 , \4171 , \4174 );
and \U$2135 ( \4176 , \2728 , \3133 );
not \U$2136 ( \4177 , \4176 );
xnor \U$2137 ( \4178 , \4177 , \3159 );
xor \U$2138 ( \4179 , 1'b0 , \4178 );
and \U$2139 ( \4180 , \2755 , \2834 );
and \U$2140 ( \4181 , \2659 , \2832 );
nor \U$2141 ( \4182 , \4180 , \4181 );
xnor \U$2142 ( \4183 , \4182 , \2839 );
xor \U$2143 ( \4184 , \4179 , \4183 );
xor \U$2144 ( \4185 , \4175 , \4184 );
xor \U$2146 ( \4186 , \4185 , 1'b1 );
and \U$2147 ( \4187 , \4116 , \4120 );
and \U$2148 ( \4188 , \4120 , \4125 );
and \U$2149 ( \4189 , \4116 , \4125 );
or \U$2150 ( \4190 , \4187 , \4188 , \4189 );
and \U$2151 ( \4191 , \4105 , \4109 );
and \U$2152 ( \4192 , \4109 , \4113 );
and \U$2153 ( \4193 , \4105 , \4113 );
or \U$2154 ( \4194 , \4191 , \4192 , \4193 );
xor \U$2155 ( \4195 , \4190 , \4194 );
xor \U$2157 ( \4196 , \4195 , 1'b0 );
xor \U$2158 ( \4197 , \4186 , \4196 );
xor \U$2159 ( \4198 , \4162 , \4197 );
xor \U$2160 ( \4199 , \4155 , \4198 );
and \U$2161 ( \4200 , \4087 , \4093 );
and \U$2162 ( \4201 , \4093 , \4138 );
and \U$2163 ( \4202 , \4087 , \4138 );
or \U$2164 ( \4203 , \4200 , \4201 , \4202 );
nor \U$2165 ( \4204 , \4199 , \4203 );
nor \U$2166 ( \4205 , \4144 , \4204 );
and \U$2167 ( \4206 , \4159 , \4161 );
and \U$2168 ( \4207 , \4161 , \4197 );
and \U$2169 ( \4208 , \4159 , \4197 );
or \U$2170 ( \4209 , \4206 , \4207 , \4208 );
and \U$2171 ( \4210 , \4190 , \4194 );
or \U$2174 ( \4211 , \4210 , 1'b0 , 1'b0 );
xor \U$2176 ( \4212 , \4211 , 1'b0 );
and \U$2177 ( \4213 , \4175 , \4184 );
xor \U$2178 ( \4214 , \4212 , \4213 );
xor \U$2179 ( \4215 , \4209 , \4214 );
and \U$2182 ( \4216 , \4150 , \4153 );
or \U$2183 ( \4217 , 1'b0 , 1'b0 , \4216 );
and \U$2184 ( \4218 , \4185 , 1'b1 );
and \U$2185 ( \4219 , 1'b1 , \4196 );
and \U$2186 ( \4220 , \4185 , \4196 );
or \U$2187 ( \4221 , \4218 , \4219 , \4220 );
xor \U$2188 ( \4222 , \4217 , \4221 );
and \U$2190 ( \4223 , \2910 , \2707 );
and \U$2191 ( \4224 , \2866 , \2705 );
nor \U$2192 ( \4225 , \4223 , \4224 );
xnor \U$2193 ( \4226 , \4225 , \2733 );
and \U$2195 ( \4227 , \3036 , \2760 );
nor \U$2196 ( \4228 , 1'b0 , \4227 );
xnor \U$2197 ( \4229 , \4228 , 1'b0 );
xor \U$2198 ( \4230 , \4226 , \4229 );
xor \U$2200 ( \4231 , \4230 , 1'b0 );
xor \U$2201 ( \4232 , 1'b0 , \4231 );
not \U$2202 ( \4233 , \3159 );
and \U$2203 ( \4234 , \2659 , \2834 );
and \U$2204 ( \4235 , \2728 , \2832 );
nor \U$2205 ( \4236 , \4234 , \4235 );
xnor \U$2206 ( \4237 , \4236 , \2839 );
xor \U$2207 ( \4238 , \4233 , \4237 );
and \U$2208 ( \4239 , \2887 , \2769 );
and \U$2209 ( \4240 , \2755 , \2767 );
nor \U$2210 ( \4241 , \4239 , \4240 );
xnor \U$2211 ( \4242 , \4241 , \2536 );
xor \U$2212 ( \4243 , \4238 , \4242 );
xor \U$2213 ( \4244 , \4232 , \4243 );
xor \U$2215 ( \4245 , \4244 , 1'b0 );
and \U$2217 ( \4246 , \4178 , \4183 );
or \U$2219 ( \4247 , 1'b0 , \4246 , 1'b0 );
and \U$2220 ( \4248 , \4166 , \4170 );
and \U$2221 ( \4249 , \4170 , \4174 );
and \U$2222 ( \4250 , \4166 , \4174 );
or \U$2223 ( \4251 , \4248 , \4249 , \4250 );
xor \U$2224 ( \4252 , \4247 , \4251 );
xor \U$2226 ( \4253 , \4252 , 1'b0 );
xor \U$2227 ( \4254 , \4245 , \4253 );
xor \U$2228 ( \4255 , \4222 , \4254 );
xor \U$2229 ( \4256 , \4215 , \4255 );
and \U$2230 ( \4257 , \4148 , \4154 );
and \U$2231 ( \4258 , \4154 , \4198 );
and \U$2232 ( \4259 , \4148 , \4198 );
or \U$2233 ( \4260 , \4257 , \4258 , \4259 );
nor \U$2234 ( \4261 , \4256 , \4260 );
and \U$2235 ( \4262 , \4217 , \4221 );
and \U$2236 ( \4263 , \4221 , \4254 );
and \U$2237 ( \4264 , \4217 , \4254 );
or \U$2238 ( \4265 , \4262 , \4263 , \4264 );
and \U$2239 ( \4266 , \4247 , \4251 );
or \U$2242 ( \4267 , \4266 , 1'b0 , 1'b0 );
xor \U$2244 ( \4268 , \4267 , 1'b0 );
and \U$2246 ( \4269 , \4231 , \4243 );
or \U$2248 ( \4270 , 1'b0 , \4269 , 1'b0 );
xor \U$2249 ( \4271 , \4268 , \4270 );
xor \U$2250 ( \4272 , \4265 , \4271 );
and \U$2253 ( \4273 , \4211 , \4213 );
or \U$2254 ( \4274 , 1'b0 , 1'b0 , \4273 );
and \U$2257 ( \4275 , \4244 , \4253 );
or \U$2258 ( \4276 , 1'b0 , 1'b0 , \4275 );
xor \U$2259 ( \4277 , \4274 , \4276 );
xor \U$2260 ( \4278 , \2890 , \2913 );
xor \U$2262 ( \4279 , \4278 , 1'b0 );
xor \U$2264 ( \4280 , 1'b0 , \2840 );
xor \U$2265 ( \4281 , \4280 , \2844 );
xor \U$2266 ( \4282 , \4279 , \4281 );
xor \U$2268 ( \4283 , \4282 , 1'b1 );
and \U$2269 ( \4284 , \4233 , \4237 );
and \U$2270 ( \4285 , \4237 , \4242 );
and \U$2271 ( \4286 , \4233 , \4242 );
or \U$2272 ( \4287 , \4284 , \4285 , \4286 );
and \U$2273 ( \4288 , \4226 , \4229 );
or \U$2276 ( \4289 , \4288 , 1'b0 , 1'b0 );
xor \U$2277 ( \4290 , \4287 , \4289 );
xor \U$2279 ( \4291 , \4290 , 1'b0 );
xor \U$2280 ( \4292 , \4283 , \4291 );
xor \U$2281 ( \4293 , \4277 , \4292 );
xor \U$2282 ( \4294 , \4272 , \4293 );
and \U$2283 ( \4295 , \4209 , \4214 );
and \U$2284 ( \4296 , \4214 , \4255 );
and \U$2285 ( \4297 , \4209 , \4255 );
or \U$2286 ( \4298 , \4295 , \4296 , \4297 );
nor \U$2287 ( \4299 , \4294 , \4298 );
nor \U$2288 ( \4300 , \4261 , \4299 );
nand \U$2289 ( \4301 , \4205 , \4300 );
and \U$2290 ( \4302 , \4274 , \4276 );
and \U$2291 ( \4303 , \4276 , \4292 );
and \U$2292 ( \4304 , \4274 , \4292 );
or \U$2293 ( \4305 , \4302 , \4303 , \4304 );
and \U$2294 ( \4306 , \4287 , \4289 );
or \U$2297 ( \4307 , \4306 , 1'b0 , 1'b0 );
xor \U$2299 ( \4308 , \4307 , 1'b0 );
and \U$2300 ( \4309 , \4279 , \4281 );
xor \U$2301 ( \4310 , \4308 , \4309 );
xor \U$2302 ( \4311 , \4305 , \4310 );
and \U$2305 ( \4312 , \4267 , \4270 );
or \U$2306 ( \4313 , 1'b0 , 1'b0 , \4312 );
and \U$2307 ( \4314 , \4282 , 1'b1 );
and \U$2308 ( \4315 , 1'b1 , \4291 );
and \U$2309 ( \4316 , \4282 , \4291 );
or \U$2310 ( \4317 , \4314 , \4315 , \4316 );
xor \U$2311 ( \4318 , \4313 , \4317 );
xor \U$2313 ( \4319 , 1'b0 , \2922 );
xor \U$2314 ( \4320 , \4319 , \2933 );
xor \U$2316 ( \4321 , \4320 , 1'b0 );
xor \U$2317 ( \4322 , \2846 , \2915 );
xor \U$2319 ( \4323 , \4322 , 1'b0 );
xor \U$2320 ( \4324 , \4321 , \4323 );
xor \U$2321 ( \4325 , \4318 , \4324 );
xor \U$2322 ( \4326 , \4311 , \4325 );
and \U$2323 ( \4327 , \4265 , \4271 );
and \U$2324 ( \4328 , \4271 , \4293 );
and \U$2325 ( \4329 , \4265 , \4293 );
or \U$2326 ( \4330 , \4327 , \4328 , \4329 );
nor \U$2327 ( \4331 , \4326 , \4330 );
and \U$2328 ( \4332 , \4313 , \4317 );
and \U$2329 ( \4333 , \4317 , \4324 );
and \U$2330 ( \4334 , \4313 , \4324 );
or \U$2331 ( \4335 , \4332 , \4333 , \4334 );
xor \U$2333 ( \4336 , \2917 , 1'b0 );
xor \U$2334 ( \4337 , \4336 , \2935 );
xor \U$2335 ( \4338 , \4335 , \4337 );
and \U$2338 ( \4339 , \4307 , \4309 );
or \U$2339 ( \4340 , 1'b0 , 1'b0 , \4339 );
and \U$2342 ( \4341 , \4320 , \4323 );
or \U$2343 ( \4342 , 1'b0 , 1'b0 , \4341 );
xor \U$2344 ( \4343 , \4340 , \4342 );
xor \U$2345 ( \4344 , \2945 , 1'b1 );
xor \U$2346 ( \4345 , \4344 , \2952 );
xor \U$2347 ( \4346 , \4343 , \4345 );
xor \U$2348 ( \4347 , \4338 , \4346 );
and \U$2349 ( \4348 , \4305 , \4310 );
and \U$2350 ( \4349 , \4310 , \4325 );
and \U$2351 ( \4350 , \4305 , \4325 );
or \U$2352 ( \4351 , \4348 , \4349 , \4350 );
nor \U$2353 ( \4352 , \4347 , \4351 );
nor \U$2354 ( \4353 , \4331 , \4352 );
and \U$2355 ( \4354 , \4340 , \4342 );
and \U$2356 ( \4355 , \4342 , \4345 );
and \U$2357 ( \4356 , \4340 , \4345 );
or \U$2358 ( \4357 , \4354 , \4355 , \4356 );
and \U$2360 ( \4358 , \2942 , \2944 );
xor \U$2361 ( \4359 , 1'b0 , \4358 );
xor \U$2362 ( \4360 , \4357 , \4359 );
xor \U$2363 ( \4361 , \2937 , \2955 );
xor \U$2364 ( \4362 , \4361 , \2958 );
xor \U$2365 ( \4363 , \4360 , \4362 );
and \U$2366 ( \4364 , \4335 , \4337 );
and \U$2367 ( \4365 , \4337 , \4346 );
and \U$2368 ( \4366 , \4335 , \4346 );
or \U$2369 ( \4367 , \4364 , \4365 , \4366 );
nor \U$2370 ( \4368 , \4363 , \4367 );
xor \U$2372 ( \4369 , \2961 , 1'b0 );
xor \U$2373 ( \4370 , \4369 , \2963 );
and \U$2374 ( \4371 , \4357 , \4359 );
and \U$2375 ( \4372 , \4359 , \4362 );
and \U$2376 ( \4373 , \4357 , \4362 );
or \U$2377 ( \4374 , \4371 , \4372 , \4373 );
nor \U$2378 ( \4375 , \4370 , \4374 );
nor \U$2379 ( \4376 , \4368 , \4375 );
nand \U$2380 ( \4377 , \4353 , \4376 );
nor \U$2381 ( \4378 , \4301 , \4377 );
nand \U$2382 ( \4379 , \4083 , \4378 );
and \U$2383 ( \4380 , \3180 , \2979 );
and \U$2384 ( \4381 , \3201 , \2976 );
nor \U$2385 ( \4382 , \4380 , \4381 );
xnor \U$2386 ( \4383 , \4382 , \2973 );
and \U$2387 ( \4384 , \3225 , \3015 );
and \U$2388 ( \4385 , \3246 , \3013 );
nor \U$2389 ( \4386 , \4384 , \4385 );
xnor \U$2390 ( \4387 , \4386 , \3041 );
and \U$2391 ( \4388 , \4383 , \4387 );
and \U$2392 ( \4389 , \3273 , \3075 );
and \U$2393 ( \4390 , \3294 , \3073 );
nor \U$2394 ( \4391 , \4389 , \4390 );
xnor \U$2395 ( \4392 , \4391 , \3101 );
and \U$2396 ( \4393 , \4387 , \4392 );
and \U$2397 ( \4394 , \4383 , \4392 );
or \U$2398 ( \4395 , \4388 , \4393 , \4394 );
and \U$2399 ( \4396 , \3294 , \3075 );
and \U$2400 ( \4397 , \3225 , \3073 );
nor \U$2401 ( \4398 , \4396 , \4397 );
xnor \U$2402 ( \4399 , \4398 , \3101 );
and \U$2403 ( \4400 , \3317 , \3133 );
and \U$2404 ( \4401 , \3273 , \3131 );
nor \U$2405 ( \4402 , \4400 , \4401 );
xnor \U$2406 ( \4403 , \4402 , \3159 );
xor \U$2407 ( \4404 , \4399 , \4403 );
nand \U$2408 ( \4405 , \3450 , \2832 );
xnor \U$2409 ( \4406 , \4405 , \2839 );
xor \U$2410 ( \4407 , \4404 , \4406 );
and \U$2411 ( \4408 , \4395 , \4407 );
and \U$2412 ( \4409 , \3201 , \2979 );
and \U$2413 ( \4410 , \3125 , \2976 );
nor \U$2414 ( \4411 , \4409 , \4410 );
xnor \U$2415 ( \4412 , \4411 , \2973 );
xor \U$2416 ( \4413 , \2839 , \4412 );
and \U$2417 ( \4414 , \3246 , \3015 );
and \U$2418 ( \4415 , \3180 , \3013 );
nor \U$2419 ( \4416 , \4414 , \4415 );
xnor \U$2420 ( \4417 , \4416 , \3041 );
xor \U$2421 ( \4418 , \4413 , \4417 );
and \U$2422 ( \4419 , \4407 , \4418 );
and \U$2423 ( \4420 , \4395 , \4418 );
or \U$2424 ( \4421 , \4408 , \4419 , \4420 );
and \U$2425 ( \4422 , \3450 , \2834 );
and \U$2426 ( \4423 , \3317 , \2832 );
nor \U$2427 ( \4424 , \4422 , \4423 );
xnor \U$2428 ( \4425 , \4424 , \2839 );
and \U$2429 ( \4426 , \3125 , \2979 );
and \U$2430 ( \4427 , \3154 , \2976 );
nor \U$2431 ( \4428 , \4426 , \4427 );
xnor \U$2432 ( \4429 , \4428 , \2973 );
and \U$2433 ( \4430 , \3180 , \3015 );
and \U$2434 ( \4431 , \3201 , \3013 );
nor \U$2435 ( \4432 , \4430 , \4431 );
xnor \U$2436 ( \4433 , \4432 , \3041 );
xor \U$2437 ( \4434 , \4429 , \4433 );
and \U$2438 ( \4435 , \3225 , \3075 );
and \U$2439 ( \4436 , \3246 , \3073 );
nor \U$2440 ( \4437 , \4435 , \4436 );
xnor \U$2441 ( \4438 , \4437 , \3101 );
xor \U$2442 ( \4439 , \4434 , \4438 );
xor \U$2443 ( \4440 , \4425 , \4439 );
xor \U$2444 ( \4441 , \4421 , \4440 );
and \U$2445 ( \4442 , \2839 , \4412 );
and \U$2446 ( \4443 , \4412 , \4417 );
and \U$2447 ( \4444 , \2839 , \4417 );
or \U$2448 ( \4445 , \4442 , \4443 , \4444 );
and \U$2449 ( \4446 , \4399 , \4403 );
and \U$2450 ( \4447 , \4403 , \4406 );
and \U$2451 ( \4448 , \4399 , \4406 );
or \U$2452 ( \4449 , \4446 , \4447 , \4448 );
xor \U$2453 ( \4450 , \4445 , \4449 );
and \U$2454 ( \4451 , \3273 , \3133 );
and \U$2455 ( \4452 , \3294 , \3131 );
nor \U$2456 ( \4453 , \4451 , \4452 );
xnor \U$2457 ( \4454 , \4453 , \3159 );
xor \U$2458 ( \4455 , \4450 , \4454 );
xor \U$2459 ( \4456 , \4441 , \4455 );
and \U$2460 ( \4457 , \3246 , \2979 );
and \U$2461 ( \4458 , \3180 , \2976 );
nor \U$2462 ( \4459 , \4457 , \4458 );
xnor \U$2463 ( \4460 , \4459 , \2973 );
and \U$2464 ( \4461 , \3159 , \4460 );
and \U$2465 ( \4462 , \3294 , \3015 );
and \U$2466 ( \4463 , \3225 , \3013 );
nor \U$2467 ( \4464 , \4462 , \4463 );
xnor \U$2468 ( \4465 , \4464 , \3041 );
and \U$2469 ( \4466 , \4460 , \4465 );
and \U$2470 ( \4467 , \3159 , \4465 );
or \U$2471 ( \4468 , \4461 , \4466 , \4467 );
and \U$2472 ( \4469 , \3317 , \3075 );
and \U$2473 ( \4470 , \3273 , \3073 );
nor \U$2474 ( \4471 , \4469 , \4470 );
xnor \U$2475 ( \4472 , \4471 , \3101 );
nand \U$2476 ( \4473 , \3450 , \3131 );
xnor \U$2477 ( \4474 , \4473 , \3159 );
and \U$2478 ( \4475 , \4472 , \4474 );
and \U$2479 ( \4476 , \4468 , \4475 );
and \U$2480 ( \4477 , \3450 , \3133 );
and \U$2481 ( \4478 , \3317 , \3131 );
nor \U$2482 ( \4479 , \4477 , \4478 );
xnor \U$2483 ( \4480 , \4479 , \3159 );
and \U$2484 ( \4481 , \4475 , \4480 );
and \U$2485 ( \4482 , \4468 , \4480 );
or \U$2486 ( \4483 , \4476 , \4481 , \4482 );
xor \U$2487 ( \4484 , \4395 , \4407 );
xor \U$2488 ( \4485 , \4484 , \4418 );
and \U$2489 ( \4486 , \4483 , \4485 );
nor \U$2490 ( \4487 , \4456 , \4486 );
and \U$2491 ( \4488 , \4429 , \4433 );
and \U$2492 ( \4489 , \4433 , \4438 );
and \U$2493 ( \4490 , \4429 , \4438 );
or \U$2494 ( \4491 , \4488 , \4489 , \4490 );
nand \U$2495 ( \4492 , \3450 , \2767 );
xnor \U$2496 ( \4493 , \4492 , \2536 );
xor \U$2497 ( \4494 , \4491 , \4493 );
and \U$2498 ( \4495 , \3246 , \3075 );
and \U$2499 ( \4496 , \3180 , \3073 );
nor \U$2500 ( \4497 , \4495 , \4496 );
xnor \U$2501 ( \4498 , \4497 , \3101 );
and \U$2502 ( \4499 , \3294 , \3133 );
and \U$2503 ( \4500 , \3225 , \3131 );
nor \U$2504 ( \4501 , \4499 , \4500 );
xnor \U$2505 ( \4502 , \4501 , \3159 );
xor \U$2506 ( \4503 , \4498 , \4502 );
and \U$2507 ( \4504 , \3317 , \2834 );
and \U$2508 ( \4505 , \3273 , \2832 );
nor \U$2509 ( \4506 , \4504 , \4505 );
xnor \U$2510 ( \4507 , \4506 , \2839 );
xor \U$2511 ( \4508 , \4503 , \4507 );
xor \U$2512 ( \4509 , \4494 , \4508 );
and \U$2513 ( \4510 , \4445 , \4449 );
and \U$2514 ( \4511 , \4449 , \4454 );
and \U$2515 ( \4512 , \4445 , \4454 );
or \U$2516 ( \4513 , \4510 , \4511 , \4512 );
and \U$2517 ( \4514 , \4425 , \4439 );
xor \U$2518 ( \4515 , \4513 , \4514 );
and \U$2519 ( \4516 , \3154 , \2979 );
and \U$2520 ( \4517 , \3063 , \2976 );
nor \U$2521 ( \4518 , \4516 , \4517 );
xnor \U$2522 ( \4519 , \4518 , \2973 );
xor \U$2523 ( \4520 , \2536 , \4519 );
and \U$2524 ( \4521 , \3201 , \3015 );
and \U$2525 ( \4522 , \3125 , \3013 );
nor \U$2526 ( \4523 , \4521 , \4522 );
xnor \U$2527 ( \4524 , \4523 , \3041 );
xor \U$2528 ( \4525 , \4520 , \4524 );
xor \U$2529 ( \4526 , \4515 , \4525 );
xor \U$2530 ( \4527 , \4509 , \4526 );
and \U$2531 ( \4528 , \4421 , \4440 );
and \U$2532 ( \4529 , \4440 , \4455 );
and \U$2533 ( \4530 , \4421 , \4455 );
or \U$2534 ( \4531 , \4528 , \4529 , \4530 );
nor \U$2535 ( \4532 , \4527 , \4531 );
nor \U$2536 ( \4533 , \4487 , \4532 );
and \U$2537 ( \4534 , \4513 , \4514 );
and \U$2538 ( \4535 , \4514 , \4525 );
and \U$2539 ( \4536 , \4513 , \4525 );
or \U$2540 ( \4537 , \4534 , \4535 , \4536 );
and \U$2541 ( \4538 , \4491 , \4493 );
and \U$2542 ( \4539 , \4493 , \4508 );
and \U$2543 ( \4540 , \4491 , \4508 );
or \U$2544 ( \4541 , \4538 , \4539 , \4540 );
and \U$2545 ( \4542 , \3063 , \2979 );
and \U$2546 ( \4543 , \3096 , \2976 );
nor \U$2547 ( \4544 , \4542 , \4543 );
xnor \U$2548 ( \4545 , \4544 , \2973 );
and \U$2549 ( \4546 , \3125 , \3015 );
and \U$2550 ( \4547 , \3154 , \3013 );
nor \U$2551 ( \4548 , \4546 , \4547 );
xnor \U$2552 ( \4549 , \4548 , \3041 );
xor \U$2553 ( \4550 , \4545 , \4549 );
and \U$2554 ( \4551 , \3180 , \3075 );
and \U$2555 ( \4552 , \3201 , \3073 );
nor \U$2556 ( \4553 , \4551 , \4552 );
xnor \U$2557 ( \4554 , \4553 , \3101 );
xor \U$2558 ( \4555 , \4550 , \4554 );
xor \U$2559 ( \4556 , \4541 , \4555 );
and \U$2560 ( \4557 , \2536 , \4519 );
and \U$2561 ( \4558 , \4519 , \4524 );
and \U$2562 ( \4559 , \2536 , \4524 );
or \U$2563 ( \4560 , \4557 , \4558 , \4559 );
and \U$2564 ( \4561 , \4498 , \4502 );
and \U$2565 ( \4562 , \4502 , \4507 );
and \U$2566 ( \4563 , \4498 , \4507 );
or \U$2567 ( \4564 , \4561 , \4562 , \4563 );
xor \U$2568 ( \4565 , \4560 , \4564 );
and \U$2569 ( \4566 , \3225 , \3133 );
and \U$2570 ( \4567 , \3246 , \3131 );
nor \U$2571 ( \4568 , \4566 , \4567 );
xnor \U$2572 ( \4569 , \4568 , \3159 );
and \U$2573 ( \4570 , \3273 , \2834 );
and \U$2574 ( \4571 , \3294 , \2832 );
nor \U$2575 ( \4572 , \4570 , \4571 );
xnor \U$2576 ( \4573 , \4572 , \2839 );
xor \U$2577 ( \4574 , \4569 , \4573 );
and \U$2578 ( \4575 , \3450 , \2769 );
and \U$2579 ( \4576 , \3317 , \2767 );
nor \U$2580 ( \4577 , \4575 , \4576 );
xnor \U$2581 ( \4578 , \4577 , \2536 );
xor \U$2582 ( \4579 , \4574 , \4578 );
xor \U$2583 ( \4580 , \4565 , \4579 );
xor \U$2584 ( \4581 , \4556 , \4580 );
xor \U$2585 ( \4582 , \4537 , \4581 );
and \U$2586 ( \4583 , \4509 , \4526 );
nor \U$2587 ( \4584 , \4582 , \4583 );
and \U$2588 ( \4585 , \4541 , \4555 );
and \U$2589 ( \4586 , \4555 , \4580 );
and \U$2590 ( \4587 , \4541 , \4580 );
or \U$2591 ( \4588 , \4585 , \4586 , \4587 );
and \U$2592 ( \4589 , \4560 , \4564 );
and \U$2593 ( \4590 , \4564 , \4579 );
and \U$2594 ( \4591 , \4560 , \4579 );
or \U$2595 ( \4592 , \4589 , \4590 , \4591 );
nand \U$2596 ( \4593 , \3450 , \2705 );
xnor \U$2597 ( \4594 , \4593 , \2733 );
and \U$2598 ( \4595 , \3201 , \3075 );
and \U$2599 ( \4596 , \3125 , \3073 );
nor \U$2600 ( \4597 , \4595 , \4596 );
xnor \U$2601 ( \4598 , \4597 , \3101 );
and \U$2602 ( \4599 , \3246 , \3133 );
and \U$2603 ( \4600 , \3180 , \3131 );
nor \U$2604 ( \4601 , \4599 , \4600 );
xnor \U$2605 ( \4602 , \4601 , \3159 );
xor \U$2606 ( \4603 , \4598 , \4602 );
and \U$2607 ( \4604 , \3294 , \2834 );
and \U$2608 ( \4605 , \3225 , \2832 );
nor \U$2609 ( \4606 , \4604 , \4605 );
xnor \U$2610 ( \4607 , \4606 , \2839 );
xor \U$2611 ( \4608 , \4603 , \4607 );
xor \U$2612 ( \4609 , \4594 , \4608 );
and \U$2613 ( \4610 , \3096 , \2979 );
and \U$2614 ( \4611 , \3003 , \2976 );
nor \U$2615 ( \4612 , \4610 , \4611 );
xnor \U$2616 ( \4613 , \4612 , \2973 );
xor \U$2617 ( \4614 , \2733 , \4613 );
and \U$2618 ( \4615 , \3154 , \3015 );
and \U$2619 ( \4616 , \3063 , \3013 );
nor \U$2620 ( \4617 , \4615 , \4616 );
xnor \U$2621 ( \4618 , \4617 , \3041 );
xor \U$2622 ( \4619 , \4614 , \4618 );
xor \U$2623 ( \4620 , \4609 , \4619 );
xor \U$2624 ( \4621 , \4592 , \4620 );
and \U$2625 ( \4622 , \4545 , \4549 );
and \U$2626 ( \4623 , \4549 , \4554 );
and \U$2627 ( \4624 , \4545 , \4554 );
or \U$2628 ( \4625 , \4622 , \4623 , \4624 );
and \U$2629 ( \4626 , \4569 , \4573 );
and \U$2630 ( \4627 , \4573 , \4578 );
and \U$2631 ( \4628 , \4569 , \4578 );
or \U$2632 ( \4629 , \4626 , \4627 , \4628 );
xor \U$2633 ( \4630 , \4625 , \4629 );
and \U$2634 ( \4631 , \3317 , \2769 );
and \U$2635 ( \4632 , \3273 , \2767 );
nor \U$2636 ( \4633 , \4631 , \4632 );
xnor \U$2637 ( \4634 , \4633 , \2536 );
xor \U$2638 ( \4635 , \4630 , \4634 );
xor \U$2639 ( \4636 , \4621 , \4635 );
xor \U$2640 ( \4637 , \4588 , \4636 );
and \U$2641 ( \4638 , \4537 , \4581 );
nor \U$2642 ( \4639 , \4637 , \4638 );
nor \U$2643 ( \4640 , \4584 , \4639 );
nand \U$2644 ( \4641 , \4533 , \4640 );
and \U$2645 ( \4642 , \4592 , \4620 );
and \U$2646 ( \4643 , \4620 , \4635 );
and \U$2647 ( \4644 , \4592 , \4635 );
or \U$2648 ( \4645 , \4642 , \4643 , \4644 );
xor \U$2649 ( \4646 , \3505 , \3509 );
xor \U$2650 ( \4647 , \4646 , \3514 );
and \U$2651 ( \4648 , \2733 , \4613 );
and \U$2652 ( \4649 , \4613 , \4618 );
and \U$2653 ( \4650 , \2733 , \4618 );
or \U$2654 ( \4651 , \4648 , \4649 , \4650 );
and \U$2655 ( \4652 , \4598 , \4602 );
and \U$2656 ( \4653 , \4602 , \4607 );
and \U$2657 ( \4654 , \4598 , \4607 );
or \U$2658 ( \4655 , \4652 , \4653 , \4654 );
xor \U$2659 ( \4656 , \4651 , \4655 );
and \U$2660 ( \4657 , \3450 , \2707 );
and \U$2661 ( \4658 , \3317 , \2705 );
nor \U$2662 ( \4659 , \4657 , \4658 );
xnor \U$2663 ( \4660 , \4659 , \2733 );
xor \U$2664 ( \4661 , \4656 , \4660 );
xor \U$2665 ( \4662 , \4647 , \4661 );
xor \U$2666 ( \4663 , \4645 , \4662 );
and \U$2667 ( \4664 , \4625 , \4629 );
and \U$2668 ( \4665 , \4629 , \4634 );
and \U$2669 ( \4666 , \4625 , \4634 );
or \U$2670 ( \4667 , \4664 , \4665 , \4666 );
and \U$2671 ( \4668 , \4594 , \4608 );
and \U$2672 ( \4669 , \4608 , \4619 );
and \U$2673 ( \4670 , \4594 , \4619 );
or \U$2674 ( \4671 , \4668 , \4669 , \4670 );
xor \U$2675 ( \4672 , \4667 , \4671 );
xor \U$2676 ( \4673 , \3521 , \3525 );
xor \U$2677 ( \4674 , \4673 , \3530 );
xor \U$2678 ( \4675 , \4672 , \4674 );
xor \U$2679 ( \4676 , \4663 , \4675 );
and \U$2680 ( \4677 , \4588 , \4636 );
nor \U$2681 ( \4678 , \4676 , \4677 );
and \U$2682 ( \4679 , \4667 , \4671 );
and \U$2683 ( \4680 , \4671 , \4674 );
and \U$2684 ( \4681 , \4667 , \4674 );
or \U$2685 ( \4682 , \4679 , \4680 , \4681 );
and \U$2686 ( \4683 , \4647 , \4661 );
xor \U$2687 ( \4684 , \4682 , \4683 );
and \U$2688 ( \4685 , \4651 , \4655 );
and \U$2689 ( \4686 , \4655 , \4660 );
and \U$2690 ( \4687 , \4651 , \4660 );
or \U$2691 ( \4688 , \4685 , \4686 , \4687 );
xor \U$2692 ( \4689 , \3541 , \3543 );
xor \U$2693 ( \4690 , \4688 , \4689 );
xor \U$2694 ( \4691 , \3517 , \3533 );
xor \U$2695 ( \4692 , \4691 , \3536 );
xor \U$2696 ( \4693 , \4690 , \4692 );
xor \U$2697 ( \4694 , \4684 , \4693 );
and \U$2698 ( \4695 , \4645 , \4662 );
and \U$2699 ( \4696 , \4662 , \4675 );
and \U$2700 ( \4697 , \4645 , \4675 );
or \U$2701 ( \4698 , \4695 , \4696 , \4697 );
nor \U$2702 ( \4699 , \4694 , \4698 );
nor \U$2703 ( \4700 , \4678 , \4699 );
and \U$2704 ( \4701 , \4688 , \4689 );
and \U$2705 ( \4702 , \4689 , \4692 );
and \U$2706 ( \4703 , \4688 , \4692 );
or \U$2707 ( \4704 , \4701 , \4702 , \4703 );
xor \U$2708 ( \4705 , \3404 , \3420 );
xor \U$2709 ( \4706 , \4705 , \3455 );
xor \U$2710 ( \4707 , \4704 , \4706 );
xor \U$2711 ( \4708 , \3539 , \3544 );
xor \U$2712 ( \4709 , \4708 , \3547 );
xor \U$2713 ( \4710 , \4707 , \4709 );
and \U$2714 ( \4711 , \4682 , \4683 );
and \U$2715 ( \4712 , \4683 , \4693 );
and \U$2716 ( \4713 , \4682 , \4693 );
or \U$2717 ( \4714 , \4711 , \4712 , \4713 );
nor \U$2718 ( \4715 , \4710 , \4714 );
xor \U$2719 ( \4716 , \3550 , \3551 );
xor \U$2720 ( \4717 , \4716 , \3554 );
and \U$2721 ( \4718 , \4704 , \4706 );
and \U$2722 ( \4719 , \4706 , \4709 );
and \U$2723 ( \4720 , \4704 , \4709 );
or \U$2724 ( \4721 , \4718 , \4719 , \4720 );
nor \U$2725 ( \4722 , \4717 , \4721 );
nor \U$2726 ( \4723 , \4715 , \4722 );
nand \U$2727 ( \4724 , \4700 , \4723 );
nor \U$2728 ( \4725 , \4641 , \4724 );
and \U$2729 ( \4726 , \3294 , \2979 );
and \U$2730 ( \4727 , \3225 , \2976 );
nor \U$2731 ( \4728 , \4726 , \4727 );
xnor \U$2732 ( \4729 , \4728 , \2973 );
and \U$2733 ( \4730 , \3101 , \4729 );
and \U$2734 ( \4731 , \3317 , \3015 );
and \U$2735 ( \4732 , \3273 , \3013 );
nor \U$2736 ( \4733 , \4731 , \4732 );
xnor \U$2737 ( \4734 , \4733 , \3041 );
and \U$2738 ( \4735 , \4729 , \4734 );
and \U$2739 ( \4736 , \3101 , \4734 );
or \U$2740 ( \4737 , \4730 , \4735 , \4736 );
and \U$2741 ( \4738 , \3225 , \2979 );
and \U$2742 ( \4739 , \3246 , \2976 );
nor \U$2743 ( \4740 , \4738 , \4739 );
xnor \U$2744 ( \4741 , \4740 , \2973 );
and \U$2745 ( \4742 , \3273 , \3015 );
and \U$2746 ( \4743 , \3294 , \3013 );
nor \U$2747 ( \4744 , \4742 , \4743 );
xnor \U$2748 ( \4745 , \4744 , \3041 );
xor \U$2749 ( \4746 , \4741 , \4745 );
and \U$2750 ( \4747 , \3450 , \3075 );
and \U$2751 ( \4748 , \3317 , \3073 );
nor \U$2752 ( \4749 , \4747 , \4748 );
xnor \U$2753 ( \4750 , \4749 , \3101 );
xor \U$2754 ( \4751 , \4746 , \4750 );
xor \U$2755 ( \4752 , \4737 , \4751 );
nand \U$2756 ( \4753 , \3450 , \3073 );
xnor \U$2757 ( \4754 , \4753 , \3101 );
xor \U$2758 ( \4755 , \3101 , \4729 );
xor \U$2759 ( \4756 , \4755 , \4734 );
and \U$2760 ( \4757 , \4754 , \4756 );
nor \U$2761 ( \4758 , \4752 , \4757 );
and \U$2762 ( \4759 , \4741 , \4745 );
and \U$2763 ( \4760 , \4745 , \4750 );
and \U$2764 ( \4761 , \4741 , \4750 );
or \U$2765 ( \4762 , \4759 , \4760 , \4761 );
xor \U$2766 ( \4763 , \4472 , \4474 );
xor \U$2767 ( \4764 , \4762 , \4763 );
xor \U$2768 ( \4765 , \3159 , \4460 );
xor \U$2769 ( \4766 , \4765 , \4465 );
xor \U$2770 ( \4767 , \4764 , \4766 );
and \U$2771 ( \4768 , \4737 , \4751 );
nor \U$2772 ( \4769 , \4767 , \4768 );
nor \U$2773 ( \4770 , \4758 , \4769 );
xor \U$2774 ( \4771 , \4383 , \4387 );
xor \U$2775 ( \4772 , \4771 , \4392 );
xor \U$2776 ( \4773 , \4468 , \4475 );
xor \U$2777 ( \4774 , \4773 , \4480 );
xor \U$2778 ( \4775 , \4772 , \4774 );
and \U$2779 ( \4776 , \4762 , \4763 );
and \U$2780 ( \4777 , \4763 , \4766 );
and \U$2781 ( \4778 , \4762 , \4766 );
or \U$2782 ( \4779 , \4776 , \4777 , \4778 );
nor \U$2783 ( \4780 , \4775 , \4779 );
xor \U$2784 ( \4781 , \4483 , \4485 );
and \U$2785 ( \4782 , \4772 , \4774 );
nor \U$2786 ( \4783 , \4781 , \4782 );
nor \U$2787 ( \4784 , \4780 , \4783 );
nand \U$2788 ( \4785 , \4770 , \4784 );
and \U$2789 ( \4786 , \3273 , \2979 );
and \U$2790 ( \4787 , \3294 , \2976 );
nor \U$2791 ( \4788 , \4786 , \4787 );
xnor \U$2792 ( \4789 , \4788 , \2973 );
and \U$2793 ( \4790 , \3450 , \3015 );
and \U$2794 ( \4791 , \3317 , \3013 );
nor \U$2795 ( \4792 , \4790 , \4791 );
xnor \U$2796 ( \4793 , \4792 , \3041 );
xor \U$2797 ( \4794 , \4789 , \4793 );
and \U$2798 ( \4795 , \3317 , \2979 );
and \U$2799 ( \4796 , \3273 , \2976 );
nor \U$2800 ( \4797 , \4795 , \4796 );
xnor \U$2801 ( \4798 , \4797 , \2973 );
and \U$2802 ( \4799 , \4798 , \3041 );
nor \U$2803 ( \4800 , \4794 , \4799 );
xor \U$2804 ( \4801 , \4754 , \4756 );
and \U$2805 ( \4802 , \4789 , \4793 );
nor \U$2806 ( \4803 , \4801 , \4802 );
nor \U$2807 ( \4804 , \4800 , \4803 );
xor \U$2808 ( \4805 , \4798 , \3041 );
nand \U$2809 ( \4806 , \3450 , \3013 );
xnor \U$2810 ( \4807 , \4806 , \3041 );
nor \U$2811 ( \4808 , \4805 , \4807 );
and \U$2812 ( \4809 , \3450 , \2979 );
and \U$2813 ( \4810 , \3317 , \2976 );
nor \U$2814 ( \4811 , \4809 , \4810 );
xnor \U$2815 ( \4812 , \4811 , \2973 );
nand \U$2816 ( \4813 , \3450 , \2976 );
xnor \U$2817 ( \4814 , \4813 , \2973 );
and \U$2818 ( \4815 , \4814 , \2973 );
nand \U$2819 ( \4816 , \4812 , \4815 );
or \U$2820 ( \4817 , \4808 , \4816 );
nand \U$2821 ( \4818 , \4805 , \4807 );
nand \U$2822 ( \4819 , \4817 , \4818 );
and \U$2823 ( \4820 , \4804 , \4819 );
nand \U$2824 ( \4821 , \4794 , \4799 );
or \U$2825 ( \4822 , \4803 , \4821 );
nand \U$2826 ( \4823 , \4801 , \4802 );
nand \U$2827 ( \4824 , \4822 , \4823 );
nor \U$2828 ( \4825 , \4820 , \4824 );
or \U$2829 ( \4826 , \4785 , \4825 );
nand \U$2830 ( \4827 , \4752 , \4757 );
or \U$2831 ( \4828 , \4769 , \4827 );
nand \U$2832 ( \4829 , \4767 , \4768 );
nand \U$2833 ( \4830 , \4828 , \4829 );
and \U$2834 ( \4831 , \4784 , \4830 );
nand \U$2835 ( \4832 , \4775 , \4779 );
or \U$2836 ( \4833 , \4783 , \4832 );
nand \U$2837 ( \4834 , \4781 , \4782 );
nand \U$2838 ( \4835 , \4833 , \4834 );
nor \U$2839 ( \4836 , \4831 , \4835 );
nand \U$2840 ( \4837 , \4826 , \4836 );
and \U$2841 ( \4838 , \4725 , \4837 );
nand \U$2842 ( \4839 , \4456 , \4486 );
or \U$2843 ( \4840 , \4532 , \4839 );
nand \U$2844 ( \4841 , \4527 , \4531 );
nand \U$2845 ( \4842 , \4840 , \4841 );
and \U$2846 ( \4843 , \4640 , \4842 );
nand \U$2847 ( \4844 , \4582 , \4583 );
or \U$2848 ( \4845 , \4639 , \4844 );
nand \U$2849 ( \4846 , \4637 , \4638 );
nand \U$2850 ( \4847 , \4845 , \4846 );
nor \U$2851 ( \4848 , \4843 , \4847 );
or \U$2852 ( \4849 , \4724 , \4848 );
nand \U$2853 ( \4850 , \4676 , \4677 );
or \U$2854 ( \4851 , \4699 , \4850 );
nand \U$2855 ( \4852 , \4694 , \4698 );
nand \U$2856 ( \4853 , \4851 , \4852 );
and \U$2857 ( \4854 , \4723 , \4853 );
nand \U$2858 ( \4855 , \4710 , \4714 );
or \U$2859 ( \4856 , \4722 , \4855 );
nand \U$2860 ( \4857 , \4717 , \4721 );
nand \U$2861 ( \4858 , \4856 , \4857 );
nor \U$2862 ( \4859 , \4854 , \4858 );
nand \U$2863 ( \4860 , \4849 , \4859 );
nor \U$2864 ( \4861 , \4838 , \4860 );
or \U$2865 ( \4862 , \4379 , \4861 );
nand \U$2866 ( \4863 , \3501 , \3557 );
or \U$2867 ( \4864 , \3633 , \4863 );
nand \U$2868 ( \4865 , \3631 , \3632 );
nand \U$2869 ( \4866 , \4864 , \4865 );
and \U$2870 ( \4867 , \3786 , \4866 );
nand \U$2871 ( \4868 , \3708 , \3709 );
or \U$2872 ( \4869 , \3785 , \4868 );
nand \U$2873 ( \4870 , \3780 , \3784 );
nand \U$2874 ( \4871 , \4869 , \4870 );
nor \U$2875 ( \4872 , \4867 , \4871 );
or \U$2876 ( \4873 , \4082 , \4872 );
nand \U$2877 ( \4874 , \3857 , \3861 );
or \U$2878 ( \4875 , \3938 , \4874 );
nand \U$2879 ( \4876 , \3933 , \3937 );
nand \U$2880 ( \4877 , \4875 , \4876 );
and \U$2881 ( \4878 , \4081 , \4877 );
nand \U$2882 ( \4879 , \4006 , \4010 );
or \U$2883 ( \4880 , \4080 , \4879 );
nand \U$2884 ( \4881 , \4075 , \4079 );
nand \U$2885 ( \4882 , \4880 , \4881 );
nor \U$2886 ( \4883 , \4878 , \4882 );
nand \U$2887 ( \4884 , \4873 , \4883 );
and \U$2888 ( \4885 , \4378 , \4884 );
nand \U$2889 ( \4886 , \4139 , \4143 );
or \U$2890 ( \4887 , \4204 , \4886 );
nand \U$2891 ( \4888 , \4199 , \4203 );
nand \U$2892 ( \4889 , \4887 , \4888 );
and \U$2893 ( \4890 , \4300 , \4889 );
nand \U$2894 ( \4891 , \4256 , \4260 );
or \U$2895 ( \4892 , \4299 , \4891 );
nand \U$2896 ( \4893 , \4294 , \4298 );
nand \U$2897 ( \4894 , \4892 , \4893 );
nor \U$2898 ( \4895 , \4890 , \4894 );
or \U$2899 ( \4896 , \4377 , \4895 );
nand \U$2900 ( \4897 , \4326 , \4330 );
or \U$2901 ( \4898 , \4352 , \4897 );
nand \U$2902 ( \4899 , \4347 , \4351 );
nand \U$2903 ( \4900 , \4898 , \4899 );
and \U$2904 ( \4901 , \4376 , \4900 );
nand \U$2905 ( \4902 , \4363 , \4367 );
or \U$2906 ( \4903 , \4375 , \4902 );
nand \U$2907 ( \4904 , \4370 , \4374 );
nand \U$2908 ( \4905 , \4903 , \4904 );
nor \U$2909 ( \4906 , \4901 , \4905 );
nand \U$2910 ( \4907 , \4896 , \4906 );
nor \U$2911 ( \4908 , \4885 , \4907 );
nand \U$2912 ( \4909 , \4862 , \4908 );
not \U$2913 ( \4910 , \4909 );
xor \U$2914 ( \4911 , \2969 , \4910 );
buf g3284_GF_PartitionCandidate( \4912_nG3284 , \4911 );
buf \U$2919 ( \4913 , RI994e3e8_15);
buf \U$2920 ( \4914 , RI994e370_16);
buf \U$2921 ( \4915 , RI994e2f8_17);
buf \U$2922 ( \4916 , RI994e280_18);
buf \U$2923 ( \4917 , RI994e208_19);
buf \U$2924 ( \4918 , RI994e190_20);
buf \U$2925 ( \4919 , RI994e118_21);
buf \U$2926 ( \4920 , RI994e0a0_22);
buf \U$2927 ( \4921 , RI994e028_23);
buf \U$2928 ( \4922 , RI994dfb0_24);
buf \U$2929 ( \4923 , RI994df38_25);
and \U$2930 ( \4924 , \4922 , \4923 );
and \U$2931 ( \4925 , \4921 , \4924 );
and \U$2932 ( \4926 , \4920 , \4925 );
and \U$2933 ( \4927 , \4919 , \4926 );
and \U$2934 ( \4928 , \4918 , \4927 );
and \U$2935 ( \4929 , \4917 , \4928 );
and \U$2936 ( \4930 , \4916 , \4929 );
and \U$2937 ( \4931 , \4915 , \4930 );
and \U$2938 ( \4932 , \4914 , \4931 );
xor \U$2939 ( \4933 , \4913 , \4932 );
buf \U$2940 ( \4934 , \4933 );
buf \U$2941 ( \4935 , \4934 );
buf \U$2942 ( \4936 , RI9921730_613);
buf \U$2943 ( \4937 , RI9921910_609);
buf \U$2944 ( \4938 , RI9921988_608);
buf \U$2945 ( \4939 , RI9921a00_607);
buf \U$2946 ( \4940 , RI9921a78_606);
buf \U$2947 ( \4941 , RI9921af0_605);
buf \U$2948 ( \4942 , RI9921b68_604);
buf \U$2949 ( \4943 , RI9921be0_603);
buf \U$2950 ( \4944 , RI9921c58_602);
buf \U$2951 ( \4945 , RI9921cd0_601);
buf \U$2952 ( \4946 , RI9921730_613);
buf \U$2953 ( \4947 , RI99217a8_612);
buf \U$2954 ( \4948 , RI9921820_611);
buf \U$2955 ( \4949 , RI9921898_610);
and \U$2956 ( \4950 , \4946 , \4947 , \4948 , \4949 );
nor \U$2957 ( \4951 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4950 );
buf \U$2958 ( \4952 , \4951 );
buf \U$2959 ( \4953 , \4952 );
xor \U$2960 ( \4954 , \4936 , \4953 );
buf \U$2961 ( \4955 , \4954 );
buf \U$2962 ( \4956 , RI99217a8_612);
and \U$2963 ( \4957 , \4936 , \4953 );
xor \U$2964 ( \4958 , \4956 , \4957 );
buf \U$2965 ( \4959 , \4958 );
buf \U$2966 ( \4960 , RI9921820_611);
and \U$2967 ( \4961 , \4956 , \4957 );
xor \U$2968 ( \4962 , \4960 , \4961 );
buf \U$2969 ( \4963 , \4962 );
buf \U$2970 ( \4964 , RI9921898_610);
and \U$2971 ( \4965 , \4960 , \4961 );
xor \U$2972 ( \4966 , \4964 , \4965 );
buf \U$2973 ( \4967 , \4966 );
buf \U$2974 ( \4968 , RI9921910_609);
and \U$2975 ( \4969 , \4964 , \4965 );
xor \U$2976 ( \4970 , \4968 , \4969 );
buf \U$2977 ( \4971 , \4970 );
not \U$2978 ( \4972 , \4971 );
buf \U$2979 ( \4973 , RI9921988_608);
and \U$2980 ( \4974 , \4968 , \4969 );
xor \U$2981 ( \4975 , \4973 , \4974 );
buf \U$2982 ( \4976 , \4975 );
buf \U$2983 ( \4977 , RI9921a00_607);
and \U$2984 ( \4978 , \4973 , \4974 );
xor \U$2985 ( \4979 , \4977 , \4978 );
buf \U$2986 ( \4980 , \4979 );
buf \U$2987 ( \4981 , RI9921a78_606);
and \U$2988 ( \4982 , \4977 , \4978 );
xor \U$2989 ( \4983 , \4981 , \4982 );
buf \U$2990 ( \4984 , \4983 );
buf \U$2991 ( \4985 , RI9921af0_605);
and \U$2992 ( \4986 , \4981 , \4982 );
xor \U$2993 ( \4987 , \4985 , \4986 );
buf \U$2994 ( \4988 , \4987 );
buf \U$2995 ( \4989 , RI9921b68_604);
and \U$2996 ( \4990 , \4985 , \4986 );
xor \U$2997 ( \4991 , \4989 , \4990 );
buf \U$2998 ( \4992 , \4991 );
buf \U$2999 ( \4993 , RI9921be0_603);
and \U$3000 ( \4994 , \4989 , \4990 );
xor \U$3001 ( \4995 , \4993 , \4994 );
buf \U$3002 ( \4996 , \4995 );
buf \U$3003 ( \4997 , RI9921c58_602);
and \U$3004 ( \4998 , \4993 , \4994 );
xor \U$3005 ( \4999 , \4997 , \4998 );
buf \U$3006 ( \5000 , \4999 );
buf \U$3007 ( \5001 , RI9921cd0_601);
and \U$3008 ( \5002 , \4997 , \4998 );
xor \U$3009 ( \5003 , \5001 , \5002 );
buf \U$3010 ( \5004 , \5003 );
nor \U$3011 ( \5005 , \4955 , \4959 , \4963 , \4967 , \4972 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3012 ( \5006 , RI995e450_236, \5005 );
not \U$3013 ( \5007 , \4955 );
not \U$3014 ( \5008 , \4959 );
not \U$3015 ( \5009 , \4963 );
not \U$3016 ( \5010 , \4967 );
nor \U$3017 ( \5011 , \5007 , \5008 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3018 ( \5012 , RI9967078_223, \5011 );
nor \U$3019 ( \5013 , \4955 , \5008 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3020 ( \5014 , RI9967690_210, \5013 );
nor \U$3021 ( \5015 , \5007 , \4959 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3022 ( \5016 , RI890fba0_197, \5015 );
nor \U$3023 ( \5017 , \4955 , \4959 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3024 ( \5018 , RI8918b88_184, \5017 );
nor \U$3025 ( \5019 , \5007 , \5008 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3026 ( \5020 , RI89253b0_171, \5019 );
nor \U$3027 ( \5021 , \4955 , \5008 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3028 ( \5022 , RI8930dc8_158, \5021 );
nor \U$3029 ( \5023 , \5007 , \4959 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3030 ( \5024 , RI8939db0_145, \5023 );
nor \U$3031 ( \5025 , \4955 , \4959 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3032 ( \5026 , RI89465d8_132, \5025 );
nor \U$3033 ( \5027 , \5007 , \5008 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3034 ( \5028 , RI89ec640_119, \5027 );
nor \U$3035 ( \5029 , \4955 , \5008 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3036 ( \5030 , RI9776f80_106, \5029 );
nor \U$3037 ( \5031 , \5007 , \4959 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3038 ( \5032 , RI9808480_93, \5031 );
nor \U$3039 ( \5033 , \4955 , \4959 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3040 ( \5034 , RI9808a98_80, \5033 );
nor \U$3041 ( \5035 , \5007 , \5008 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3042 ( \5036 , RI9819730_67, \5035 );
nor \U$3043 ( \5037 , \4955 , \5008 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3044 ( \5038 , RI98abc38_54, \5037 );
nor \U$3045 ( \5039 , \5007 , \4959 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3046 ( \5040 , RI98bc8d0_41, \5039 );
nor \U$3047 ( \5041 , \4955 , \4959 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$3048 ( \5042 , RI994ddd0_28, \5041 );
or \U$3049 ( \5043 , \5006 , \5012 , \5014 , \5016 , \5018 , \5020 , \5022 , \5024 , \5026 , \5028 , \5030 , \5032 , \5034 , \5036 , \5038 , \5040 , \5042 );
buf \U$3050 ( \5044 , \4976 );
buf \U$3051 ( \5045 , \4980 );
buf \U$3052 ( \5046 , \4984 );
buf \U$3053 ( \5047 , \4988 );
buf \U$3054 ( \5048 , \4992 );
buf \U$3055 ( \5049 , \4996 );
buf \U$3056 ( \5050 , \5000 );
buf \U$3057 ( \5051 , \5004 );
buf \U$3058 ( \5052 , \4971 );
buf \U$3059 ( \5053 , \4955 );
buf \U$3060 ( \5054 , \4959 );
buf \U$3061 ( \5055 , \4963 );
buf \U$3062 ( \5056 , \4967 );
or \U$3063 ( \5057 , \5053 , \5054 , \5055 , \5056 );
and \U$3064 ( \5058 , \5052 , \5057 );
or \U$3065 ( \5059 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5058 );
buf \U$3066 ( \5060 , \5059 );
_DC g2232 ( \5061_nG2232 , \5043 , \5060 );
buf \U$3067 ( \5062 , \5061_nG2232 );
not \U$3068 ( \5063 , \5062 );
xor \U$3069 ( \5064 , \4935 , \5063 );
xor \U$3070 ( \5065 , \4914 , \4931 );
buf \U$3071 ( \5066 , \5065 );
buf \U$3072 ( \5067 , \5066 );
and \U$3073 ( \5068 , RI995e3d8_237, \5005 );
and \U$3074 ( \5069 , RI99669e8_224, \5011 );
and \U$3075 ( \5070 , RI9967618_211, \5013 );
and \U$3076 ( \5071 , RI890fb28_198, \5015 );
and \U$3077 ( \5072 , RI8918b10_185, \5017 );
and \U$3078 ( \5073 , RI8925338_172, \5019 );
and \U$3079 ( \5074 , RI8930d50_159, \5021 );
and \U$3080 ( \5075 , RI8939d38_146, \5023 );
and \U$3081 ( \5076 , RI8946560_133, \5025 );
and \U$3082 ( \5077 , RI89ec5c8_120, \5027 );
and \U$3083 ( \5078 , RI9776f08_107, \5029 );
and \U$3084 ( \5079 , RI9808408_94, \5031 );
and \U$3085 ( \5080 , RI9808a20_81, \5033 );
and \U$3086 ( \5081 , RI98196b8_68, \5035 );
and \U$3087 ( \5082 , RI98abbc0_55, \5037 );
and \U$3088 ( \5083 , RI98bc858_42, \5039 );
and \U$3089 ( \5084 , RI994dd58_29, \5041 );
or \U$3090 ( \5085 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 );
_DC g220e ( \5086_nG220e , \5085 , \5060 );
buf \U$3091 ( \5087 , \5086_nG220e );
not \U$3092 ( \5088 , \5087 );
and \U$3093 ( \5089 , \5067 , \5088 );
xor \U$3094 ( \5090 , \4915 , \4930 );
buf \U$3095 ( \5091 , \5090 );
buf \U$3096 ( \5092 , \5091 );
and \U$3097 ( \5093 , RI9959fe0_238, \5005 );
and \U$3098 ( \5094 , RI995e978_225, \5011 );
and \U$3099 ( \5095 , RI99675a0_212, \5013 );
and \U$3100 ( \5096 , RI890fab0_199, \5015 );
and \U$3101 ( \5097 , RI8918a98_186, \5017 );
and \U$3102 ( \5098 , RI89252c0_173, \5019 );
and \U$3103 ( \5099 , RI8930cd8_160, \5021 );
and \U$3104 ( \5100 , RI8939cc0_147, \5023 );
and \U$3105 ( \5101 , RI89464e8_134, \5025 );
and \U$3106 ( \5102 , RI89ec550_121, \5027 );
and \U$3107 ( \5103 , RI9776e90_108, \5029 );
and \U$3108 ( \5104 , RI9808390_95, \5031 );
and \U$3109 ( \5105 , RI98089a8_82, \5033 );
and \U$3110 ( \5106 , RI9819640_69, \5035 );
and \U$3111 ( \5107 , RI98abb48_56, \5037 );
and \U$3112 ( \5108 , RI98bc7e0_43, \5039 );
and \U$3113 ( \5109 , RI994dce0_30, \5041 );
or \U$3114 ( \5110 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 );
_DC g207b ( \5111_nG207b , \5110 , \5060 );
buf \U$3115 ( \5112 , \5111_nG207b );
not \U$3116 ( \5113 , \5112 );
and \U$3117 ( \5114 , \5092 , \5113 );
xor \U$3118 ( \5115 , \4916 , \4929 );
buf \U$3119 ( \5116 , \5115 );
buf \U$3120 ( \5117 , \5116 );
and \U$3121 ( \5118 , RI9959f68_239, \5005 );
and \U$3122 ( \5119 , RI995e900_226, \5011 );
and \U$3123 ( \5120 , RI9967528_213, \5013 );
and \U$3124 ( \5121 , RI890fa38_200, \5015 );
and \U$3125 ( \5122 , RI8918a20_187, \5017 );
and \U$3126 ( \5123 , RI8925248_174, \5019 );
and \U$3127 ( \5124 , RI8930c60_161, \5021 );
and \U$3128 ( \5125 , RI8939c48_148, \5023 );
and \U$3129 ( \5126 , RI8946470_135, \5025 );
and \U$3130 ( \5127 , RI89ec4d8_122, \5027 );
and \U$3131 ( \5128 , RI9776e18_109, \5029 );
and \U$3132 ( \5129 , RI9808318_96, \5031 );
and \U$3133 ( \5130 , RI9808930_83, \5033 );
and \U$3134 ( \5131 , RI98195c8_70, \5035 );
and \U$3135 ( \5132 , RI98abad0_57, \5037 );
and \U$3136 ( \5133 , RI98bc768_44, \5039 );
and \U$3137 ( \5134 , RI994dc68_31, \5041 );
or \U$3138 ( \5135 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 );
_DC g2057 ( \5136_nG2057 , \5135 , \5060 );
buf \U$3139 ( \5137 , \5136_nG2057 );
not \U$3140 ( \5138 , \5137 );
and \U$3141 ( \5139 , \5117 , \5138 );
xor \U$3142 ( \5140 , \4917 , \4928 );
buf \U$3143 ( \5141 , \5140 );
buf \U$3144 ( \5142 , \5141 );
and \U$3145 ( \5143 , RI9959860_240, \5005 );
and \U$3146 ( \5144 , RI995e888_227, \5011 );
and \U$3147 ( \5145 , RI99674b0_214, \5013 );
and \U$3148 ( \5146 , RI890f9c0_201, \5015 );
and \U$3149 ( \5147 , RI89189a8_188, \5017 );
and \U$3150 ( \5148 , RI89251d0_175, \5019 );
and \U$3151 ( \5149 , RI8930be8_162, \5021 );
and \U$3152 ( \5150 , RI8939bd0_149, \5023 );
and \U$3153 ( \5151 , RI89463f8_136, \5025 );
and \U$3154 ( \5152 , RI89ec460_123, \5027 );
and \U$3155 ( \5153 , RI9776da0_110, \5029 );
and \U$3156 ( \5154 , RI98082a0_97, \5031 );
and \U$3157 ( \5155 , RI98088b8_84, \5033 );
and \U$3158 ( \5156 , RI9819550_71, \5035 );
and \U$3159 ( \5157 , RI98aba58_58, \5037 );
and \U$3160 ( \5158 , RI98bc6f0_45, \5039 );
and \U$3161 ( \5159 , RI994dbf0_32, \5041 );
or \U$3162 ( \5160 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 );
_DC g1ed8 ( \5161_nG1ed8 , \5160 , \5060 );
buf \U$3163 ( \5162 , \5161_nG1ed8 );
not \U$3164 ( \5163 , \5162 );
and \U$3165 ( \5164 , \5142 , \5163 );
xor \U$3166 ( \5165 , \4918 , \4927 );
buf \U$3167 ( \5166 , \5165 );
buf \U$3168 ( \5167 , \5166 );
and \U$3169 ( \5168 , RI994d998_241, \5005 );
and \U$3170 ( \5169 , RI995e810_228, \5011 );
and \U$3171 ( \5170 , RI9967438_215, \5013 );
and \U$3172 ( \5171 , RI890f948_202, \5015 );
and \U$3173 ( \5172 , RI8918930_189, \5017 );
and \U$3174 ( \5173 , RI8925158_176, \5019 );
and \U$3175 ( \5174 , RI8930b70_163, \5021 );
and \U$3176 ( \5175 , RI8939b58_150, \5023 );
and \U$3177 ( \5176 , RI8946380_137, \5025 );
and \U$3178 ( \5177 , RI89ec3e8_124, \5027 );
and \U$3179 ( \5178 , RI9776d28_111, \5029 );
and \U$3180 ( \5179 , RI9808228_98, \5031 );
and \U$3181 ( \5180 , RI9808840_85, \5033 );
and \U$3182 ( \5181 , RI98194d8_72, \5035 );
and \U$3183 ( \5182 , RI98ab9e0_59, \5037 );
and \U$3184 ( \5183 , RI98abff8_46, \5039 );
and \U$3185 ( \5184 , RI98bcc90_33, \5041 );
or \U$3186 ( \5185 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 );
_DC g1eb4 ( \5186_nG1eb4 , \5185 , \5060 );
buf \U$3187 ( \5187 , \5186_nG1eb4 );
not \U$3188 ( \5188 , \5187 );
and \U$3189 ( \5189 , \5167 , \5188 );
xor \U$3190 ( \5190 , \4919 , \4926 );
buf \U$3191 ( \5191 , \5190 );
buf \U$3192 ( \5192 , \5191 );
and \U$3193 ( \5193 , RI994d920_242, \5005 );
and \U$3194 ( \5194 , RI995e798_229, \5011 );
and \U$3195 ( \5195 , RI99673c0_216, \5013 );
and \U$3196 ( \5196 , RI890f8d0_203, \5015 );
and \U$3197 ( \5197 , RI89188b8_190, \5017 );
and \U$3198 ( \5198 , RI89250e0_177, \5019 );
and \U$3199 ( \5199 , RI8930af8_164, \5021 );
and \U$3200 ( \5200 , RI8939ae0_151, \5023 );
and \U$3201 ( \5201 , RI8946308_138, \5025 );
and \U$3202 ( \5202 , RI89ec370_125, \5027 );
and \U$3203 ( \5203 , RI89ec988_112, \5029 );
and \U$3204 ( \5204 , RI97772c8_99, \5031 );
and \U$3205 ( \5205 , RI98087c8_86, \5033 );
and \U$3206 ( \5206 , RI9819460_73, \5035 );
and \U$3207 ( \5207 , RI98ab968_60, \5037 );
and \U$3208 ( \5208 , RI98abf80_47, \5039 );
and \U$3209 ( \5209 , RI98bcc18_34, \5041 );
or \U$3210 ( \5210 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 );
_DC g1d69 ( \5211_nG1d69 , \5210 , \5060 );
buf \U$3211 ( \5212 , \5211_nG1d69 );
not \U$3212 ( \5213 , \5212 );
and \U$3213 ( \5214 , \5192 , \5213 );
xor \U$3214 ( \5215 , \4920 , \4925 );
buf \U$3215 ( \5216 , \5215 );
buf \U$3216 ( \5217 , \5216 );
and \U$3217 ( \5218 , RI994d8a8_243, \5005 );
and \U$3218 ( \5219 , RI995e720_230, \5011 );
and \U$3219 ( \5220 , RI9967348_217, \5013 );
and \U$3220 ( \5221 , RI890f858_204, \5015 );
and \U$3221 ( \5222 , RI8918840_191, \5017 );
and \U$3222 ( \5223 , RI8925068_178, \5019 );
and \U$3223 ( \5224 , RI8930a80_165, \5021 );
and \U$3224 ( \5225 , RI8939a68_152, \5023 );
and \U$3225 ( \5226 , RI8946290_139, \5025 );
and \U$3226 ( \5227 , RI89ec2f8_126, \5027 );
and \U$3227 ( \5228 , RI89ec910_113, \5029 );
and \U$3228 ( \5229 , RI9777250_100, \5031 );
and \U$3229 ( \5230 , RI9808750_87, \5033 );
and \U$3230 ( \5231 , RI98193e8_74, \5035 );
and \U$3231 ( \5232 , RI98ab8f0_61, \5037 );
and \U$3232 ( \5233 , RI98abf08_48, \5039 );
and \U$3233 ( \5234 , RI98bcba0_35, \5041 );
or \U$3234 ( \5235 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 );
_DC g1d45 ( \5236_nG1d45 , \5235 , \5060 );
buf \U$3235 ( \5237 , \5236_nG1d45 );
not \U$3236 ( \5238 , \5237 );
and \U$3237 ( \5239 , \5217 , \5238 );
xor \U$3238 ( \5240 , \4921 , \4924 );
buf \U$3239 ( \5241 , \5240 );
buf \U$3240 ( \5242 , \5241 );
and \U$3241 ( \5243 , RI994d830_244, \5005 );
and \U$3242 ( \5244 , RI995e6a8_231, \5011 );
and \U$3243 ( \5245 , RI99672d0_218, \5013 );
and \U$3244 ( \5246 , RI890f7e0_205, \5015 );
and \U$3245 ( \5247 , RI89187c8_192, \5017 );
and \U$3246 ( \5248 , RI8924ff0_179, \5019 );
and \U$3247 ( \5249 , RI8930a08_166, \5021 );
and \U$3248 ( \5250 , RI89399f0_153, \5023 );
and \U$3249 ( \5251 , RI8946218_140, \5025 );
and \U$3250 ( \5252 , RI89ec280_127, \5027 );
and \U$3251 ( \5253 , RI89ec898_114, \5029 );
and \U$3252 ( \5254 , RI97771d8_101, \5031 );
and \U$3253 ( \5255 , RI98086d8_88, \5033 );
and \U$3254 ( \5256 , RI9819370_75, \5035 );
and \U$3255 ( \5257 , RI98ab878_62, \5037 );
and \U$3256 ( \5258 , RI98abe90_49, \5039 );
and \U$3257 ( \5259 , RI98bcb28_36, \5041 );
or \U$3258 ( \5260 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 );
_DC g1c2a ( \5261_nG1c2a , \5260 , \5060 );
buf \U$3259 ( \5262 , \5261_nG1c2a );
not \U$3260 ( \5263 , \5262 );
and \U$3261 ( \5264 , \5242 , \5263 );
xor \U$3262 ( \5265 , \4922 , \4923 );
buf \U$3263 ( \5266 , \5265 );
buf \U$3264 ( \5267 , \5266 );
and \U$3265 ( \5268 , RI994d7b8_245, \5005 );
and \U$3266 ( \5269 , RI995e630_232, \5011 );
and \U$3267 ( \5270 , RI9967258_219, \5013 );
and \U$3268 ( \5271 , RI890f768_206, \5015 );
and \U$3269 ( \5272 , RI8918750_193, \5017 );
and \U$3270 ( \5273 , RI8924f78_180, \5019 );
and \U$3271 ( \5274 , RI8930990_167, \5021 );
and \U$3272 ( \5275 , RI8939978_154, \5023 );
and \U$3273 ( \5276 , RI89461a0_141, \5025 );
and \U$3274 ( \5277 , RI89ec208_128, \5027 );
and \U$3275 ( \5278 , RI89ec820_115, \5029 );
and \U$3276 ( \5279 , RI9777160_102, \5031 );
and \U$3277 ( \5280 , RI9808660_89, \5033 );
and \U$3278 ( \5281 , RI98192f8_76, \5035 );
and \U$3279 ( \5282 , RI98ab800_63, \5037 );
and \U$3280 ( \5283 , RI98abe18_50, \5039 );
and \U$3281 ( \5284 , RI98bcab0_37, \5041 );
or \U$3282 ( \5285 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 );
_DC g1c43 ( \5286_nG1c43 , \5285 , \5060 );
buf \U$3283 ( \5287 , \5286_nG1c43 );
not \U$3284 ( \5288 , \5287 );
and \U$3285 ( \5289 , \5267 , \5288 );
not \U$3286 ( \5290 , \4923 );
buf \U$3287 ( \5291 , \5290 );
buf \U$3288 ( \5292 , \5291 );
and \U$3289 ( \5293 , RI994d740_246, \5005 );
and \U$3290 ( \5294 , RI995e5b8_233, \5011 );
and \U$3291 ( \5295 , RI99671e0_220, \5013 );
and \U$3292 ( \5296 , RI890f6f0_207, \5015 );
and \U$3293 ( \5297 , RI89186d8_194, \5017 );
and \U$3294 ( \5298 , RI8924f00_181, \5019 );
and \U$3295 ( \5299 , RI8930918_168, \5021 );
and \U$3296 ( \5300 , RI8939900_155, \5023 );
and \U$3297 ( \5301 , RI8946128_142, \5025 );
and \U$3298 ( \5302 , RI89ec190_129, \5027 );
and \U$3299 ( \5303 , RI89ec7a8_116, \5029 );
and \U$3300 ( \5304 , RI97770e8_103, \5031 );
and \U$3301 ( \5305 , RI98085e8_90, \5033 );
and \U$3302 ( \5306 , RI9819280_77, \5035 );
and \U$3303 ( \5307 , RI98ab788_64, \5037 );
and \U$3304 ( \5308 , RI98abda0_51, \5039 );
and \U$3305 ( \5309 , RI98bca38_38, \5041 );
or \U$3306 ( \5310 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 );
_DC g1b40 ( \5311_nG1b40 , \5310 , \5060 );
buf \U$3307 ( \5312 , \5311_nG1b40 );
not \U$3308 ( \5313 , \5312 );
and \U$3309 ( \5314 , \5292 , \5313 );
buf \U$3310 ( \5315 , RI994dec0_26);
buf \U$3313 ( \5316 , \5315 );
and \U$3314 ( \5317 , RI994d6c8_247, \5005 );
and \U$3315 ( \5318 , RI995e540_234, \5011 );
and \U$3316 ( \5319 , RI9967168_221, \5013 );
and \U$3317 ( \5320 , RI890f678_208, \5015 );
and \U$3318 ( \5321 , RI8918660_195, \5017 );
and \U$3319 ( \5322 , RI8924e88_182, \5019 );
and \U$3320 ( \5323 , RI89308a0_169, \5021 );
and \U$3321 ( \5324 , RI8939888_156, \5023 );
and \U$3322 ( \5325 , RI89460b0_143, \5025 );
and \U$3323 ( \5326 , RI89ec118_130, \5027 );
and \U$3324 ( \5327 , RI89ec730_117, \5029 );
and \U$3325 ( \5328 , RI9777070_104, \5031 );
and \U$3326 ( \5329 , RI9808570_91, \5033 );
and \U$3327 ( \5330 , RI9819208_78, \5035 );
and \U$3328 ( \5331 , RI98ab710_65, \5037 );
and \U$3329 ( \5332 , RI98abd28_52, \5039 );
and \U$3330 ( \5333 , RI98bc9c0_39, \5041 );
or \U$3331 ( \5334 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 );
_DC g1b24 ( \5335_nG1b24 , \5334 , \5060 );
buf \U$3332 ( \5336 , \5335_nG1b24 );
not \U$3333 ( \5337 , \5336 );
or \U$3334 ( \5338 , \5316 , \5337 );
and \U$3335 ( \5339 , \5313 , \5338 );
and \U$3336 ( \5340 , \5292 , \5338 );
or \U$3337 ( \5341 , \5314 , \5339 , \5340 );
and \U$3338 ( \5342 , \5288 , \5341 );
and \U$3339 ( \5343 , \5267 , \5341 );
or \U$3340 ( \5344 , \5289 , \5342 , \5343 );
and \U$3341 ( \5345 , \5263 , \5344 );
and \U$3342 ( \5346 , \5242 , \5344 );
or \U$3343 ( \5347 , \5264 , \5345 , \5346 );
and \U$3344 ( \5348 , \5238 , \5347 );
and \U$3345 ( \5349 , \5217 , \5347 );
or \U$3346 ( \5350 , \5239 , \5348 , \5349 );
and \U$3347 ( \5351 , \5213 , \5350 );
and \U$3348 ( \5352 , \5192 , \5350 );
or \U$3349 ( \5353 , \5214 , \5351 , \5352 );
and \U$3350 ( \5354 , \5188 , \5353 );
and \U$3351 ( \5355 , \5167 , \5353 );
or \U$3352 ( \5356 , \5189 , \5354 , \5355 );
and \U$3353 ( \5357 , \5163 , \5356 );
and \U$3354 ( \5358 , \5142 , \5356 );
or \U$3355 ( \5359 , \5164 , \5357 , \5358 );
and \U$3356 ( \5360 , \5138 , \5359 );
and \U$3357 ( \5361 , \5117 , \5359 );
or \U$3358 ( \5362 , \5139 , \5360 , \5361 );
and \U$3359 ( \5363 , \5113 , \5362 );
and \U$3360 ( \5364 , \5092 , \5362 );
or \U$3361 ( \5365 , \5114 , \5363 , \5364 );
and \U$3362 ( \5366 , \5088 , \5365 );
and \U$3363 ( \5367 , \5067 , \5365 );
or \U$3364 ( \5368 , \5089 , \5366 , \5367 );
xor \U$3365 ( \5369 , \5064 , \5368 );
buf g223b_GF_PartitionCandidate( \5370_nG223b , \5369 );
buf \U$3366 ( \5371 , \5370_nG223b );
xor \U$3367 ( \5372 , \5067 , \5088 );
xor \U$3368 ( \5373 , \5372 , \5365 );
buf g2217_GF_PartitionCandidate( \5374_nG2217 , \5373 );
buf \U$3369 ( \5375 , \5374_nG2217 );
xor \U$3370 ( \5376 , \5092 , \5113 );
xor \U$3371 ( \5377 , \5376 , \5362 );
buf g2084_GF_PartitionCandidate( \5378_nG2084 , \5377 );
buf \U$3372 ( \5379 , \5378_nG2084 );
and \U$3373 ( \5380 , \5375 , \5379 );
not \U$3374 ( \5381 , \5380 );
and \U$3375 ( \5382 , \5371 , \5381 );
not \U$3376 ( \5383 , \5382 );
buf \U$3377 ( \5384 , \4955 );
buf \U$3378 ( \5385 , \4976 );
buf \U$3379 ( \5386 , \4980 );
buf \U$3380 ( \5387 , \4984 );
buf \U$3381 ( \5388 , \4988 );
buf \U$3382 ( \5389 , \4992 );
buf \U$3383 ( \5390 , \4996 );
buf \U$3384 ( \5391 , \5000 );
buf \U$3385 ( \5392 , \5004 );
buf \U$3386 ( \5393 , \4971 );
nor \U$3387 ( \5394 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 );
buf \U$3388 ( \5395 , \5394 );
buf \U$3389 ( \5396 , \5395 );
xor \U$3390 ( \5397 , \5384 , \5396 );
buf \U$3391 ( \5398 , \5397 );
buf \U$3392 ( \5399 , \4959 );
and \U$3393 ( \5400 , \5384 , \5396 );
xor \U$3394 ( \5401 , \5399 , \5400 );
buf \U$3395 ( \5402 , \5401 );
buf \U$3396 ( \5403 , \4963 );
and \U$3397 ( \5404 , \5399 , \5400 );
xor \U$3398 ( \5405 , \5403 , \5404 );
buf \U$3399 ( \5406 , \5405 );
buf \U$3400 ( \5407 , \4967 );
and \U$3401 ( \5408 , \5403 , \5404 );
xor \U$3402 ( \5409 , \5407 , \5408 );
buf \U$3403 ( \5410 , \5409 );
buf \U$3404 ( \5411 , \4971 );
and \U$3405 ( \5412 , \5407 , \5408 );
xor \U$3406 ( \5413 , \5411 , \5412 );
buf \U$3407 ( \5414 , \5413 );
not \U$3408 ( \5415 , \5414 );
buf \U$3409 ( \5416 , \4976 );
and \U$3410 ( \5417 , \5411 , \5412 );
xor \U$3411 ( \5418 , \5416 , \5417 );
buf \U$3412 ( \5419 , \5418 );
buf \U$3413 ( \5420 , \4980 );
and \U$3414 ( \5421 , \5416 , \5417 );
xor \U$3415 ( \5422 , \5420 , \5421 );
buf \U$3416 ( \5423 , \5422 );
buf \U$3417 ( \5424 , \4984 );
and \U$3418 ( \5425 , \5420 , \5421 );
xor \U$3419 ( \5426 , \5424 , \5425 );
buf \U$3420 ( \5427 , \5426 );
buf \U$3421 ( \5428 , \4988 );
and \U$3422 ( \5429 , \5424 , \5425 );
xor \U$3423 ( \5430 , \5428 , \5429 );
buf \U$3424 ( \5431 , \5430 );
buf \U$3425 ( \5432 , \4992 );
and \U$3426 ( \5433 , \5428 , \5429 );
xor \U$3427 ( \5434 , \5432 , \5433 );
buf \U$3428 ( \5435 , \5434 );
buf \U$3429 ( \5436 , \4996 );
and \U$3430 ( \5437 , \5432 , \5433 );
xor \U$3431 ( \5438 , \5436 , \5437 );
buf \U$3432 ( \5439 , \5438 );
buf \U$3433 ( \5440 , \5000 );
and \U$3434 ( \5441 , \5436 , \5437 );
xor \U$3435 ( \5442 , \5440 , \5441 );
buf \U$3436 ( \5443 , \5442 );
buf \U$3437 ( \5444 , \5004 );
and \U$3438 ( \5445 , \5440 , \5441 );
xor \U$3439 ( \5446 , \5444 , \5445 );
buf \U$3440 ( \5447 , \5446 );
nor \U$3441 ( \5448 , \5398 , \5402 , \5406 , \5410 , \5415 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3442 ( \5449 , RI9922bd0_569, \5448 );
not \U$3443 ( \5450 , \5398 );
not \U$3444 ( \5451 , \5402 );
not \U$3445 ( \5452 , \5406 );
not \U$3446 ( \5453 , \5410 );
nor \U$3447 ( \5454 , \5450 , \5451 , \5452 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3448 ( \5455 , RI9923800_549, \5454 );
nor \U$3449 ( \5456 , \5398 , \5451 , \5452 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3450 ( \5457 , RI9924160_529, \5456 );
nor \U$3451 ( \5458 , \5450 , \5402 , \5452 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3452 ( \5459 , RI9924ac0_509, \5458 );
nor \U$3453 ( \5460 , \5398 , \5402 , \5452 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3454 ( \5461 , RI9925ab0_489, \5460 );
nor \U$3455 ( \5462 , \5450 , \5451 , \5406 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3456 ( \5463 , RI9926410_469, \5462 );
nor \U$3457 ( \5464 , \5398 , \5451 , \5406 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3458 ( \5465 , RI9926d70_449, \5464 );
nor \U$3459 ( \5466 , \5450 , \5402 , \5406 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3460 ( \5467 , RI9928120_429, \5466 );
nor \U$3461 ( \5468 , \5398 , \5402 , \5406 , \5453 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3462 ( \5469 , RI9928a80_409, \5468 );
nor \U$3463 ( \5470 , \5450 , \5451 , \5452 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3464 ( \5471 , RI992a1f0_389, \5470 );
nor \U$3465 ( \5472 , \5398 , \5451 , \5452 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3466 ( \5473 , RI992ab50_369, \5472 );
nor \U$3467 ( \5474 , \5450 , \5402 , \5452 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3468 ( \5475 , RI992b4b0_349, \5474 );
nor \U$3469 ( \5476 , \5398 , \5402 , \5452 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3470 ( \5477 , RI992cfe0_329, \5476 );
nor \U$3471 ( \5478 , \5450 , \5451 , \5406 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3472 ( \5479 , RI992eed0_309, \5478 );
nor \U$3473 ( \5480 , \5398 , \5451 , \5406 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3474 ( \5481 , RI992f830_289, \5480 );
nor \U$3475 ( \5482 , \5450 , \5402 , \5406 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3476 ( \5483 , RI9931ae0_269, \5482 );
nor \U$3477 ( \5484 , \5398 , \5402 , \5406 , \5410 , \5414 , \5419 , \5423 , \5427 , \5431 , \5435 , \5439 , \5443 , \5447 );
and \U$3478 ( \5485 , RI994d5d8_249, \5484 );
or \U$3479 ( \5486 , \5449 , \5455 , \5457 , \5459 , \5461 , \5463 , \5465 , \5467 , \5469 , \5471 , \5473 , \5475 , \5477 , \5479 , \5481 , \5483 , \5485 );
buf \U$3480 ( \5487 , \5419 );
buf \U$3481 ( \5488 , \5423 );
buf \U$3482 ( \5489 , \5427 );
buf \U$3483 ( \5490 , \5431 );
buf \U$3484 ( \5491 , \5435 );
buf \U$3485 ( \5492 , \5439 );
buf \U$3486 ( \5493 , \5443 );
buf \U$3487 ( \5494 , \5447 );
buf \U$3488 ( \5495 , \5414 );
buf \U$3489 ( \5496 , \5398 );
buf \U$3490 ( \5497 , \5402 );
buf \U$3491 ( \5498 , \5406 );
buf \U$3492 ( \5499 , \5410 );
or \U$3493 ( \5500 , \5496 , \5497 , \5498 , \5499 );
and \U$3494 ( \5501 , \5495 , \5500 );
or \U$3495 ( \5502 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5501 );
buf \U$3496 ( \5503 , \5502 );
_DC g290c ( \5504_nG290c , \5486 , \5503 );
buf \U$3497 ( \5505 , \5504_nG290c );
buf \U$3498 ( \5506 , RI994e460_14);
and \U$3499 ( \5507 , \4913 , \4932 );
and \U$3500 ( \5508 , \5506 , \5507 );
buf \U$3501 ( \5509 , \5508 );
buf \U$3502 ( \5510 , \5509 );
xor \U$3503 ( \5511 , \5506 , \5507 );
buf \U$3504 ( \5512 , \5511 );
buf \U$3505 ( \5513 , \5512 );
and \U$3506 ( \5514 , RI995e4c8_235, \5005 );
and \U$3507 ( \5515 , RI99670f0_222, \5011 );
and \U$3508 ( \5516 , RI890f600_209, \5013 );
and \U$3509 ( \5517 , RI89185e8_196, \5015 );
and \U$3510 ( \5518 , RI8924e10_183, \5017 );
and \U$3511 ( \5519 , RI8930828_170, \5019 );
and \U$3512 ( \5520 , RI8939810_157, \5021 );
and \U$3513 ( \5521 , RI8946038_144, \5023 );
and \U$3514 ( \5522 , RI89ec0a0_131, \5025 );
and \U$3515 ( \5523 , RI89ec6b8_118, \5027 );
and \U$3516 ( \5524 , RI9776ff8_105, \5029 );
and \U$3517 ( \5525 , RI98084f8_92, \5031 );
and \U$3518 ( \5526 , RI9808b10_79, \5033 );
and \U$3519 ( \5527 , RI98197a8_66, \5035 );
and \U$3520 ( \5528 , RI98abcb0_53, \5037 );
and \U$3521 ( \5529 , RI98bc948_40, \5039 );
and \U$3522 ( \5530 , RI994de48_27, \5041 );
or \U$3523 ( \5531 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 );
_DC g23ed ( \5532_nG23ed , \5531 , \5060 );
buf \U$3524 ( \5533 , \5532_nG23ed );
not \U$3525 ( \5534 , \5533 );
and \U$3526 ( \5535 , \5513 , \5534 );
and \U$3527 ( \5536 , \4935 , \5063 );
and \U$3528 ( \5537 , \5063 , \5368 );
and \U$3529 ( \5538 , \4935 , \5368 );
or \U$3530 ( \5539 , \5536 , \5537 , \5538 );
and \U$3531 ( \5540 , \5534 , \5539 );
and \U$3532 ( \5541 , \5513 , \5539 );
or \U$3533 ( \5542 , \5535 , \5540 , \5541 );
xnor \U$3534 ( \5543 , \5510 , \5542 );
buf g2402_GF_PartitionCandidate( \5544_nG2402 , \5543 );
buf \U$3535 ( \5545 , \5544_nG2402 );
xor \U$3536 ( \5546 , \5513 , \5534 );
xor \U$3537 ( \5547 , \5546 , \5539 );
buf g23f6_GF_PartitionCandidate( \5548_nG23f6 , \5547 );
buf \U$3538 ( \5549 , \5548_nG23f6 );
xor \U$3539 ( \5550 , \5545 , \5549 );
xor \U$3540 ( \5551 , \5549 , \5371 );
not \U$3541 ( \5552 , \5551 );
and \U$3542 ( \5553 , \5550 , \5552 );
and \U$3543 ( \5554 , \5505 , \5553 );
and \U$3544 ( \5555 , RI9922f18_568, \5448 );
and \U$3545 ( \5556 , RI9923878_548, \5454 );
and \U$3546 ( \5557 , RI99241d8_528, \5456 );
and \U$3547 ( \5558 , RI9924b38_508, \5458 );
and \U$3548 ( \5559 , RI9925b28_488, \5460 );
and \U$3549 ( \5560 , RI9926488_468, \5462 );
and \U$3550 ( \5561 , RI9926de8_448, \5464 );
and \U$3551 ( \5562 , RI9928198_428, \5466 );
and \U$3552 ( \5563 , RI9928af8_408, \5468 );
and \U$3553 ( \5564 , RI992a268_388, \5470 );
and \U$3554 ( \5565 , RI992abc8_368, \5472 );
and \U$3555 ( \5566 , RI992c6f8_348, \5474 );
and \U$3556 ( \5567 , RI992d058_328, \5476 );
and \U$3557 ( \5568 , RI992ef48_308, \5478 );
and \U$3558 ( \5569 , RI992f8a8_288, \5480 );
and \U$3559 ( \5570 , RI9931b58_268, \5482 );
and \U$3560 ( \5571 , RI994d650_248, \5484 );
or \U$3561 ( \5572 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 );
_DC g2a01 ( \5573_nG2a01 , \5572 , \5503 );
buf \U$3562 ( \5574 , \5573_nG2a01 );
and \U$3563 ( \5575 , \5574 , \5551 );
nor \U$3564 ( \5576 , \5554 , \5575 );
and \U$3565 ( \5577 , \5549 , \5371 );
not \U$3566 ( \5578 , \5577 );
and \U$3567 ( \5579 , \5545 , \5578 );
xnor \U$3568 ( \5580 , \5576 , \5579 );
xor \U$3569 ( \5581 , \5383 , \5580 );
and \U$3571 ( \5582 , RI9922b58_570, \5448 );
and \U$3572 ( \5583 , RI9923788_550, \5454 );
and \U$3573 ( \5584 , RI99240e8_530, \5456 );
and \U$3574 ( \5585 , RI9924a48_510, \5458 );
and \U$3575 ( \5586 , RI9925a38_490, \5460 );
and \U$3576 ( \5587 , RI9926398_470, \5462 );
and \U$3577 ( \5588 , RI9926cf8_450, \5464 );
and \U$3578 ( \5589 , RI99280a8_430, \5466 );
and \U$3579 ( \5590 , RI9928a08_410, \5468 );
and \U$3580 ( \5591 , RI992a178_390, \5470 );
and \U$3581 ( \5592 , RI992aad8_370, \5472 );
and \U$3582 ( \5593 , RI992b438_350, \5474 );
and \U$3583 ( \5594 , RI992cf68_330, \5476 );
and \U$3584 ( \5595 , RI992ee58_310, \5478 );
and \U$3585 ( \5596 , RI992f7b8_290, \5480 );
and \U$3586 ( \5597 , RI9931a68_270, \5482 );
and \U$3587 ( \5598 , RI994d560_250, \5484 );
or \U$3588 ( \5599 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 );
_DC g2843 ( \5600_nG2843 , \5599 , \5503 );
buf \U$3589 ( \5601 , \5600_nG2843 );
or \U$3590 ( \5602 , \5510 , \5542 );
not \U$3591 ( \5603 , \5602 );
buf g25dc_GF_PartitionCandidate( \5604_nG25dc , \5603 );
buf \U$3592 ( \5605 , \5604_nG25dc );
xor \U$3593 ( \5606 , \5605 , \5545 );
and \U$3594 ( \5607 , \5601 , \5606 );
nor \U$3595 ( \5608 , 1'b0 , \5607 );
xnor \U$3597 ( \5609 , \5608 , 1'b0 );
xor \U$3598 ( \5610 , \5581 , \5609 );
xor \U$3599 ( \5611 , 1'b0 , \5610 );
xor \U$3601 ( \5612 , \5371 , \5375 );
xor \U$3602 ( \5613 , \5375 , \5379 );
not \U$3603 ( \5614 , \5613 );
and \U$3604 ( \5615 , \5612 , \5614 );
and \U$3605 ( \5616 , \5574 , \5615 );
not \U$3606 ( \5617 , \5616 );
xnor \U$3607 ( \5618 , \5617 , \5382 );
and \U$3608 ( \5619 , \5601 , \5553 );
and \U$3609 ( \5620 , \5505 , \5551 );
nor \U$3610 ( \5621 , \5619 , \5620 );
xnor \U$3611 ( \5622 , \5621 , \5579 );
and \U$3612 ( \5623 , \5618 , \5622 );
or \U$3614 ( \5624 , 1'b0 , \5623 , 1'b0 );
xor \U$3616 ( \5625 , \5624 , 1'b0 );
xor \U$3618 ( \5626 , \5625 , 1'b0 );
and \U$3619 ( \5627 , \5611 , \5626 );
or \U$3620 ( \5628 , 1'b0 , 1'b0 , \5627 );
and \U$3623 ( \5629 , \5574 , \5553 );
not \U$3624 ( \5630 , \5629 );
xnor \U$3625 ( \5631 , \5630 , \5579 );
xor \U$3626 ( \5632 , 1'b0 , \5631 );
and \U$3628 ( \5633 , \5505 , \5606 );
nor \U$3629 ( \5634 , 1'b0 , \5633 );
xnor \U$3630 ( \5635 , \5634 , 1'b0 );
xor \U$3631 ( \5636 , \5632 , \5635 );
xor \U$3632 ( \5637 , 1'b0 , \5636 );
xor \U$3634 ( \5638 , \5637 , 1'b1 );
and \U$3635 ( \5639 , \5383 , \5580 );
and \U$3636 ( \5640 , \5580 , \5609 );
and \U$3637 ( \5641 , \5383 , \5609 );
or \U$3638 ( \5642 , \5639 , \5640 , \5641 );
xor \U$3640 ( \5643 , \5642 , 1'b0 );
xor \U$3642 ( \5644 , \5643 , 1'b0 );
xor \U$3643 ( \5645 , \5638 , \5644 );
and \U$3644 ( \5646 , \5628 , \5645 );
or \U$3646 ( \5647 , 1'b0 , \5646 , 1'b0 );
xor \U$3648 ( \5648 , \5647 , 1'b0 );
and \U$3650 ( \5649 , \5637 , 1'b1 );
and \U$3651 ( \5650 , 1'b1 , \5644 );
and \U$3652 ( \5651 , \5637 , \5644 );
or \U$3653 ( \5652 , \5649 , \5650 , \5651 );
xor \U$3654 ( \5653 , 1'b0 , \5652 );
not \U$3656 ( \5654 , \5579 );
and \U$3658 ( \5655 , \5574 , \5606 );
nor \U$3659 ( \5656 , 1'b0 , \5655 );
xnor \U$3660 ( \5657 , \5656 , 1'b0 );
xor \U$3661 ( \5658 , \5654 , \5657 );
xor \U$3663 ( \5659 , \5658 , 1'b0 );
xor \U$3664 ( \5660 , 1'b0 , \5659 );
xor \U$3666 ( \5661 , \5660 , 1'b0 );
and \U$3668 ( \5662 , \5631 , \5635 );
or \U$3670 ( \5663 , 1'b0 , \5662 , 1'b0 );
xor \U$3672 ( \5664 , \5663 , 1'b0 );
xor \U$3674 ( \5665 , \5664 , 1'b0 );
xor \U$3675 ( \5666 , \5661 , \5665 );
xor \U$3676 ( \5667 , \5653 , \5666 );
xor \U$3677 ( \5668 , \5648 , \5667 );
xor \U$3683 ( \5669 , \5117 , \5138 );
xor \U$3684 ( \5670 , \5669 , \5359 );
buf g2060_GF_PartitionCandidate( \5671_nG2060 , \5670 );
buf \U$3685 ( \5672 , \5671_nG2060 );
xor \U$3686 ( \5673 , \5379 , \5672 );
xor \U$3687 ( \5674 , \5142 , \5163 );
xor \U$3688 ( \5675 , \5674 , \5356 );
buf g1ee1_GF_PartitionCandidate( \5676_nG1ee1 , \5675 );
buf \U$3689 ( \5677 , \5676_nG1ee1 );
xor \U$3690 ( \5678 , \5672 , \5677 );
not \U$3691 ( \5679 , \5678 );
and \U$3692 ( \5680 , \5673 , \5679 );
and \U$3693 ( \5681 , \5574 , \5680 );
not \U$3694 ( \5682 , \5681 );
and \U$3695 ( \5683 , \5672 , \5677 );
not \U$3696 ( \5684 , \5683 );
and \U$3697 ( \5685 , \5379 , \5684 );
xnor \U$3698 ( \5686 , \5682 , \5685 );
and \U$3699 ( \5687 , \5601 , \5615 );
and \U$3700 ( \5688 , \5505 , \5613 );
nor \U$3701 ( \5689 , \5687 , \5688 );
xnor \U$3702 ( \5690 , \5689 , \5382 );
and \U$3703 ( \5691 , \5686 , \5690 );
or \U$3705 ( \5692 , 1'b0 , \5691 , 1'b0 );
and \U$3706 ( \5693 , RI9922a68_572, \5448 );
and \U$3707 ( \5694 , RI9923698_552, \5454 );
and \U$3708 ( \5695 , RI9923ff8_532, \5456 );
and \U$3709 ( \5696 , RI9924958_512, \5458 );
and \U$3710 ( \5697 , RI9925948_492, \5460 );
and \U$3711 ( \5698 , RI99262a8_472, \5462 );
and \U$3712 ( \5699 , RI9926c08_452, \5464 );
and \U$3713 ( \5700 , RI9927fb8_432, \5466 );
and \U$3714 ( \5701 , RI9928918_412, \5468 );
and \U$3715 ( \5702 , RI9929278_392, \5470 );
and \U$3716 ( \5703 , RI992a9e8_372, \5472 );
and \U$3717 ( \5704 , RI992b348_352, \5474 );
and \U$3718 ( \5705 , RI992ce78_332, \5476 );
and \U$3719 ( \5706 , RI992ed68_312, \5478 );
and \U$3720 ( \5707 , RI992f6c8_292, \5480 );
and \U$3721 ( \5708 , RI9931978_272, \5482 );
and \U$3722 ( \5709 , RI994d470_252, \5484 );
or \U$3723 ( \5710 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 );
_DC g26a4 ( \5711_nG26a4 , \5710 , \5503 );
buf \U$3724 ( \5712 , \5711_nG26a4 );
and \U$3725 ( \5713 , \5712 , \5553 );
and \U$3726 ( \5714 , RI9922ae0_571, \5448 );
and \U$3727 ( \5715 , RI9923710_551, \5454 );
and \U$3728 ( \5716 , RI9924070_531, \5456 );
and \U$3729 ( \5717 , RI99249d0_511, \5458 );
and \U$3730 ( \5718 , RI99259c0_491, \5460 );
and \U$3731 ( \5719 , RI9926320_471, \5462 );
and \U$3732 ( \5720 , RI9926c80_451, \5464 );
and \U$3733 ( \5721 , RI9928030_431, \5466 );
and \U$3734 ( \5722 , RI9928990_411, \5468 );
and \U$3735 ( \5723 , RI992a100_391, \5470 );
and \U$3736 ( \5724 , RI992aa60_371, \5472 );
and \U$3737 ( \5725 , RI992b3c0_351, \5474 );
and \U$3738 ( \5726 , RI992cef0_331, \5476 );
and \U$3739 ( \5727 , RI992ede0_311, \5478 );
and \U$3740 ( \5728 , RI992f740_291, \5480 );
and \U$3741 ( \5729 , RI99319f0_271, \5482 );
and \U$3742 ( \5730 , RI994d4e8_251, \5484 );
or \U$3743 ( \5731 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 );
_DC g2782 ( \5732_nG2782 , \5731 , \5503 );
buf \U$3744 ( \5733 , \5732_nG2782 );
and \U$3745 ( \5734 , \5733 , \5551 );
nor \U$3746 ( \5735 , \5713 , \5734 );
xnor \U$3747 ( \5736 , \5735 , \5579 );
and \U$3749 ( \5737 , RI99229f0_573, \5448 );
and \U$3750 ( \5738 , RI9923620_553, \5454 );
and \U$3751 ( \5739 , RI9923f80_533, \5456 );
and \U$3752 ( \5740 , RI99248e0_513, \5458 );
and \U$3753 ( \5741 , RI99258d0_493, \5460 );
and \U$3754 ( \5742 , RI9926230_473, \5462 );
and \U$3755 ( \5743 , RI9926b90_453, \5464 );
and \U$3756 ( \5744 , RI9927f40_433, \5466 );
and \U$3757 ( \5745 , RI99288a0_413, \5468 );
and \U$3758 ( \5746 , RI9929200_393, \5470 );
and \U$3759 ( \5747 , RI992a970_373, \5472 );
and \U$3760 ( \5748 , RI992b2d0_353, \5474 );
and \U$3761 ( \5749 , RI992ce00_333, \5476 );
and \U$3762 ( \5750 , RI992ecf0_313, \5478 );
and \U$3763 ( \5751 , RI992f650_293, \5480 );
and \U$3764 ( \5752 , RI9931900_273, \5482 );
and \U$3765 ( \5753 , RI994d3f8_253, \5484 );
or \U$3766 ( \5754 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 );
_DC g25bb ( \5755_nG25bb , \5754 , \5503 );
buf \U$3767 ( \5756 , \5755_nG25bb );
and \U$3768 ( \5757 , \5756 , \5606 );
nor \U$3769 ( \5758 , 1'b0 , \5757 );
xnor \U$3770 ( \5759 , \5758 , 1'b0 );
and \U$3771 ( \5760 , \5736 , \5759 );
or \U$3774 ( \5761 , \5760 , 1'b0 , 1'b0 );
and \U$3775 ( \5762 , \5692 , \5761 );
or \U$3778 ( \5763 , \5762 , 1'b0 , 1'b0 );
and \U$3781 ( \5764 , \5712 , \5606 );
nor \U$3782 ( \5765 , 1'b0 , \5764 );
xnor \U$3783 ( \5766 , \5765 , 1'b0 );
xor \U$3785 ( \5767 , \5766 , 1'b0 );
xor \U$3787 ( \5768 , \5767 , 1'b0 );
not \U$3788 ( \5769 , \5685 );
and \U$3789 ( \5770 , \5505 , \5615 );
and \U$3790 ( \5771 , \5574 , \5613 );
nor \U$3791 ( \5772 , \5770 , \5771 );
xnor \U$3792 ( \5773 , \5772 , \5382 );
xor \U$3793 ( \5774 , \5769 , \5773 );
and \U$3794 ( \5775 , \5733 , \5553 );
and \U$3795 ( \5776 , \5601 , \5551 );
nor \U$3796 ( \5777 , \5775 , \5776 );
xnor \U$3797 ( \5778 , \5777 , \5579 );
xor \U$3798 ( \5779 , \5774 , \5778 );
and \U$3799 ( \5780 , \5768 , \5779 );
or \U$3801 ( \5781 , 1'b0 , \5780 , 1'b0 );
and \U$3802 ( \5782 , \5763 , \5781 );
or \U$3803 ( \5783 , 1'b0 , 1'b0 , \5782 );
and \U$3805 ( \5784 , \5733 , \5606 );
nor \U$3806 ( \5785 , 1'b0 , \5784 );
xnor \U$3807 ( \5786 , \5785 , 1'b0 );
xor \U$3809 ( \5787 , \5786 , 1'b0 );
xor \U$3811 ( \5788 , \5787 , 1'b0 );
xor \U$3813 ( \5789 , 1'b0 , \5618 );
xor \U$3814 ( \5790 , \5789 , \5622 );
xor \U$3815 ( \5791 , \5788 , \5790 );
and \U$3817 ( \5792 , \5791 , 1'b1 );
and \U$3818 ( \5793 , \5769 , \5773 );
and \U$3819 ( \5794 , \5773 , \5778 );
and \U$3820 ( \5795 , \5769 , \5778 );
or \U$3821 ( \5796 , \5793 , \5794 , \5795 );
xor \U$3823 ( \5797 , \5796 , 1'b0 );
xor \U$3825 ( \5798 , \5797 , 1'b0 );
and \U$3826 ( \5799 , 1'b1 , \5798 );
and \U$3827 ( \5800 , \5791 , \5798 );
or \U$3828 ( \5801 , \5792 , \5799 , \5800 );
and \U$3829 ( \5802 , \5783 , \5801 );
xor \U$3831 ( \5803 , \5611 , 1'b0 );
xor \U$3832 ( \5804 , \5803 , \5626 );
and \U$3833 ( \5805 , \5801 , \5804 );
and \U$3834 ( \5806 , \5783 , \5804 );
or \U$3835 ( \5807 , \5802 , \5805 , \5806 );
xor \U$3837 ( \5808 , 1'b0 , \5628 );
xor \U$3838 ( \5809 , \5808 , \5645 );
and \U$3839 ( \5810 , \5807 , \5809 );
or \U$3840 ( \5811 , 1'b0 , 1'b0 , \5810 );
nand \U$3841 ( \5812 , \5668 , \5811 );
nor \U$3842 ( \5813 , \5668 , \5811 );
not \U$3843 ( \5814 , \5813 );
nand \U$3844 ( \5815 , \5812 , \5814 );
xor \U$3845 ( \5816 , \5292 , \5313 );
xor \U$3846 ( \5817 , \5816 , \5338 );
buf g1b47_GF_PartitionCandidate( \5818_nG1b47 , \5817 );
buf \U$3847 ( \5819 , \5818_nG1b47 );
xor \U$3848 ( \5820 , \5316 , \5336 );
buf g1b27_GF_PartitionCandidate( \5821_nG1b27 , \5820 );
buf \U$3849 ( \5822 , \5821_nG1b27 );
xor \U$3850 ( \5823 , \5819 , \5822 );
not \U$3851 ( \5824 , \5822 );
and \U$3852 ( \5825 , \5823 , \5824 );
and \U$3853 ( \5826 , \5756 , \5825 );
and \U$3854 ( \5827 , \5712 , \5822 );
nor \U$3855 ( \5828 , \5826 , \5827 );
xnor \U$3856 ( \5829 , \5828 , \5819 );
and \U$3857 ( \5830 , RI9922900_575, \5448 );
and \U$3858 ( \5831 , RI9923530_555, \5454 );
and \U$3859 ( \5832 , RI9923e90_535, \5456 );
and \U$3860 ( \5833 , RI99247f0_515, \5458 );
and \U$3861 ( \5834 , RI99257e0_495, \5460 );
and \U$3862 ( \5835 , RI9926140_475, \5462 );
and \U$3863 ( \5836 , RI9926aa0_455, \5464 );
and \U$3864 ( \5837 , RI9927e50_435, \5466 );
and \U$3865 ( \5838 , RI99287b0_415, \5468 );
and \U$3866 ( \5839 , RI9929110_395, \5470 );
and \U$3867 ( \5840 , RI992a880_375, \5472 );
and \U$3868 ( \5841 , RI992b1e0_355, \5474 );
and \U$3869 ( \5842 , RI992cd10_335, \5476 );
and \U$3870 ( \5843 , RI992d670_315, \5478 );
and \U$3871 ( \5844 , RI992f560_295, \5480 );
and \U$3872 ( \5845 , RI9931810_275, \5482 );
and \U$3873 ( \5846 , RI9935f50_255, \5484 );
or \U$3874 ( \5847 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 );
_DC g242a ( \5848_nG242a , \5847 , \5503 );
buf \U$3875 ( \5849 , \5848_nG242a );
xor \U$3876 ( \5850 , \5242 , \5263 );
xor \U$3877 ( \5851 , \5850 , \5344 );
buf g1c4f_GF_PartitionCandidate( \5852_nG1c4f , \5851 );
buf \U$3878 ( \5853 , \5852_nG1c4f );
xor \U$3879 ( \5854 , \5267 , \5288 );
xor \U$3880 ( \5855 , \5854 , \5341 );
buf g1c53_GF_PartitionCandidate( \5856_nG1c53 , \5855 );
buf \U$3881 ( \5857 , \5856_nG1c53 );
xor \U$3882 ( \5858 , \5853 , \5857 );
xor \U$3883 ( \5859 , \5857 , \5819 );
not \U$3884 ( \5860 , \5859 );
and \U$3885 ( \5861 , \5858 , \5860 );
and \U$3886 ( \5862 , \5849 , \5861 );
and \U$3887 ( \5863 , RI9922978_574, \5448 );
and \U$3888 ( \5864 , RI99235a8_554, \5454 );
and \U$3889 ( \5865 , RI9923f08_534, \5456 );
and \U$3890 ( \5866 , RI9924868_514, \5458 );
and \U$3891 ( \5867 , RI9925858_494, \5460 );
and \U$3892 ( \5868 , RI99261b8_474, \5462 );
and \U$3893 ( \5869 , RI9926b18_454, \5464 );
and \U$3894 ( \5870 , RI9927ec8_434, \5466 );
and \U$3895 ( \5871 , RI9928828_414, \5468 );
and \U$3896 ( \5872 , RI9929188_394, \5470 );
and \U$3897 ( \5873 , RI992a8f8_374, \5472 );
and \U$3898 ( \5874 , RI992b258_354, \5474 );
and \U$3899 ( \5875 , RI992cd88_334, \5476 );
and \U$3900 ( \5876 , RI992d6e8_314, \5478 );
and \U$3901 ( \5877 , RI992f5d8_294, \5480 );
and \U$3902 ( \5878 , RI9931888_274, \5482 );
and \U$3903 ( \5879 , RI9935fc8_254, \5484 );
or \U$3904 ( \5880 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 );
_DC g24d7 ( \5881_nG24d7 , \5880 , \5503 );
buf \U$3905 ( \5882 , \5881_nG24d7 );
and \U$3906 ( \5883 , \5882 , \5859 );
nor \U$3907 ( \5884 , \5862 , \5883 );
and \U$3908 ( \5885 , \5857 , \5819 );
not \U$3909 ( \5886 , \5885 );
and \U$3910 ( \5887 , \5853 , \5886 );
xnor \U$3911 ( \5888 , \5884 , \5887 );
and \U$3912 ( \5889 , \5829 , \5888 );
and \U$3913 ( \5890 , RI9922810_577, \5448 );
and \U$3914 ( \5891 , RI9923440_557, \5454 );
and \U$3915 ( \5892 , RI9923da0_537, \5456 );
and \U$3916 ( \5893 , RI9924700_517, \5458 );
and \U$3917 ( \5894 , RI99256f0_497, \5460 );
and \U$3918 ( \5895 , RI9926050_477, \5462 );
and \U$3919 ( \5896 , RI99269b0_457, \5464 );
and \U$3920 ( \5897 , RI9927d60_437, \5466 );
and \U$3921 ( \5898 , RI99286c0_417, \5468 );
and \U$3922 ( \5899 , RI9929020_397, \5470 );
and \U$3923 ( \5900 , RI992a790_377, \5472 );
and \U$3924 ( \5901 , RI992b0f0_357, \5474 );
and \U$3925 ( \5902 , RI992cc20_337, \5476 );
and \U$3926 ( \5903 , RI992d580_317, \5478 );
and \U$3927 ( \5904 , RI992f470_297, \5480 );
and \U$3928 ( \5905 , RI9931720_277, \5482 );
and \U$3929 ( \5906 , RI9933d90_257, \5484 );
or \U$3930 ( \5907 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 );
_DC g226a ( \5908_nG226a , \5907 , \5503 );
buf \U$3931 ( \5909 , \5908_nG226a );
xor \U$3932 ( \5910 , \5192 , \5213 );
xor \U$3933 ( \5911 , \5910 , \5350 );
buf g1d72_GF_PartitionCandidate( \5912_nG1d72 , \5911 );
buf \U$3934 ( \5913 , \5912_nG1d72 );
xor \U$3935 ( \5914 , \5217 , \5238 );
xor \U$3936 ( \5915 , \5914 , \5347 );
buf g1d4e_GF_PartitionCandidate( \5916_nG1d4e , \5915 );
buf \U$3937 ( \5917 , \5916_nG1d4e );
xor \U$3938 ( \5918 , \5913 , \5917 );
xor \U$3939 ( \5919 , \5917 , \5853 );
not \U$3940 ( \5920 , \5919 );
and \U$3941 ( \5921 , \5918 , \5920 );
and \U$3942 ( \5922 , \5909 , \5921 );
and \U$3943 ( \5923 , RI9922888_576, \5448 );
and \U$3944 ( \5924 , RI99234b8_556, \5454 );
and \U$3945 ( \5925 , RI9923e18_536, \5456 );
and \U$3946 ( \5926 , RI9924778_516, \5458 );
and \U$3947 ( \5927 , RI9925768_496, \5460 );
and \U$3948 ( \5928 , RI99260c8_476, \5462 );
and \U$3949 ( \5929 , RI9926a28_456, \5464 );
and \U$3950 ( \5930 , RI9927dd8_436, \5466 );
and \U$3951 ( \5931 , RI9928738_416, \5468 );
and \U$3952 ( \5932 , RI9929098_396, \5470 );
and \U$3953 ( \5933 , RI992a808_376, \5472 );
and \U$3954 ( \5934 , RI992b168_356, \5474 );
and \U$3955 ( \5935 , RI992cc98_336, \5476 );
and \U$3956 ( \5936 , RI992d5f8_316, \5478 );
and \U$3957 ( \5937 , RI992f4e8_296, \5480 );
and \U$3958 ( \5938 , RI9931798_276, \5482 );
and \U$3959 ( \5939 , RI9935ed8_256, \5484 );
or \U$3960 ( \5940 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 );
_DC g2302 ( \5941_nG2302 , \5940 , \5503 );
buf \U$3961 ( \5942 , \5941_nG2302 );
and \U$3962 ( \5943 , \5942 , \5919 );
nor \U$3963 ( \5944 , \5922 , \5943 );
and \U$3964 ( \5945 , \5917 , \5853 );
not \U$3965 ( \5946 , \5945 );
and \U$3966 ( \5947 , \5913 , \5946 );
xnor \U$3967 ( \5948 , \5944 , \5947 );
and \U$3968 ( \5949 , \5888 , \5948 );
and \U$3969 ( \5950 , \5829 , \5948 );
or \U$3970 ( \5951 , \5889 , \5949 , \5950 );
and \U$3971 ( \5952 , RI9922720_579, \5448 );
and \U$3972 ( \5953 , RI9923350_559, \5454 );
and \U$3973 ( \5954 , RI9923cb0_539, \5456 );
and \U$3974 ( \5955 , RI9924610_519, \5458 );
and \U$3975 ( \5956 , RI9925600_499, \5460 );
and \U$3976 ( \5957 , RI9925f60_479, \5462 );
and \U$3977 ( \5958 , RI99268c0_459, \5464 );
and \U$3978 ( \5959 , RI9927c70_439, \5466 );
and \U$3979 ( \5960 , RI99285d0_419, \5468 );
and \U$3980 ( \5961 , RI9928f30_399, \5470 );
and \U$3981 ( \5962 , RI992a6a0_379, \5472 );
and \U$3982 ( \5963 , RI992b000_359, \5474 );
and \U$3983 ( \5964 , RI992cb30_339, \5476 );
and \U$3984 ( \5965 , RI992d490_319, \5478 );
and \U$3985 ( \5966 , RI992f380_299, \5480 );
and \U$3986 ( \5967 , RI9931630_279, \5482 );
and \U$3987 ( \5968 , RI9933ca0_259, \5484 );
or \U$3988 ( \5969 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 );
_DC g209f ( \5970_nG209f , \5969 , \5503 );
buf \U$3989 ( \5971 , \5970_nG209f );
xor \U$3990 ( \5972 , \5167 , \5188 );
xor \U$3991 ( \5973 , \5972 , \5353 );
buf g1ebd_GF_PartitionCandidate( \5974_nG1ebd , \5973 );
buf \U$3992 ( \5975 , \5974_nG1ebd );
xor \U$3993 ( \5976 , \5677 , \5975 );
xor \U$3994 ( \5977 , \5975 , \5913 );
not \U$3995 ( \5978 , \5977 );
and \U$3996 ( \5979 , \5976 , \5978 );
and \U$3997 ( \5980 , \5971 , \5979 );
and \U$3998 ( \5981 , RI9922798_578, \5448 );
and \U$3999 ( \5982 , RI99233c8_558, \5454 );
and \U$4000 ( \5983 , RI9923d28_538, \5456 );
and \U$4001 ( \5984 , RI9924688_518, \5458 );
and \U$4002 ( \5985 , RI9925678_498, \5460 );
and \U$4003 ( \5986 , RI9925fd8_478, \5462 );
and \U$4004 ( \5987 , RI9926938_458, \5464 );
and \U$4005 ( \5988 , RI9927ce8_438, \5466 );
and \U$4006 ( \5989 , RI9928648_418, \5468 );
and \U$4007 ( \5990 , RI9928fa8_398, \5470 );
and \U$4008 ( \5991 , RI992a718_378, \5472 );
and \U$4009 ( \5992 , RI992b078_358, \5474 );
and \U$4010 ( \5993 , RI992cba8_338, \5476 );
and \U$4011 ( \5994 , RI992d508_318, \5478 );
and \U$4012 ( \5995 , RI992f3f8_298, \5480 );
and \U$4013 ( \5996 , RI99316a8_278, \5482 );
and \U$4014 ( \5997 , RI9933d18_258, \5484 );
or \U$4015 ( \5998 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 );
_DC g2129 ( \5999_nG2129 , \5998 , \5503 );
buf \U$4016 ( \6000 , \5999_nG2129 );
and \U$4017 ( \6001 , \6000 , \5977 );
nor \U$4018 ( \6002 , \5980 , \6001 );
and \U$4019 ( \6003 , \5975 , \5913 );
not \U$4020 ( \6004 , \6003 );
and \U$4021 ( \6005 , \5677 , \6004 );
xnor \U$4022 ( \6006 , \6002 , \6005 );
and \U$4023 ( \6007 , RI9922630_581, \5448 );
and \U$4024 ( \6008 , RI9923260_561, \5454 );
and \U$4025 ( \6009 , RI9923bc0_541, \5456 );
and \U$4026 ( \6010 , RI9924520_521, \5458 );
and \U$4027 ( \6011 , RI9925510_501, \5460 );
and \U$4028 ( \6012 , RI9925e70_481, \5462 );
and \U$4029 ( \6013 , RI99267d0_461, \5464 );
and \U$4030 ( \6014 , RI9927b80_441, \5466 );
and \U$4031 ( \6015 , RI99284e0_421, \5468 );
and \U$4032 ( \6016 , RI9928e40_401, \5470 );
and \U$4033 ( \6017 , RI992a5b0_381, \5472 );
and \U$4034 ( \6018 , RI992af10_361, \5474 );
and \U$4035 ( \6019 , RI992ca40_341, \5476 );
and \U$4036 ( \6020 , RI992d3a0_321, \5478 );
and \U$4037 ( \6021 , RI992f290_301, \5480 );
and \U$4038 ( \6022 , RI9931540_281, \5482 );
and \U$4039 ( \6023 , RI9933bb0_261, \5484 );
or \U$4040 ( \6024 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 );
_DC g1efc ( \6025_nG1efc , \6024 , \5503 );
buf \U$4041 ( \6026 , \6025_nG1efc );
and \U$4042 ( \6027 , \6026 , \5680 );
and \U$4043 ( \6028 , RI99226a8_580, \5448 );
and \U$4044 ( \6029 , RI99232d8_560, \5454 );
and \U$4045 ( \6030 , RI9923c38_540, \5456 );
and \U$4046 ( \6031 , RI9924598_520, \5458 );
and \U$4047 ( \6032 , RI9925588_500, \5460 );
and \U$4048 ( \6033 , RI9925ee8_480, \5462 );
and \U$4049 ( \6034 , RI9926848_460, \5464 );
and \U$4050 ( \6035 , RI9927bf8_440, \5466 );
and \U$4051 ( \6036 , RI9928558_420, \5468 );
and \U$4052 ( \6037 , RI9928eb8_400, \5470 );
and \U$4053 ( \6038 , RI992a628_380, \5472 );
and \U$4054 ( \6039 , RI992af88_360, \5474 );
and \U$4055 ( \6040 , RI992cab8_340, \5476 );
and \U$4056 ( \6041 , RI992d418_320, \5478 );
and \U$4057 ( \6042 , RI992f308_300, \5480 );
and \U$4058 ( \6043 , RI99315b8_280, \5482 );
and \U$4059 ( \6044 , RI9933c28_260, \5484 );
or \U$4060 ( \6045 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 );
_DC g1f70 ( \6046_nG1f70 , \6045 , \5503 );
buf \U$4061 ( \6047 , \6046_nG1f70 );
and \U$4062 ( \6048 , \6047 , \5678 );
nor \U$4063 ( \6049 , \6027 , \6048 );
xnor \U$4064 ( \6050 , \6049 , \5685 );
and \U$4065 ( \6051 , \6006 , \6050 );
and \U$4066 ( \6052 , RI9922540_583, \5448 );
and \U$4067 ( \6053 , RI9923170_563, \5454 );
and \U$4068 ( \6054 , RI9923ad0_543, \5456 );
and \U$4069 ( \6055 , RI9924430_523, \5458 );
and \U$4070 ( \6056 , RI9924d90_503, \5460 );
and \U$4071 ( \6057 , RI9925d80_483, \5462 );
and \U$4072 ( \6058 , RI99266e0_463, \5464 );
and \U$4073 ( \6059 , RI9927040_443, \5466 );
and \U$4074 ( \6060 , RI99283f0_423, \5468 );
and \U$4075 ( \6061 , RI9928d50_403, \5470 );
and \U$4076 ( \6062 , RI992a4c0_383, \5472 );
and \U$4077 ( \6063 , RI992ae20_363, \5474 );
and \U$4078 ( \6064 , RI992c950_343, \5476 );
and \U$4079 ( \6065 , RI992d2b0_323, \5478 );
and \U$4080 ( \6066 , RI992f1a0_303, \5480 );
and \U$4081 ( \6067 , RI9931450_283, \5482 );
and \U$4082 ( \6068 , RI9933ac0_263, \5484 );
or \U$4083 ( \6069 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 );
_DC g1d8b ( \6070_nG1d8b , \6069 , \5503 );
buf \U$4084 ( \6071 , \6070_nG1d8b );
and \U$4085 ( \6072 , \6071 , \5615 );
and \U$4086 ( \6073 , RI99225b8_582, \5448 );
and \U$4087 ( \6074 , RI99231e8_562, \5454 );
and \U$4088 ( \6075 , RI9923b48_542, \5456 );
and \U$4089 ( \6076 , RI99244a8_522, \5458 );
and \U$4090 ( \6077 , RI9924e08_502, \5460 );
and \U$4091 ( \6078 , RI9925df8_482, \5462 );
and \U$4092 ( \6079 , RI9926758_462, \5464 );
and \U$4093 ( \6080 , RI9927b08_442, \5466 );
and \U$4094 ( \6081 , RI9928468_422, \5468 );
and \U$4095 ( \6082 , RI9928dc8_402, \5470 );
and \U$4096 ( \6083 , RI992a538_382, \5472 );
and \U$4097 ( \6084 , RI992ae98_362, \5474 );
and \U$4098 ( \6085 , RI992c9c8_342, \5476 );
and \U$4099 ( \6086 , RI992d328_322, \5478 );
and \U$4100 ( \6087 , RI992f218_302, \5480 );
and \U$4101 ( \6088 , RI99314c8_282, \5482 );
and \U$4102 ( \6089 , RI9933b38_262, \5484 );
or \U$4103 ( \6090 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 );
_DC g1df2 ( \6091_nG1df2 , \6090 , \5503 );
buf \U$4104 ( \6092 , \6091_nG1df2 );
and \U$4105 ( \6093 , \6092 , \5613 );
nor \U$4106 ( \6094 , \6072 , \6093 );
xnor \U$4107 ( \6095 , \6094 , \5382 );
and \U$4108 ( \6096 , \6050 , \6095 );
and \U$4109 ( \6097 , \6006 , \6095 );
or \U$4110 ( \6098 , \6051 , \6096 , \6097 );
and \U$4111 ( \6099 , \5951 , \6098 );
and \U$4112 ( \6100 , RI9922450_585, \5448 );
and \U$4113 ( \6101 , RI9923080_565, \5454 );
and \U$4114 ( \6102 , RI99239e0_545, \5456 );
and \U$4115 ( \6103 , RI9924340_525, \5458 );
and \U$4116 ( \6104 , RI9924ca0_505, \5460 );
and \U$4117 ( \6105 , RI9925c90_485, \5462 );
and \U$4118 ( \6106 , RI99265f0_465, \5464 );
and \U$4119 ( \6107 , RI9926f50_445, \5466 );
and \U$4120 ( \6108 , RI9928300_425, \5468 );
and \U$4121 ( \6109 , RI9928c60_405, \5470 );
and \U$4122 ( \6110 , RI992a3d0_385, \5472 );
and \U$4123 ( \6111 , RI992ad30_365, \5474 );
and \U$4124 ( \6112 , RI992c860_345, \5476 );
and \U$4125 ( \6113 , RI992d1c0_325, \5478 );
and \U$4126 ( \6114 , RI992f0b0_305, \5480 );
and \U$4127 ( \6115 , RI9931360_285, \5482 );
and \U$4128 ( \6116 , RI99339d0_265, \5484 );
or \U$4129 ( \6117 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 );
_DC g1c0d ( \6118_nG1c0d , \6117 , \5503 );
buf \U$4130 ( \6119 , \6118_nG1c0d );
and \U$4131 ( \6120 , \6119 , \5553 );
and \U$4132 ( \6121 , RI99224c8_584, \5448 );
and \U$4133 ( \6122 , RI99230f8_564, \5454 );
and \U$4134 ( \6123 , RI9923a58_544, \5456 );
and \U$4135 ( \6124 , RI99243b8_524, \5458 );
and \U$4136 ( \6125 , RI9924d18_504, \5460 );
and \U$4137 ( \6126 , RI9925d08_484, \5462 );
and \U$4138 ( \6127 , RI9926668_464, \5464 );
and \U$4139 ( \6128 , RI9926fc8_444, \5466 );
and \U$4140 ( \6129 , RI9928378_424, \5468 );
and \U$4141 ( \6130 , RI9928cd8_404, \5470 );
and \U$4142 ( \6131 , RI992a448_384, \5472 );
and \U$4143 ( \6132 , RI992ada8_364, \5474 );
and \U$4144 ( \6133 , RI992c8d8_344, \5476 );
and \U$4145 ( \6134 , RI992d238_324, \5478 );
and \U$4146 ( \6135 , RI992f128_304, \5480 );
and \U$4147 ( \6136 , RI99313d8_284, \5482 );
and \U$4148 ( \6137 , RI9933a48_264, \5484 );
or \U$4149 ( \6138 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 );
_DC g1ca0 ( \6139_nG1ca0 , \6138 , \5503 );
buf \U$4150 ( \6140 , \6139_nG1ca0 );
and \U$4151 ( \6141 , \6140 , \5551 );
nor \U$4152 ( \6142 , \6120 , \6141 );
xnor \U$4153 ( \6143 , \6142 , \5579 );
and \U$4155 ( \6144 , RI99223d8_586, \5448 );
and \U$4156 ( \6145 , RI9923008_566, \5454 );
and \U$4157 ( \6146 , RI9923968_546, \5456 );
and \U$4158 ( \6147 , RI99242c8_526, \5458 );
and \U$4159 ( \6148 , RI9924c28_506, \5460 );
and \U$4160 ( \6149 , RI9925c18_486, \5462 );
and \U$4161 ( \6150 , RI9926578_466, \5464 );
and \U$4162 ( \6151 , RI9926ed8_446, \5466 );
and \U$4163 ( \6152 , RI9928288_426, \5468 );
and \U$4164 ( \6153 , RI9928be8_406, \5470 );
and \U$4165 ( \6154 , RI992a358_386, \5472 );
and \U$4166 ( \6155 , RI992acb8_366, \5474 );
and \U$4167 ( \6156 , RI992c7e8_346, \5476 );
and \U$4168 ( \6157 , RI992d148_326, \5478 );
and \U$4169 ( \6158 , RI992f038_306, \5480 );
and \U$4170 ( \6159 , RI99312e8_286, \5482 );
and \U$4171 ( \6160 , RI9933958_266, \5484 );
or \U$4172 ( \6161 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 );
_DC g1b85 ( \6162_nG1b85 , \6161 , \5503 );
buf \U$4173 ( \6163 , \6162_nG1b85 );
and \U$4174 ( \6164 , \6163 , \5606 );
nor \U$4175 ( \6165 , 1'b0 , \6164 );
xnor \U$4176 ( \6166 , \6165 , 1'b0 );
and \U$4177 ( \6167 , \6143 , \6166 );
and \U$4178 ( \6168 , \6098 , \6167 );
and \U$4179 ( \6169 , \5951 , \6167 );
or \U$4180 ( \6170 , \6099 , \6168 , \6169 );
and \U$4182 ( \6171 , \6092 , \5615 );
and \U$4183 ( \6172 , \6026 , \5613 );
nor \U$4184 ( \6173 , \6171 , \6172 );
xnor \U$4185 ( \6174 , \6173 , \5382 );
and \U$4186 ( \6175 , \6140 , \5553 );
and \U$4187 ( \6176 , \6071 , \5551 );
nor \U$4188 ( \6177 , \6175 , \6176 );
xnor \U$4189 ( \6178 , \6177 , \5579 );
xor \U$4190 ( \6179 , \6174 , \6178 );
and \U$4192 ( \6180 , \6119 , \5606 );
nor \U$4193 ( \6181 , 1'b0 , \6180 );
xnor \U$4194 ( \6182 , \6181 , 1'b0 );
xor \U$4195 ( \6183 , \6179 , \6182 );
and \U$4196 ( \6184 , \5942 , \5921 );
and \U$4197 ( \6185 , \5849 , \5919 );
nor \U$4198 ( \6186 , \6184 , \6185 );
xnor \U$4199 ( \6187 , \6186 , \5947 );
and \U$4200 ( \6188 , \6000 , \5979 );
and \U$4201 ( \6189 , \5909 , \5977 );
nor \U$4202 ( \6190 , \6188 , \6189 );
xnor \U$4203 ( \6191 , \6190 , \6005 );
xor \U$4204 ( \6192 , \6187 , \6191 );
and \U$4205 ( \6193 , \6047 , \5680 );
and \U$4206 ( \6194 , \5971 , \5678 );
nor \U$4207 ( \6195 , \6193 , \6194 );
xnor \U$4208 ( \6196 , \6195 , \5685 );
xor \U$4209 ( \6197 , \6192 , \6196 );
and \U$4210 ( \6198 , \6183 , \6197 );
or \U$4212 ( \6199 , 1'b0 , \6198 , 1'b0 );
xor \U$4213 ( \6200 , \6170 , \6199 );
and \U$4214 ( \6201 , \6071 , \5553 );
and \U$4215 ( \6202 , \6092 , \5551 );
nor \U$4216 ( \6203 , \6201 , \6202 );
xnor \U$4217 ( \6204 , \6203 , \5579 );
and \U$4219 ( \6205 , \6140 , \5606 );
nor \U$4220 ( \6206 , 1'b0 , \6205 );
xnor \U$4221 ( \6207 , \6206 , 1'b0 );
xor \U$4222 ( \6208 , \6204 , \6207 );
xor \U$4224 ( \6209 , \6208 , 1'b0 );
and \U$4225 ( \6210 , \5909 , \5979 );
and \U$4226 ( \6211 , \5942 , \5977 );
nor \U$4227 ( \6212 , \6210 , \6211 );
xnor \U$4228 ( \6213 , \6212 , \6005 );
and \U$4229 ( \6214 , \5971 , \5680 );
and \U$4230 ( \6215 , \6000 , \5678 );
nor \U$4231 ( \6216 , \6214 , \6215 );
xnor \U$4232 ( \6217 , \6216 , \5685 );
xor \U$4233 ( \6218 , \6213 , \6217 );
and \U$4234 ( \6219 , \6026 , \5615 );
and \U$4235 ( \6220 , \6047 , \5613 );
nor \U$4236 ( \6221 , \6219 , \6220 );
xnor \U$4237 ( \6222 , \6221 , \5382 );
xor \U$4238 ( \6223 , \6218 , \6222 );
xor \U$4239 ( \6224 , \6209 , \6223 );
and \U$4240 ( \6225 , \5733 , \5825 );
and \U$4241 ( \6226 , \5601 , \5822 );
nor \U$4242 ( \6227 , \6225 , \6226 );
xnor \U$4243 ( \6228 , \6227 , \5819 );
and \U$4244 ( \6229 , \5756 , \5861 );
and \U$4245 ( \6230 , \5712 , \5859 );
nor \U$4246 ( \6231 , \6229 , \6230 );
xnor \U$4247 ( \6232 , \6231 , \5887 );
xor \U$4248 ( \6233 , \6228 , \6232 );
and \U$4249 ( \6234 , \5849 , \5921 );
and \U$4250 ( \6235 , \5882 , \5919 );
nor \U$4251 ( \6236 , \6234 , \6235 );
xnor \U$4252 ( \6237 , \6236 , \5947 );
xor \U$4253 ( \6238 , \6233 , \6237 );
xor \U$4254 ( \6239 , \6224 , \6238 );
xor \U$4255 ( \6240 , \6200 , \6239 );
and \U$4257 ( \6241 , \5882 , \5825 );
and \U$4258 ( \6242 , \5756 , \5822 );
nor \U$4259 ( \6243 , \6241 , \6242 );
xnor \U$4260 ( \6244 , \6243 , \5819 );
and \U$4261 ( \6245 , \5942 , \5861 );
and \U$4262 ( \6246 , \5849 , \5859 );
nor \U$4263 ( \6247 , \6245 , \6246 );
xnor \U$4264 ( \6248 , \6247 , \5887 );
and \U$4265 ( \6249 , \6244 , \6248 );
or \U$4267 ( \6250 , 1'b0 , \6249 , 1'b0 );
and \U$4268 ( \6251 , \6000 , \5921 );
and \U$4269 ( \6252 , \5909 , \5919 );
nor \U$4270 ( \6253 , \6251 , \6252 );
xnor \U$4271 ( \6254 , \6253 , \5947 );
and \U$4272 ( \6255 , \6047 , \5979 );
and \U$4273 ( \6256 , \5971 , \5977 );
nor \U$4274 ( \6257 , \6255 , \6256 );
xnor \U$4275 ( \6258 , \6257 , \6005 );
and \U$4276 ( \6259 , \6254 , \6258 );
and \U$4277 ( \6260 , \6092 , \5680 );
and \U$4278 ( \6261 , \6026 , \5678 );
nor \U$4279 ( \6262 , \6260 , \6261 );
xnor \U$4280 ( \6263 , \6262 , \5685 );
and \U$4281 ( \6264 , \6258 , \6263 );
and \U$4282 ( \6265 , \6254 , \6263 );
or \U$4283 ( \6266 , \6259 , \6264 , \6265 );
and \U$4284 ( \6267 , \6250 , \6266 );
and \U$4285 ( \6268 , \6140 , \5615 );
and \U$4286 ( \6269 , \6071 , \5613 );
nor \U$4287 ( \6270 , \6268 , \6269 );
xnor \U$4288 ( \6271 , \6270 , \5382 );
and \U$4289 ( \6272 , \6163 , \5553 );
and \U$4290 ( \6273 , \6119 , \5551 );
nor \U$4291 ( \6274 , \6272 , \6273 );
xnor \U$4292 ( \6275 , \6274 , \5579 );
and \U$4293 ( \6276 , \6271 , \6275 );
and \U$4294 ( \6277 , RI9922360_587, \5448 );
and \U$4295 ( \6278 , RI9922f90_567, \5454 );
and \U$4296 ( \6279 , RI99238f0_547, \5456 );
and \U$4297 ( \6280 , RI9924250_527, \5458 );
and \U$4298 ( \6281 , RI9924bb0_507, \5460 );
and \U$4299 ( \6282 , RI9925ba0_487, \5462 );
and \U$4300 ( \6283 , RI9926500_467, \5464 );
and \U$4301 ( \6284 , RI9926e60_447, \5466 );
and \U$4302 ( \6285 , RI9928210_427, \5468 );
and \U$4303 ( \6286 , RI9928b70_407, \5470 );
and \U$4304 ( \6287 , RI992a2e0_387, \5472 );
and \U$4305 ( \6288 , RI992ac40_367, \5474 );
and \U$4306 ( \6289 , RI992c770_347, \5476 );
and \U$4307 ( \6290 , RI992d0d0_327, \5478 );
and \U$4308 ( \6291 , RI992efc0_307, \5480 );
and \U$4309 ( \6292 , RI992f920_287, \5482 );
and \U$4310 ( \6293 , RI99338e0_267, \5484 );
or \U$4311 ( \6294 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 );
_DC g1aea ( \6295_nG1aea , \6294 , \5503 );
buf \U$4312 ( \6296 , \6295_nG1aea );
nand \U$4313 ( \6297 , \6296 , \5606 );
xnor \U$4314 ( \6298 , \6297 , 1'b0 );
and \U$4315 ( \6299 , \6275 , \6298 );
and \U$4316 ( \6300 , \6271 , \6298 );
or \U$4317 ( \6301 , \6276 , \6299 , \6300 );
and \U$4318 ( \6302 , \6266 , \6301 );
and \U$4319 ( \6303 , \6250 , \6301 );
or \U$4320 ( \6304 , \6267 , \6302 , \6303 );
xor \U$4321 ( \6305 , \6143 , \6166 );
xor \U$4322 ( \6306 , \6006 , \6050 );
xor \U$4323 ( \6307 , \6306 , \6095 );
and \U$4324 ( \6308 , \6305 , \6307 );
xor \U$4325 ( \6309 , \5829 , \5888 );
xor \U$4326 ( \6310 , \6309 , \5948 );
and \U$4327 ( \6311 , \6307 , \6310 );
and \U$4328 ( \6312 , \6305 , \6310 );
or \U$4329 ( \6313 , \6308 , \6311 , \6312 );
and \U$4330 ( \6314 , \6304 , \6313 );
and \U$4332 ( \6315 , \5712 , \5825 );
and \U$4333 ( \6316 , \5733 , \5822 );
nor \U$4334 ( \6317 , \6315 , \6316 );
xnor \U$4335 ( \6318 , \6317 , \5819 );
xor \U$4336 ( \6319 , 1'b0 , \6318 );
and \U$4337 ( \6320 , \5882 , \5861 );
and \U$4338 ( \6321 , \5756 , \5859 );
nor \U$4339 ( \6322 , \6320 , \6321 );
xnor \U$4340 ( \6323 , \6322 , \5887 );
xor \U$4341 ( \6324 , \6319 , \6323 );
and \U$4342 ( \6325 , \6313 , \6324 );
and \U$4343 ( \6326 , \6304 , \6324 );
or \U$4344 ( \6327 , \6314 , \6325 , \6326 );
xor \U$4346 ( \6328 , 1'b0 , \6183 );
xor \U$4347 ( \6329 , \6328 , \6197 );
xor \U$4348 ( \6330 , \5951 , \6098 );
xor \U$4349 ( \6331 , \6330 , \6167 );
and \U$4350 ( \6332 , \6329 , \6331 );
xor \U$4351 ( \6333 , \6327 , \6332 );
and \U$4353 ( \6334 , \6318 , \6323 );
or \U$4355 ( \6335 , 1'b0 , \6334 , 1'b0 );
and \U$4356 ( \6336 , \6187 , \6191 );
and \U$4357 ( \6337 , \6191 , \6196 );
and \U$4358 ( \6338 , \6187 , \6196 );
or \U$4359 ( \6339 , \6336 , \6337 , \6338 );
xor \U$4360 ( \6340 , \6335 , \6339 );
and \U$4361 ( \6341 , \6174 , \6178 );
and \U$4362 ( \6342 , \6178 , \6182 );
and \U$4363 ( \6343 , \6174 , \6182 );
or \U$4364 ( \6344 , \6341 , \6342 , \6343 );
xor \U$4365 ( \6345 , \6340 , \6344 );
xor \U$4366 ( \6346 , \6333 , \6345 );
xor \U$4367 ( \6347 , \6240 , \6346 );
and \U$4368 ( \6348 , \5849 , \5825 );
and \U$4369 ( \6349 , \5882 , \5822 );
nor \U$4370 ( \6350 , \6348 , \6349 );
xnor \U$4371 ( \6351 , \6350 , \5819 );
and \U$4372 ( \6352 , \5909 , \5861 );
and \U$4373 ( \6353 , \5942 , \5859 );
nor \U$4374 ( \6354 , \6352 , \6353 );
xnor \U$4375 ( \6355 , \6354 , \5887 );
and \U$4376 ( \6356 , \6351 , \6355 );
and \U$4377 ( \6357 , \5971 , \5921 );
and \U$4378 ( \6358 , \6000 , \5919 );
nor \U$4379 ( \6359 , \6357 , \6358 );
xnor \U$4380 ( \6360 , \6359 , \5947 );
and \U$4381 ( \6361 , \6355 , \6360 );
and \U$4382 ( \6362 , \6351 , \6360 );
or \U$4383 ( \6363 , \6356 , \6361 , \6362 );
and \U$4384 ( \6364 , \6026 , \5979 );
and \U$4385 ( \6365 , \6047 , \5977 );
nor \U$4386 ( \6366 , \6364 , \6365 );
xnor \U$4387 ( \6367 , \6366 , \6005 );
and \U$4388 ( \6368 , \6071 , \5680 );
and \U$4389 ( \6369 , \6092 , \5678 );
nor \U$4390 ( \6370 , \6368 , \6369 );
xnor \U$4391 ( \6371 , \6370 , \5685 );
and \U$4392 ( \6372 , \6367 , \6371 );
and \U$4393 ( \6373 , \6119 , \5615 );
and \U$4394 ( \6374 , \6140 , \5613 );
nor \U$4395 ( \6375 , \6373 , \6374 );
xnor \U$4396 ( \6376 , \6375 , \5382 );
and \U$4397 ( \6377 , \6371 , \6376 );
and \U$4398 ( \6378 , \6367 , \6376 );
or \U$4399 ( \6379 , \6372 , \6377 , \6378 );
and \U$4400 ( \6380 , \6363 , \6379 );
xor \U$4401 ( \6381 , \6271 , \6275 );
xor \U$4402 ( \6382 , \6381 , \6298 );
and \U$4403 ( \6383 , \6379 , \6382 );
and \U$4404 ( \6384 , \6363 , \6382 );
or \U$4405 ( \6385 , \6380 , \6383 , \6384 );
xor \U$4406 ( \6386 , \6254 , \6258 );
xor \U$4407 ( \6387 , \6386 , \6263 );
xor \U$4408 ( \6388 , 1'b0 , \6244 );
xor \U$4409 ( \6389 , \6388 , \6248 );
and \U$4410 ( \6390 , \6387 , \6389 );
and \U$4411 ( \6391 , \6385 , \6390 );
xor \U$4412 ( \6392 , \6305 , \6307 );
xor \U$4413 ( \6393 , \6392 , \6310 );
and \U$4414 ( \6394 , \6390 , \6393 );
and \U$4415 ( \6395 , \6385 , \6393 );
or \U$4416 ( \6396 , \6391 , \6394 , \6395 );
xor \U$4417 ( \6397 , \6329 , \6331 );
and \U$4418 ( \6398 , \6396 , \6397 );
xor \U$4419 ( \6399 , \6304 , \6313 );
xor \U$4420 ( \6400 , \6399 , \6324 );
and \U$4421 ( \6401 , \6397 , \6400 );
and \U$4422 ( \6402 , \6396 , \6400 );
or \U$4423 ( \6403 , \6398 , \6401 , \6402 );
nor \U$4424 ( \6404 , \6347 , \6403 );
and \U$4425 ( \6405 , \6327 , \6332 );
and \U$4426 ( \6406 , \6332 , \6345 );
and \U$4427 ( \6407 , \6327 , \6345 );
or \U$4428 ( \6408 , \6405 , \6406 , \6407 );
and \U$4429 ( \6409 , \6170 , \6199 );
and \U$4430 ( \6410 , \6199 , \6239 );
and \U$4431 ( \6411 , \6170 , \6239 );
or \U$4432 ( \6412 , \6409 , \6410 , \6411 );
and \U$4434 ( \6413 , \5601 , \5825 );
and \U$4435 ( \6414 , \5505 , \5822 );
nor \U$4436 ( \6415 , \6413 , \6414 );
xnor \U$4437 ( \6416 , \6415 , \5819 );
xor \U$4438 ( \6417 , 1'b0 , \6416 );
and \U$4439 ( \6418 , \5712 , \5861 );
and \U$4440 ( \6419 , \5733 , \5859 );
nor \U$4441 ( \6420 , \6418 , \6419 );
xnor \U$4442 ( \6421 , \6420 , \5887 );
xor \U$4443 ( \6422 , \6417 , \6421 );
and \U$4445 ( \6423 , \6047 , \5615 );
and \U$4446 ( \6424 , \5971 , \5613 );
nor \U$4447 ( \6425 , \6423 , \6424 );
xnor \U$4448 ( \6426 , \6425 , \5382 );
and \U$4449 ( \6427 , \6092 , \5553 );
and \U$4450 ( \6428 , \6026 , \5551 );
nor \U$4451 ( \6429 , \6427 , \6428 );
xnor \U$4452 ( \6430 , \6429 , \5579 );
xor \U$4453 ( \6431 , \6426 , \6430 );
and \U$4455 ( \6432 , \6071 , \5606 );
nor \U$4456 ( \6433 , 1'b0 , \6432 );
xnor \U$4457 ( \6434 , \6433 , 1'b0 );
xor \U$4458 ( \6435 , \6431 , \6434 );
xor \U$4459 ( \6436 , 1'b0 , \6435 );
xor \U$4460 ( \6437 , \6422 , \6436 );
and \U$4461 ( \6438 , \6228 , \6232 );
and \U$4462 ( \6439 , \6232 , \6237 );
and \U$4463 ( \6440 , \6228 , \6237 );
or \U$4464 ( \6441 , \6438 , \6439 , \6440 );
and \U$4465 ( \6442 , \6213 , \6217 );
and \U$4466 ( \6443 , \6217 , \6222 );
and \U$4467 ( \6444 , \6213 , \6222 );
or \U$4468 ( \6445 , \6442 , \6443 , \6444 );
xor \U$4469 ( \6446 , \6441 , \6445 );
and \U$4470 ( \6447 , \6204 , \6207 );
or \U$4473 ( \6448 , \6447 , 1'b0 , 1'b0 );
xor \U$4474 ( \6449 , \6446 , \6448 );
xor \U$4475 ( \6450 , \6437 , \6449 );
xor \U$4476 ( \6451 , \6412 , \6450 );
and \U$4477 ( \6452 , \6335 , \6339 );
and \U$4478 ( \6453 , \6339 , \6344 );
and \U$4479 ( \6454 , \6335 , \6344 );
or \U$4480 ( \6455 , \6452 , \6453 , \6454 );
and \U$4481 ( \6456 , \6209 , \6223 );
and \U$4482 ( \6457 , \6223 , \6238 );
and \U$4483 ( \6458 , \6209 , \6238 );
or \U$4484 ( \6459 , \6456 , \6457 , \6458 );
xor \U$4485 ( \6460 , \6455 , \6459 );
and \U$4486 ( \6461 , \5882 , \5921 );
and \U$4487 ( \6462 , \5756 , \5919 );
nor \U$4488 ( \6463 , \6461 , \6462 );
xnor \U$4489 ( \6464 , \6463 , \5947 );
and \U$4490 ( \6465 , \5942 , \5979 );
and \U$4491 ( \6466 , \5849 , \5977 );
nor \U$4492 ( \6467 , \6465 , \6466 );
xnor \U$4493 ( \6468 , \6467 , \6005 );
xor \U$4494 ( \6469 , \6464 , \6468 );
and \U$4495 ( \6470 , \6000 , \5680 );
and \U$4496 ( \6471 , \5909 , \5678 );
nor \U$4497 ( \6472 , \6470 , \6471 );
xnor \U$4498 ( \6473 , \6472 , \5685 );
xor \U$4499 ( \6474 , \6469 , \6473 );
xor \U$4500 ( \6475 , \6460 , \6474 );
xor \U$4501 ( \6476 , \6451 , \6475 );
xor \U$4502 ( \6477 , \6408 , \6476 );
and \U$4503 ( \6478 , \6240 , \6346 );
nor \U$4504 ( \6479 , \6477 , \6478 );
nor \U$4505 ( \6480 , \6404 , \6479 );
and \U$4506 ( \6481 , \6412 , \6450 );
and \U$4507 ( \6482 , \6450 , \6475 );
and \U$4508 ( \6483 , \6412 , \6475 );
or \U$4509 ( \6484 , \6481 , \6482 , \6483 );
and \U$4511 ( \6485 , \6416 , \6421 );
or \U$4513 ( \6486 , 1'b0 , \6485 , 1'b0 );
and \U$4514 ( \6487 , \6464 , \6468 );
and \U$4515 ( \6488 , \6468 , \6473 );
and \U$4516 ( \6489 , \6464 , \6473 );
or \U$4517 ( \6490 , \6487 , \6488 , \6489 );
xor \U$4518 ( \6491 , \6486 , \6490 );
and \U$4519 ( \6492 , \6426 , \6430 );
and \U$4520 ( \6493 , \6430 , \6434 );
and \U$4521 ( \6494 , \6426 , \6434 );
or \U$4522 ( \6495 , \6492 , \6493 , \6494 );
xor \U$4523 ( \6496 , \6491 , \6495 );
and \U$4524 ( \6497 , \6441 , \6445 );
and \U$4525 ( \6498 , \6445 , \6448 );
and \U$4526 ( \6499 , \6441 , \6448 );
or \U$4527 ( \6500 , \6497 , \6498 , \6499 );
xor \U$4529 ( \6501 , \6500 , 1'b0 );
and \U$4530 ( \6502 , \5505 , \5825 );
and \U$4531 ( \6503 , \5574 , \5822 );
nor \U$4532 ( \6504 , \6502 , \6503 );
xnor \U$4533 ( \6505 , \6504 , \5819 );
and \U$4534 ( \6506 , \5733 , \5861 );
and \U$4535 ( \6507 , \5601 , \5859 );
nor \U$4536 ( \6508 , \6506 , \6507 );
xnor \U$4537 ( \6509 , \6508 , \5887 );
xor \U$4538 ( \6510 , \6505 , \6509 );
and \U$4539 ( \6511 , \5756 , \5921 );
and \U$4540 ( \6512 , \5712 , \5919 );
nor \U$4541 ( \6513 , \6511 , \6512 );
xnor \U$4542 ( \6514 , \6513 , \5947 );
xor \U$4543 ( \6515 , \6510 , \6514 );
xor \U$4544 ( \6516 , \6501 , \6515 );
xor \U$4545 ( \6517 , \6496 , \6516 );
xor \U$4546 ( \6518 , \6484 , \6517 );
and \U$4547 ( \6519 , \6455 , \6459 );
and \U$4548 ( \6520 , \6459 , \6474 );
and \U$4549 ( \6521 , \6455 , \6474 );
or \U$4550 ( \6522 , \6519 , \6520 , \6521 );
and \U$4551 ( \6523 , \6422 , \6436 );
and \U$4552 ( \6524 , \6436 , \6449 );
and \U$4553 ( \6525 , \6422 , \6449 );
or \U$4554 ( \6526 , \6523 , \6524 , \6525 );
xor \U$4555 ( \6527 , \6522 , \6526 );
and \U$4557 ( \6528 , \6026 , \5553 );
and \U$4558 ( \6529 , \6047 , \5551 );
nor \U$4559 ( \6530 , \6528 , \6529 );
xnor \U$4560 ( \6531 , \6530 , \5579 );
and \U$4562 ( \6532 , \6092 , \5606 );
nor \U$4563 ( \6533 , 1'b0 , \6532 );
xnor \U$4564 ( \6534 , \6533 , 1'b0 );
xor \U$4565 ( \6535 , \6531 , \6534 );
xor \U$4567 ( \6536 , \6535 , 1'b0 );
xor \U$4568 ( \6537 , 1'b0 , \6536 );
and \U$4569 ( \6538 , \5849 , \5979 );
and \U$4570 ( \6539 , \5882 , \5977 );
nor \U$4571 ( \6540 , \6538 , \6539 );
xnor \U$4572 ( \6541 , \6540 , \6005 );
and \U$4573 ( \6542 , \5909 , \5680 );
and \U$4574 ( \6543 , \5942 , \5678 );
nor \U$4575 ( \6544 , \6542 , \6543 );
xnor \U$4576 ( \6545 , \6544 , \5685 );
xor \U$4577 ( \6546 , \6541 , \6545 );
and \U$4578 ( \6547 , \5971 , \5615 );
and \U$4579 ( \6548 , \6000 , \5613 );
nor \U$4580 ( \6549 , \6547 , \6548 );
xnor \U$4581 ( \6550 , \6549 , \5382 );
xor \U$4582 ( \6551 , \6546 , \6550 );
xor \U$4583 ( \6552 , \6537 , \6551 );
xor \U$4584 ( \6553 , \6527 , \6552 );
xor \U$4585 ( \6554 , \6518 , \6553 );
and \U$4586 ( \6555 , \6408 , \6476 );
nor \U$4587 ( \6556 , \6554 , \6555 );
and \U$4588 ( \6557 , \6522 , \6526 );
and \U$4589 ( \6558 , \6526 , \6552 );
and \U$4590 ( \6559 , \6522 , \6552 );
or \U$4591 ( \6560 , \6557 , \6558 , \6559 );
and \U$4592 ( \6561 , \6496 , \6516 );
xor \U$4593 ( \6562 , \6560 , \6561 );
and \U$4596 ( \6563 , \6500 , \6515 );
or \U$4597 ( \6564 , 1'b0 , 1'b0 , \6563 );
and \U$4599 ( \6565 , \6000 , \5615 );
and \U$4600 ( \6566 , \5909 , \5613 );
nor \U$4601 ( \6567 , \6565 , \6566 );
xnor \U$4602 ( \6568 , \6567 , \5382 );
and \U$4603 ( \6569 , \6047 , \5553 );
and \U$4604 ( \6570 , \5971 , \5551 );
nor \U$4605 ( \6571 , \6569 , \6570 );
xnor \U$4606 ( \6572 , \6571 , \5579 );
xor \U$4607 ( \6573 , \6568 , \6572 );
and \U$4609 ( \6574 , \6026 , \5606 );
nor \U$4610 ( \6575 , 1'b0 , \6574 );
xnor \U$4611 ( \6576 , \6575 , 1'b0 );
xor \U$4612 ( \6577 , \6573 , \6576 );
xor \U$4613 ( \6578 , 1'b0 , \6577 );
and \U$4614 ( \6579 , \5712 , \5921 );
and \U$4615 ( \6580 , \5733 , \5919 );
nor \U$4616 ( \6581 , \6579 , \6580 );
xnor \U$4617 ( \6582 , \6581 , \5947 );
and \U$4618 ( \6583 , \5882 , \5979 );
and \U$4619 ( \6584 , \5756 , \5977 );
nor \U$4620 ( \6585 , \6583 , \6584 );
xnor \U$4621 ( \6586 , \6585 , \6005 );
xor \U$4622 ( \6587 , \6582 , \6586 );
and \U$4623 ( \6588 , \5942 , \5680 );
and \U$4624 ( \6589 , \5849 , \5678 );
nor \U$4625 ( \6590 , \6588 , \6589 );
xnor \U$4626 ( \6591 , \6590 , \5685 );
xor \U$4627 ( \6592 , \6587 , \6591 );
xor \U$4628 ( \6593 , \6578 , \6592 );
and \U$4629 ( \6594 , \6505 , \6509 );
and \U$4630 ( \6595 , \6509 , \6514 );
and \U$4631 ( \6596 , \6505 , \6514 );
or \U$4632 ( \6597 , \6594 , \6595 , \6596 );
and \U$4633 ( \6598 , \6541 , \6545 );
and \U$4634 ( \6599 , \6545 , \6550 );
and \U$4635 ( \6600 , \6541 , \6550 );
or \U$4636 ( \6601 , \6598 , \6599 , \6600 );
xor \U$4637 ( \6602 , \6597 , \6601 );
and \U$4638 ( \6603 , \6531 , \6534 );
or \U$4641 ( \6604 , \6603 , 1'b0 , 1'b0 );
xor \U$4642 ( \6605 , \6602 , \6604 );
xor \U$4643 ( \6606 , \6593 , \6605 );
xor \U$4644 ( \6607 , \6564 , \6606 );
and \U$4645 ( \6608 , \6486 , \6490 );
and \U$4646 ( \6609 , \6490 , \6495 );
and \U$4647 ( \6610 , \6486 , \6495 );
or \U$4648 ( \6611 , \6608 , \6609 , \6610 );
and \U$4650 ( \6612 , \6536 , \6551 );
or \U$4652 ( \6613 , 1'b0 , \6612 , 1'b0 );
xor \U$4653 ( \6614 , \6611 , \6613 );
and \U$4655 ( \6615 , \5574 , \5825 );
not \U$4656 ( \6616 , \6615 );
xnor \U$4657 ( \6617 , \6616 , \5819 );
xor \U$4658 ( \6618 , 1'b0 , \6617 );
and \U$4659 ( \6619 , \5601 , \5861 );
and \U$4660 ( \6620 , \5505 , \5859 );
nor \U$4661 ( \6621 , \6619 , \6620 );
xnor \U$4662 ( \6622 , \6621 , \5887 );
xor \U$4663 ( \6623 , \6618 , \6622 );
xor \U$4664 ( \6624 , \6614 , \6623 );
xor \U$4665 ( \6625 , \6607 , \6624 );
xor \U$4666 ( \6626 , \6562 , \6625 );
and \U$4667 ( \6627 , \6484 , \6517 );
and \U$4668 ( \6628 , \6517 , \6553 );
and \U$4669 ( \6629 , \6484 , \6553 );
or \U$4670 ( \6630 , \6627 , \6628 , \6629 );
nor \U$4671 ( \6631 , \6626 , \6630 );
nor \U$4672 ( \6632 , \6556 , \6631 );
nand \U$4673 ( \6633 , \6480 , \6632 );
and \U$4674 ( \6634 , \6564 , \6606 );
and \U$4675 ( \6635 , \6606 , \6624 );
and \U$4676 ( \6636 , \6564 , \6624 );
or \U$4677 ( \6637 , \6634 , \6635 , \6636 );
and \U$4678 ( \6638 , \6597 , \6601 );
and \U$4679 ( \6639 , \6601 , \6604 );
and \U$4680 ( \6640 , \6597 , \6604 );
or \U$4681 ( \6641 , \6638 , \6639 , \6640 );
and \U$4683 ( \6642 , \6577 , \6592 );
or \U$4685 ( \6643 , 1'b0 , \6642 , 1'b0 );
xor \U$4686 ( \6644 , \6641 , \6643 );
and \U$4687 ( \6645 , \5756 , \5979 );
and \U$4688 ( \6646 , \5712 , \5977 );
nor \U$4689 ( \6647 , \6645 , \6646 );
xnor \U$4690 ( \6648 , \6647 , \6005 );
and \U$4691 ( \6649 , \5849 , \5680 );
and \U$4692 ( \6650 , \5882 , \5678 );
nor \U$4693 ( \6651 , \6649 , \6650 );
xnor \U$4694 ( \6652 , \6651 , \5685 );
xor \U$4695 ( \6653 , \6648 , \6652 );
and \U$4696 ( \6654 , \5909 , \5615 );
and \U$4697 ( \6655 , \5942 , \5613 );
nor \U$4698 ( \6656 , \6654 , \6655 );
xnor \U$4699 ( \6657 , \6656 , \5382 );
xor \U$4700 ( \6658 , \6653 , \6657 );
xor \U$4701 ( \6659 , \6644 , \6658 );
xor \U$4702 ( \6660 , \6637 , \6659 );
and \U$4703 ( \6661 , \6611 , \6613 );
and \U$4704 ( \6662 , \6613 , \6623 );
and \U$4705 ( \6663 , \6611 , \6623 );
or \U$4706 ( \6664 , \6661 , \6662 , \6663 );
and \U$4707 ( \6665 , \6593 , \6605 );
xor \U$4708 ( \6666 , \6664 , \6665 );
not \U$4709 ( \6667 , \5819 );
and \U$4710 ( \6668 , \5505 , \5861 );
and \U$4711 ( \6669 , \5574 , \5859 );
nor \U$4712 ( \6670 , \6668 , \6669 );
xnor \U$4713 ( \6671 , \6670 , \5887 );
xor \U$4714 ( \6672 , \6667 , \6671 );
and \U$4715 ( \6673 , \5733 , \5921 );
and \U$4716 ( \6674 , \5601 , \5919 );
nor \U$4717 ( \6675 , \6673 , \6674 );
xnor \U$4718 ( \6676 , \6675 , \5947 );
xor \U$4719 ( \6677 , \6672 , \6676 );
and \U$4721 ( \6678 , \5971 , \5553 );
and \U$4722 ( \6679 , \6000 , \5551 );
nor \U$4723 ( \6680 , \6678 , \6679 );
xnor \U$4724 ( \6681 , \6680 , \5579 );
and \U$4726 ( \6682 , \6047 , \5606 );
nor \U$4727 ( \6683 , 1'b0 , \6682 );
xnor \U$4728 ( \6684 , \6683 , 1'b0 );
xor \U$4729 ( \6685 , \6681 , \6684 );
xor \U$4731 ( \6686 , \6685 , 1'b0 );
xor \U$4732 ( \6687 , 1'b1 , \6686 );
xor \U$4733 ( \6688 , \6677 , \6687 );
and \U$4735 ( \6689 , \6617 , \6622 );
or \U$4737 ( \6690 , 1'b0 , \6689 , 1'b0 );
and \U$4738 ( \6691 , \6582 , \6586 );
and \U$4739 ( \6692 , \6586 , \6591 );
and \U$4740 ( \6693 , \6582 , \6591 );
or \U$4741 ( \6694 , \6691 , \6692 , \6693 );
xor \U$4742 ( \6695 , \6690 , \6694 );
and \U$4743 ( \6696 , \6568 , \6572 );
and \U$4744 ( \6697 , \6572 , \6576 );
and \U$4745 ( \6698 , \6568 , \6576 );
or \U$4746 ( \6699 , \6696 , \6697 , \6698 );
xor \U$4747 ( \6700 , \6695 , \6699 );
xor \U$4748 ( \6701 , \6688 , \6700 );
xor \U$4749 ( \6702 , \6666 , \6701 );
xor \U$4750 ( \6703 , \6660 , \6702 );
and \U$4751 ( \6704 , \6560 , \6561 );
and \U$4752 ( \6705 , \6561 , \6625 );
and \U$4753 ( \6706 , \6560 , \6625 );
or \U$4754 ( \6707 , \6704 , \6705 , \6706 );
nor \U$4755 ( \6708 , \6703 , \6707 );
and \U$4756 ( \6709 , \6664 , \6665 );
and \U$4757 ( \6710 , \6665 , \6701 );
and \U$4758 ( \6711 , \6664 , \6701 );
or \U$4759 ( \6712 , \6709 , \6710 , \6711 );
and \U$4760 ( \6713 , \6667 , \6671 );
and \U$4761 ( \6714 , \6671 , \6676 );
and \U$4762 ( \6715 , \6667 , \6676 );
or \U$4763 ( \6716 , \6713 , \6714 , \6715 );
and \U$4764 ( \6717 , \6648 , \6652 );
and \U$4765 ( \6718 , \6652 , \6657 );
and \U$4766 ( \6719 , \6648 , \6657 );
or \U$4767 ( \6720 , \6717 , \6718 , \6719 );
xor \U$4768 ( \6721 , \6716 , \6720 );
and \U$4769 ( \6722 , \6681 , \6684 );
or \U$4772 ( \6723 , \6722 , 1'b0 , 1'b0 );
xor \U$4773 ( \6724 , \6721 , \6723 );
and \U$4774 ( \6725 , \6690 , \6694 );
and \U$4775 ( \6726 , \6694 , \6699 );
and \U$4776 ( \6727 , \6690 , \6699 );
or \U$4777 ( \6728 , \6725 , \6726 , \6727 );
and \U$4780 ( \6729 , 1'b1 , \6686 );
or \U$4782 ( \6730 , 1'b0 , \6729 , 1'b0 );
xor \U$4783 ( \6731 , \6728 , \6730 );
and \U$4784 ( \6732 , \6000 , \5553 );
and \U$4785 ( \6733 , \5909 , \5551 );
nor \U$4786 ( \6734 , \6732 , \6733 );
xnor \U$4787 ( \6735 , \6734 , \5579 );
and \U$4789 ( \6736 , \5971 , \5606 );
nor \U$4790 ( \6737 , 1'b0 , \6736 );
xnor \U$4791 ( \6738 , \6737 , 1'b0 );
xor \U$4792 ( \6739 , \6735 , \6738 );
xor \U$4794 ( \6740 , \6739 , 1'b0 );
and \U$4795 ( \6741 , \5712 , \5979 );
and \U$4796 ( \6742 , \5733 , \5977 );
nor \U$4797 ( \6743 , \6741 , \6742 );
xnor \U$4798 ( \6744 , \6743 , \6005 );
and \U$4799 ( \6745 , \5882 , \5680 );
and \U$4800 ( \6746 , \5756 , \5678 );
nor \U$4801 ( \6747 , \6745 , \6746 );
xnor \U$4802 ( \6748 , \6747 , \5685 );
xor \U$4803 ( \6749 , \6744 , \6748 );
and \U$4804 ( \6750 , \5942 , \5615 );
and \U$4805 ( \6751 , \5849 , \5613 );
nor \U$4806 ( \6752 , \6750 , \6751 );
xnor \U$4807 ( \6753 , \6752 , \5382 );
xor \U$4808 ( \6754 , \6749 , \6753 );
xor \U$4809 ( \6755 , \6740 , \6754 );
and \U$4811 ( \6756 , \5574 , \5861 );
not \U$4812 ( \6757 , \6756 );
xnor \U$4813 ( \6758 , \6757 , \5887 );
xor \U$4814 ( \6759 , 1'b0 , \6758 );
and \U$4815 ( \6760 , \5601 , \5921 );
and \U$4816 ( \6761 , \5505 , \5919 );
nor \U$4817 ( \6762 , \6760 , \6761 );
xnor \U$4818 ( \6763 , \6762 , \5947 );
xor \U$4819 ( \6764 , \6759 , \6763 );
xor \U$4820 ( \6765 , \6755 , \6764 );
xor \U$4821 ( \6766 , \6731 , \6765 );
xor \U$4822 ( \6767 , \6724 , \6766 );
xor \U$4823 ( \6768 , \6712 , \6767 );
and \U$4824 ( \6769 , \6641 , \6643 );
and \U$4825 ( \6770 , \6643 , \6658 );
and \U$4826 ( \6771 , \6641 , \6658 );
or \U$4827 ( \6772 , \6769 , \6770 , \6771 );
and \U$4828 ( \6773 , \6677 , \6687 );
and \U$4829 ( \6774 , \6687 , \6700 );
and \U$4830 ( \6775 , \6677 , \6700 );
or \U$4831 ( \6776 , \6773 , \6774 , \6775 );
xor \U$4832 ( \6777 , \6772 , \6776 );
xor \U$4834 ( \6778 , \6777 , 1'b1 );
xor \U$4835 ( \6779 , \6768 , \6778 );
and \U$4836 ( \6780 , \6637 , \6659 );
and \U$4837 ( \6781 , \6659 , \6702 );
and \U$4838 ( \6782 , \6637 , \6702 );
or \U$4839 ( \6783 , \6780 , \6781 , \6782 );
nor \U$4840 ( \6784 , \6779 , \6783 );
nor \U$4841 ( \6785 , \6708 , \6784 );
and \U$4842 ( \6786 , \6772 , \6776 );
and \U$4843 ( \6787 , \6776 , 1'b1 );
and \U$4844 ( \6788 , \6772 , 1'b1 );
or \U$4845 ( \6789 , \6786 , \6787 , \6788 );
and \U$4846 ( \6790 , \6724 , \6766 );
xor \U$4847 ( \6791 , \6789 , \6790 );
and \U$4848 ( \6792 , \6728 , \6730 );
and \U$4849 ( \6793 , \6730 , \6765 );
and \U$4850 ( \6794 , \6728 , \6765 );
or \U$4851 ( \6795 , \6792 , \6793 , \6794 );
and \U$4853 ( \6796 , \6000 , \5606 );
nor \U$4854 ( \6797 , 1'b0 , \6796 );
xnor \U$4855 ( \6798 , \6797 , 1'b0 );
xor \U$4857 ( \6799 , \6798 , 1'b0 );
xor \U$4859 ( \6800 , \6799 , 1'b0 );
and \U$4860 ( \6801 , \5756 , \5680 );
and \U$4861 ( \6802 , \5712 , \5678 );
nor \U$4862 ( \6803 , \6801 , \6802 );
xnor \U$4863 ( \6804 , \6803 , \5685 );
and \U$4864 ( \6805 , \5849 , \5615 );
and \U$4865 ( \6806 , \5882 , \5613 );
nor \U$4866 ( \6807 , \6805 , \6806 );
xnor \U$4867 ( \6808 , \6807 , \5382 );
xor \U$4868 ( \6809 , \6804 , \6808 );
and \U$4869 ( \6810 , \5909 , \5553 );
and \U$4870 ( \6811 , \5942 , \5551 );
nor \U$4871 ( \6812 , \6810 , \6811 );
xnor \U$4872 ( \6813 , \6812 , \5579 );
xor \U$4873 ( \6814 , \6809 , \6813 );
xor \U$4874 ( \6815 , \6800 , \6814 );
not \U$4875 ( \6816 , \5887 );
and \U$4876 ( \6817 , \5505 , \5921 );
and \U$4877 ( \6818 , \5574 , \5919 );
nor \U$4878 ( \6819 , \6817 , \6818 );
xnor \U$4879 ( \6820 , \6819 , \5947 );
xor \U$4880 ( \6821 , \6816 , \6820 );
and \U$4881 ( \6822 , \5733 , \5979 );
and \U$4882 ( \6823 , \5601 , \5977 );
nor \U$4883 ( \6824 , \6822 , \6823 );
xnor \U$4884 ( \6825 , \6824 , \6005 );
xor \U$4885 ( \6826 , \6821 , \6825 );
xor \U$4886 ( \6827 , \6815 , \6826 );
xor \U$4888 ( \6828 , \6827 , 1'b0 );
and \U$4890 ( \6829 , \6758 , \6763 );
or \U$4892 ( \6830 , 1'b0 , \6829 , 1'b0 );
and \U$4893 ( \6831 , \6744 , \6748 );
and \U$4894 ( \6832 , \6748 , \6753 );
and \U$4895 ( \6833 , \6744 , \6753 );
or \U$4896 ( \6834 , \6831 , \6832 , \6833 );
xor \U$4897 ( \6835 , \6830 , \6834 );
and \U$4898 ( \6836 , \6735 , \6738 );
or \U$4901 ( \6837 , \6836 , 1'b0 , 1'b0 );
xor \U$4902 ( \6838 , \6835 , \6837 );
xor \U$4903 ( \6839 , \6828 , \6838 );
xor \U$4904 ( \6840 , \6795 , \6839 );
and \U$4905 ( \6841 , \6716 , \6720 );
and \U$4906 ( \6842 , \6720 , \6723 );
and \U$4907 ( \6843 , \6716 , \6723 );
or \U$4908 ( \6844 , \6841 , \6842 , \6843 );
xor \U$4910 ( \6845 , \6844 , 1'b0 );
and \U$4911 ( \6846 , \6740 , \6754 );
and \U$4912 ( \6847 , \6754 , \6764 );
and \U$4913 ( \6848 , \6740 , \6764 );
or \U$4914 ( \6849 , \6846 , \6847 , \6848 );
xor \U$4915 ( \6850 , \6845 , \6849 );
xor \U$4916 ( \6851 , \6840 , \6850 );
xor \U$4917 ( \6852 , \6791 , \6851 );
and \U$4918 ( \6853 , \6712 , \6767 );
and \U$4919 ( \6854 , \6767 , \6778 );
and \U$4920 ( \6855 , \6712 , \6778 );
or \U$4921 ( \6856 , \6853 , \6854 , \6855 );
nor \U$4922 ( \6857 , \6852 , \6856 );
and \U$4923 ( \6858 , \6795 , \6839 );
and \U$4924 ( \6859 , \6839 , \6850 );
and \U$4925 ( \6860 , \6795 , \6850 );
or \U$4926 ( \6861 , \6858 , \6859 , \6860 );
and \U$4927 ( \6862 , \6830 , \6834 );
and \U$4928 ( \6863 , \6834 , \6837 );
and \U$4929 ( \6864 , \6830 , \6837 );
or \U$4930 ( \6865 , \6862 , \6863 , \6864 );
xor \U$4932 ( \6866 , \6865 , 1'b0 );
and \U$4933 ( \6867 , \6800 , \6814 );
and \U$4934 ( \6868 , \6814 , \6826 );
and \U$4935 ( \6869 , \6800 , \6826 );
or \U$4936 ( \6870 , \6867 , \6868 , \6869 );
xor \U$4937 ( \6871 , \6866 , \6870 );
xor \U$4938 ( \6872 , \6861 , \6871 );
and \U$4941 ( \6873 , \6844 , \6849 );
or \U$4942 ( \6874 , 1'b0 , 1'b0 , \6873 );
and \U$4945 ( \6875 , \6827 , \6838 );
or \U$4946 ( \6876 , 1'b0 , 1'b0 , \6875 );
xor \U$4947 ( \6877 , \6874 , \6876 );
and \U$4948 ( \6878 , \5712 , \5680 );
and \U$4949 ( \6879 , \5733 , \5678 );
nor \U$4950 ( \6880 , \6878 , \6879 );
xnor \U$4951 ( \6881 , \6880 , \5685 );
and \U$4952 ( \6882 , \5882 , \5615 );
and \U$4953 ( \6883 , \5756 , \5613 );
nor \U$4954 ( \6884 , \6882 , \6883 );
xnor \U$4955 ( \6885 , \6884 , \5382 );
xor \U$4956 ( \6886 , \6881 , \6885 );
and \U$4957 ( \6887 , \5942 , \5553 );
and \U$4958 ( \6888 , \5849 , \5551 );
nor \U$4959 ( \6889 , \6887 , \6888 );
xnor \U$4960 ( \6890 , \6889 , \5579 );
xor \U$4961 ( \6891 , \6886 , \6890 );
and \U$4963 ( \6892 , \5574 , \5921 );
not \U$4964 ( \6893 , \6892 );
xnor \U$4965 ( \6894 , \6893 , \5947 );
xor \U$4966 ( \6895 , 1'b0 , \6894 );
and \U$4967 ( \6896 , \5601 , \5979 );
and \U$4968 ( \6897 , \5505 , \5977 );
nor \U$4969 ( \6898 , \6896 , \6897 );
xnor \U$4970 ( \6899 , \6898 , \6005 );
xor \U$4971 ( \6900 , \6895 , \6899 );
xor \U$4972 ( \6901 , \6891 , \6900 );
and \U$4975 ( \6902 , \5909 , \5606 );
nor \U$4976 ( \6903 , 1'b0 , \6902 );
xnor \U$4977 ( \6904 , \6903 , 1'b0 );
xor \U$4979 ( \6905 , \6904 , 1'b0 );
xor \U$4981 ( \6906 , \6905 , 1'b0 );
xnor \U$4982 ( \6907 , 1'b0 , \6906 );
xor \U$4983 ( \6908 , \6901 , \6907 );
and \U$4984 ( \6909 , \6816 , \6820 );
and \U$4985 ( \6910 , \6820 , \6825 );
and \U$4986 ( \6911 , \6816 , \6825 );
or \U$4987 ( \6912 , \6909 , \6910 , \6911 );
and \U$4988 ( \6913 , \6804 , \6808 );
and \U$4989 ( \6914 , \6808 , \6813 );
and \U$4990 ( \6915 , \6804 , \6813 );
or \U$4991 ( \6916 , \6913 , \6914 , \6915 );
xor \U$4992 ( \6917 , \6912 , \6916 );
xor \U$4994 ( \6918 , \6917 , 1'b0 );
xor \U$4995 ( \6919 , \6908 , \6918 );
xor \U$4996 ( \6920 , \6877 , \6919 );
xor \U$4997 ( \6921 , \6872 , \6920 );
and \U$4998 ( \6922 , \6789 , \6790 );
and \U$4999 ( \6923 , \6790 , \6851 );
and \U$5000 ( \6924 , \6789 , \6851 );
or \U$5001 ( \6925 , \6922 , \6923 , \6924 );
nor \U$5002 ( \6926 , \6921 , \6925 );
nor \U$5003 ( \6927 , \6857 , \6926 );
nand \U$5004 ( \6928 , \6785 , \6927 );
nor \U$5005 ( \6929 , \6633 , \6928 );
and \U$5006 ( \6930 , \6874 , \6876 );
and \U$5007 ( \6931 , \6876 , \6919 );
and \U$5008 ( \6932 , \6874 , \6919 );
or \U$5009 ( \6933 , \6930 , \6931 , \6932 );
and \U$5010 ( \6934 , \6912 , \6916 );
or \U$5013 ( \6935 , \6934 , 1'b0 , 1'b0 );
or \U$5014 ( \6936 , 1'b0 , \6906 );
xor \U$5015 ( \6937 , \6935 , \6936 );
and \U$5016 ( \6938 , \6891 , \6900 );
xor \U$5017 ( \6939 , \6937 , \6938 );
xor \U$5018 ( \6940 , \6933 , \6939 );
and \U$5021 ( \6941 , \6865 , \6870 );
or \U$5022 ( \6942 , 1'b0 , 1'b0 , \6941 );
and \U$5023 ( \6943 , \6901 , \6907 );
and \U$5024 ( \6944 , \6907 , \6918 );
and \U$5025 ( \6945 , \6901 , \6918 );
or \U$5026 ( \6946 , \6943 , \6944 , \6945 );
xor \U$5027 ( \6947 , \6942 , \6946 );
and \U$5029 ( \6948 , \5756 , \5615 );
and \U$5030 ( \6949 , \5712 , \5613 );
nor \U$5031 ( \6950 , \6948 , \6949 );
xnor \U$5032 ( \6951 , \6950 , \5382 );
and \U$5033 ( \6952 , \5849 , \5553 );
and \U$5034 ( \6953 , \5882 , \5551 );
nor \U$5035 ( \6954 , \6952 , \6953 );
xnor \U$5036 ( \6955 , \6954 , \5579 );
xor \U$5037 ( \6956 , \6951 , \6955 );
and \U$5039 ( \6957 , \5942 , \5606 );
nor \U$5040 ( \6958 , 1'b0 , \6957 );
xnor \U$5041 ( \6959 , \6958 , 1'b0 );
xor \U$5042 ( \6960 , \6956 , \6959 );
xor \U$5043 ( \6961 , 1'b0 , \6960 );
not \U$5044 ( \6962 , \5947 );
and \U$5045 ( \6963 , \5505 , \5979 );
and \U$5046 ( \6964 , \5574 , \5977 );
nor \U$5047 ( \6965 , \6963 , \6964 );
xnor \U$5048 ( \6966 , \6965 , \6005 );
xor \U$5049 ( \6967 , \6962 , \6966 );
and \U$5050 ( \6968 , \5733 , \5680 );
and \U$5051 ( \6969 , \5601 , \5678 );
nor \U$5052 ( \6970 , \6968 , \6969 );
xnor \U$5053 ( \6971 , \6970 , \5685 );
xor \U$5054 ( \6972 , \6967 , \6971 );
xor \U$5055 ( \6973 , \6961 , \6972 );
xor \U$5057 ( \6974 , \6973 , 1'b0 );
and \U$5059 ( \6975 , \6894 , \6899 );
or \U$5061 ( \6976 , 1'b0 , \6975 , 1'b0 );
and \U$5062 ( \6977 , \6881 , \6885 );
and \U$5063 ( \6978 , \6885 , \6890 );
and \U$5064 ( \6979 , \6881 , \6890 );
or \U$5065 ( \6980 , \6977 , \6978 , \6979 );
xor \U$5066 ( \6981 , \6976 , \6980 );
xor \U$5068 ( \6982 , \6981 , 1'b0 );
xor \U$5069 ( \6983 , \6974 , \6982 );
xor \U$5070 ( \6984 , \6947 , \6983 );
xor \U$5071 ( \6985 , \6940 , \6984 );
and \U$5072 ( \6986 , \6861 , \6871 );
and \U$5073 ( \6987 , \6871 , \6920 );
and \U$5074 ( \6988 , \6861 , \6920 );
or \U$5075 ( \6989 , \6986 , \6987 , \6988 );
nor \U$5076 ( \6990 , \6985 , \6989 );
and \U$5077 ( \6991 , \6942 , \6946 );
and \U$5078 ( \6992 , \6946 , \6983 );
and \U$5079 ( \6993 , \6942 , \6983 );
or \U$5080 ( \6994 , \6991 , \6992 , \6993 );
and \U$5081 ( \6995 , \6976 , \6980 );
or \U$5084 ( \6996 , \6995 , 1'b0 , 1'b0 );
xor \U$5086 ( \6997 , \6996 , 1'b0 );
and \U$5088 ( \6998 , \6960 , \6972 );
or \U$5090 ( \6999 , 1'b0 , \6998 , 1'b0 );
xor \U$5091 ( \7000 , \6997 , \6999 );
xor \U$5092 ( \7001 , \6994 , \7000 );
and \U$5093 ( \7002 , \6935 , \6936 );
and \U$5094 ( \7003 , \6936 , \6938 );
and \U$5095 ( \7004 , \6935 , \6938 );
or \U$5096 ( \7005 , \7002 , \7003 , \7004 );
and \U$5099 ( \7006 , \6973 , \6982 );
or \U$5100 ( \7007 , 1'b0 , 1'b0 , \7006 );
xor \U$5101 ( \7008 , \7005 , \7007 );
and \U$5102 ( \7009 , \5712 , \5615 );
and \U$5103 ( \7010 , \5733 , \5613 );
nor \U$5104 ( \7011 , \7009 , \7010 );
xnor \U$5105 ( \7012 , \7011 , \5382 );
and \U$5106 ( \7013 , \5882 , \5553 );
and \U$5107 ( \7014 , \5756 , \5551 );
nor \U$5108 ( \7015 , \7013 , \7014 );
xnor \U$5109 ( \7016 , \7015 , \5579 );
xor \U$5110 ( \7017 , \7012 , \7016 );
and \U$5112 ( \7018 , \5849 , \5606 );
nor \U$5113 ( \7019 , 1'b0 , \7018 );
xnor \U$5114 ( \7020 , \7019 , 1'b0 );
xor \U$5115 ( \7021 , \7017 , \7020 );
and \U$5117 ( \7022 , \5574 , \5979 );
not \U$5118 ( \7023 , \7022 );
xnor \U$5119 ( \7024 , \7023 , \6005 );
xor \U$5120 ( \7025 , 1'b0 , \7024 );
and \U$5121 ( \7026 , \5601 , \5680 );
and \U$5122 ( \7027 , \5505 , \5678 );
nor \U$5123 ( \7028 , \7026 , \7027 );
xnor \U$5124 ( \7029 , \7028 , \5685 );
xor \U$5125 ( \7030 , \7025 , \7029 );
xor \U$5126 ( \7031 , \7021 , \7030 );
xor \U$5128 ( \7032 , \7031 , 1'b1 );
and \U$5129 ( \7033 , \6962 , \6966 );
and \U$5130 ( \7034 , \6966 , \6971 );
and \U$5131 ( \7035 , \6962 , \6971 );
or \U$5132 ( \7036 , \7033 , \7034 , \7035 );
and \U$5133 ( \7037 , \6951 , \6955 );
and \U$5134 ( \7038 , \6955 , \6959 );
and \U$5135 ( \7039 , \6951 , \6959 );
or \U$5136 ( \7040 , \7037 , \7038 , \7039 );
xor \U$5137 ( \7041 , \7036 , \7040 );
xor \U$5139 ( \7042 , \7041 , 1'b0 );
xor \U$5140 ( \7043 , \7032 , \7042 );
xor \U$5141 ( \7044 , \7008 , \7043 );
xor \U$5142 ( \7045 , \7001 , \7044 );
and \U$5143 ( \7046 , \6933 , \6939 );
and \U$5144 ( \7047 , \6939 , \6984 );
and \U$5145 ( \7048 , \6933 , \6984 );
or \U$5146 ( \7049 , \7046 , \7047 , \7048 );
nor \U$5147 ( \7050 , \7045 , \7049 );
nor \U$5148 ( \7051 , \6990 , \7050 );
and \U$5149 ( \7052 , \7005 , \7007 );
and \U$5150 ( \7053 , \7007 , \7043 );
and \U$5151 ( \7054 , \7005 , \7043 );
or \U$5152 ( \7055 , \7052 , \7053 , \7054 );
and \U$5153 ( \7056 , \7036 , \7040 );
or \U$5156 ( \7057 , \7056 , 1'b0 , 1'b0 );
xor \U$5158 ( \7058 , \7057 , 1'b0 );
and \U$5159 ( \7059 , \7021 , \7030 );
xor \U$5160 ( \7060 , \7058 , \7059 );
xor \U$5161 ( \7061 , \7055 , \7060 );
and \U$5164 ( \7062 , \6996 , \6999 );
or \U$5165 ( \7063 , 1'b0 , 1'b0 , \7062 );
and \U$5166 ( \7064 , \7031 , 1'b1 );
and \U$5167 ( \7065 , 1'b1 , \7042 );
and \U$5168 ( \7066 , \7031 , \7042 );
or \U$5169 ( \7067 , \7064 , \7065 , \7066 );
xor \U$5170 ( \7068 , \7063 , \7067 );
and \U$5172 ( \7069 , \5756 , \5553 );
and \U$5173 ( \7070 , \5712 , \5551 );
nor \U$5174 ( \7071 , \7069 , \7070 );
xnor \U$5175 ( \7072 , \7071 , \5579 );
and \U$5177 ( \7073 , \5882 , \5606 );
nor \U$5178 ( \7074 , 1'b0 , \7073 );
xnor \U$5179 ( \7075 , \7074 , 1'b0 );
xor \U$5180 ( \7076 , \7072 , \7075 );
xor \U$5182 ( \7077 , \7076 , 1'b0 );
xor \U$5183 ( \7078 , 1'b0 , \7077 );
not \U$5184 ( \7079 , \6005 );
and \U$5185 ( \7080 , \5505 , \5680 );
and \U$5186 ( \7081 , \5574 , \5678 );
nor \U$5187 ( \7082 , \7080 , \7081 );
xnor \U$5188 ( \7083 , \7082 , \5685 );
xor \U$5189 ( \7084 , \7079 , \7083 );
and \U$5190 ( \7085 , \5733 , \5615 );
and \U$5191 ( \7086 , \5601 , \5613 );
nor \U$5192 ( \7087 , \7085 , \7086 );
xnor \U$5193 ( \7088 , \7087 , \5382 );
xor \U$5194 ( \7089 , \7084 , \7088 );
xor \U$5195 ( \7090 , \7078 , \7089 );
xor \U$5197 ( \7091 , \7090 , 1'b0 );
and \U$5199 ( \7092 , \7024 , \7029 );
or \U$5201 ( \7093 , 1'b0 , \7092 , 1'b0 );
and \U$5202 ( \7094 , \7012 , \7016 );
and \U$5203 ( \7095 , \7016 , \7020 );
and \U$5204 ( \7096 , \7012 , \7020 );
or \U$5205 ( \7097 , \7094 , \7095 , \7096 );
xor \U$5206 ( \7098 , \7093 , \7097 );
xor \U$5208 ( \7099 , \7098 , 1'b0 );
xor \U$5209 ( \7100 , \7091 , \7099 );
xor \U$5210 ( \7101 , \7068 , \7100 );
xor \U$5211 ( \7102 , \7061 , \7101 );
and \U$5212 ( \7103 , \6994 , \7000 );
and \U$5213 ( \7104 , \7000 , \7044 );
and \U$5214 ( \7105 , \6994 , \7044 );
or \U$5215 ( \7106 , \7103 , \7104 , \7105 );
nor \U$5216 ( \7107 , \7102 , \7106 );
and \U$5217 ( \7108 , \7063 , \7067 );
and \U$5218 ( \7109 , \7067 , \7100 );
and \U$5219 ( \7110 , \7063 , \7100 );
or \U$5220 ( \7111 , \7108 , \7109 , \7110 );
and \U$5221 ( \7112 , \7093 , \7097 );
or \U$5224 ( \7113 , \7112 , 1'b0 , 1'b0 );
xor \U$5226 ( \7114 , \7113 , 1'b0 );
and \U$5228 ( \7115 , \7077 , \7089 );
or \U$5230 ( \7116 , 1'b0 , \7115 , 1'b0 );
xor \U$5231 ( \7117 , \7114 , \7116 );
xor \U$5232 ( \7118 , \7111 , \7117 );
and \U$5235 ( \7119 , \7057 , \7059 );
or \U$5236 ( \7120 , 1'b0 , 1'b0 , \7119 );
and \U$5239 ( \7121 , \7090 , \7099 );
or \U$5240 ( \7122 , 1'b0 , 1'b0 , \7121 );
xor \U$5241 ( \7123 , \7120 , \7122 );
xor \U$5242 ( \7124 , \5736 , \5759 );
xor \U$5244 ( \7125 , \7124 , 1'b0 );
xor \U$5246 ( \7126 , 1'b0 , \5686 );
xor \U$5247 ( \7127 , \7126 , \5690 );
xor \U$5248 ( \7128 , \7125 , \7127 );
xor \U$5250 ( \7129 , \7128 , 1'b1 );
and \U$5251 ( \7130 , \7079 , \7083 );
and \U$5252 ( \7131 , \7083 , \7088 );
and \U$5253 ( \7132 , \7079 , \7088 );
or \U$5254 ( \7133 , \7130 , \7131 , \7132 );
and \U$5255 ( \7134 , \7072 , \7075 );
or \U$5258 ( \7135 , \7134 , 1'b0 , 1'b0 );
xor \U$5259 ( \7136 , \7133 , \7135 );
xor \U$5261 ( \7137 , \7136 , 1'b0 );
xor \U$5262 ( \7138 , \7129 , \7137 );
xor \U$5263 ( \7139 , \7123 , \7138 );
xor \U$5264 ( \7140 , \7118 , \7139 );
and \U$5265 ( \7141 , \7055 , \7060 );
and \U$5266 ( \7142 , \7060 , \7101 );
and \U$5267 ( \7143 , \7055 , \7101 );
or \U$5268 ( \7144 , \7141 , \7142 , \7143 );
nor \U$5269 ( \7145 , \7140 , \7144 );
nor \U$5270 ( \7146 , \7107 , \7145 );
nand \U$5271 ( \7147 , \7051 , \7146 );
and \U$5272 ( \7148 , \7120 , \7122 );
and \U$5273 ( \7149 , \7122 , \7138 );
and \U$5274 ( \7150 , \7120 , \7138 );
or \U$5275 ( \7151 , \7148 , \7149 , \7150 );
and \U$5276 ( \7152 , \7133 , \7135 );
or \U$5279 ( \7153 , \7152 , 1'b0 , 1'b0 );
xor \U$5281 ( \7154 , \7153 , 1'b0 );
and \U$5282 ( \7155 , \7125 , \7127 );
xor \U$5283 ( \7156 , \7154 , \7155 );
xor \U$5284 ( \7157 , \7151 , \7156 );
and \U$5287 ( \7158 , \7113 , \7116 );
or \U$5288 ( \7159 , 1'b0 , 1'b0 , \7158 );
and \U$5289 ( \7160 , \7128 , 1'b1 );
and \U$5290 ( \7161 , 1'b1 , \7137 );
and \U$5291 ( \7162 , \7128 , \7137 );
or \U$5292 ( \7163 , \7160 , \7161 , \7162 );
xor \U$5293 ( \7164 , \7159 , \7163 );
xor \U$5295 ( \7165 , 1'b0 , \5768 );
xor \U$5296 ( \7166 , \7165 , \5779 );
xor \U$5298 ( \7167 , \7166 , 1'b0 );
xor \U$5299 ( \7168 , \5692 , \5761 );
xor \U$5301 ( \7169 , \7168 , 1'b0 );
xor \U$5302 ( \7170 , \7167 , \7169 );
xor \U$5303 ( \7171 , \7164 , \7170 );
xor \U$5304 ( \7172 , \7157 , \7171 );
and \U$5305 ( \7173 , \7111 , \7117 );
and \U$5306 ( \7174 , \7117 , \7139 );
and \U$5307 ( \7175 , \7111 , \7139 );
or \U$5308 ( \7176 , \7173 , \7174 , \7175 );
nor \U$5309 ( \7177 , \7172 , \7176 );
and \U$5310 ( \7178 , \7159 , \7163 );
and \U$5311 ( \7179 , \7163 , \7170 );
and \U$5312 ( \7180 , \7159 , \7170 );
or \U$5313 ( \7181 , \7178 , \7179 , \7180 );
xor \U$5315 ( \7182 , \5763 , 1'b0 );
xor \U$5316 ( \7183 , \7182 , \5781 );
xor \U$5317 ( \7184 , \7181 , \7183 );
and \U$5320 ( \7185 , \7153 , \7155 );
or \U$5321 ( \7186 , 1'b0 , 1'b0 , \7185 );
and \U$5324 ( \7187 , \7166 , \7169 );
or \U$5325 ( \7188 , 1'b0 , 1'b0 , \7187 );
xor \U$5326 ( \7189 , \7186 , \7188 );
xor \U$5327 ( \7190 , \5791 , 1'b1 );
xor \U$5328 ( \7191 , \7190 , \5798 );
xor \U$5329 ( \7192 , \7189 , \7191 );
xor \U$5330 ( \7193 , \7184 , \7192 );
and \U$5331 ( \7194 , \7151 , \7156 );
and \U$5332 ( \7195 , \7156 , \7171 );
and \U$5333 ( \7196 , \7151 , \7171 );
or \U$5334 ( \7197 , \7194 , \7195 , \7196 );
nor \U$5335 ( \7198 , \7193 , \7197 );
nor \U$5336 ( \7199 , \7177 , \7198 );
and \U$5337 ( \7200 , \7186 , \7188 );
and \U$5338 ( \7201 , \7188 , \7191 );
and \U$5339 ( \7202 , \7186 , \7191 );
or \U$5340 ( \7203 , \7200 , \7201 , \7202 );
and \U$5342 ( \7204 , \5788 , \5790 );
xor \U$5343 ( \7205 , 1'b0 , \7204 );
xor \U$5344 ( \7206 , \7203 , \7205 );
xor \U$5345 ( \7207 , \5783 , \5801 );
xor \U$5346 ( \7208 , \7207 , \5804 );
xor \U$5347 ( \7209 , \7206 , \7208 );
and \U$5348 ( \7210 , \7181 , \7183 );
and \U$5349 ( \7211 , \7183 , \7192 );
and \U$5350 ( \7212 , \7181 , \7192 );
or \U$5351 ( \7213 , \7210 , \7211 , \7212 );
nor \U$5352 ( \7214 , \7209 , \7213 );
xor \U$5354 ( \7215 , \5807 , 1'b0 );
xor \U$5355 ( \7216 , \7215 , \5809 );
and \U$5356 ( \7217 , \7203 , \7205 );
and \U$5357 ( \7218 , \7205 , \7208 );
and \U$5358 ( \7219 , \7203 , \7208 );
or \U$5359 ( \7220 , \7217 , \7218 , \7219 );
nor \U$5360 ( \7221 , \7216 , \7220 );
nor \U$5361 ( \7222 , \7214 , \7221 );
nand \U$5362 ( \7223 , \7199 , \7222 );
nor \U$5363 ( \7224 , \7147 , \7223 );
nand \U$5364 ( \7225 , \6929 , \7224 );
and \U$5365 ( \7226 , \6026 , \5825 );
and \U$5366 ( \7227 , \6047 , \5822 );
nor \U$5367 ( \7228 , \7226 , \7227 );
xnor \U$5368 ( \7229 , \7228 , \5819 );
and \U$5369 ( \7230 , \6071 , \5861 );
and \U$5370 ( \7231 , \6092 , \5859 );
nor \U$5371 ( \7232 , \7230 , \7231 );
xnor \U$5372 ( \7233 , \7232 , \5887 );
and \U$5373 ( \7234 , \7229 , \7233 );
and \U$5374 ( \7235 , \6119 , \5921 );
and \U$5375 ( \7236 , \6140 , \5919 );
nor \U$5376 ( \7237 , \7235 , \7236 );
xnor \U$5377 ( \7238 , \7237 , \5947 );
and \U$5378 ( \7239 , \7233 , \7238 );
and \U$5379 ( \7240 , \7229 , \7238 );
or \U$5380 ( \7241 , \7234 , \7239 , \7240 );
and \U$5381 ( \7242 , \6140 , \5921 );
and \U$5382 ( \7243 , \6071 , \5919 );
nor \U$5383 ( \7244 , \7242 , \7243 );
xnor \U$5384 ( \7245 , \7244 , \5947 );
and \U$5385 ( \7246 , \6163 , \5979 );
and \U$5386 ( \7247 , \6119 , \5977 );
nor \U$5387 ( \7248 , \7246 , \7247 );
xnor \U$5388 ( \7249 , \7248 , \6005 );
xor \U$5389 ( \7250 , \7245 , \7249 );
nand \U$5390 ( \7251 , \6296 , \5678 );
xnor \U$5391 ( \7252 , \7251 , \5685 );
xor \U$5392 ( \7253 , \7250 , \7252 );
and \U$5393 ( \7254 , \7241 , \7253 );
and \U$5394 ( \7255 , \6047 , \5825 );
and \U$5395 ( \7256 , \5971 , \5822 );
nor \U$5396 ( \7257 , \7255 , \7256 );
xnor \U$5397 ( \7258 , \7257 , \5819 );
xor \U$5398 ( \7259 , \5685 , \7258 );
and \U$5399 ( \7260 , \6092 , \5861 );
and \U$5400 ( \7261 , \6026 , \5859 );
nor \U$5401 ( \7262 , \7260 , \7261 );
xnor \U$5402 ( \7263 , \7262 , \5887 );
xor \U$5403 ( \7264 , \7259 , \7263 );
and \U$5404 ( \7265 , \7253 , \7264 );
and \U$5405 ( \7266 , \7241 , \7264 );
or \U$5406 ( \7267 , \7254 , \7265 , \7266 );
and \U$5407 ( \7268 , \6296 , \5680 );
and \U$5408 ( \7269 , \6163 , \5678 );
nor \U$5409 ( \7270 , \7268 , \7269 );
xnor \U$5410 ( \7271 , \7270 , \5685 );
and \U$5411 ( \7272 , \5971 , \5825 );
and \U$5412 ( \7273 , \6000 , \5822 );
nor \U$5413 ( \7274 , \7272 , \7273 );
xnor \U$5414 ( \7275 , \7274 , \5819 );
and \U$5415 ( \7276 , \6026 , \5861 );
and \U$5416 ( \7277 , \6047 , \5859 );
nor \U$5417 ( \7278 , \7276 , \7277 );
xnor \U$5418 ( \7279 , \7278 , \5887 );
xor \U$5419 ( \7280 , \7275 , \7279 );
and \U$5420 ( \7281 , \6071 , \5921 );
and \U$5421 ( \7282 , \6092 , \5919 );
nor \U$5422 ( \7283 , \7281 , \7282 );
xnor \U$5423 ( \7284 , \7283 , \5947 );
xor \U$5424 ( \7285 , \7280 , \7284 );
xor \U$5425 ( \7286 , \7271 , \7285 );
xor \U$5426 ( \7287 , \7267 , \7286 );
and \U$5427 ( \7288 , \5685 , \7258 );
and \U$5428 ( \7289 , \7258 , \7263 );
and \U$5429 ( \7290 , \5685 , \7263 );
or \U$5430 ( \7291 , \7288 , \7289 , \7290 );
and \U$5431 ( \7292 , \7245 , \7249 );
and \U$5432 ( \7293 , \7249 , \7252 );
and \U$5433 ( \7294 , \7245 , \7252 );
or \U$5434 ( \7295 , \7292 , \7293 , \7294 );
xor \U$5435 ( \7296 , \7291 , \7295 );
and \U$5436 ( \7297 , \6119 , \5979 );
and \U$5437 ( \7298 , \6140 , \5977 );
nor \U$5438 ( \7299 , \7297 , \7298 );
xnor \U$5439 ( \7300 , \7299 , \6005 );
xor \U$5440 ( \7301 , \7296 , \7300 );
xor \U$5441 ( \7302 , \7287 , \7301 );
and \U$5442 ( \7303 , \6092 , \5825 );
and \U$5443 ( \7304 , \6026 , \5822 );
nor \U$5444 ( \7305 , \7303 , \7304 );
xnor \U$5445 ( \7306 , \7305 , \5819 );
and \U$5446 ( \7307 , \6005 , \7306 );
and \U$5447 ( \7308 , \6140 , \5861 );
and \U$5448 ( \7309 , \6071 , \5859 );
nor \U$5449 ( \7310 , \7308 , \7309 );
xnor \U$5450 ( \7311 , \7310 , \5887 );
and \U$5451 ( \7312 , \7306 , \7311 );
and \U$5452 ( \7313 , \6005 , \7311 );
or \U$5453 ( \7314 , \7307 , \7312 , \7313 );
and \U$5454 ( \7315 , \6163 , \5921 );
and \U$5455 ( \7316 , \6119 , \5919 );
nor \U$5456 ( \7317 , \7315 , \7316 );
xnor \U$5457 ( \7318 , \7317 , \5947 );
nand \U$5458 ( \7319 , \6296 , \5977 );
xnor \U$5459 ( \7320 , \7319 , \6005 );
and \U$5460 ( \7321 , \7318 , \7320 );
and \U$5461 ( \7322 , \7314 , \7321 );
and \U$5462 ( \7323 , \6296 , \5979 );
and \U$5463 ( \7324 , \6163 , \5977 );
nor \U$5464 ( \7325 , \7323 , \7324 );
xnor \U$5465 ( \7326 , \7325 , \6005 );
and \U$5466 ( \7327 , \7321 , \7326 );
and \U$5467 ( \7328 , \7314 , \7326 );
or \U$5468 ( \7329 , \7322 , \7327 , \7328 );
xor \U$5469 ( \7330 , \7241 , \7253 );
xor \U$5470 ( \7331 , \7330 , \7264 );
and \U$5471 ( \7332 , \7329 , \7331 );
nor \U$5472 ( \7333 , \7302 , \7332 );
and \U$5473 ( \7334 , \7275 , \7279 );
and \U$5474 ( \7335 , \7279 , \7284 );
and \U$5475 ( \7336 , \7275 , \7284 );
or \U$5476 ( \7337 , \7334 , \7335 , \7336 );
nand \U$5477 ( \7338 , \6296 , \5613 );
xnor \U$5478 ( \7339 , \7338 , \5382 );
xor \U$5479 ( \7340 , \7337 , \7339 );
and \U$5480 ( \7341 , \6092 , \5921 );
and \U$5481 ( \7342 , \6026 , \5919 );
nor \U$5482 ( \7343 , \7341 , \7342 );
xnor \U$5483 ( \7344 , \7343 , \5947 );
and \U$5484 ( \7345 , \6140 , \5979 );
and \U$5485 ( \7346 , \6071 , \5977 );
nor \U$5486 ( \7347 , \7345 , \7346 );
xnor \U$5487 ( \7348 , \7347 , \6005 );
xor \U$5488 ( \7349 , \7344 , \7348 );
and \U$5489 ( \7350 , \6163 , \5680 );
and \U$5490 ( \7351 , \6119 , \5678 );
nor \U$5491 ( \7352 , \7350 , \7351 );
xnor \U$5492 ( \7353 , \7352 , \5685 );
xor \U$5493 ( \7354 , \7349 , \7353 );
xor \U$5494 ( \7355 , \7340 , \7354 );
and \U$5495 ( \7356 , \7291 , \7295 );
and \U$5496 ( \7357 , \7295 , \7300 );
and \U$5497 ( \7358 , \7291 , \7300 );
or \U$5498 ( \7359 , \7356 , \7357 , \7358 );
and \U$5499 ( \7360 , \7271 , \7285 );
xor \U$5500 ( \7361 , \7359 , \7360 );
and \U$5501 ( \7362 , \6000 , \5825 );
and \U$5502 ( \7363 , \5909 , \5822 );
nor \U$5503 ( \7364 , \7362 , \7363 );
xnor \U$5504 ( \7365 , \7364 , \5819 );
xor \U$5505 ( \7366 , \5382 , \7365 );
and \U$5506 ( \7367 , \6047 , \5861 );
and \U$5507 ( \7368 , \5971 , \5859 );
nor \U$5508 ( \7369 , \7367 , \7368 );
xnor \U$5509 ( \7370 , \7369 , \5887 );
xor \U$5510 ( \7371 , \7366 , \7370 );
xor \U$5511 ( \7372 , \7361 , \7371 );
xor \U$5512 ( \7373 , \7355 , \7372 );
and \U$5513 ( \7374 , \7267 , \7286 );
and \U$5514 ( \7375 , \7286 , \7301 );
and \U$5515 ( \7376 , \7267 , \7301 );
or \U$5516 ( \7377 , \7374 , \7375 , \7376 );
nor \U$5517 ( \7378 , \7373 , \7377 );
nor \U$5518 ( \7379 , \7333 , \7378 );
and \U$5519 ( \7380 , \7359 , \7360 );
and \U$5520 ( \7381 , \7360 , \7371 );
and \U$5521 ( \7382 , \7359 , \7371 );
or \U$5522 ( \7383 , \7380 , \7381 , \7382 );
and \U$5523 ( \7384 , \7337 , \7339 );
and \U$5524 ( \7385 , \7339 , \7354 );
and \U$5525 ( \7386 , \7337 , \7354 );
or \U$5526 ( \7387 , \7384 , \7385 , \7386 );
and \U$5527 ( \7388 , \5909 , \5825 );
and \U$5528 ( \7389 , \5942 , \5822 );
nor \U$5529 ( \7390 , \7388 , \7389 );
xnor \U$5530 ( \7391 , \7390 , \5819 );
and \U$5531 ( \7392 , \5971 , \5861 );
and \U$5532 ( \7393 , \6000 , \5859 );
nor \U$5533 ( \7394 , \7392 , \7393 );
xnor \U$5534 ( \7395 , \7394 , \5887 );
xor \U$5535 ( \7396 , \7391 , \7395 );
and \U$5536 ( \7397 , \6026 , \5921 );
and \U$5537 ( \7398 , \6047 , \5919 );
nor \U$5538 ( \7399 , \7397 , \7398 );
xnor \U$5539 ( \7400 , \7399 , \5947 );
xor \U$5540 ( \7401 , \7396 , \7400 );
xor \U$5541 ( \7402 , \7387 , \7401 );
and \U$5542 ( \7403 , \5382 , \7365 );
and \U$5543 ( \7404 , \7365 , \7370 );
and \U$5544 ( \7405 , \5382 , \7370 );
or \U$5545 ( \7406 , \7403 , \7404 , \7405 );
and \U$5546 ( \7407 , \7344 , \7348 );
and \U$5547 ( \7408 , \7348 , \7353 );
and \U$5548 ( \7409 , \7344 , \7353 );
or \U$5549 ( \7410 , \7407 , \7408 , \7409 );
xor \U$5550 ( \7411 , \7406 , \7410 );
and \U$5551 ( \7412 , \6071 , \5979 );
and \U$5552 ( \7413 , \6092 , \5977 );
nor \U$5553 ( \7414 , \7412 , \7413 );
xnor \U$5554 ( \7415 , \7414 , \6005 );
and \U$5555 ( \7416 , \6119 , \5680 );
and \U$5556 ( \7417 , \6140 , \5678 );
nor \U$5557 ( \7418 , \7416 , \7417 );
xnor \U$5558 ( \7419 , \7418 , \5685 );
xor \U$5559 ( \7420 , \7415 , \7419 );
and \U$5560 ( \7421 , \6296 , \5615 );
and \U$5561 ( \7422 , \6163 , \5613 );
nor \U$5562 ( \7423 , \7421 , \7422 );
xnor \U$5563 ( \7424 , \7423 , \5382 );
xor \U$5564 ( \7425 , \7420 , \7424 );
xor \U$5565 ( \7426 , \7411 , \7425 );
xor \U$5566 ( \7427 , \7402 , \7426 );
xor \U$5567 ( \7428 , \7383 , \7427 );
and \U$5568 ( \7429 , \7355 , \7372 );
nor \U$5569 ( \7430 , \7428 , \7429 );
and \U$5570 ( \7431 , \7387 , \7401 );
and \U$5571 ( \7432 , \7401 , \7426 );
and \U$5572 ( \7433 , \7387 , \7426 );
or \U$5573 ( \7434 , \7431 , \7432 , \7433 );
and \U$5574 ( \7435 , \7406 , \7410 );
and \U$5575 ( \7436 , \7410 , \7425 );
and \U$5576 ( \7437 , \7406 , \7425 );
or \U$5577 ( \7438 , \7435 , \7436 , \7437 );
nand \U$5578 ( \7439 , \6296 , \5551 );
xnor \U$5579 ( \7440 , \7439 , \5579 );
and \U$5580 ( \7441 , \6047 , \5921 );
and \U$5581 ( \7442 , \5971 , \5919 );
nor \U$5582 ( \7443 , \7441 , \7442 );
xnor \U$5583 ( \7444 , \7443 , \5947 );
and \U$5584 ( \7445 , \6092 , \5979 );
and \U$5585 ( \7446 , \6026 , \5977 );
nor \U$5586 ( \7447 , \7445 , \7446 );
xnor \U$5587 ( \7448 , \7447 , \6005 );
xor \U$5588 ( \7449 , \7444 , \7448 );
and \U$5589 ( \7450 , \6140 , \5680 );
and \U$5590 ( \7451 , \6071 , \5678 );
nor \U$5591 ( \7452 , \7450 , \7451 );
xnor \U$5592 ( \7453 , \7452 , \5685 );
xor \U$5593 ( \7454 , \7449 , \7453 );
xor \U$5594 ( \7455 , \7440 , \7454 );
and \U$5595 ( \7456 , \5942 , \5825 );
and \U$5596 ( \7457 , \5849 , \5822 );
nor \U$5597 ( \7458 , \7456 , \7457 );
xnor \U$5598 ( \7459 , \7458 , \5819 );
xor \U$5599 ( \7460 , \5579 , \7459 );
and \U$5600 ( \7461 , \6000 , \5861 );
and \U$5601 ( \7462 , \5909 , \5859 );
nor \U$5602 ( \7463 , \7461 , \7462 );
xnor \U$5603 ( \7464 , \7463 , \5887 );
xor \U$5604 ( \7465 , \7460 , \7464 );
xor \U$5605 ( \7466 , \7455 , \7465 );
xor \U$5606 ( \7467 , \7438 , \7466 );
and \U$5607 ( \7468 , \7391 , \7395 );
and \U$5608 ( \7469 , \7395 , \7400 );
and \U$5609 ( \7470 , \7391 , \7400 );
or \U$5610 ( \7471 , \7468 , \7469 , \7470 );
and \U$5611 ( \7472 , \7415 , \7419 );
and \U$5612 ( \7473 , \7419 , \7424 );
and \U$5613 ( \7474 , \7415 , \7424 );
or \U$5614 ( \7475 , \7472 , \7473 , \7474 );
xor \U$5615 ( \7476 , \7471 , \7475 );
and \U$5616 ( \7477 , \6163 , \5615 );
and \U$5617 ( \7478 , \6119 , \5613 );
nor \U$5618 ( \7479 , \7477 , \7478 );
xnor \U$5619 ( \7480 , \7479 , \5382 );
xor \U$5620 ( \7481 , \7476 , \7480 );
xor \U$5621 ( \7482 , \7467 , \7481 );
xor \U$5622 ( \7483 , \7434 , \7482 );
and \U$5623 ( \7484 , \7383 , \7427 );
nor \U$5624 ( \7485 , \7483 , \7484 );
nor \U$5625 ( \7486 , \7430 , \7485 );
nand \U$5626 ( \7487 , \7379 , \7486 );
and \U$5627 ( \7488 , \7438 , \7466 );
and \U$5628 ( \7489 , \7466 , \7481 );
and \U$5629 ( \7490 , \7438 , \7481 );
or \U$5630 ( \7491 , \7488 , \7489 , \7490 );
xor \U$5631 ( \7492 , \6351 , \6355 );
xor \U$5632 ( \7493 , \7492 , \6360 );
and \U$5633 ( \7494 , \5579 , \7459 );
and \U$5634 ( \7495 , \7459 , \7464 );
and \U$5635 ( \7496 , \5579 , \7464 );
or \U$5636 ( \7497 , \7494 , \7495 , \7496 );
and \U$5637 ( \7498 , \7444 , \7448 );
and \U$5638 ( \7499 , \7448 , \7453 );
and \U$5639 ( \7500 , \7444 , \7453 );
or \U$5640 ( \7501 , \7498 , \7499 , \7500 );
xor \U$5641 ( \7502 , \7497 , \7501 );
and \U$5642 ( \7503 , \6296 , \5553 );
and \U$5643 ( \7504 , \6163 , \5551 );
nor \U$5644 ( \7505 , \7503 , \7504 );
xnor \U$5645 ( \7506 , \7505 , \5579 );
xor \U$5646 ( \7507 , \7502 , \7506 );
xor \U$5647 ( \7508 , \7493 , \7507 );
xor \U$5648 ( \7509 , \7491 , \7508 );
and \U$5649 ( \7510 , \7471 , \7475 );
and \U$5650 ( \7511 , \7475 , \7480 );
and \U$5651 ( \7512 , \7471 , \7480 );
or \U$5652 ( \7513 , \7510 , \7511 , \7512 );
and \U$5653 ( \7514 , \7440 , \7454 );
and \U$5654 ( \7515 , \7454 , \7465 );
and \U$5655 ( \7516 , \7440 , \7465 );
or \U$5656 ( \7517 , \7514 , \7515 , \7516 );
xor \U$5657 ( \7518 , \7513 , \7517 );
xor \U$5658 ( \7519 , \6367 , \6371 );
xor \U$5659 ( \7520 , \7519 , \6376 );
xor \U$5660 ( \7521 , \7518 , \7520 );
xor \U$5661 ( \7522 , \7509 , \7521 );
and \U$5662 ( \7523 , \7434 , \7482 );
nor \U$5663 ( \7524 , \7522 , \7523 );
and \U$5664 ( \7525 , \7513 , \7517 );
and \U$5665 ( \7526 , \7517 , \7520 );
and \U$5666 ( \7527 , \7513 , \7520 );
or \U$5667 ( \7528 , \7525 , \7526 , \7527 );
and \U$5668 ( \7529 , \7493 , \7507 );
xor \U$5669 ( \7530 , \7528 , \7529 );
and \U$5670 ( \7531 , \7497 , \7501 );
and \U$5671 ( \7532 , \7501 , \7506 );
and \U$5672 ( \7533 , \7497 , \7506 );
or \U$5673 ( \7534 , \7531 , \7532 , \7533 );
xor \U$5674 ( \7535 , \6387 , \6389 );
xor \U$5675 ( \7536 , \7534 , \7535 );
xor \U$5676 ( \7537 , \6363 , \6379 );
xor \U$5677 ( \7538 , \7537 , \6382 );
xor \U$5678 ( \7539 , \7536 , \7538 );
xor \U$5679 ( \7540 , \7530 , \7539 );
and \U$5680 ( \7541 , \7491 , \7508 );
and \U$5681 ( \7542 , \7508 , \7521 );
and \U$5682 ( \7543 , \7491 , \7521 );
or \U$5683 ( \7544 , \7541 , \7542 , \7543 );
nor \U$5684 ( \7545 , \7540 , \7544 );
nor \U$5685 ( \7546 , \7524 , \7545 );
and \U$5686 ( \7547 , \7534 , \7535 );
and \U$5687 ( \7548 , \7535 , \7538 );
and \U$5688 ( \7549 , \7534 , \7538 );
or \U$5689 ( \7550 , \7547 , \7548 , \7549 );
xor \U$5690 ( \7551 , \6250 , \6266 );
xor \U$5691 ( \7552 , \7551 , \6301 );
xor \U$5692 ( \7553 , \7550 , \7552 );
xor \U$5693 ( \7554 , \6385 , \6390 );
xor \U$5694 ( \7555 , \7554 , \6393 );
xor \U$5695 ( \7556 , \7553 , \7555 );
and \U$5696 ( \7557 , \7528 , \7529 );
and \U$5697 ( \7558 , \7529 , \7539 );
and \U$5698 ( \7559 , \7528 , \7539 );
or \U$5699 ( \7560 , \7557 , \7558 , \7559 );
nor \U$5700 ( \7561 , \7556 , \7560 );
xor \U$5701 ( \7562 , \6396 , \6397 );
xor \U$5702 ( \7563 , \7562 , \6400 );
and \U$5703 ( \7564 , \7550 , \7552 );
and \U$5704 ( \7565 , \7552 , \7555 );
and \U$5705 ( \7566 , \7550 , \7555 );
or \U$5706 ( \7567 , \7564 , \7565 , \7566 );
nor \U$5707 ( \7568 , \7563 , \7567 );
nor \U$5708 ( \7569 , \7561 , \7568 );
nand \U$5709 ( \7570 , \7546 , \7569 );
nor \U$5710 ( \7571 , \7487 , \7570 );
and \U$5711 ( \7572 , \6140 , \5825 );
and \U$5712 ( \7573 , \6071 , \5822 );
nor \U$5713 ( \7574 , \7572 , \7573 );
xnor \U$5714 ( \7575 , \7574 , \5819 );
and \U$5715 ( \7576 , \5947 , \7575 );
and \U$5716 ( \7577 , \6163 , \5861 );
and \U$5717 ( \7578 , \6119 , \5859 );
nor \U$5718 ( \7579 , \7577 , \7578 );
xnor \U$5719 ( \7580 , \7579 , \5887 );
and \U$5720 ( \7581 , \7575 , \7580 );
and \U$5721 ( \7582 , \5947 , \7580 );
or \U$5722 ( \7583 , \7576 , \7581 , \7582 );
and \U$5723 ( \7584 , \6071 , \5825 );
and \U$5724 ( \7585 , \6092 , \5822 );
nor \U$5725 ( \7586 , \7584 , \7585 );
xnor \U$5726 ( \7587 , \7586 , \5819 );
and \U$5727 ( \7588 , \6119 , \5861 );
and \U$5728 ( \7589 , \6140 , \5859 );
nor \U$5729 ( \7590 , \7588 , \7589 );
xnor \U$5730 ( \7591 , \7590 , \5887 );
xor \U$5731 ( \7592 , \7587 , \7591 );
and \U$5732 ( \7593 , \6296 , \5921 );
and \U$5733 ( \7594 , \6163 , \5919 );
nor \U$5734 ( \7595 , \7593 , \7594 );
xnor \U$5735 ( \7596 , \7595 , \5947 );
xor \U$5736 ( \7597 , \7592 , \7596 );
xor \U$5737 ( \7598 , \7583 , \7597 );
nand \U$5738 ( \7599 , \6296 , \5919 );
xnor \U$5739 ( \7600 , \7599 , \5947 );
xor \U$5740 ( \7601 , \5947 , \7575 );
xor \U$5741 ( \7602 , \7601 , \7580 );
and \U$5742 ( \7603 , \7600 , \7602 );
nor \U$5743 ( \7604 , \7598 , \7603 );
and \U$5744 ( \7605 , \7587 , \7591 );
and \U$5745 ( \7606 , \7591 , \7596 );
and \U$5746 ( \7607 , \7587 , \7596 );
or \U$5747 ( \7608 , \7605 , \7606 , \7607 );
xor \U$5748 ( \7609 , \7318 , \7320 );
xor \U$5749 ( \7610 , \7608 , \7609 );
xor \U$5750 ( \7611 , \6005 , \7306 );
xor \U$5751 ( \7612 , \7611 , \7311 );
xor \U$5752 ( \7613 , \7610 , \7612 );
and \U$5753 ( \7614 , \7583 , \7597 );
nor \U$5754 ( \7615 , \7613 , \7614 );
nor \U$5755 ( \7616 , \7604 , \7615 );
xor \U$5756 ( \7617 , \7229 , \7233 );
xor \U$5757 ( \7618 , \7617 , \7238 );
xor \U$5758 ( \7619 , \7314 , \7321 );
xor \U$5759 ( \7620 , \7619 , \7326 );
xor \U$5760 ( \7621 , \7618 , \7620 );
and \U$5761 ( \7622 , \7608 , \7609 );
and \U$5762 ( \7623 , \7609 , \7612 );
and \U$5763 ( \7624 , \7608 , \7612 );
or \U$5764 ( \7625 , \7622 , \7623 , \7624 );
nor \U$5765 ( \7626 , \7621 , \7625 );
xor \U$5766 ( \7627 , \7329 , \7331 );
and \U$5767 ( \7628 , \7618 , \7620 );
nor \U$5768 ( \7629 , \7627 , \7628 );
nor \U$5769 ( \7630 , \7626 , \7629 );
nand \U$5770 ( \7631 , \7616 , \7630 );
and \U$5771 ( \7632 , \6119 , \5825 );
and \U$5772 ( \7633 , \6140 , \5822 );
nor \U$5773 ( \7634 , \7632 , \7633 );
xnor \U$5774 ( \7635 , \7634 , \5819 );
and \U$5775 ( \7636 , \6296 , \5861 );
and \U$5776 ( \7637 , \6163 , \5859 );
nor \U$5777 ( \7638 , \7636 , \7637 );
xnor \U$5778 ( \7639 , \7638 , \5887 );
xor \U$5779 ( \7640 , \7635 , \7639 );
and \U$5780 ( \7641 , \6163 , \5825 );
and \U$5781 ( \7642 , \6119 , \5822 );
nor \U$5782 ( \7643 , \7641 , \7642 );
xnor \U$5783 ( \7644 , \7643 , \5819 );
and \U$5784 ( \7645 , \7644 , \5887 );
nor \U$5785 ( \7646 , \7640 , \7645 );
xor \U$5786 ( \7647 , \7600 , \7602 );
and \U$5787 ( \7648 , \7635 , \7639 );
nor \U$5788 ( \7649 , \7647 , \7648 );
nor \U$5789 ( \7650 , \7646 , \7649 );
xor \U$5790 ( \7651 , \7644 , \5887 );
nand \U$5791 ( \7652 , \6296 , \5859 );
xnor \U$5792 ( \7653 , \7652 , \5887 );
nor \U$5793 ( \7654 , \7651 , \7653 );
and \U$5794 ( \7655 , \6296 , \5825 );
and \U$5795 ( \7656 , \6163 , \5822 );
nor \U$5796 ( \7657 , \7655 , \7656 );
xnor \U$5797 ( \7658 , \7657 , \5819 );
nand \U$5798 ( \7659 , \6296 , \5822 );
xnor \U$5799 ( \7660 , \7659 , \5819 );
and \U$5800 ( \7661 , \7660 , \5819 );
nand \U$5801 ( \7662 , \7658 , \7661 );
or \U$5802 ( \7663 , \7654 , \7662 );
nand \U$5803 ( \7664 , \7651 , \7653 );
nand \U$5804 ( \7665 , \7663 , \7664 );
and \U$5805 ( \7666 , \7650 , \7665 );
nand \U$5806 ( \7667 , \7640 , \7645 );
or \U$5807 ( \7668 , \7649 , \7667 );
nand \U$5808 ( \7669 , \7647 , \7648 );
nand \U$5809 ( \7670 , \7668 , \7669 );
nor \U$5810 ( \7671 , \7666 , \7670 );
or \U$5811 ( \7672 , \7631 , \7671 );
nand \U$5812 ( \7673 , \7598 , \7603 );
or \U$5813 ( \7674 , \7615 , \7673 );
nand \U$5814 ( \7675 , \7613 , \7614 );
nand \U$5815 ( \7676 , \7674 , \7675 );
and \U$5816 ( \7677 , \7630 , \7676 );
nand \U$5817 ( \7678 , \7621 , \7625 );
or \U$5818 ( \7679 , \7629 , \7678 );
nand \U$5819 ( \7680 , \7627 , \7628 );
nand \U$5820 ( \7681 , \7679 , \7680 );
nor \U$5821 ( \7682 , \7677 , \7681 );
nand \U$5822 ( \7683 , \7672 , \7682 );
and \U$5823 ( \7684 , \7571 , \7683 );
nand \U$5824 ( \7685 , \7302 , \7332 );
or \U$5825 ( \7686 , \7378 , \7685 );
nand \U$5826 ( \7687 , \7373 , \7377 );
nand \U$5827 ( \7688 , \7686 , \7687 );
and \U$5828 ( \7689 , \7486 , \7688 );
nand \U$5829 ( \7690 , \7428 , \7429 );
or \U$5830 ( \7691 , \7485 , \7690 );
nand \U$5831 ( \7692 , \7483 , \7484 );
nand \U$5832 ( \7693 , \7691 , \7692 );
nor \U$5833 ( \7694 , \7689 , \7693 );
or \U$5834 ( \7695 , \7570 , \7694 );
nand \U$5835 ( \7696 , \7522 , \7523 );
or \U$5836 ( \7697 , \7545 , \7696 );
nand \U$5837 ( \7698 , \7540 , \7544 );
nand \U$5838 ( \7699 , \7697 , \7698 );
and \U$5839 ( \7700 , \7569 , \7699 );
nand \U$5840 ( \7701 , \7556 , \7560 );
or \U$5841 ( \7702 , \7568 , \7701 );
nand \U$5842 ( \7703 , \7563 , \7567 );
nand \U$5843 ( \7704 , \7702 , \7703 );
nor \U$5844 ( \7705 , \7700 , \7704 );
nand \U$5845 ( \7706 , \7695 , \7705 );
nor \U$5846 ( \7707 , \7684 , \7706 );
or \U$5847 ( \7708 , \7225 , \7707 );
nand \U$5848 ( \7709 , \6347 , \6403 );
or \U$5849 ( \7710 , \6479 , \7709 );
nand \U$5850 ( \7711 , \6477 , \6478 );
nand \U$5851 ( \7712 , \7710 , \7711 );
and \U$5852 ( \7713 , \6632 , \7712 );
nand \U$5853 ( \7714 , \6554 , \6555 );
or \U$5854 ( \7715 , \6631 , \7714 );
nand \U$5855 ( \7716 , \6626 , \6630 );
nand \U$5856 ( \7717 , \7715 , \7716 );
nor \U$5857 ( \7718 , \7713 , \7717 );
or \U$5858 ( \7719 , \6928 , \7718 );
nand \U$5859 ( \7720 , \6703 , \6707 );
or \U$5860 ( \7721 , \6784 , \7720 );
nand \U$5861 ( \7722 , \6779 , \6783 );
nand \U$5862 ( \7723 , \7721 , \7722 );
and \U$5863 ( \7724 , \6927 , \7723 );
nand \U$5864 ( \7725 , \6852 , \6856 );
or \U$5865 ( \7726 , \6926 , \7725 );
nand \U$5866 ( \7727 , \6921 , \6925 );
nand \U$5867 ( \7728 , \7726 , \7727 );
nor \U$5868 ( \7729 , \7724 , \7728 );
nand \U$5869 ( \7730 , \7719 , \7729 );
and \U$5870 ( \7731 , \7224 , \7730 );
nand \U$5871 ( \7732 , \6985 , \6989 );
or \U$5872 ( \7733 , \7050 , \7732 );
nand \U$5873 ( \7734 , \7045 , \7049 );
nand \U$5874 ( \7735 , \7733 , \7734 );
and \U$5875 ( \7736 , \7146 , \7735 );
nand \U$5876 ( \7737 , \7102 , \7106 );
or \U$5877 ( \7738 , \7145 , \7737 );
nand \U$5878 ( \7739 , \7140 , \7144 );
nand \U$5879 ( \7740 , \7738 , \7739 );
nor \U$5880 ( \7741 , \7736 , \7740 );
or \U$5881 ( \7742 , \7223 , \7741 );
nand \U$5882 ( \7743 , \7172 , \7176 );
or \U$5883 ( \7744 , \7198 , \7743 );
nand \U$5884 ( \7745 , \7193 , \7197 );
nand \U$5885 ( \7746 , \7744 , \7745 );
and \U$5886 ( \7747 , \7222 , \7746 );
nand \U$5887 ( \7748 , \7209 , \7213 );
or \U$5888 ( \7749 , \7221 , \7748 );
nand \U$5889 ( \7750 , \7216 , \7220 );
nand \U$5890 ( \7751 , \7749 , \7750 );
nor \U$5891 ( \7752 , \7747 , \7751 );
nand \U$5892 ( \7753 , \7742 , \7752 );
nor \U$5893 ( \7754 , \7731 , \7753 );
nand \U$5894 ( \7755 , \7708 , \7754 );
not \U$5895 ( \7756 , \7755 );
xor \U$5896 ( \7757 , \5815 , \7756 );
buf g32b2_GF_PartitionCandidate( \7758_nG32b2 , \7757 );
buf \U$5897 ( \7759 , RI994e460_14);
buf \U$5898 ( \7760 , RI994e3e8_15);
buf \U$5899 ( \7761 , RI994e370_16);
buf \U$5900 ( \7762 , RI994e2f8_17);
buf \U$5901 ( \7763 , RI994e280_18);
buf \U$5902 ( \7764 , RI994e208_19);
buf \U$5903 ( \7765 , RI994e190_20);
buf \U$5904 ( \7766 , RI994e118_21);
buf \U$5905 ( \7767 , RI994e0a0_22);
buf \U$5906 ( \7768 , RI994e028_23);
buf \U$5907 ( \7769 , RI994dfb0_24);
buf \U$5908 ( \7770 , RI994df38_25);
not \U$5909 ( \7771 , RI99216b8_614);
buf \U$5910 ( \7772 , \7771 );
and \U$5911 ( \7773 , \7770 , \7772 );
and \U$5912 ( \7774 , \7769 , \7773 );
and \U$5913 ( \7775 , \7768 , \7774 );
and \U$5914 ( \7776 , \7767 , \7775 );
and \U$5915 ( \7777 , \7766 , \7776 );
and \U$5916 ( \7778 , \7765 , \7777 );
and \U$5917 ( \7779 , \7764 , \7778 );
and \U$5918 ( \7780 , \7763 , \7779 );
and \U$5919 ( \7781 , \7762 , \7780 );
and \U$5920 ( \7782 , \7761 , \7781 );
and \U$5921 ( \7783 , \7760 , \7782 );
xor \U$5922 ( \7784 , \7759 , \7783 );
buf \U$5923 ( \7785 , \7784 );
buf \U$5924 ( \7786 , \7785 );
not \U$5925 ( \7787 , \7786 );
nor \U$5926 ( \7788 , \4955 , \4959 , \4963 , \4967 , \4972 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5927 ( \7789 , RI995e4c8_235, \7788 );
nor \U$5928 ( \7790 , \5007 , \5008 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5929 ( \7791 , RI99670f0_222, \7790 );
nor \U$5930 ( \7792 , \4955 , \5008 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5931 ( \7793 , RI890f600_209, \7792 );
nor \U$5932 ( \7794 , \5007 , \4959 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5933 ( \7795 , RI89185e8_196, \7794 );
nor \U$5934 ( \7796 , \4955 , \4959 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5935 ( \7797 , RI8924e10_183, \7796 );
nor \U$5936 ( \7798 , \5007 , \5008 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5937 ( \7799 , RI8930828_170, \7798 );
nor \U$5938 ( \7800 , \4955 , \5008 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5939 ( \7801 , RI8939810_157, \7800 );
nor \U$5940 ( \7802 , \5007 , \4959 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5941 ( \7803 , RI8946038_144, \7802 );
nor \U$5942 ( \7804 , \4955 , \4959 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5943 ( \7805 , RI89ec0a0_131, \7804 );
nor \U$5944 ( \7806 , \5007 , \5008 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5945 ( \7807 , RI89ec6b8_118, \7806 );
nor \U$5946 ( \7808 , \4955 , \5008 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5947 ( \7809 , RI9776ff8_105, \7808 );
nor \U$5948 ( \7810 , \5007 , \4959 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5949 ( \7811 , RI98084f8_92, \7810 );
nor \U$5950 ( \7812 , \4955 , \4959 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5951 ( \7813 , RI9808b10_79, \7812 );
nor \U$5952 ( \7814 , \5007 , \5008 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5953 ( \7815 , RI98197a8_66, \7814 );
nor \U$5954 ( \7816 , \4955 , \5008 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5955 ( \7817 , RI98abcb0_53, \7816 );
nor \U$5956 ( \7818 , \5007 , \4959 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5957 ( \7819 , RI98bc948_40, \7818 );
nor \U$5958 ( \7820 , \4955 , \4959 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$5959 ( \7821 , RI994de48_27, \7820 );
or \U$5960 ( \7822 , \7789 , \7791 , \7793 , \7795 , \7797 , \7799 , \7801 , \7803 , \7805 , \7807 , \7809 , \7811 , \7813 , \7815 , \7817 , \7819 , \7821 );
buf \U$5961 ( \7823 , \4976 );
buf \U$5962 ( \7824 , \4980 );
buf \U$5963 ( \7825 , \4984 );
buf \U$5964 ( \7826 , \4988 );
buf \U$5965 ( \7827 , \4992 );
buf \U$5966 ( \7828 , \4996 );
buf \U$5967 ( \7829 , \5000 );
buf \U$5968 ( \7830 , \5004 );
buf \U$5969 ( \7831 , \4971 );
buf \U$5970 ( \7832 , \4955 );
buf \U$5971 ( \7833 , \4959 );
buf \U$5972 ( \7834 , \4963 );
buf \U$5973 ( \7835 , \4967 );
or \U$5974 ( \7836 , \7832 , \7833 , \7834 , \7835 );
and \U$5975 ( \7837 , \7831 , \7836 );
or \U$5976 ( \7838 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7837 );
buf \U$5977 ( \7839 , \7838 );
_DC g1080 ( \7840_nG1080 , \7822 , \7839 );
buf \U$5978 ( \7841 , \7840_nG1080 );
and \U$5979 ( \7842 , \7787 , \7841 );
xor \U$5980 ( \7843 , \7760 , \7782 );
buf \U$5981 ( \7844 , \7843 );
buf \U$5982 ( \7845 , \7844 );
not \U$5983 ( \7846 , \7845 );
and \U$5984 ( \7847 , RI995e450_236, \7788 );
and \U$5985 ( \7848 , RI9967078_223, \7790 );
and \U$5986 ( \7849 , RI9967690_210, \7792 );
and \U$5987 ( \7850 , RI890fba0_197, \7794 );
and \U$5988 ( \7851 , RI8918b88_184, \7796 );
and \U$5989 ( \7852 , RI89253b0_171, \7798 );
and \U$5990 ( \7853 , RI8930dc8_158, \7800 );
and \U$5991 ( \7854 , RI8939db0_145, \7802 );
and \U$5992 ( \7855 , RI89465d8_132, \7804 );
and \U$5993 ( \7856 , RI89ec640_119, \7806 );
and \U$5994 ( \7857 , RI9776f80_106, \7808 );
and \U$5995 ( \7858 , RI9808480_93, \7810 );
and \U$5996 ( \7859 , RI9808a98_80, \7812 );
and \U$5997 ( \7860 , RI9819730_67, \7814 );
and \U$5998 ( \7861 , RI98abc38_54, \7816 );
and \U$5999 ( \7862 , RI98bc8d0_41, \7818 );
and \U$6000 ( \7863 , RI994ddd0_28, \7820 );
or \U$6001 ( \7864 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 );
_DC g1099 ( \7865_nG1099 , \7864 , \7839 );
buf \U$6002 ( \7866 , \7865_nG1099 );
and \U$6003 ( \7867 , \7846 , \7866 );
xor \U$6004 ( \7868 , \7761 , \7781 );
buf \U$6005 ( \7869 , \7868 );
buf \U$6006 ( \7870 , \7869 );
not \U$6007 ( \7871 , \7870 );
and \U$6008 ( \7872 , RI995e3d8_237, \7788 );
and \U$6009 ( \7873 , RI99669e8_224, \7790 );
and \U$6010 ( \7874 , RI9967618_211, \7792 );
and \U$6011 ( \7875 , RI890fb28_198, \7794 );
and \U$6012 ( \7876 , RI8918b10_185, \7796 );
and \U$6013 ( \7877 , RI8925338_172, \7798 );
and \U$6014 ( \7878 , RI8930d50_159, \7800 );
and \U$6015 ( \7879 , RI8939d38_146, \7802 );
and \U$6016 ( \7880 , RI8946560_133, \7804 );
and \U$6017 ( \7881 , RI89ec5c8_120, \7806 );
and \U$6018 ( \7882 , RI9776f08_107, \7808 );
and \U$6019 ( \7883 , RI9808408_94, \7810 );
and \U$6020 ( \7884 , RI9808a20_81, \7812 );
and \U$6021 ( \7885 , RI98196b8_68, \7814 );
and \U$6022 ( \7886 , RI98abbc0_55, \7816 );
and \U$6023 ( \7887 , RI98bc858_42, \7818 );
and \U$6024 ( \7888 , RI994dd58_29, \7820 );
or \U$6025 ( \7889 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 );
_DC g10b2 ( \7890_nG10b2 , \7889 , \7839 );
buf \U$6026 ( \7891 , \7890_nG10b2 );
and \U$6027 ( \7892 , \7871 , \7891 );
xor \U$6028 ( \7893 , \7762 , \7780 );
buf \U$6029 ( \7894 , \7893 );
buf \U$6030 ( \7895 , \7894 );
not \U$6031 ( \7896 , \7895 );
and \U$6032 ( \7897 , RI9959fe0_238, \7788 );
and \U$6033 ( \7898 , RI995e978_225, \7790 );
and \U$6034 ( \7899 , RI99675a0_212, \7792 );
and \U$6035 ( \7900 , RI890fab0_199, \7794 );
and \U$6036 ( \7901 , RI8918a98_186, \7796 );
and \U$6037 ( \7902 , RI89252c0_173, \7798 );
and \U$6038 ( \7903 , RI8930cd8_160, \7800 );
and \U$6039 ( \7904 , RI8939cc0_147, \7802 );
and \U$6040 ( \7905 , RI89464e8_134, \7804 );
and \U$6041 ( \7906 , RI89ec550_121, \7806 );
and \U$6042 ( \7907 , RI9776e90_108, \7808 );
and \U$6043 ( \7908 , RI9808390_95, \7810 );
and \U$6044 ( \7909 , RI98089a8_82, \7812 );
and \U$6045 ( \7910 , RI9819640_69, \7814 );
and \U$6046 ( \7911 , RI98abb48_56, \7816 );
and \U$6047 ( \7912 , RI98bc7e0_43, \7818 );
and \U$6048 ( \7913 , RI994dce0_30, \7820 );
or \U$6049 ( \7914 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 );
_DC g10cb ( \7915_nG10cb , \7914 , \7839 );
buf \U$6050 ( \7916 , \7915_nG10cb );
and \U$6051 ( \7917 , \7896 , \7916 );
xor \U$6052 ( \7918 , \7763 , \7779 );
buf \U$6053 ( \7919 , \7918 );
buf \U$6054 ( \7920 , \7919 );
not \U$6055 ( \7921 , \7920 );
and \U$6056 ( \7922 , RI9959f68_239, \7788 );
and \U$6057 ( \7923 , RI995e900_226, \7790 );
and \U$6058 ( \7924 , RI9967528_213, \7792 );
and \U$6059 ( \7925 , RI890fa38_200, \7794 );
and \U$6060 ( \7926 , RI8918a20_187, \7796 );
and \U$6061 ( \7927 , RI8925248_174, \7798 );
and \U$6062 ( \7928 , RI8930c60_161, \7800 );
and \U$6063 ( \7929 , RI8939c48_148, \7802 );
and \U$6064 ( \7930 , RI8946470_135, \7804 );
and \U$6065 ( \7931 , RI89ec4d8_122, \7806 );
and \U$6066 ( \7932 , RI9776e18_109, \7808 );
and \U$6067 ( \7933 , RI9808318_96, \7810 );
and \U$6068 ( \7934 , RI9808930_83, \7812 );
and \U$6069 ( \7935 , RI98195c8_70, \7814 );
and \U$6070 ( \7936 , RI98abad0_57, \7816 );
and \U$6071 ( \7937 , RI98bc768_44, \7818 );
and \U$6072 ( \7938 , RI994dc68_31, \7820 );
or \U$6073 ( \7939 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 );
_DC g10e4 ( \7940_nG10e4 , \7939 , \7839 );
buf \U$6074 ( \7941 , \7940_nG10e4 );
and \U$6075 ( \7942 , \7921 , \7941 );
xor \U$6076 ( \7943 , \7764 , \7778 );
buf \U$6077 ( \7944 , \7943 );
buf \U$6078 ( \7945 , \7944 );
not \U$6079 ( \7946 , \7945 );
and \U$6080 ( \7947 , RI9959860_240, \7788 );
and \U$6081 ( \7948 , RI995e888_227, \7790 );
and \U$6082 ( \7949 , RI99674b0_214, \7792 );
and \U$6083 ( \7950 , RI890f9c0_201, \7794 );
and \U$6084 ( \7951 , RI89189a8_188, \7796 );
and \U$6085 ( \7952 , RI89251d0_175, \7798 );
and \U$6086 ( \7953 , RI8930be8_162, \7800 );
and \U$6087 ( \7954 , RI8939bd0_149, \7802 );
and \U$6088 ( \7955 , RI89463f8_136, \7804 );
and \U$6089 ( \7956 , RI89ec460_123, \7806 );
and \U$6090 ( \7957 , RI9776da0_110, \7808 );
and \U$6091 ( \7958 , RI98082a0_97, \7810 );
and \U$6092 ( \7959 , RI98088b8_84, \7812 );
and \U$6093 ( \7960 , RI9819550_71, \7814 );
and \U$6094 ( \7961 , RI98aba58_58, \7816 );
and \U$6095 ( \7962 , RI98bc6f0_45, \7818 );
and \U$6096 ( \7963 , RI994dbf0_32, \7820 );
or \U$6097 ( \7964 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 );
_DC g10fd ( \7965_nG10fd , \7964 , \7839 );
buf \U$6098 ( \7966 , \7965_nG10fd );
and \U$6099 ( \7967 , \7946 , \7966 );
xor \U$6100 ( \7968 , \7765 , \7777 );
buf \U$6101 ( \7969 , \7968 );
buf \U$6102 ( \7970 , \7969 );
not \U$6103 ( \7971 , \7970 );
and \U$6104 ( \7972 , RI994d998_241, \7788 );
and \U$6105 ( \7973 , RI995e810_228, \7790 );
and \U$6106 ( \7974 , RI9967438_215, \7792 );
and \U$6107 ( \7975 , RI890f948_202, \7794 );
and \U$6108 ( \7976 , RI8918930_189, \7796 );
and \U$6109 ( \7977 , RI8925158_176, \7798 );
and \U$6110 ( \7978 , RI8930b70_163, \7800 );
and \U$6111 ( \7979 , RI8939b58_150, \7802 );
and \U$6112 ( \7980 , RI8946380_137, \7804 );
and \U$6113 ( \7981 , RI89ec3e8_124, \7806 );
and \U$6114 ( \7982 , RI9776d28_111, \7808 );
and \U$6115 ( \7983 , RI9808228_98, \7810 );
and \U$6116 ( \7984 , RI9808840_85, \7812 );
and \U$6117 ( \7985 , RI98194d8_72, \7814 );
and \U$6118 ( \7986 , RI98ab9e0_59, \7816 );
and \U$6119 ( \7987 , RI98abff8_46, \7818 );
and \U$6120 ( \7988 , RI98bcc90_33, \7820 );
or \U$6121 ( \7989 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 );
_DC g1116 ( \7990_nG1116 , \7989 , \7839 );
buf \U$6122 ( \7991 , \7990_nG1116 );
and \U$6123 ( \7992 , \7971 , \7991 );
xor \U$6124 ( \7993 , \7766 , \7776 );
buf \U$6125 ( \7994 , \7993 );
buf \U$6126 ( \7995 , \7994 );
not \U$6127 ( \7996 , \7995 );
and \U$6128 ( \7997 , RI994d920_242, \7788 );
and \U$6129 ( \7998 , RI995e798_229, \7790 );
and \U$6130 ( \7999 , RI99673c0_216, \7792 );
and \U$6131 ( \8000 , RI890f8d0_203, \7794 );
and \U$6132 ( \8001 , RI89188b8_190, \7796 );
and \U$6133 ( \8002 , RI89250e0_177, \7798 );
and \U$6134 ( \8003 , RI8930af8_164, \7800 );
and \U$6135 ( \8004 , RI8939ae0_151, \7802 );
and \U$6136 ( \8005 , RI8946308_138, \7804 );
and \U$6137 ( \8006 , RI89ec370_125, \7806 );
and \U$6138 ( \8007 , RI89ec988_112, \7808 );
and \U$6139 ( \8008 , RI97772c8_99, \7810 );
and \U$6140 ( \8009 , RI98087c8_86, \7812 );
and \U$6141 ( \8010 , RI9819460_73, \7814 );
and \U$6142 ( \8011 , RI98ab968_60, \7816 );
and \U$6143 ( \8012 , RI98abf80_47, \7818 );
and \U$6144 ( \8013 , RI98bcc18_34, \7820 );
or \U$6145 ( \8014 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 );
_DC g112f ( \8015_nG112f , \8014 , \7839 );
buf \U$6146 ( \8016 , \8015_nG112f );
and \U$6147 ( \8017 , \7996 , \8016 );
xor \U$6148 ( \8018 , \7767 , \7775 );
buf \U$6149 ( \8019 , \8018 );
buf \U$6150 ( \8020 , \8019 );
not \U$6151 ( \8021 , \8020 );
and \U$6152 ( \8022 , RI994d8a8_243, \7788 );
and \U$6153 ( \8023 , RI995e720_230, \7790 );
and \U$6154 ( \8024 , RI9967348_217, \7792 );
and \U$6155 ( \8025 , RI890f858_204, \7794 );
and \U$6156 ( \8026 , RI8918840_191, \7796 );
and \U$6157 ( \8027 , RI8925068_178, \7798 );
and \U$6158 ( \8028 , RI8930a80_165, \7800 );
and \U$6159 ( \8029 , RI8939a68_152, \7802 );
and \U$6160 ( \8030 , RI8946290_139, \7804 );
and \U$6161 ( \8031 , RI89ec2f8_126, \7806 );
and \U$6162 ( \8032 , RI89ec910_113, \7808 );
and \U$6163 ( \8033 , RI9777250_100, \7810 );
and \U$6164 ( \8034 , RI9808750_87, \7812 );
and \U$6165 ( \8035 , RI98193e8_74, \7814 );
and \U$6166 ( \8036 , RI98ab8f0_61, \7816 );
and \U$6167 ( \8037 , RI98abf08_48, \7818 );
and \U$6168 ( \8038 , RI98bcba0_35, \7820 );
or \U$6169 ( \8039 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 );
_DC g1148 ( \8040_nG1148 , \8039 , \7839 );
buf \U$6170 ( \8041 , \8040_nG1148 );
and \U$6171 ( \8042 , \8021 , \8041 );
xor \U$6172 ( \8043 , \7768 , \7774 );
buf \U$6173 ( \8044 , \8043 );
buf \U$6174 ( \8045 , \8044 );
not \U$6175 ( \8046 , \8045 );
and \U$6176 ( \8047 , RI994d830_244, \7788 );
and \U$6177 ( \8048 , RI995e6a8_231, \7790 );
and \U$6178 ( \8049 , RI99672d0_218, \7792 );
and \U$6179 ( \8050 , RI890f7e0_205, \7794 );
and \U$6180 ( \8051 , RI89187c8_192, \7796 );
and \U$6181 ( \8052 , RI8924ff0_179, \7798 );
and \U$6182 ( \8053 , RI8930a08_166, \7800 );
and \U$6183 ( \8054 , RI89399f0_153, \7802 );
and \U$6184 ( \8055 , RI8946218_140, \7804 );
and \U$6185 ( \8056 , RI89ec280_127, \7806 );
and \U$6186 ( \8057 , RI89ec898_114, \7808 );
and \U$6187 ( \8058 , RI97771d8_101, \7810 );
and \U$6188 ( \8059 , RI98086d8_88, \7812 );
and \U$6189 ( \8060 , RI9819370_75, \7814 );
and \U$6190 ( \8061 , RI98ab878_62, \7816 );
and \U$6191 ( \8062 , RI98abe90_49, \7818 );
and \U$6192 ( \8063 , RI98bcb28_36, \7820 );
or \U$6193 ( \8064 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 );
_DC g1161 ( \8065_nG1161 , \8064 , \7839 );
buf \U$6194 ( \8066 , \8065_nG1161 );
and \U$6195 ( \8067 , \8046 , \8066 );
xor \U$6196 ( \8068 , \7769 , \7773 );
buf \U$6197 ( \8069 , \8068 );
buf \U$6198 ( \8070 , \8069 );
not \U$6199 ( \8071 , \8070 );
and \U$6200 ( \8072 , RI994d7b8_245, \7788 );
and \U$6201 ( \8073 , RI995e630_232, \7790 );
and \U$6202 ( \8074 , RI9967258_219, \7792 );
and \U$6203 ( \8075 , RI890f768_206, \7794 );
and \U$6204 ( \8076 , RI8918750_193, \7796 );
and \U$6205 ( \8077 , RI8924f78_180, \7798 );
and \U$6206 ( \8078 , RI8930990_167, \7800 );
and \U$6207 ( \8079 , RI8939978_154, \7802 );
and \U$6208 ( \8080 , RI89461a0_141, \7804 );
and \U$6209 ( \8081 , RI89ec208_128, \7806 );
and \U$6210 ( \8082 , RI89ec820_115, \7808 );
and \U$6211 ( \8083 , RI9777160_102, \7810 );
and \U$6212 ( \8084 , RI9808660_89, \7812 );
and \U$6213 ( \8085 , RI98192f8_76, \7814 );
and \U$6214 ( \8086 , RI98ab800_63, \7816 );
and \U$6215 ( \8087 , RI98abe18_50, \7818 );
and \U$6216 ( \8088 , RI98bcab0_37, \7820 );
or \U$6217 ( \8089 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 );
_DC g117a ( \8090_nG117a , \8089 , \7839 );
buf \U$6218 ( \8091 , \8090_nG117a );
and \U$6219 ( \8092 , \8071 , \8091 );
xor \U$6220 ( \8093 , \7770 , \7772 );
buf \U$6221 ( \8094 , \8093 );
buf \U$6222 ( \8095 , \8094 );
not \U$6223 ( \8096 , \8095 );
and \U$6224 ( \8097 , RI994d740_246, \7788 );
and \U$6225 ( \8098 , RI995e5b8_233, \7790 );
and \U$6226 ( \8099 , RI99671e0_220, \7792 );
and \U$6227 ( \8100 , RI890f6f0_207, \7794 );
and \U$6228 ( \8101 , RI89186d8_194, \7796 );
and \U$6229 ( \8102 , RI8924f00_181, \7798 );
and \U$6230 ( \8103 , RI8930918_168, \7800 );
and \U$6231 ( \8104 , RI8939900_155, \7802 );
and \U$6232 ( \8105 , RI8946128_142, \7804 );
and \U$6233 ( \8106 , RI89ec190_129, \7806 );
and \U$6234 ( \8107 , RI89ec7a8_116, \7808 );
and \U$6235 ( \8108 , RI97770e8_103, \7810 );
and \U$6236 ( \8109 , RI98085e8_90, \7812 );
and \U$6237 ( \8110 , RI9819280_77, \7814 );
and \U$6238 ( \8111 , RI98ab788_64, \7816 );
and \U$6239 ( \8112 , RI98abda0_51, \7818 );
and \U$6240 ( \8113 , RI98bca38_38, \7820 );
or \U$6241 ( \8114 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 );
_DC g1193 ( \8115_nG1193 , \8114 , \7839 );
buf \U$6242 ( \8116 , \8115_nG1193 );
and \U$6243 ( \8117 , \8096 , \8116 );
buf \U$6244 ( \8118 , RI994dec0_26);
buf \U$6247 ( \8119 , \8118 );
not \U$6248 ( \8120 , \8119 );
and \U$6249 ( \8121 , RI994d6c8_247, \7788 );
and \U$6250 ( \8122 , RI995e540_234, \7790 );
and \U$6251 ( \8123 , RI9967168_221, \7792 );
and \U$6252 ( \8124 , RI890f678_208, \7794 );
and \U$6253 ( \8125 , RI8918660_195, \7796 );
and \U$6254 ( \8126 , RI8924e88_182, \7798 );
and \U$6255 ( \8127 , RI89308a0_169, \7800 );
and \U$6256 ( \8128 , RI8939888_156, \7802 );
and \U$6257 ( \8129 , RI89460b0_143, \7804 );
and \U$6258 ( \8130 , RI89ec118_130, \7806 );
and \U$6259 ( \8131 , RI89ec730_117, \7808 );
and \U$6260 ( \8132 , RI9777070_104, \7810 );
and \U$6261 ( \8133 , RI9808570_91, \7812 );
and \U$6262 ( \8134 , RI9819208_78, \7814 );
and \U$6263 ( \8135 , RI98ab710_65, \7816 );
and \U$6264 ( \8136 , RI98abd28_52, \7818 );
and \U$6265 ( \8137 , RI98bc9c0_39, \7820 );
or \U$6266 ( \8138 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 );
_DC g11ad ( \8139_nG11ad , \8138 , \7839 );
buf \U$6267 ( \8140 , \8139_nG11ad );
and \U$6268 ( \8141 , \8120 , \8140 );
xnor \U$6269 ( \8142 , \8095 , \8116 );
and \U$6270 ( \8143 , \8141 , \8142 );
or \U$6271 ( \8144 , \8117 , \8143 );
xnor \U$6272 ( \8145 , \8070 , \8091 );
and \U$6273 ( \8146 , \8144 , \8145 );
or \U$6274 ( \8147 , \8092 , \8146 );
xnor \U$6275 ( \8148 , \8045 , \8066 );
and \U$6276 ( \8149 , \8147 , \8148 );
or \U$6277 ( \8150 , \8067 , \8149 );
xnor \U$6278 ( \8151 , \8020 , \8041 );
and \U$6279 ( \8152 , \8150 , \8151 );
or \U$6280 ( \8153 , \8042 , \8152 );
xnor \U$6281 ( \8154 , \7995 , \8016 );
and \U$6282 ( \8155 , \8153 , \8154 );
or \U$6283 ( \8156 , \8017 , \8155 );
xnor \U$6284 ( \8157 , \7970 , \7991 );
and \U$6285 ( \8158 , \8156 , \8157 );
or \U$6286 ( \8159 , \7992 , \8158 );
xnor \U$6287 ( \8160 , \7945 , \7966 );
and \U$6288 ( \8161 , \8159 , \8160 );
or \U$6289 ( \8162 , \7967 , \8161 );
xnor \U$6290 ( \8163 , \7920 , \7941 );
and \U$6291 ( \8164 , \8162 , \8163 );
or \U$6292 ( \8165 , \7942 , \8164 );
xnor \U$6293 ( \8166 , \7895 , \7916 );
and \U$6294 ( \8167 , \8165 , \8166 );
or \U$6295 ( \8168 , \7917 , \8167 );
xnor \U$6296 ( \8169 , \7870 , \7891 );
and \U$6297 ( \8170 , \8168 , \8169 );
or \U$6298 ( \8171 , \7892 , \8170 );
xnor \U$6299 ( \8172 , \7845 , \7866 );
and \U$6300 ( \8173 , \8171 , \8172 );
or \U$6301 ( \8174 , \7867 , \8173 );
xnor \U$6302 ( \8175 , \7786 , \7841 );
and \U$6303 ( \8176 , \8174 , \8175 );
or \U$6304 ( \8177 , \7842 , \8176 );
not \U$6305 ( \8178 , \8177 );
buf \U$6306 ( \8179 , \8178 );
buf \U$6307 ( \8180 , RI9921910_609);
buf \U$6308 ( \8181 , RI9921988_608);
buf \U$6309 ( \8182 , RI9921a00_607);
buf \U$6310 ( \8183 , RI9921a78_606);
buf \U$6311 ( \8184 , RI9921af0_605);
buf \U$6312 ( \8185 , RI9921b68_604);
buf \U$6313 ( \8186 , RI9921be0_603);
buf \U$6314 ( \8187 , RI9921c58_602);
buf \U$6315 ( \8188 , RI9921cd0_601);
buf \U$6316 ( \8189 , RI9921730_613);
buf \U$6317 ( \8190 , RI99217a8_612);
buf \U$6318 ( \8191 , RI9921820_611);
buf \U$6319 ( \8192 , RI9921898_610);
and \U$6320 ( \8193 , \8189 , \8190 , \8191 , \8192 );
nor \U$6321 ( \8194 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8193 );
buf \U$6322 ( \8195 , \8194 );
and \U$6323 ( \8196 , \8179 , \8195 );
nor \U$6324 ( \8197 , RI9921730_613, RI99217a8_612, RI9921820_611, RI9921898_610, \2158 , RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6325 ( \8198 , RI995e4c8_235, \8197 );
nor \U$6326 ( \8199 , \2161 , \2162 , \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6327 ( \8200 , RI99670f0_222, \8199 );
nor \U$6328 ( \8201 , RI9921730_613, \2162 , \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6329 ( \8202 , RI890f600_209, \8201 );
nor \U$6330 ( \8203 , \2161 , RI99217a8_612, \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6331 ( \8204 , RI89185e8_196, \8203 );
nor \U$6332 ( \8205 , RI9921730_613, RI99217a8_612, \2163 , \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6333 ( \8206 , RI8924e10_183, \8205 );
nor \U$6334 ( \8207 , \2161 , \2162 , RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6335 ( \8208 , RI8930828_170, \8207 );
nor \U$6336 ( \8209 , RI9921730_613, \2162 , RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6337 ( \8210 , RI8939810_157, \8209 );
nor \U$6338 ( \8211 , \2161 , RI99217a8_612, RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6339 ( \8212 , RI8946038_144, \8211 );
nor \U$6340 ( \8213 , RI9921730_613, RI99217a8_612, RI9921820_611, \2164 , RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6341 ( \8214 , RI89ec0a0_131, \8213 );
nor \U$6342 ( \8215 , \2161 , \2162 , \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6343 ( \8216 , RI89ec6b8_118, \8215 );
nor \U$6344 ( \8217 , RI9921730_613, \2162 , \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6345 ( \8218 , RI9776ff8_105, \8217 );
nor \U$6346 ( \8219 , \2161 , RI99217a8_612, \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6347 ( \8220 , RI98084f8_92, \8219 );
nor \U$6348 ( \8221 , RI9921730_613, RI99217a8_612, \2163 , RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6349 ( \8222 , RI9808b10_79, \8221 );
nor \U$6350 ( \8223 , \2161 , \2162 , RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6351 ( \8224 , RI98197a8_66, \8223 );
nor \U$6352 ( \8225 , RI9921730_613, \2162 , RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6353 ( \8226 , RI98abcb0_53, \8225 );
nor \U$6354 ( \8227 , \2161 , RI99217a8_612, RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6355 ( \8228 , RI98bc948_40, \8227 );
nor \U$6356 ( \8229 , RI9921730_613, RI99217a8_612, RI9921820_611, RI9921898_610, RI9921910_609, RI9921988_608, RI9921a00_607, RI9921a78_606, RI9921af0_605, RI9921b68_604, RI9921be0_603, RI9921c58_602, RI9921cd0_601);
and \U$6357 ( \8230 , RI994de48_27, \8229 );
or \U$6358 ( \8231 , \8198 , \8200 , \8202 , \8204 , \8206 , \8208 , \8210 , \8212 , \8214 , \8216 , \8218 , \8220 , \8222 , \8224 , \8226 , \8228 , \8230 );
buf \U$6359 ( \8232 , RI9921988_608);
buf \U$6360 ( \8233 , RI9921a00_607);
buf \U$6361 ( \8234 , RI9921a78_606);
buf \U$6362 ( \8235 , RI9921af0_605);
buf \U$6363 ( \8236 , RI9921b68_604);
buf \U$6364 ( \8237 , RI9921be0_603);
buf \U$6365 ( \8238 , RI9921c58_602);
buf \U$6366 ( \8239 , RI9921cd0_601);
buf \U$6367 ( \8240 , RI9921910_609);
buf \U$6368 ( \8241 , RI9921730_613);
buf \U$6369 ( \8242 , RI99217a8_612);
buf \U$6370 ( \8243 , RI9921820_611);
buf \U$6371 ( \8244 , RI9921898_610);
or \U$6372 ( \8245 , \8241 , \8242 , \8243 , \8244 );
and \U$6373 ( \8246 , \8240 , \8245 );
or \U$6374 ( \8247 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8246 );
buf \U$6375 ( \8248 , \8247 );
_DC g1220 ( \8249_nG1220 , \8231 , \8248 );
buf \U$6376 ( \8250 , \8249_nG1220 );
not \U$6377 ( \8251 , \8250 );
nor \U$6378 ( \8252 , \4955 , \4959 , \4963 , \4967 , \4972 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6379 ( \8253 , RI995e4c8_235, \8252 );
nor \U$6380 ( \8254 , \5007 , \5008 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6381 ( \8255 , RI99670f0_222, \8254 );
nor \U$6382 ( \8256 , \4955 , \5008 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6383 ( \8257 , RI890f600_209, \8256 );
nor \U$6384 ( \8258 , \5007 , \4959 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6385 ( \8259 , RI89185e8_196, \8258 );
nor \U$6386 ( \8260 , \4955 , \4959 , \5009 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6387 ( \8261 , RI8924e10_183, \8260 );
nor \U$6388 ( \8262 , \5007 , \5008 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6389 ( \8263 , RI8930828_170, \8262 );
nor \U$6390 ( \8264 , \4955 , \5008 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6391 ( \8265 , RI8939810_157, \8264 );
nor \U$6392 ( \8266 , \5007 , \4959 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6393 ( \8267 , RI8946038_144, \8266 );
nor \U$6394 ( \8268 , \4955 , \4959 , \4963 , \5010 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6395 ( \8269 , RI89ec0a0_131, \8268 );
nor \U$6396 ( \8270 , \5007 , \5008 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6397 ( \8271 , RI89ec6b8_118, \8270 );
nor \U$6398 ( \8272 , \4955 , \5008 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6399 ( \8273 , RI9776ff8_105, \8272 );
nor \U$6400 ( \8274 , \5007 , \4959 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6401 ( \8275 , RI98084f8_92, \8274 );
nor \U$6402 ( \8276 , \4955 , \4959 , \5009 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6403 ( \8277 , RI9808b10_79, \8276 );
nor \U$6404 ( \8278 , \5007 , \5008 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6405 ( \8279 , RI98197a8_66, \8278 );
nor \U$6406 ( \8280 , \4955 , \5008 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6407 ( \8281 , RI98abcb0_53, \8280 );
nor \U$6408 ( \8282 , \5007 , \4959 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6409 ( \8283 , RI98bc948_40, \8282 );
nor \U$6410 ( \8284 , \4955 , \4959 , \4963 , \4967 , \4971 , \4976 , \4980 , \4984 , \4988 , \4992 , \4996 , \5000 , \5004 );
and \U$6411 ( \8285 , RI994de48_27, \8284 );
or \U$6412 ( \8286 , \8253 , \8255 , \8257 , \8259 , \8261 , \8263 , \8265 , \8267 , \8269 , \8271 , \8273 , \8275 , \8277 , \8279 , \8281 , \8283 , \8285 );
buf \U$6413 ( \8287 , \4976 );
buf \U$6414 ( \8288 , \4980 );
buf \U$6415 ( \8289 , \4984 );
buf \U$6416 ( \8290 , \4988 );
buf \U$6417 ( \8291 , \4992 );
buf \U$6418 ( \8292 , \4996 );
buf \U$6419 ( \8293 , \5000 );
buf \U$6420 ( \8294 , \5004 );
buf \U$6421 ( \8295 , \4971 );
buf \U$6422 ( \8296 , \4955 );
buf \U$6423 ( \8297 , \4959 );
buf \U$6424 ( \8298 , \4963 );
buf \U$6425 ( \8299 , \4967 );
or \U$6426 ( \8300 , \8296 , \8297 , \8298 , \8299 );
and \U$6427 ( \8301 , \8295 , \8300 );
or \U$6428 ( \8302 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8301 );
buf \U$6429 ( \8303 , \8302 );
_DC g1257 ( \8304_nG1257 , \8286 , \8303 );
buf \U$6430 ( \8305 , \8304_nG1257 );
and \U$6431 ( \8306 , \8251 , \8305 );
and \U$6432 ( \8307 , RI995e450_236, \8197 );
and \U$6433 ( \8308 , RI9967078_223, \8199 );
and \U$6434 ( \8309 , RI9967690_210, \8201 );
and \U$6435 ( \8310 , RI890fba0_197, \8203 );
and \U$6436 ( \8311 , RI8918b88_184, \8205 );
and \U$6437 ( \8312 , RI89253b0_171, \8207 );
and \U$6438 ( \8313 , RI8930dc8_158, \8209 );
and \U$6439 ( \8314 , RI8939db0_145, \8211 );
and \U$6440 ( \8315 , RI89465d8_132, \8213 );
and \U$6441 ( \8316 , RI89ec640_119, \8215 );
and \U$6442 ( \8317 , RI9776f80_106, \8217 );
and \U$6443 ( \8318 , RI9808480_93, \8219 );
and \U$6444 ( \8319 , RI9808a98_80, \8221 );
and \U$6445 ( \8320 , RI9819730_67, \8223 );
and \U$6446 ( \8321 , RI98abc38_54, \8225 );
and \U$6447 ( \8322 , RI98bc8d0_41, \8227 );
and \U$6448 ( \8323 , RI994ddd0_28, \8229 );
or \U$6449 ( \8324 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 );
_DC g126c ( \8325_nG126c , \8324 , \8248 );
buf \U$6450 ( \8326 , \8325_nG126c );
not \U$6451 ( \8327 , \8326 );
and \U$6452 ( \8328 , RI995e450_236, \8252 );
and \U$6453 ( \8329 , RI9967078_223, \8254 );
and \U$6454 ( \8330 , RI9967690_210, \8256 );
and \U$6455 ( \8331 , RI890fba0_197, \8258 );
and \U$6456 ( \8332 , RI8918b88_184, \8260 );
and \U$6457 ( \8333 , RI89253b0_171, \8262 );
and \U$6458 ( \8334 , RI8930dc8_158, \8264 );
and \U$6459 ( \8335 , RI8939db0_145, \8266 );
and \U$6460 ( \8336 , RI89465d8_132, \8268 );
and \U$6461 ( \8337 , RI89ec640_119, \8270 );
and \U$6462 ( \8338 , RI9776f80_106, \8272 );
and \U$6463 ( \8339 , RI9808480_93, \8274 );
and \U$6464 ( \8340 , RI9808a98_80, \8276 );
and \U$6465 ( \8341 , RI9819730_67, \8278 );
and \U$6466 ( \8342 , RI98abc38_54, \8280 );
and \U$6467 ( \8343 , RI98bc8d0_41, \8282 );
and \U$6468 ( \8344 , RI994ddd0_28, \8284 );
or \U$6469 ( \8345 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 );
_DC g1281 ( \8346_nG1281 , \8345 , \8303 );
buf \U$6470 ( \8347 , \8346_nG1281 );
and \U$6471 ( \8348 , \8327 , \8347 );
and \U$6472 ( \8349 , RI995e3d8_237, \8197 );
and \U$6473 ( \8350 , RI99669e8_224, \8199 );
and \U$6474 ( \8351 , RI9967618_211, \8201 );
and \U$6475 ( \8352 , RI890fb28_198, \8203 );
and \U$6476 ( \8353 , RI8918b10_185, \8205 );
and \U$6477 ( \8354 , RI8925338_172, \8207 );
and \U$6478 ( \8355 , RI8930d50_159, \8209 );
and \U$6479 ( \8356 , RI8939d38_146, \8211 );
and \U$6480 ( \8357 , RI8946560_133, \8213 );
and \U$6481 ( \8358 , RI89ec5c8_120, \8215 );
and \U$6482 ( \8359 , RI9776f08_107, \8217 );
and \U$6483 ( \8360 , RI9808408_94, \8219 );
and \U$6484 ( \8361 , RI9808a20_81, \8221 );
and \U$6485 ( \8362 , RI98196b8_68, \8223 );
and \U$6486 ( \8363 , RI98abbc0_55, \8225 );
and \U$6487 ( \8364 , RI98bc858_42, \8227 );
and \U$6488 ( \8365 , RI994dd58_29, \8229 );
or \U$6489 ( \8366 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 );
_DC g1296 ( \8367_nG1296 , \8366 , \8248 );
buf \U$6490 ( \8368 , \8367_nG1296 );
not \U$6491 ( \8369 , \8368 );
and \U$6492 ( \8370 , RI995e3d8_237, \8252 );
and \U$6493 ( \8371 , RI99669e8_224, \8254 );
and \U$6494 ( \8372 , RI9967618_211, \8256 );
and \U$6495 ( \8373 , RI890fb28_198, \8258 );
and \U$6496 ( \8374 , RI8918b10_185, \8260 );
and \U$6497 ( \8375 , RI8925338_172, \8262 );
and \U$6498 ( \8376 , RI8930d50_159, \8264 );
and \U$6499 ( \8377 , RI8939d38_146, \8266 );
and \U$6500 ( \8378 , RI8946560_133, \8268 );
and \U$6501 ( \8379 , RI89ec5c8_120, \8270 );
and \U$6502 ( \8380 , RI9776f08_107, \8272 );
and \U$6503 ( \8381 , RI9808408_94, \8274 );
and \U$6504 ( \8382 , RI9808a20_81, \8276 );
and \U$6505 ( \8383 , RI98196b8_68, \8278 );
and \U$6506 ( \8384 , RI98abbc0_55, \8280 );
and \U$6507 ( \8385 , RI98bc858_42, \8282 );
and \U$6508 ( \8386 , RI994dd58_29, \8284 );
or \U$6509 ( \8387 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 );
_DC g12ab ( \8388_nG12ab , \8387 , \8303 );
buf \U$6510 ( \8389 , \8388_nG12ab );
and \U$6511 ( \8390 , \8369 , \8389 );
and \U$6512 ( \8391 , RI9959fe0_238, \8197 );
and \U$6513 ( \8392 , RI995e978_225, \8199 );
and \U$6514 ( \8393 , RI99675a0_212, \8201 );
and \U$6515 ( \8394 , RI890fab0_199, \8203 );
and \U$6516 ( \8395 , RI8918a98_186, \8205 );
and \U$6517 ( \8396 , RI89252c0_173, \8207 );
and \U$6518 ( \8397 , RI8930cd8_160, \8209 );
and \U$6519 ( \8398 , RI8939cc0_147, \8211 );
and \U$6520 ( \8399 , RI89464e8_134, \8213 );
and \U$6521 ( \8400 , RI89ec550_121, \8215 );
and \U$6522 ( \8401 , RI9776e90_108, \8217 );
and \U$6523 ( \8402 , RI9808390_95, \8219 );
and \U$6524 ( \8403 , RI98089a8_82, \8221 );
and \U$6525 ( \8404 , RI9819640_69, \8223 );
and \U$6526 ( \8405 , RI98abb48_56, \8225 );
and \U$6527 ( \8406 , RI98bc7e0_43, \8227 );
and \U$6528 ( \8407 , RI994dce0_30, \8229 );
or \U$6529 ( \8408 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 );
_DC g12c0 ( \8409_nG12c0 , \8408 , \8248 );
buf \U$6530 ( \8410 , \8409_nG12c0 );
not \U$6531 ( \8411 , \8410 );
and \U$6532 ( \8412 , RI9959fe0_238, \8252 );
and \U$6533 ( \8413 , RI995e978_225, \8254 );
and \U$6534 ( \8414 , RI99675a0_212, \8256 );
and \U$6535 ( \8415 , RI890fab0_199, \8258 );
and \U$6536 ( \8416 , RI8918a98_186, \8260 );
and \U$6537 ( \8417 , RI89252c0_173, \8262 );
and \U$6538 ( \8418 , RI8930cd8_160, \8264 );
and \U$6539 ( \8419 , RI8939cc0_147, \8266 );
and \U$6540 ( \8420 , RI89464e8_134, \8268 );
and \U$6541 ( \8421 , RI89ec550_121, \8270 );
and \U$6542 ( \8422 , RI9776e90_108, \8272 );
and \U$6543 ( \8423 , RI9808390_95, \8274 );
and \U$6544 ( \8424 , RI98089a8_82, \8276 );
and \U$6545 ( \8425 , RI9819640_69, \8278 );
and \U$6546 ( \8426 , RI98abb48_56, \8280 );
and \U$6547 ( \8427 , RI98bc7e0_43, \8282 );
and \U$6548 ( \8428 , RI994dce0_30, \8284 );
or \U$6549 ( \8429 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 );
_DC g12d5 ( \8430_nG12d5 , \8429 , \8303 );
buf \U$6550 ( \8431 , \8430_nG12d5 );
and \U$6551 ( \8432 , \8411 , \8431 );
and \U$6552 ( \8433 , RI9959f68_239, \8197 );
and \U$6553 ( \8434 , RI995e900_226, \8199 );
and \U$6554 ( \8435 , RI9967528_213, \8201 );
and \U$6555 ( \8436 , RI890fa38_200, \8203 );
and \U$6556 ( \8437 , RI8918a20_187, \8205 );
and \U$6557 ( \8438 , RI8925248_174, \8207 );
and \U$6558 ( \8439 , RI8930c60_161, \8209 );
and \U$6559 ( \8440 , RI8939c48_148, \8211 );
and \U$6560 ( \8441 , RI8946470_135, \8213 );
and \U$6561 ( \8442 , RI89ec4d8_122, \8215 );
and \U$6562 ( \8443 , RI9776e18_109, \8217 );
and \U$6563 ( \8444 , RI9808318_96, \8219 );
and \U$6564 ( \8445 , RI9808930_83, \8221 );
and \U$6565 ( \8446 , RI98195c8_70, \8223 );
and \U$6566 ( \8447 , RI98abad0_57, \8225 );
and \U$6567 ( \8448 , RI98bc768_44, \8227 );
and \U$6568 ( \8449 , RI994dc68_31, \8229 );
or \U$6569 ( \8450 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 );
_DC g12ea ( \8451_nG12ea , \8450 , \8248 );
buf \U$6570 ( \8452 , \8451_nG12ea );
not \U$6571 ( \8453 , \8452 );
and \U$6572 ( \8454 , RI9959f68_239, \8252 );
and \U$6573 ( \8455 , RI995e900_226, \8254 );
and \U$6574 ( \8456 , RI9967528_213, \8256 );
and \U$6575 ( \8457 , RI890fa38_200, \8258 );
and \U$6576 ( \8458 , RI8918a20_187, \8260 );
and \U$6577 ( \8459 , RI8925248_174, \8262 );
and \U$6578 ( \8460 , RI8930c60_161, \8264 );
and \U$6579 ( \8461 , RI8939c48_148, \8266 );
and \U$6580 ( \8462 , RI8946470_135, \8268 );
and \U$6581 ( \8463 , RI89ec4d8_122, \8270 );
and \U$6582 ( \8464 , RI9776e18_109, \8272 );
and \U$6583 ( \8465 , RI9808318_96, \8274 );
and \U$6584 ( \8466 , RI9808930_83, \8276 );
and \U$6585 ( \8467 , RI98195c8_70, \8278 );
and \U$6586 ( \8468 , RI98abad0_57, \8280 );
and \U$6587 ( \8469 , RI98bc768_44, \8282 );
and \U$6588 ( \8470 , RI994dc68_31, \8284 );
or \U$6589 ( \8471 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 );
_DC g12ff ( \8472_nG12ff , \8471 , \8303 );
buf \U$6590 ( \8473 , \8472_nG12ff );
and \U$6591 ( \8474 , \8453 , \8473 );
and \U$6592 ( \8475 , RI9959860_240, \8197 );
and \U$6593 ( \8476 , RI995e888_227, \8199 );
and \U$6594 ( \8477 , RI99674b0_214, \8201 );
and \U$6595 ( \8478 , RI890f9c0_201, \8203 );
and \U$6596 ( \8479 , RI89189a8_188, \8205 );
and \U$6597 ( \8480 , RI89251d0_175, \8207 );
and \U$6598 ( \8481 , RI8930be8_162, \8209 );
and \U$6599 ( \8482 , RI8939bd0_149, \8211 );
and \U$6600 ( \8483 , RI89463f8_136, \8213 );
and \U$6601 ( \8484 , RI89ec460_123, \8215 );
and \U$6602 ( \8485 , RI9776da0_110, \8217 );
and \U$6603 ( \8486 , RI98082a0_97, \8219 );
and \U$6604 ( \8487 , RI98088b8_84, \8221 );
and \U$6605 ( \8488 , RI9819550_71, \8223 );
and \U$6606 ( \8489 , RI98aba58_58, \8225 );
and \U$6607 ( \8490 , RI98bc6f0_45, \8227 );
and \U$6608 ( \8491 , RI994dbf0_32, \8229 );
or \U$6609 ( \8492 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 );
_DC g1314 ( \8493_nG1314 , \8492 , \8248 );
buf \U$6610 ( \8494 , \8493_nG1314 );
not \U$6611 ( \8495 , \8494 );
and \U$6612 ( \8496 , RI9959860_240, \8252 );
and \U$6613 ( \8497 , RI995e888_227, \8254 );
and \U$6614 ( \8498 , RI99674b0_214, \8256 );
and \U$6615 ( \8499 , RI890f9c0_201, \8258 );
and \U$6616 ( \8500 , RI89189a8_188, \8260 );
and \U$6617 ( \8501 , RI89251d0_175, \8262 );
and \U$6618 ( \8502 , RI8930be8_162, \8264 );
and \U$6619 ( \8503 , RI8939bd0_149, \8266 );
and \U$6620 ( \8504 , RI89463f8_136, \8268 );
and \U$6621 ( \8505 , RI89ec460_123, \8270 );
and \U$6622 ( \8506 , RI9776da0_110, \8272 );
and \U$6623 ( \8507 , RI98082a0_97, \8274 );
and \U$6624 ( \8508 , RI98088b8_84, \8276 );
and \U$6625 ( \8509 , RI9819550_71, \8278 );
and \U$6626 ( \8510 , RI98aba58_58, \8280 );
and \U$6627 ( \8511 , RI98bc6f0_45, \8282 );
and \U$6628 ( \8512 , RI994dbf0_32, \8284 );
or \U$6629 ( \8513 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 );
_DC g1329 ( \8514_nG1329 , \8513 , \8303 );
buf \U$6630 ( \8515 , \8514_nG1329 );
and \U$6631 ( \8516 , \8495 , \8515 );
and \U$6632 ( \8517 , RI994d998_241, \8197 );
and \U$6633 ( \8518 , RI995e810_228, \8199 );
and \U$6634 ( \8519 , RI9967438_215, \8201 );
and \U$6635 ( \8520 , RI890f948_202, \8203 );
and \U$6636 ( \8521 , RI8918930_189, \8205 );
and \U$6637 ( \8522 , RI8925158_176, \8207 );
and \U$6638 ( \8523 , RI8930b70_163, \8209 );
and \U$6639 ( \8524 , RI8939b58_150, \8211 );
and \U$6640 ( \8525 , RI8946380_137, \8213 );
and \U$6641 ( \8526 , RI89ec3e8_124, \8215 );
and \U$6642 ( \8527 , RI9776d28_111, \8217 );
and \U$6643 ( \8528 , RI9808228_98, \8219 );
and \U$6644 ( \8529 , RI9808840_85, \8221 );
and \U$6645 ( \8530 , RI98194d8_72, \8223 );
and \U$6646 ( \8531 , RI98ab9e0_59, \8225 );
and \U$6647 ( \8532 , RI98abff8_46, \8227 );
and \U$6648 ( \8533 , RI98bcc90_33, \8229 );
or \U$6649 ( \8534 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 );
_DC g133e ( \8535_nG133e , \8534 , \8248 );
buf \U$6650 ( \8536 , \8535_nG133e );
not \U$6651 ( \8537 , \8536 );
and \U$6652 ( \8538 , RI994d998_241, \8252 );
and \U$6653 ( \8539 , RI995e810_228, \8254 );
and \U$6654 ( \8540 , RI9967438_215, \8256 );
and \U$6655 ( \8541 , RI890f948_202, \8258 );
and \U$6656 ( \8542 , RI8918930_189, \8260 );
and \U$6657 ( \8543 , RI8925158_176, \8262 );
and \U$6658 ( \8544 , RI8930b70_163, \8264 );
and \U$6659 ( \8545 , RI8939b58_150, \8266 );
and \U$6660 ( \8546 , RI8946380_137, \8268 );
and \U$6661 ( \8547 , RI89ec3e8_124, \8270 );
and \U$6662 ( \8548 , RI9776d28_111, \8272 );
and \U$6663 ( \8549 , RI9808228_98, \8274 );
and \U$6664 ( \8550 , RI9808840_85, \8276 );
and \U$6665 ( \8551 , RI98194d8_72, \8278 );
and \U$6666 ( \8552 , RI98ab9e0_59, \8280 );
and \U$6667 ( \8553 , RI98abff8_46, \8282 );
and \U$6668 ( \8554 , RI98bcc90_33, \8284 );
or \U$6669 ( \8555 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 );
_DC g1353 ( \8556_nG1353 , \8555 , \8303 );
buf \U$6670 ( \8557 , \8556_nG1353 );
and \U$6671 ( \8558 , \8537 , \8557 );
and \U$6672 ( \8559 , RI994d920_242, \8197 );
and \U$6673 ( \8560 , RI995e798_229, \8199 );
and \U$6674 ( \8561 , RI99673c0_216, \8201 );
and \U$6675 ( \8562 , RI890f8d0_203, \8203 );
and \U$6676 ( \8563 , RI89188b8_190, \8205 );
and \U$6677 ( \8564 , RI89250e0_177, \8207 );
and \U$6678 ( \8565 , RI8930af8_164, \8209 );
and \U$6679 ( \8566 , RI8939ae0_151, \8211 );
and \U$6680 ( \8567 , RI8946308_138, \8213 );
and \U$6681 ( \8568 , RI89ec370_125, \8215 );
and \U$6682 ( \8569 , RI89ec988_112, \8217 );
and \U$6683 ( \8570 , RI97772c8_99, \8219 );
and \U$6684 ( \8571 , RI98087c8_86, \8221 );
and \U$6685 ( \8572 , RI9819460_73, \8223 );
and \U$6686 ( \8573 , RI98ab968_60, \8225 );
and \U$6687 ( \8574 , RI98abf80_47, \8227 );
and \U$6688 ( \8575 , RI98bcc18_34, \8229 );
or \U$6689 ( \8576 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 );
_DC g1368 ( \8577_nG1368 , \8576 , \8248 );
buf \U$6690 ( \8578 , \8577_nG1368 );
not \U$6691 ( \8579 , \8578 );
and \U$6692 ( \8580 , RI994d920_242, \8252 );
and \U$6693 ( \8581 , RI995e798_229, \8254 );
and \U$6694 ( \8582 , RI99673c0_216, \8256 );
and \U$6695 ( \8583 , RI890f8d0_203, \8258 );
and \U$6696 ( \8584 , RI89188b8_190, \8260 );
and \U$6697 ( \8585 , RI89250e0_177, \8262 );
and \U$6698 ( \8586 , RI8930af8_164, \8264 );
and \U$6699 ( \8587 , RI8939ae0_151, \8266 );
and \U$6700 ( \8588 , RI8946308_138, \8268 );
and \U$6701 ( \8589 , RI89ec370_125, \8270 );
and \U$6702 ( \8590 , RI89ec988_112, \8272 );
and \U$6703 ( \8591 , RI97772c8_99, \8274 );
and \U$6704 ( \8592 , RI98087c8_86, \8276 );
and \U$6705 ( \8593 , RI9819460_73, \8278 );
and \U$6706 ( \8594 , RI98ab968_60, \8280 );
and \U$6707 ( \8595 , RI98abf80_47, \8282 );
and \U$6708 ( \8596 , RI98bcc18_34, \8284 );
or \U$6709 ( \8597 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 );
_DC g137d ( \8598_nG137d , \8597 , \8303 );
buf \U$6710 ( \8599 , \8598_nG137d );
and \U$6711 ( \8600 , \8579 , \8599 );
and \U$6712 ( \8601 , RI994d8a8_243, \8197 );
and \U$6713 ( \8602 , RI995e720_230, \8199 );
and \U$6714 ( \8603 , RI9967348_217, \8201 );
and \U$6715 ( \8604 , RI890f858_204, \8203 );
and \U$6716 ( \8605 , RI8918840_191, \8205 );
and \U$6717 ( \8606 , RI8925068_178, \8207 );
and \U$6718 ( \8607 , RI8930a80_165, \8209 );
and \U$6719 ( \8608 , RI8939a68_152, \8211 );
and \U$6720 ( \8609 , RI8946290_139, \8213 );
and \U$6721 ( \8610 , RI89ec2f8_126, \8215 );
and \U$6722 ( \8611 , RI89ec910_113, \8217 );
and \U$6723 ( \8612 , RI9777250_100, \8219 );
and \U$6724 ( \8613 , RI9808750_87, \8221 );
and \U$6725 ( \8614 , RI98193e8_74, \8223 );
and \U$6726 ( \8615 , RI98ab8f0_61, \8225 );
and \U$6727 ( \8616 , RI98abf08_48, \8227 );
and \U$6728 ( \8617 , RI98bcba0_35, \8229 );
or \U$6729 ( \8618 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 );
_DC g1392 ( \8619_nG1392 , \8618 , \8248 );
buf \U$6730 ( \8620 , \8619_nG1392 );
not \U$6731 ( \8621 , \8620 );
and \U$6732 ( \8622 , RI994d8a8_243, \8252 );
and \U$6733 ( \8623 , RI995e720_230, \8254 );
and \U$6734 ( \8624 , RI9967348_217, \8256 );
and \U$6735 ( \8625 , RI890f858_204, \8258 );
and \U$6736 ( \8626 , RI8918840_191, \8260 );
and \U$6737 ( \8627 , RI8925068_178, \8262 );
and \U$6738 ( \8628 , RI8930a80_165, \8264 );
and \U$6739 ( \8629 , RI8939a68_152, \8266 );
and \U$6740 ( \8630 , RI8946290_139, \8268 );
and \U$6741 ( \8631 , RI89ec2f8_126, \8270 );
and \U$6742 ( \8632 , RI89ec910_113, \8272 );
and \U$6743 ( \8633 , RI9777250_100, \8274 );
and \U$6744 ( \8634 , RI9808750_87, \8276 );
and \U$6745 ( \8635 , RI98193e8_74, \8278 );
and \U$6746 ( \8636 , RI98ab8f0_61, \8280 );
and \U$6747 ( \8637 , RI98abf08_48, \8282 );
and \U$6748 ( \8638 , RI98bcba0_35, \8284 );
or \U$6749 ( \8639 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 );
_DC g13a7 ( \8640_nG13a7 , \8639 , \8303 );
buf \U$6750 ( \8641 , \8640_nG13a7 );
and \U$6751 ( \8642 , \8621 , \8641 );
and \U$6752 ( \8643 , RI994d830_244, \8197 );
and \U$6753 ( \8644 , RI995e6a8_231, \8199 );
and \U$6754 ( \8645 , RI99672d0_218, \8201 );
and \U$6755 ( \8646 , RI890f7e0_205, \8203 );
and \U$6756 ( \8647 , RI89187c8_192, \8205 );
and \U$6757 ( \8648 , RI8924ff0_179, \8207 );
and \U$6758 ( \8649 , RI8930a08_166, \8209 );
and \U$6759 ( \8650 , RI89399f0_153, \8211 );
and \U$6760 ( \8651 , RI8946218_140, \8213 );
and \U$6761 ( \8652 , RI89ec280_127, \8215 );
and \U$6762 ( \8653 , RI89ec898_114, \8217 );
and \U$6763 ( \8654 , RI97771d8_101, \8219 );
and \U$6764 ( \8655 , RI98086d8_88, \8221 );
and \U$6765 ( \8656 , RI9819370_75, \8223 );
and \U$6766 ( \8657 , RI98ab878_62, \8225 );
and \U$6767 ( \8658 , RI98abe90_49, \8227 );
and \U$6768 ( \8659 , RI98bcb28_36, \8229 );
or \U$6769 ( \8660 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 );
_DC g13bc ( \8661_nG13bc , \8660 , \8248 );
buf \U$6770 ( \8662 , \8661_nG13bc );
not \U$6771 ( \8663 , \8662 );
and \U$6772 ( \8664 , RI994d830_244, \8252 );
and \U$6773 ( \8665 , RI995e6a8_231, \8254 );
and \U$6774 ( \8666 , RI99672d0_218, \8256 );
and \U$6775 ( \8667 , RI890f7e0_205, \8258 );
and \U$6776 ( \8668 , RI89187c8_192, \8260 );
and \U$6777 ( \8669 , RI8924ff0_179, \8262 );
and \U$6778 ( \8670 , RI8930a08_166, \8264 );
and \U$6779 ( \8671 , RI89399f0_153, \8266 );
and \U$6780 ( \8672 , RI8946218_140, \8268 );
and \U$6781 ( \8673 , RI89ec280_127, \8270 );
and \U$6782 ( \8674 , RI89ec898_114, \8272 );
and \U$6783 ( \8675 , RI97771d8_101, \8274 );
and \U$6784 ( \8676 , RI98086d8_88, \8276 );
and \U$6785 ( \8677 , RI9819370_75, \8278 );
and \U$6786 ( \8678 , RI98ab878_62, \8280 );
and \U$6787 ( \8679 , RI98abe90_49, \8282 );
and \U$6788 ( \8680 , RI98bcb28_36, \8284 );
or \U$6789 ( \8681 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 );
_DC g13d1 ( \8682_nG13d1 , \8681 , \8303 );
buf \U$6790 ( \8683 , \8682_nG13d1 );
and \U$6791 ( \8684 , \8663 , \8683 );
and \U$6792 ( \8685 , RI994d7b8_245, \8197 );
and \U$6793 ( \8686 , RI995e630_232, \8199 );
and \U$6794 ( \8687 , RI9967258_219, \8201 );
and \U$6795 ( \8688 , RI890f768_206, \8203 );
and \U$6796 ( \8689 , RI8918750_193, \8205 );
and \U$6797 ( \8690 , RI8924f78_180, \8207 );
and \U$6798 ( \8691 , RI8930990_167, \8209 );
and \U$6799 ( \8692 , RI8939978_154, \8211 );
and \U$6800 ( \8693 , RI89461a0_141, \8213 );
and \U$6801 ( \8694 , RI89ec208_128, \8215 );
and \U$6802 ( \8695 , RI89ec820_115, \8217 );
and \U$6803 ( \8696 , RI9777160_102, \8219 );
and \U$6804 ( \8697 , RI9808660_89, \8221 );
and \U$6805 ( \8698 , RI98192f8_76, \8223 );
and \U$6806 ( \8699 , RI98ab800_63, \8225 );
and \U$6807 ( \8700 , RI98abe18_50, \8227 );
and \U$6808 ( \8701 , RI98bcab0_37, \8229 );
or \U$6809 ( \8702 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 );
_DC g13e6 ( \8703_nG13e6 , \8702 , \8248 );
buf \U$6810 ( \8704 , \8703_nG13e6 );
not \U$6811 ( \8705 , \8704 );
and \U$6812 ( \8706 , RI994d7b8_245, \8252 );
and \U$6813 ( \8707 , RI995e630_232, \8254 );
and \U$6814 ( \8708 , RI9967258_219, \8256 );
and \U$6815 ( \8709 , RI890f768_206, \8258 );
and \U$6816 ( \8710 , RI8918750_193, \8260 );
and \U$6817 ( \8711 , RI8924f78_180, \8262 );
and \U$6818 ( \8712 , RI8930990_167, \8264 );
and \U$6819 ( \8713 , RI8939978_154, \8266 );
and \U$6820 ( \8714 , RI89461a0_141, \8268 );
and \U$6821 ( \8715 , RI89ec208_128, \8270 );
and \U$6822 ( \8716 , RI89ec820_115, \8272 );
and \U$6823 ( \8717 , RI9777160_102, \8274 );
and \U$6824 ( \8718 , RI9808660_89, \8276 );
and \U$6825 ( \8719 , RI98192f8_76, \8278 );
and \U$6826 ( \8720 , RI98ab800_63, \8280 );
and \U$6827 ( \8721 , RI98abe18_50, \8282 );
and \U$6828 ( \8722 , RI98bcab0_37, \8284 );
or \U$6829 ( \8723 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 );
_DC g13fb ( \8724_nG13fb , \8723 , \8303 );
buf \U$6830 ( \8725 , \8724_nG13fb );
and \U$6831 ( \8726 , \8705 , \8725 );
and \U$6832 ( \8727 , RI994d740_246, \8197 );
and \U$6833 ( \8728 , RI995e5b8_233, \8199 );
and \U$6834 ( \8729 , RI99671e0_220, \8201 );
and \U$6835 ( \8730 , RI890f6f0_207, \8203 );
and \U$6836 ( \8731 , RI89186d8_194, \8205 );
and \U$6837 ( \8732 , RI8924f00_181, \8207 );
and \U$6838 ( \8733 , RI8930918_168, \8209 );
and \U$6839 ( \8734 , RI8939900_155, \8211 );
and \U$6840 ( \8735 , RI8946128_142, \8213 );
and \U$6841 ( \8736 , RI89ec190_129, \8215 );
and \U$6842 ( \8737 , RI89ec7a8_116, \8217 );
and \U$6843 ( \8738 , RI97770e8_103, \8219 );
and \U$6844 ( \8739 , RI98085e8_90, \8221 );
and \U$6845 ( \8740 , RI9819280_77, \8223 );
and \U$6846 ( \8741 , RI98ab788_64, \8225 );
and \U$6847 ( \8742 , RI98abda0_51, \8227 );
and \U$6848 ( \8743 , RI98bca38_38, \8229 );
or \U$6849 ( \8744 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 );
_DC g1410 ( \8745_nG1410 , \8744 , \8248 );
buf \U$6850 ( \8746 , \8745_nG1410 );
not \U$6851 ( \8747 , \8746 );
and \U$6852 ( \8748 , RI994d740_246, \8252 );
and \U$6853 ( \8749 , RI995e5b8_233, \8254 );
and \U$6854 ( \8750 , RI99671e0_220, \8256 );
and \U$6855 ( \8751 , RI890f6f0_207, \8258 );
and \U$6856 ( \8752 , RI89186d8_194, \8260 );
and \U$6857 ( \8753 , RI8924f00_181, \8262 );
and \U$6858 ( \8754 , RI8930918_168, \8264 );
and \U$6859 ( \8755 , RI8939900_155, \8266 );
and \U$6860 ( \8756 , RI8946128_142, \8268 );
and \U$6861 ( \8757 , RI89ec190_129, \8270 );
and \U$6862 ( \8758 , RI89ec7a8_116, \8272 );
and \U$6863 ( \8759 , RI97770e8_103, \8274 );
and \U$6864 ( \8760 , RI98085e8_90, \8276 );
and \U$6865 ( \8761 , RI9819280_77, \8278 );
and \U$6866 ( \8762 , RI98ab788_64, \8280 );
and \U$6867 ( \8763 , RI98abda0_51, \8282 );
and \U$6868 ( \8764 , RI98bca38_38, \8284 );
or \U$6869 ( \8765 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 );
_DC g1425 ( \8766_nG1425 , \8765 , \8303 );
buf \U$6870 ( \8767 , \8766_nG1425 );
and \U$6871 ( \8768 , \8747 , \8767 );
and \U$6872 ( \8769 , RI994d6c8_247, \8197 );
and \U$6873 ( \8770 , RI995e540_234, \8199 );
and \U$6874 ( \8771 , RI9967168_221, \8201 );
and \U$6875 ( \8772 , RI890f678_208, \8203 );
and \U$6876 ( \8773 , RI8918660_195, \8205 );
and \U$6877 ( \8774 , RI8924e88_182, \8207 );
and \U$6878 ( \8775 , RI89308a0_169, \8209 );
and \U$6879 ( \8776 , RI8939888_156, \8211 );
and \U$6880 ( \8777 , RI89460b0_143, \8213 );
and \U$6881 ( \8778 , RI89ec118_130, \8215 );
and \U$6882 ( \8779 , RI89ec730_117, \8217 );
and \U$6883 ( \8780 , RI9777070_104, \8219 );
and \U$6884 ( \8781 , RI9808570_91, \8221 );
and \U$6885 ( \8782 , RI9819208_78, \8223 );
and \U$6886 ( \8783 , RI98ab710_65, \8225 );
and \U$6887 ( \8784 , RI98abd28_52, \8227 );
and \U$6888 ( \8785 , RI98bc9c0_39, \8229 );
or \U$6889 ( \8786 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 );
_DC g143a ( \8787_nG143a , \8786 , \8248 );
buf \U$6890 ( \8788 , \8787_nG143a );
not \U$6891 ( \8789 , \8788 );
and \U$6892 ( \8790 , RI994d6c8_247, \8252 );
and \U$6893 ( \8791 , RI995e540_234, \8254 );
and \U$6894 ( \8792 , RI9967168_221, \8256 );
and \U$6895 ( \8793 , RI890f678_208, \8258 );
and \U$6896 ( \8794 , RI8918660_195, \8260 );
and \U$6897 ( \8795 , RI8924e88_182, \8262 );
and \U$6898 ( \8796 , RI89308a0_169, \8264 );
and \U$6899 ( \8797 , RI8939888_156, \8266 );
and \U$6900 ( \8798 , RI89460b0_143, \8268 );
and \U$6901 ( \8799 , RI89ec118_130, \8270 );
and \U$6902 ( \8800 , RI89ec730_117, \8272 );
and \U$6903 ( \8801 , RI9777070_104, \8274 );
and \U$6904 ( \8802 , RI9808570_91, \8276 );
and \U$6905 ( \8803 , RI9819208_78, \8278 );
and \U$6906 ( \8804 , RI98ab710_65, \8280 );
and \U$6907 ( \8805 , RI98abd28_52, \8282 );
and \U$6908 ( \8806 , RI98bc9c0_39, \8284 );
or \U$6909 ( \8807 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 );
_DC g144f ( \8808_nG144f , \8807 , \8303 );
buf \U$6910 ( \8809 , \8808_nG144f );
and \U$6911 ( \8810 , \8789 , \8809 );
xnor \U$6912 ( \8811 , \8767 , \8746 );
and \U$6913 ( \8812 , \8810 , \8811 );
or \U$6914 ( \8813 , \8768 , \8812 );
xnor \U$6915 ( \8814 , \8725 , \8704 );
and \U$6916 ( \8815 , \8813 , \8814 );
or \U$6917 ( \8816 , \8726 , \8815 );
xnor \U$6918 ( \8817 , \8683 , \8662 );
and \U$6919 ( \8818 , \8816 , \8817 );
or \U$6920 ( \8819 , \8684 , \8818 );
xnor \U$6921 ( \8820 , \8641 , \8620 );
and \U$6922 ( \8821 , \8819 , \8820 );
or \U$6923 ( \8822 , \8642 , \8821 );
xnor \U$6924 ( \8823 , \8599 , \8578 );
and \U$6925 ( \8824 , \8822 , \8823 );
or \U$6926 ( \8825 , \8600 , \8824 );
xnor \U$6927 ( \8826 , \8557 , \8536 );
and \U$6928 ( \8827 , \8825 , \8826 );
or \U$6929 ( \8828 , \8558 , \8827 );
xnor \U$6930 ( \8829 , \8515 , \8494 );
and \U$6931 ( \8830 , \8828 , \8829 );
or \U$6932 ( \8831 , \8516 , \8830 );
xnor \U$6933 ( \8832 , \8473 , \8452 );
and \U$6934 ( \8833 , \8831 , \8832 );
or \U$6935 ( \8834 , \8474 , \8833 );
xnor \U$6936 ( \8835 , \8431 , \8410 );
and \U$6937 ( \8836 , \8834 , \8835 );
or \U$6938 ( \8837 , \8432 , \8836 );
xnor \U$6939 ( \8838 , \8389 , \8368 );
and \U$6940 ( \8839 , \8837 , \8838 );
or \U$6941 ( \8840 , \8390 , \8839 );
xnor \U$6942 ( \8841 , \8347 , \8326 );
and \U$6943 ( \8842 , \8840 , \8841 );
or \U$6944 ( \8843 , \8348 , \8842 );
xnor \U$6945 ( \8844 , \8305 , \8250 );
and \U$6946 ( \8845 , \8843 , \8844 );
or \U$6947 ( \8846 , \8306 , \8845 );
buf \U$6948 ( \8847 , \8846 );
and \U$6949 ( \8848 , \8196 , \8847 );
_HMUX g32b3_GF_PartitionCandidate ( \8849_nG32b3 , \4912_nG3284 , \7758_nG32b2 , \8848 );
buf \U$6950 ( \8850 , \8849_nG32b3 );
not \U$6951 ( \8851 , \4375 );
nand \U$6952 ( \8852 , \4904 , \8851 );
nor \U$6953 ( \8853 , \4722 , \3558 );
nor \U$6954 ( \8854 , \3633 , \3710 );
nand \U$6955 ( \8855 , \8853 , \8854 );
nor \U$6956 ( \8856 , \3785 , \3862 );
nor \U$6957 ( \8857 , \3938 , \4011 );
nand \U$6958 ( \8858 , \8856 , \8857 );
nor \U$6959 ( \8859 , \8855 , \8858 );
nor \U$6960 ( \8860 , \4080 , \4144 );
nor \U$6961 ( \8861 , \4204 , \4261 );
nand \U$6962 ( \8862 , \8860 , \8861 );
nor \U$6963 ( \8863 , \4299 , \4331 );
nor \U$6964 ( \8864 , \4352 , \4368 );
nand \U$6965 ( \8865 , \8863 , \8864 );
nor \U$6966 ( \8866 , \8862 , \8865 );
nand \U$6967 ( \8867 , \8859 , \8866 );
nor \U$6968 ( \8868 , \4783 , \4487 );
nor \U$6969 ( \8869 , \4532 , \4584 );
nand \U$6970 ( \8870 , \8868 , \8869 );
nor \U$6971 ( \8871 , \4639 , \4678 );
nor \U$6972 ( \8872 , \4699 , \4715 );
nand \U$6973 ( \8873 , \8871 , \8872 );
nor \U$6974 ( \8874 , \8870 , \8873 );
nor \U$6975 ( \8875 , \4803 , \4758 );
nor \U$6976 ( \8876 , \4769 , \4780 );
nand \U$6977 ( \8877 , \8875 , \8876 );
nor \U$6978 ( \8878 , \4808 , \4800 );
not \U$6979 ( \8879 , \4816 );
and \U$6980 ( \8880 , \8878 , \8879 );
or \U$6981 ( \8881 , \4800 , \4818 );
nand \U$6982 ( \8882 , \8881 , \4821 );
nor \U$6983 ( \8883 , \8880 , \8882 );
or \U$6984 ( \8884 , \8877 , \8883 );
or \U$6985 ( \8885 , \4758 , \4823 );
nand \U$6986 ( \8886 , \8885 , \4827 );
and \U$6987 ( \8887 , \8876 , \8886 );
or \U$6988 ( \8888 , \4780 , \4829 );
nand \U$6989 ( \8889 , \8888 , \4832 );
nor \U$6990 ( \8890 , \8887 , \8889 );
nand \U$6991 ( \8891 , \8884 , \8890 );
and \U$6992 ( \8892 , \8874 , \8891 );
or \U$6993 ( \8893 , \4487 , \4834 );
nand \U$6994 ( \8894 , \8893 , \4839 );
and \U$6995 ( \8895 , \8869 , \8894 );
or \U$6996 ( \8896 , \4584 , \4841 );
nand \U$6997 ( \8897 , \8896 , \4844 );
nor \U$6998 ( \8898 , \8895 , \8897 );
or \U$6999 ( \8899 , \8873 , \8898 );
or \U$7000 ( \8900 , \4678 , \4846 );
nand \U$7001 ( \8901 , \8900 , \4850 );
and \U$7002 ( \8902 , \8872 , \8901 );
or \U$7003 ( \8903 , \4715 , \4852 );
nand \U$7004 ( \8904 , \8903 , \4855 );
nor \U$7005 ( \8905 , \8902 , \8904 );
nand \U$7006 ( \8906 , \8899 , \8905 );
nor \U$7007 ( \8907 , \8892 , \8906 );
or \U$7008 ( \8908 , \8867 , \8907 );
or \U$7009 ( \8909 , \3558 , \4857 );
nand \U$7010 ( \8910 , \8909 , \4863 );
and \U$7011 ( \8911 , \8854 , \8910 );
or \U$7012 ( \8912 , \3710 , \4865 );
nand \U$7013 ( \8913 , \8912 , \4868 );
nor \U$7014 ( \8914 , \8911 , \8913 );
or \U$7015 ( \8915 , \8858 , \8914 );
or \U$7016 ( \8916 , \3862 , \4870 );
nand \U$7017 ( \8917 , \8916 , \4874 );
and \U$7018 ( \8918 , \8857 , \8917 );
or \U$7019 ( \8919 , \4011 , \4876 );
nand \U$7020 ( \8920 , \8919 , \4879 );
nor \U$7021 ( \8921 , \8918 , \8920 );
nand \U$7022 ( \8922 , \8915 , \8921 );
and \U$7023 ( \8923 , \8866 , \8922 );
or \U$7024 ( \8924 , \4144 , \4881 );
nand \U$7025 ( \8925 , \8924 , \4886 );
and \U$7026 ( \8926 , \8861 , \8925 );
or \U$7027 ( \8927 , \4261 , \4888 );
nand \U$7028 ( \8928 , \8927 , \4891 );
nor \U$7029 ( \8929 , \8926 , \8928 );
or \U$7030 ( \8930 , \8865 , \8929 );
or \U$7031 ( \8931 , \4331 , \4893 );
nand \U$7032 ( \8932 , \8931 , \4897 );
and \U$7033 ( \8933 , \8864 , \8932 );
or \U$7034 ( \8934 , \4368 , \4899 );
nand \U$7035 ( \8935 , \8934 , \4902 );
nor \U$7036 ( \8936 , \8933 , \8935 );
nand \U$7037 ( \8937 , \8930 , \8936 );
nor \U$7038 ( \8938 , \8923 , \8937 );
nand \U$7039 ( \8939 , \8908 , \8938 );
not \U$7040 ( \8940 , \8939 );
xor \U$7041 ( \8941 , \8852 , \8940 );
buf g3221_GF_PartitionCandidate( \8942_nG3221 , \8941 );
not \U$7042 ( \8943 , \7221 );
nand \U$7043 ( \8944 , \7750 , \8943 );
nor \U$7044 ( \8945 , \7568 , \6404 );
nor \U$7045 ( \8946 , \6479 , \6556 );
nand \U$7046 ( \8947 , \8945 , \8946 );
nor \U$7047 ( \8948 , \6631 , \6708 );
nor \U$7048 ( \8949 , \6784 , \6857 );
nand \U$7049 ( \8950 , \8948 , \8949 );
nor \U$7050 ( \8951 , \8947 , \8950 );
nor \U$7051 ( \8952 , \6926 , \6990 );
nor \U$7052 ( \8953 , \7050 , \7107 );
nand \U$7053 ( \8954 , \8952 , \8953 );
nor \U$7054 ( \8955 , \7145 , \7177 );
nor \U$7055 ( \8956 , \7198 , \7214 );
nand \U$7056 ( \8957 , \8955 , \8956 );
nor \U$7057 ( \8958 , \8954 , \8957 );
nand \U$7058 ( \8959 , \8951 , \8958 );
nor \U$7059 ( \8960 , \7629 , \7333 );
nor \U$7060 ( \8961 , \7378 , \7430 );
nand \U$7061 ( \8962 , \8960 , \8961 );
nor \U$7062 ( \8963 , \7485 , \7524 );
nor \U$7063 ( \8964 , \7545 , \7561 );
nand \U$7064 ( \8965 , \8963 , \8964 );
nor \U$7065 ( \8966 , \8962 , \8965 );
nor \U$7066 ( \8967 , \7649 , \7604 );
nor \U$7067 ( \8968 , \7615 , \7626 );
nand \U$7068 ( \8969 , \8967 , \8968 );
nor \U$7069 ( \8970 , \7654 , \7646 );
not \U$7070 ( \8971 , \7662 );
and \U$7071 ( \8972 , \8970 , \8971 );
or \U$7072 ( \8973 , \7646 , \7664 );
nand \U$7073 ( \8974 , \8973 , \7667 );
nor \U$7074 ( \8975 , \8972 , \8974 );
or \U$7075 ( \8976 , \8969 , \8975 );
or \U$7076 ( \8977 , \7604 , \7669 );
nand \U$7077 ( \8978 , \8977 , \7673 );
and \U$7078 ( \8979 , \8968 , \8978 );
or \U$7079 ( \8980 , \7626 , \7675 );
nand \U$7080 ( \8981 , \8980 , \7678 );
nor \U$7081 ( \8982 , \8979 , \8981 );
nand \U$7082 ( \8983 , \8976 , \8982 );
and \U$7083 ( \8984 , \8966 , \8983 );
or \U$7084 ( \8985 , \7333 , \7680 );
nand \U$7085 ( \8986 , \8985 , \7685 );
and \U$7086 ( \8987 , \8961 , \8986 );
or \U$7087 ( \8988 , \7430 , \7687 );
nand \U$7088 ( \8989 , \8988 , \7690 );
nor \U$7089 ( \8990 , \8987 , \8989 );
or \U$7090 ( \8991 , \8965 , \8990 );
or \U$7091 ( \8992 , \7524 , \7692 );
nand \U$7092 ( \8993 , \8992 , \7696 );
and \U$7093 ( \8994 , \8964 , \8993 );
or \U$7094 ( \8995 , \7561 , \7698 );
nand \U$7095 ( \8996 , \8995 , \7701 );
nor \U$7096 ( \8997 , \8994 , \8996 );
nand \U$7097 ( \8998 , \8991 , \8997 );
nor \U$7098 ( \8999 , \8984 , \8998 );
or \U$7099 ( \9000 , \8959 , \8999 );
or \U$7100 ( \9001 , \6404 , \7703 );
nand \U$7101 ( \9002 , \9001 , \7709 );
and \U$7102 ( \9003 , \8946 , \9002 );
or \U$7103 ( \9004 , \6556 , \7711 );
nand \U$7104 ( \9005 , \9004 , \7714 );
nor \U$7105 ( \9006 , \9003 , \9005 );
or \U$7106 ( \9007 , \8950 , \9006 );
or \U$7107 ( \9008 , \6708 , \7716 );
nand \U$7108 ( \9009 , \9008 , \7720 );
and \U$7109 ( \9010 , \8949 , \9009 );
or \U$7110 ( \9011 , \6857 , \7722 );
nand \U$7111 ( \9012 , \9011 , \7725 );
nor \U$7112 ( \9013 , \9010 , \9012 );
nand \U$7113 ( \9014 , \9007 , \9013 );
and \U$7114 ( \9015 , \8958 , \9014 );
or \U$7115 ( \9016 , \6990 , \7727 );
nand \U$7116 ( \9017 , \9016 , \7732 );
and \U$7117 ( \9018 , \8953 , \9017 );
or \U$7118 ( \9019 , \7107 , \7734 );
nand \U$7119 ( \9020 , \9019 , \7737 );
nor \U$7120 ( \9021 , \9018 , \9020 );
or \U$7121 ( \9022 , \8957 , \9021 );
or \U$7122 ( \9023 , \7177 , \7739 );
nand \U$7123 ( \9024 , \9023 , \7743 );
and \U$7124 ( \9025 , \8956 , \9024 );
or \U$7125 ( \9026 , \7214 , \7745 );
nand \U$7126 ( \9027 , \9026 , \7748 );
nor \U$7127 ( \9028 , \9025 , \9027 );
nand \U$7128 ( \9029 , \9022 , \9028 );
nor \U$7129 ( \9030 , \9015 , \9029 );
nand \U$7130 ( \9031 , \9000 , \9030 );
not \U$7131 ( \9032 , \9031 );
xor \U$7132 ( \9033 , \8944 , \9032 );
buf g3255_GF_PartitionCandidate( \9034_nG3255 , \9033 );
_HMUX g3256_GF_PartitionCandidate ( \9035_nG3256 , \8942_nG3221 , \9034_nG3255 , \8848 );
buf \U$7133 ( \9036 , \9035_nG3256 );
not \U$7134 ( \9037 , \4368 );
nand \U$7135 ( \9038 , \4902 , \9037 );
nand \U$7136 ( \9039 , \4723 , \3634 );
nand \U$7137 ( \9040 , \3786 , \3939 );
nor \U$7138 ( \9041 , \9039 , \9040 );
nand \U$7139 ( \9042 , \4081 , \4205 );
nand \U$7140 ( \9043 , \4300 , \4353 );
nor \U$7141 ( \9044 , \9042 , \9043 );
nand \U$7142 ( \9045 , \9041 , \9044 );
nand \U$7143 ( \9046 , \4784 , \4533 );
nand \U$7144 ( \9047 , \4640 , \4700 );
nor \U$7145 ( \9048 , \9046 , \9047 );
nand \U$7146 ( \9049 , \4804 , \4770 );
not \U$7147 ( \9050 , \4819 );
or \U$7148 ( \9051 , \9049 , \9050 );
and \U$7149 ( \9052 , \4770 , \4824 );
nor \U$7150 ( \9053 , \9052 , \4830 );
nand \U$7151 ( \9054 , \9051 , \9053 );
and \U$7152 ( \9055 , \9048 , \9054 );
and \U$7153 ( \9056 , \4533 , \4835 );
nor \U$7154 ( \9057 , \9056 , \4842 );
or \U$7155 ( \9058 , \9047 , \9057 );
and \U$7156 ( \9059 , \4700 , \4847 );
nor \U$7157 ( \9060 , \9059 , \4853 );
nand \U$7158 ( \9061 , \9058 , \9060 );
nor \U$7159 ( \9062 , \9055 , \9061 );
or \U$7160 ( \9063 , \9045 , \9062 );
and \U$7161 ( \9064 , \3634 , \4858 );
nor \U$7162 ( \9065 , \9064 , \4866 );
or \U$7163 ( \9066 , \9040 , \9065 );
and \U$7164 ( \9067 , \3939 , \4871 );
nor \U$7165 ( \9068 , \9067 , \4877 );
nand \U$7166 ( \9069 , \9066 , \9068 );
and \U$7167 ( \9070 , \9044 , \9069 );
and \U$7168 ( \9071 , \4205 , \4882 );
nor \U$7169 ( \9072 , \9071 , \4889 );
or \U$7170 ( \9073 , \9043 , \9072 );
and \U$7171 ( \9074 , \4353 , \4894 );
nor \U$7172 ( \9075 , \9074 , \4900 );
nand \U$7173 ( \9076 , \9073 , \9075 );
nor \U$7174 ( \9077 , \9070 , \9076 );
nand \U$7175 ( \9078 , \9063 , \9077 );
not \U$7176 ( \9079 , \9078 );
xor \U$7177 ( \9080 , \9038 , \9079 );
buf g31b2_GF_PartitionCandidate( \9081_nG31b2 , \9080 );
not \U$7178 ( \9082 , \7214 );
nand \U$7179 ( \9083 , \7748 , \9082 );
nand \U$7180 ( \9084 , \7569 , \6480 );
nand \U$7181 ( \9085 , \6632 , \6785 );
nor \U$7182 ( \9086 , \9084 , \9085 );
nand \U$7183 ( \9087 , \6927 , \7051 );
nand \U$7184 ( \9088 , \7146 , \7199 );
nor \U$7185 ( \9089 , \9087 , \9088 );
nand \U$7186 ( \9090 , \9086 , \9089 );
nand \U$7187 ( \9091 , \7630 , \7379 );
nand \U$7188 ( \9092 , \7486 , \7546 );
nor \U$7189 ( \9093 , \9091 , \9092 );
nand \U$7190 ( \9094 , \7650 , \7616 );
not \U$7191 ( \9095 , \7665 );
or \U$7192 ( \9096 , \9094 , \9095 );
and \U$7193 ( \9097 , \7616 , \7670 );
nor \U$7194 ( \9098 , \9097 , \7676 );
nand \U$7195 ( \9099 , \9096 , \9098 );
and \U$7196 ( \9100 , \9093 , \9099 );
and \U$7197 ( \9101 , \7379 , \7681 );
nor \U$7198 ( \9102 , \9101 , \7688 );
or \U$7199 ( \9103 , \9092 , \9102 );
and \U$7200 ( \9104 , \7546 , \7693 );
nor \U$7201 ( \9105 , \9104 , \7699 );
nand \U$7202 ( \9106 , \9103 , \9105 );
nor \U$7203 ( \9107 , \9100 , \9106 );
or \U$7204 ( \9108 , \9090 , \9107 );
and \U$7205 ( \9109 , \6480 , \7704 );
nor \U$7206 ( \9110 , \9109 , \7712 );
or \U$7207 ( \9111 , \9085 , \9110 );
and \U$7208 ( \9112 , \6785 , \7717 );
nor \U$7209 ( \9113 , \9112 , \7723 );
nand \U$7210 ( \9114 , \9111 , \9113 );
and \U$7211 ( \9115 , \9089 , \9114 );
and \U$7212 ( \9116 , \7051 , \7728 );
nor \U$7213 ( \9117 , \9116 , \7735 );
or \U$7214 ( \9118 , \9088 , \9117 );
and \U$7215 ( \9119 , \7199 , \7740 );
nor \U$7216 ( \9120 , \9119 , \7746 );
nand \U$7217 ( \9121 , \9118 , \9120 );
nor \U$7218 ( \9122 , \9115 , \9121 );
nand \U$7219 ( \9123 , \9108 , \9122 );
not \U$7220 ( \9124 , \9123 );
xor \U$7221 ( \9125 , \9083 , \9124 );
buf g31ec_GF_PartitionCandidate( \9126_nG31ec , \9125 );
_HMUX g31ed_GF_PartitionCandidate ( \9127_nG31ed , \9081_nG31b2 , \9126_nG31ec , \8848 );
buf \U$7222 ( \9128 , \9127_nG31ed );
not \U$7223 ( \9129 , \4352 );
nand \U$7224 ( \9130 , \4899 , \9129 );
nand \U$7225 ( \9131 , \8872 , \8853 );
nand \U$7226 ( \9132 , \8854 , \8856 );
nor \U$7227 ( \9133 , \9131 , \9132 );
nand \U$7228 ( \9134 , \8857 , \8860 );
nand \U$7229 ( \9135 , \8861 , \8863 );
nor \U$7230 ( \9136 , \9134 , \9135 );
nand \U$7231 ( \9137 , \9133 , \9136 );
nand \U$7232 ( \9138 , \8876 , \8868 );
nand \U$7233 ( \9139 , \8869 , \8871 );
nor \U$7234 ( \9140 , \9138 , \9139 );
nand \U$7235 ( \9141 , \8878 , \8875 );
or \U$7236 ( \9142 , \9141 , \4816 );
and \U$7237 ( \9143 , \8875 , \8882 );
nor \U$7238 ( \9144 , \9143 , \8886 );
nand \U$7239 ( \9145 , \9142 , \9144 );
and \U$7240 ( \9146 , \9140 , \9145 );
and \U$7241 ( \9147 , \8868 , \8889 );
nor \U$7242 ( \9148 , \9147 , \8894 );
or \U$7243 ( \9149 , \9139 , \9148 );
and \U$7244 ( \9150 , \8871 , \8897 );
nor \U$7245 ( \9151 , \9150 , \8901 );
nand \U$7246 ( \9152 , \9149 , \9151 );
nor \U$7247 ( \9153 , \9146 , \9152 );
or \U$7248 ( \9154 , \9137 , \9153 );
and \U$7249 ( \9155 , \8853 , \8904 );
nor \U$7250 ( \9156 , \9155 , \8910 );
or \U$7251 ( \9157 , \9132 , \9156 );
and \U$7252 ( \9158 , \8856 , \8913 );
nor \U$7253 ( \9159 , \9158 , \8917 );
nand \U$7254 ( \9160 , \9157 , \9159 );
and \U$7255 ( \9161 , \9136 , \9160 );
and \U$7256 ( \9162 , \8860 , \8920 );
nor \U$7257 ( \9163 , \9162 , \8925 );
or \U$7258 ( \9164 , \9135 , \9163 );
and \U$7259 ( \9165 , \8863 , \8928 );
nor \U$7260 ( \9166 , \9165 , \8932 );
nand \U$7261 ( \9167 , \9164 , \9166 );
nor \U$7262 ( \9168 , \9161 , \9167 );
nand \U$7263 ( \9169 , \9154 , \9168 );
not \U$7264 ( \9170 , \9169 );
xor \U$7265 ( \9171 , \9130 , \9170 );
buf g3135_GF_PartitionCandidate( \9172_nG3135 , \9171 );
not \U$7266 ( \9173 , \7198 );
nand \U$7267 ( \9174 , \7745 , \9173 );
nand \U$7268 ( \9175 , \8964 , \8945 );
nand \U$7269 ( \9176 , \8946 , \8948 );
nor \U$7270 ( \9177 , \9175 , \9176 );
nand \U$7271 ( \9178 , \8949 , \8952 );
nand \U$7272 ( \9179 , \8953 , \8955 );
nor \U$7273 ( \9180 , \9178 , \9179 );
nand \U$7274 ( \9181 , \9177 , \9180 );
nand \U$7275 ( \9182 , \8968 , \8960 );
nand \U$7276 ( \9183 , \8961 , \8963 );
nor \U$7277 ( \9184 , \9182 , \9183 );
nand \U$7278 ( \9185 , \8970 , \8967 );
or \U$7279 ( \9186 , \9185 , \7662 );
and \U$7280 ( \9187 , \8967 , \8974 );
nor \U$7281 ( \9188 , \9187 , \8978 );
nand \U$7282 ( \9189 , \9186 , \9188 );
and \U$7283 ( \9190 , \9184 , \9189 );
and \U$7284 ( \9191 , \8960 , \8981 );
nor \U$7285 ( \9192 , \9191 , \8986 );
or \U$7286 ( \9193 , \9183 , \9192 );
and \U$7287 ( \9194 , \8963 , \8989 );
nor \U$7288 ( \9195 , \9194 , \8993 );
nand \U$7289 ( \9196 , \9193 , \9195 );
nor \U$7290 ( \9197 , \9190 , \9196 );
or \U$7291 ( \9198 , \9181 , \9197 );
and \U$7292 ( \9199 , \8945 , \8996 );
nor \U$7293 ( \9200 , \9199 , \9002 );
or \U$7294 ( \9201 , \9176 , \9200 );
and \U$7295 ( \9202 , \8948 , \9005 );
nor \U$7296 ( \9203 , \9202 , \9009 );
nand \U$7297 ( \9204 , \9201 , \9203 );
and \U$7298 ( \9205 , \9180 , \9204 );
and \U$7299 ( \9206 , \8952 , \9012 );
nor \U$7300 ( \9207 , \9206 , \9017 );
or \U$7301 ( \9208 , \9179 , \9207 );
and \U$7302 ( \9209 , \8955 , \9020 );
nor \U$7303 ( \9210 , \9209 , \9024 );
nand \U$7304 ( \9211 , \9208 , \9210 );
nor \U$7305 ( \9212 , \9205 , \9211 );
nand \U$7306 ( \9213 , \9198 , \9212 );
not \U$7307 ( \9214 , \9213 );
xor \U$7308 ( \9215 , \9174 , \9214 );
buf g3177_GF_PartitionCandidate( \9216_nG3177 , \9215 );
_HMUX g3178_GF_PartitionCandidate ( \9217_nG3178 , \9172_nG3135 , \9216_nG3177 , \8848 );
buf \U$7309 ( \9218 , \9217_nG3178 );
not \U$7310 ( \9219 , \4331 );
nand \U$7311 ( \9220 , \4897 , \9219 );
nor \U$7312 ( \9221 , \4724 , \3787 );
nor \U$7313 ( \9222 , \4082 , \4301 );
nand \U$7314 ( \9223 , \9221 , \9222 );
nor \U$7315 ( \9224 , \4785 , \4641 );
not \U$7316 ( \9225 , \4825 );
and \U$7317 ( \9226 , \9224 , \9225 );
or \U$7318 ( \9227 , \4641 , \4836 );
nand \U$7319 ( \9228 , \9227 , \4848 );
nor \U$7320 ( \9229 , \9226 , \9228 );
or \U$7321 ( \9230 , \9223 , \9229 );
or \U$7322 ( \9231 , \3787 , \4859 );
nand \U$7323 ( \9232 , \9231 , \4872 );
and \U$7324 ( \9233 , \9222 , \9232 );
or \U$7325 ( \9234 , \4301 , \4883 );
nand \U$7326 ( \9235 , \9234 , \4895 );
nor \U$7327 ( \9236 , \9233 , \9235 );
nand \U$7328 ( \9237 , \9230 , \9236 );
not \U$7329 ( \9238 , \9237 );
xor \U$7330 ( \9239 , \9220 , \9238 );
buf g30ac_GF_PartitionCandidate( \9240_nG30ac , \9239 );
not \U$7331 ( \9241 , \7177 );
nand \U$7332 ( \9242 , \7743 , \9241 );
nor \U$7333 ( \9243 , \7570 , \6633 );
nor \U$7334 ( \9244 , \6928 , \7147 );
nand \U$7335 ( \9245 , \9243 , \9244 );
nor \U$7336 ( \9246 , \7631 , \7487 );
not \U$7337 ( \9247 , \7671 );
and \U$7338 ( \9248 , \9246 , \9247 );
or \U$7339 ( \9249 , \7487 , \7682 );
nand \U$7340 ( \9250 , \9249 , \7694 );
nor \U$7341 ( \9251 , \9248 , \9250 );
or \U$7342 ( \9252 , \9245 , \9251 );
or \U$7343 ( \9253 , \6633 , \7705 );
nand \U$7344 ( \9254 , \9253 , \7718 );
and \U$7345 ( \9255 , \9244 , \9254 );
or \U$7346 ( \9256 , \7147 , \7729 );
nand \U$7347 ( \9257 , \9256 , \7741 );
nor \U$7348 ( \9258 , \9255 , \9257 );
nand \U$7349 ( \9259 , \9252 , \9258 );
not \U$7350 ( \9260 , \9259 );
xor \U$7351 ( \9261 , \9242 , \9260 );
buf g30f2_GF_PartitionCandidate( \9262_nG30f2 , \9261 );
_HMUX g30f3_GF_PartitionCandidate ( \9263_nG30f3 , \9240_nG30ac , \9262_nG30f2 , \8848 );
buf \U$7352 ( \9264 , \9263_nG30f3 );
not \U$7353 ( \9265 , \4299 );
nand \U$7354 ( \9266 , \4893 , \9265 );
nor \U$7355 ( \9267 , \8873 , \8855 );
nor \U$7356 ( \9268 , \8858 , \8862 );
nand \U$7357 ( \9269 , \9267 , \9268 );
nor \U$7358 ( \9270 , \8877 , \8870 );
not \U$7359 ( \9271 , \8883 );
and \U$7360 ( \9272 , \9270 , \9271 );
or \U$7361 ( \9273 , \8870 , \8890 );
nand \U$7362 ( \9274 , \9273 , \8898 );
nor \U$7363 ( \9275 , \9272 , \9274 );
or \U$7364 ( \9276 , \9269 , \9275 );
or \U$7365 ( \9277 , \8855 , \8905 );
nand \U$7366 ( \9278 , \9277 , \8914 );
and \U$7367 ( \9279 , \9268 , \9278 );
or \U$7368 ( \9280 , \8862 , \8921 );
nand \U$7369 ( \9281 , \9280 , \8929 );
nor \U$7370 ( \9282 , \9279 , \9281 );
nand \U$7371 ( \9283 , \9276 , \9282 );
not \U$7372 ( \9284 , \9283 );
xor \U$7373 ( \9285 , \9266 , \9284 );
buf g301d_GF_PartitionCandidate( \9286_nG301d , \9285 );
not \U$7374 ( \9287 , \7145 );
nand \U$7375 ( \9288 , \7739 , \9287 );
nor \U$7376 ( \9289 , \8965 , \8947 );
nor \U$7377 ( \9290 , \8950 , \8954 );
nand \U$7378 ( \9291 , \9289 , \9290 );
nor \U$7379 ( \9292 , \8969 , \8962 );
not \U$7380 ( \9293 , \8975 );
and \U$7381 ( \9294 , \9292 , \9293 );
or \U$7382 ( \9295 , \8962 , \8982 );
nand \U$7383 ( \9296 , \9295 , \8990 );
nor \U$7384 ( \9297 , \9294 , \9296 );
or \U$7385 ( \9298 , \9291 , \9297 );
or \U$7386 ( \9299 , \8947 , \8997 );
nand \U$7387 ( \9300 , \9299 , \9006 );
and \U$7388 ( \9301 , \9290 , \9300 );
or \U$7389 ( \9302 , \8954 , \9013 );
nand \U$7390 ( \9303 , \9302 , \9021 );
nor \U$7391 ( \9304 , \9301 , \9303 );
nand \U$7392 ( \9305 , \9298 , \9304 );
not \U$7393 ( \9306 , \9305 );
xor \U$7394 ( \9307 , \9288 , \9306 );
buf g3065_GF_PartitionCandidate( \9308_nG3065 , \9307 );
_HMUX g3066_GF_PartitionCandidate ( \9309_nG3066 , \9286_nG301d , \9308_nG3065 , \8848 );
buf \U$7395 ( \9310 , \9309_nG3066 );
not \U$7396 ( \9311 , \4261 );
nand \U$7397 ( \9312 , \4891 , \9311 );
nor \U$7398 ( \9313 , \9047 , \9039 );
nor \U$7399 ( \9314 , \9040 , \9042 );
nand \U$7400 ( \9315 , \9313 , \9314 );
nor \U$7401 ( \9316 , \9049 , \9046 );
and \U$7402 ( \9317 , \9316 , \4819 );
or \U$7403 ( \9318 , \9046 , \9053 );
nand \U$7404 ( \9319 , \9318 , \9057 );
nor \U$7405 ( \9320 , \9317 , \9319 );
or \U$7406 ( \9321 , \9315 , \9320 );
or \U$7407 ( \9322 , \9039 , \9060 );
nand \U$7408 ( \9323 , \9322 , \9065 );
and \U$7409 ( \9324 , \9314 , \9323 );
or \U$7410 ( \9325 , \9042 , \9068 );
nand \U$7411 ( \9326 , \9325 , \9072 );
nor \U$7412 ( \9327 , \9324 , \9326 );
nand \U$7413 ( \9328 , \9321 , \9327 );
not \U$7414 ( \9329 , \9328 );
xor \U$7415 ( \9330 , \9312 , \9329 );
buf g2f88_GF_PartitionCandidate( \9331_nG2f88 , \9330 );
not \U$7416 ( \9332 , \7107 );
nand \U$7417 ( \9333 , \7737 , \9332 );
nor \U$7418 ( \9334 , \9092 , \9084 );
nor \U$7419 ( \9335 , \9085 , \9087 );
nand \U$7420 ( \9336 , \9334 , \9335 );
nor \U$7421 ( \9337 , \9094 , \9091 );
and \U$7422 ( \9338 , \9337 , \7665 );
or \U$7423 ( \9339 , \9091 , \9098 );
nand \U$7424 ( \9340 , \9339 , \9102 );
nor \U$7425 ( \9341 , \9338 , \9340 );
or \U$7426 ( \9342 , \9336 , \9341 );
or \U$7427 ( \9343 , \9084 , \9105 );
nand \U$7428 ( \9344 , \9343 , \9110 );
and \U$7429 ( \9345 , \9335 , \9344 );
or \U$7430 ( \9346 , \9087 , \9113 );
nand \U$7431 ( \9347 , \9346 , \9117 );
nor \U$7432 ( \9348 , \9345 , \9347 );
nand \U$7433 ( \9349 , \9342 , \9348 );
not \U$7434 ( \9350 , \9349 );
xor \U$7435 ( \9351 , \9333 , \9350 );
buf g2fd4_GF_PartitionCandidate( \9352_nG2fd4 , \9351 );
_HMUX g2fd5_GF_PartitionCandidate ( \9353_nG2fd5 , \9331_nG2f88 , \9352_nG2fd4 , \8848 );
buf \U$7436 ( \9354 , \9353_nG2fd5 );
not \U$7437 ( \9355 , \4204 );
nand \U$7438 ( \9356 , \4888 , \9355 );
nor \U$7439 ( \9357 , \9139 , \9131 );
nor \U$7440 ( \9358 , \9132 , \9134 );
nand \U$7441 ( \9359 , \9357 , \9358 );
nor \U$7442 ( \9360 , \9141 , \9138 );
and \U$7443 ( \9361 , \9360 , \8879 );
or \U$7444 ( \9362 , \9138 , \9144 );
nand \U$7445 ( \9363 , \9362 , \9148 );
nor \U$7446 ( \9364 , \9361 , \9363 );
or \U$7447 ( \9365 , \9359 , \9364 );
or \U$7448 ( \9366 , \9131 , \9151 );
nand \U$7449 ( \9367 , \9366 , \9156 );
and \U$7450 ( \9368 , \9358 , \9367 );
or \U$7451 ( \9369 , \9134 , \9159 );
nand \U$7452 ( \9370 , \9369 , \9163 );
nor \U$7453 ( \9371 , \9368 , \9370 );
nand \U$7454 ( \9372 , \9365 , \9371 );
not \U$7455 ( \9373 , \9372 );
xor \U$7456 ( \9374 , \9356 , \9373 );
buf g2eeb_GF_PartitionCandidate( \9375_nG2eeb , \9374 );
not \U$7457 ( \9376 , \7050 );
nand \U$7458 ( \9377 , \7734 , \9376 );
nor \U$7459 ( \9378 , \9183 , \9175 );
nor \U$7460 ( \9379 , \9176 , \9178 );
nand \U$7461 ( \9380 , \9378 , \9379 );
nor \U$7462 ( \9381 , \9185 , \9182 );
and \U$7463 ( \9382 , \9381 , \8971 );
or \U$7464 ( \9383 , \9182 , \9188 );
nand \U$7465 ( \9384 , \9383 , \9192 );
nor \U$7466 ( \9385 , \9382 , \9384 );
or \U$7467 ( \9386 , \9380 , \9385 );
or \U$7468 ( \9387 , \9175 , \9195 );
nand \U$7469 ( \9388 , \9387 , \9200 );
and \U$7470 ( \9389 , \9379 , \9388 );
or \U$7471 ( \9390 , \9178 , \9203 );
nand \U$7472 ( \9391 , \9390 , \9207 );
nor \U$7473 ( \9392 , \9389 , \9391 );
nand \U$7474 ( \9393 , \9386 , \9392 );
not \U$7475 ( \9394 , \9393 );
xor \U$7476 ( \9395 , \9377 , \9394 );
buf g2f3b_GF_PartitionCandidate( \9396_nG2f3b , \9395 );
_HMUX g2f3c_GF_PartitionCandidate ( \9397_nG2f3c , \9375_nG2eeb , \9396_nG2f3b , \8848 );
buf \U$7477 ( \9398 , \9397_nG2f3c );
not \U$7478 ( \9399 , \4144 );
nand \U$7479 ( \9400 , \4886 , \9399 );
nand \U$7480 ( \9401 , \4725 , \4083 );
not \U$7481 ( \9402 , \4837 );
or \U$7482 ( \9403 , \9401 , \9402 );
and \U$7483 ( \9404 , \4083 , \4860 );
nor \U$7484 ( \9405 , \9404 , \4884 );
nand \U$7485 ( \9406 , \9403 , \9405 );
not \U$7486 ( \9407 , \9406 );
xor \U$7487 ( \9408 , \9400 , \9407 );
buf g2e49_GF_PartitionCandidate( \9409_nG2e49 , \9408 );
not \U$7488 ( \9410 , \6990 );
nand \U$7489 ( \9411 , \7732 , \9410 );
nand \U$7490 ( \9412 , \7571 , \6929 );
not \U$7491 ( \9413 , \7683 );
or \U$7492 ( \9414 , \9412 , \9413 );
and \U$7493 ( \9415 , \6929 , \7706 );
nor \U$7494 ( \9416 , \9415 , \7730 );
nand \U$7495 ( \9417 , \9414 , \9416 );
not \U$7496 ( \9418 , \9417 );
xor \U$7497 ( \9419 , \9411 , \9418 );
buf g2e9a_GF_PartitionCandidate( \9420_nG2e9a , \9419 );
_HMUX g2e9b_GF_PartitionCandidate ( \9421_nG2e9b , \9409_nG2e49 , \9420_nG2e9a , \8848 );
buf \U$7498 ( \9422 , \9421_nG2e9b );
not \U$7499 ( \9423 , \4080 );
nand \U$7500 ( \9424 , \4881 , \9423 );
nand \U$7501 ( \9425 , \8874 , \8859 );
not \U$7502 ( \9426 , \8891 );
or \U$7503 ( \9427 , \9425 , \9426 );
and \U$7504 ( \9428 , \8859 , \8906 );
nor \U$7505 ( \9429 , \9428 , \8922 );
nand \U$7506 ( \9430 , \9427 , \9429 );
not \U$7507 ( \9431 , \9430 );
xor \U$7508 ( \9432 , \9424 , \9431 );
buf g2d9e_GF_PartitionCandidate( \9433_nG2d9e , \9432 );
not \U$7509 ( \9434 , \6926 );
nand \U$7510 ( \9435 , \7727 , \9434 );
nand \U$7511 ( \9436 , \8966 , \8951 );
not \U$7512 ( \9437 , \8983 );
or \U$7513 ( \9438 , \9436 , \9437 );
and \U$7514 ( \9439 , \8951 , \8998 );
nor \U$7515 ( \9440 , \9439 , \9014 );
nand \U$7516 ( \9441 , \9438 , \9440 );
not \U$7517 ( \9442 , \9441 );
xor \U$7518 ( \9443 , \9435 , \9442 );
buf g2df7_GF_PartitionCandidate( \9444_nG2df7 , \9443 );
_HMUX g2df8_GF_PartitionCandidate ( \9445_nG2df8 , \9433_nG2d9e , \9444_nG2df7 , \8848 );
buf \U$7519 ( \9446 , \9445_nG2df8 );
not \U$7520 ( \9447 , \4011 );
nand \U$7521 ( \9448 , \4879 , \9447 );
nand \U$7522 ( \9449 , \9048 , \9041 );
not \U$7523 ( \9450 , \9054 );
or \U$7524 ( \9451 , \9449 , \9450 );
and \U$7525 ( \9452 , \9041 , \9061 );
nor \U$7526 ( \9453 , \9452 , \9069 );
nand \U$7527 ( \9454 , \9451 , \9453 );
not \U$7528 ( \9455 , \9454 );
xor \U$7529 ( \9456 , \9448 , \9455 );
buf g2ce8_GF_PartitionCandidate( \9457_nG2ce8 , \9456 );
not \U$7530 ( \9458 , \6857 );
nand \U$7531 ( \9459 , \7725 , \9458 );
nand \U$7532 ( \9460 , \9093 , \9086 );
not \U$7533 ( \9461 , \9099 );
or \U$7534 ( \9462 , \9460 , \9461 );
and \U$7535 ( \9463 , \9086 , \9106 );
nor \U$7536 ( \9464 , \9463 , \9114 );
nand \U$7537 ( \9465 , \9462 , \9464 );
not \U$7538 ( \9466 , \9465 );
xor \U$7539 ( \9467 , \9459 , \9466 );
buf g2d44_GF_PartitionCandidate( \9468_nG2d44 , \9467 );
_HMUX g2d45_GF_PartitionCandidate ( \9469_nG2d45 , \9457_nG2ce8 , \9468_nG2d44 , \8848 );
buf \U$7540 ( \9470 , \9469_nG2d45 );
not \U$7541 ( \9471 , \3938 );
nand \U$7542 ( \9472 , \4876 , \9471 );
nand \U$7543 ( \9473 , \9140 , \9133 );
not \U$7544 ( \9474 , \9145 );
or \U$7545 ( \9475 , \9473 , \9474 );
and \U$7546 ( \9476 , \9133 , \9152 );
nor \U$7547 ( \9477 , \9476 , \9160 );
nand \U$7548 ( \9478 , \9475 , \9477 );
not \U$7549 ( \9479 , \9478 );
xor \U$7550 ( \9480 , \9472 , \9479 );
buf g2c2b_GF_PartitionCandidate( \9481_nG2c2b , \9480 );
not \U$7551 ( \9482 , \6784 );
nand \U$7552 ( \9483 , \7722 , \9482 );
nand \U$7553 ( \9484 , \9184 , \9177 );
not \U$7554 ( \9485 , \9189 );
or \U$7555 ( \9486 , \9484 , \9485 );
and \U$7556 ( \9487 , \9177 , \9196 );
nor \U$7557 ( \9488 , \9487 , \9204 );
nand \U$7558 ( \9489 , \9486 , \9488 );
not \U$7559 ( \9490 , \9489 );
xor \U$7560 ( \9491 , \9483 , \9490 );
buf g2c8b_GF_PartitionCandidate( \9492_nG2c8b , \9491 );
_HMUX g2c8c_GF_PartitionCandidate ( \9493_nG2c8c , \9481_nG2c2b , \9492_nG2c8b , \8848 );
buf \U$7561 ( \9494 , \9493_nG2c8c );
not \U$7562 ( \9495 , \3862 );
nand \U$7563 ( \9496 , \4874 , \9495 );
nand \U$7564 ( \9497 , \9224 , \9221 );
or \U$7565 ( \9498 , \9497 , \4825 );
and \U$7566 ( \9499 , \9221 , \9228 );
nor \U$7567 ( \9500 , \9499 , \9232 );
nand \U$7568 ( \9501 , \9498 , \9500 );
not \U$7569 ( \9502 , \9501 );
xor \U$7570 ( \9503 , \9496 , \9502 );
buf g2b6b_GF_PartitionCandidate( \9504_nG2b6b , \9503 );
not \U$7571 ( \9505 , \6708 );
nand \U$7572 ( \9506 , \7720 , \9505 );
nand \U$7573 ( \9507 , \9246 , \9243 );
or \U$7574 ( \9508 , \9507 , \7671 );
and \U$7575 ( \9509 , \9243 , \9250 );
nor \U$7576 ( \9510 , \9509 , \9254 );
nand \U$7577 ( \9511 , \9508 , \9510 );
not \U$7578 ( \9512 , \9511 );
xor \U$7579 ( \9513 , \9506 , \9512 );
buf g2bca_GF_PartitionCandidate( \9514_nG2bca , \9513 );
_HMUX g2bcb_GF_PartitionCandidate ( \9515_nG2bcb , \9504_nG2b6b , \9514_nG2bca , \8848 );
buf \U$7580 ( \9516 , \9515_nG2bcb );
not \U$7581 ( \9517 , \3785 );
nand \U$7582 ( \9518 , \4870 , \9517 );
nand \U$7583 ( \9519 , \9270 , \9267 );
or \U$7584 ( \9520 , \9519 , \8883 );
and \U$7585 ( \9521 , \9267 , \9274 );
nor \U$7586 ( \9522 , \9521 , \9278 );
nand \U$7587 ( \9523 , \9520 , \9522 );
not \U$7588 ( \9524 , \9523 );
xor \U$7589 ( \9525 , \9518 , \9524 );
buf g2aac_GF_PartitionCandidate( \9526_nG2aac , \9525 );
not \U$7590 ( \9527 , \6631 );
nand \U$7591 ( \9528 , \7716 , \9527 );
nand \U$7592 ( \9529 , \9292 , \9289 );
or \U$7593 ( \9530 , \9529 , \8975 );
and \U$7594 ( \9531 , \9289 , \9296 );
nor \U$7595 ( \9532 , \9531 , \9300 );
nand \U$7596 ( \9533 , \9530 , \9532 );
not \U$7597 ( \9534 , \9533 );
xor \U$7598 ( \9535 , \9528 , \9534 );
buf g2b0b_GF_PartitionCandidate( \9536_nG2b0b , \9535 );
_HMUX g2b0c_GF_PartitionCandidate ( \9537_nG2b0c , \9526_nG2aac , \9536_nG2b0b , \8848 );
buf \U$7599 ( \9538 , \9537_nG2b0c );
not \U$7600 ( \9539 , \3710 );
nand \U$7601 ( \9540 , \4868 , \9539 );
nand \U$7602 ( \9541 , \9316 , \9313 );
or \U$7603 ( \9542 , \9541 , \9050 );
and \U$7604 ( \9543 , \9313 , \9319 );
nor \U$7605 ( \9544 , \9543 , \9323 );
nand \U$7606 ( \9545 , \9542 , \9544 );
not \U$7607 ( \9546 , \9545 );
xor \U$7608 ( \9547 , \9540 , \9546 );
buf g29d8_GF_PartitionCandidate( \9548_nG29d8 , \9547 );
not \U$7609 ( \9549 , \6556 );
nand \U$7610 ( \9550 , \7714 , \9549 );
nand \U$7611 ( \9551 , \9337 , \9334 );
or \U$7612 ( \9552 , \9551 , \9095 );
and \U$7613 ( \9553 , \9334 , \9340 );
nor \U$7614 ( \9554 , \9553 , \9344 );
nand \U$7615 ( \9555 , \9552 , \9554 );
not \U$7616 ( \9556 , \9555 );
xor \U$7617 ( \9557 , \9550 , \9556 );
buf g2a4c_GF_PartitionCandidate( \9558_nG2a4c , \9557 );
_HMUX g2a4d_GF_PartitionCandidate ( \9559_nG2a4d , \9548_nG29d8 , \9558_nG2a4c , \8848 );
buf \U$7618 ( \9560 , \9559_nG2a4d );
not \U$7619 ( \9561 , \3633 );
nand \U$7620 ( \9562 , \4865 , \9561 );
nand \U$7621 ( \9563 , \9360 , \9357 );
or \U$7622 ( \9564 , \9563 , \4816 );
and \U$7623 ( \9565 , \9357 , \9363 );
nor \U$7624 ( \9566 , \9565 , \9367 );
nand \U$7625 ( \9567 , \9564 , \9566 );
not \U$7626 ( \9568 , \9567 );
xor \U$7627 ( \9569 , \9562 , \9568 );
buf g28f0_GF_PartitionCandidate( \9570_nG28f0 , \9569 );
not \U$7628 ( \9571 , \6479 );
nand \U$7629 ( \9572 , \7711 , \9571 );
nand \U$7630 ( \9573 , \9381 , \9378 );
or \U$7631 ( \9574 , \9573 , \7662 );
and \U$7632 ( \9575 , \9378 , \9384 );
nor \U$7633 ( \9576 , \9575 , \9388 );
nand \U$7634 ( \9577 , \9574 , \9576 );
not \U$7635 ( \9578 , \9577 );
xor \U$7636 ( \9579 , \9572 , \9578 );
buf g2963_GF_PartitionCandidate( \9580_nG2963 , \9579 );
_HMUX g2964_GF_PartitionCandidate ( \9581_nG2964 , \9570_nG28f0 , \9580_nG2963 , \8848 );
buf \U$7637 ( \9582 , \9581_nG2964 );
not \U$7638 ( \9583 , \3558 );
nand \U$7639 ( \9584 , \4863 , \9583 );
xor \U$7640 ( \9585 , \9584 , \4861 );
buf g2810_GF_PartitionCandidate( \9586_nG2810 , \9585 );
not \U$7641 ( \9587 , \6404 );
nand \U$7642 ( \9588 , \7709 , \9587 );
xor \U$7643 ( \9589 , \9588 , \7707 );
buf g287c_GF_PartitionCandidate( \9590_nG287c , \9589 );
_HMUX g287d_GF_PartitionCandidate ( \9591_nG287d , \9586_nG2810 , \9590_nG287c , \8848 );
buf \U$7644 ( \9592 , \9591_nG287d );
not \U$7645 ( \9593 , \4722 );
nand \U$7646 ( \9594 , \4857 , \9593 );
xor \U$7647 ( \9595 , \9594 , \8907 );
buf g2737_GF_PartitionCandidate( \9596_nG2737 , \9595 );
not \U$7648 ( \9597 , \7568 );
nand \U$7649 ( \9598 , \7703 , \9597 );
xor \U$7650 ( \9599 , \9598 , \8999 );
buf g27a3_GF_PartitionCandidate( \9600_nG27a3 , \9599 );
_HMUX g27a4_GF_PartitionCandidate ( \9601_nG27a4 , \9596_nG2737 , \9600_nG27a3 , \8848 );
buf \U$7651 ( \9602 , \9601_nG27a4 );
not \U$7652 ( \9603 , \4715 );
nand \U$7653 ( \9604 , \4855 , \9603 );
xor \U$7654 ( \9605 , \9604 , \9062 );
buf g2662_GF_PartitionCandidate( \9606_nG2662 , \9605 );
not \U$7655 ( \9607 , \7561 );
nand \U$7656 ( \9608 , \7701 , \9607 );
xor \U$7657 ( \9609 , \9608 , \9107 );
buf g26ca_GF_PartitionCandidate( \9610_nG26ca , \9609 );
_HMUX g26cb_GF_PartitionCandidate ( \9611_nG26cb , \9606_nG2662 , \9610_nG26ca , \8848 );
buf \U$7658 ( \9612 , \9611_nG26cb );
not \U$7659 ( \9613 , \4699 );
nand \U$7660 ( \9614 , \4852 , \9613 );
xor \U$7661 ( \9615 , \9614 , \9153 );
buf g258f_GF_PartitionCandidate( \9616_nG258f , \9615 );
not \U$7662 ( \9617 , \7545 );
nand \U$7663 ( \9618 , \7698 , \9617 );
xor \U$7664 ( \9619 , \9618 , \9197 );
buf g25f9_GF_PartitionCandidate( \9620_nG25f9 , \9619 );
_HMUX g25fa_GF_PartitionCandidate ( \9621_nG25fa , \9616_nG258f , \9620_nG25f9 , \8848 );
buf \U$7665 ( \9622 , \9621_nG25fa );
not \U$7666 ( \9623 , \4678 );
nand \U$7667 ( \9624 , \4850 , \9623 );
xor \U$7668 ( \9625 , \9624 , \9229 );
buf g24bf_GF_PartitionCandidate( \9626_nG24bf , \9625 );
not \U$7669 ( \9627 , \7524 );
nand \U$7670 ( \9628 , \7696 , \9627 );
xor \U$7671 ( \9629 , \9628 , \9251 );
buf g2524_GF_PartitionCandidate( \9630_nG2524 , \9629 );
_HMUX g2525_GF_PartitionCandidate ( \9631_nG2525 , \9626_nG24bf , \9630_nG2524 , \8848 );
buf \U$7672 ( \9632 , \9631_nG2525 );
not \U$7673 ( \9633 , \4639 );
nand \U$7674 ( \9634 , \4846 , \9633 );
xor \U$7675 ( \9635 , \9634 , \9275 );
buf g23cd_GF_PartitionCandidate( \9636_nG23cd , \9635 );
not \U$7676 ( \9637 , \7485 );
nand \U$7677 ( \9638 , \7692 , \9637 );
xor \U$7678 ( \9639 , \9638 , \9297 );
buf g2459_GF_PartitionCandidate( \9640_nG2459 , \9639 );
_HMUX g245a_GF_PartitionCandidate ( \9641_nG245a , \9636_nG23cd , \9640_nG2459 , \8848 );
buf \U$7679 ( \9642 , \9641_nG245a );
not \U$7680 ( \9643 , \4584 );
nand \U$7681 ( \9644 , \4844 , \9643 );
xor \U$7682 ( \9645 , \9644 , \9320 );
buf g22e6_GF_PartitionCandidate( \9646_nG22e6 , \9645 );
not \U$7683 ( \9647 , \7430 );
nand \U$7684 ( \9648 , \7690 , \9647 );
xor \U$7685 ( \9649 , \9648 , \9341 );
buf g2340_GF_PartitionCandidate( \9650_nG2340 , \9649 );
_HMUX g2341_GF_PartitionCandidate ( \9651_nG2341 , \9646_nG22e6 , \9650_nG2340 , \8848 );
buf \U$7686 ( \9652 , \9651_nG2341 );
not \U$7687 ( \9653 , \4532 );
nand \U$7688 ( \9654 , \4841 , \9653 );
xor \U$7689 ( \9655 , \9654 , \9364 );
buf g21f2_GF_PartitionCandidate( \9656_nG21f2 , \9655 );
not \U$7690 ( \9657 , \7378 );
nand \U$7691 ( \9658 , \7687 , \9657 );
xor \U$7692 ( \9659 , \9658 , \9385 );
buf g228b_GF_PartitionCandidate( \9660_nG228b , \9659 );
_HMUX g228c_GF_PartitionCandidate ( \9661_nG228c , \9656_nG21f2 , \9660_nG228b , \8848 );
buf \U$7693 ( \9662 , \9661_nG228c );
not \U$7694 ( \9663 , \4487 );
nand \U$7695 ( \9664 , \4839 , \9663 );
xor \U$7696 ( \9665 , \9664 , \9402 );
buf g210a_GF_PartitionCandidate( \9666_nG210a , \9665 );
not \U$7697 ( \9667 , \7333 );
nand \U$7698 ( \9668 , \7685 , \9667 );
xor \U$7699 ( \9669 , \9668 , \9413 );
buf g2158_GF_PartitionCandidate( \9670_nG2158 , \9669 );
_HMUX g2159_GF_PartitionCandidate ( \9671_nG2159 , \9666_nG210a , \9670_nG2158 , \8848 );
buf \U$7700 ( \9672 , \9671_nG2159 );
not \U$7701 ( \9673 , \4783 );
nand \U$7702 ( \9674 , \4834 , \9673 );
xor \U$7703 ( \9675 , \9674 , \9426 );
buf g202e_GF_PartitionCandidate( \9676_nG202e , \9675 );
not \U$7704 ( \9677 , \7629 );
nand \U$7705 ( \9678 , \7680 , \9677 );
xor \U$7706 ( \9679 , \9678 , \9437 );
buf g20bb_GF_PartitionCandidate( \9680_nG20bb , \9679 );
_HMUX g20bc_GF_PartitionCandidate ( \9681_nG20bc , \9676_nG202e , \9680_nG20bb , \8848 );
buf \U$7707 ( \9682 , \9681_nG20bc );
not \U$7708 ( \9683 , \4780 );
nand \U$7709 ( \9684 , \4832 , \9683 );
xor \U$7710 ( \9685 , \9684 , \9450 );
buf g1f5c_GF_PartitionCandidate( \9686_nG1f5c , \9685 );
not \U$7711 ( \9687 , \7626 );
nand \U$7712 ( \9688 , \7678 , \9687 );
xor \U$7713 ( \9689 , \9688 , \9461 );
buf g1fa0_GF_PartitionCandidate( \9690_nG1fa0 , \9689 );
_HMUX g1fa1_GF_PartitionCandidate ( \9691_nG1fa1 , \9686_nG1f5c , \9690_nG1fa0 , \8848 );
buf \U$7714 ( \9692 , \9691_nG1fa1 );
buf \U$7719 ( \9693 , RI995f080_2);
buf \U$7720 ( \9694 , RI995f008_3);
buf \U$7721 ( \9695 , RI995ef90_4);
buf \U$7722 ( \9696 , RI995ef18_5);
buf \U$7723 ( \9697 , RI995eea0_6);
buf \U$7724 ( \9698 , RI995ee28_7);
buf \U$7725 ( \9699 , RI995edb0_8);
buf \U$7726 ( \9700 , RI995ed38_9);
buf \U$7727 ( \9701 , RI995ecc0_10);
buf \U$7728 ( \9702 , RI995ec48_11);
buf \U$7729 ( \9703 , RI995ebd0_12);
and \U$7730 ( \9704 , \9702 , \9703 );
and \U$7731 ( \9705 , \9701 , \9704 );
and \U$7732 ( \9706 , \9700 , \9705 );
and \U$7733 ( \9707 , \9699 , \9706 );
and \U$7734 ( \9708 , \9698 , \9707 );
and \U$7735 ( \9709 , \9697 , \9708 );
and \U$7736 ( \9710 , \9696 , \9709 );
and \U$7737 ( \9711 , \9695 , \9710 );
and \U$7738 ( \9712 , \9694 , \9711 );
xor \U$7739 ( \9713 , \9693 , \9712 );
buf \U$7740 ( \9714 , \9713 );
buf \U$7741 ( \9715 , \9714 );
not \U$7742 ( \9716 , RI9921f28_596);
nor \U$7743 ( \9717 , RI9921d48_600, RI9921dc0_599, RI9921e38_598, RI9921eb0_597, \9716 , RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7744 ( \9718 , RI995e450_236, \9717 );
not \U$7745 ( \9719 , RI9921d48_600);
not \U$7746 ( \9720 , RI9921dc0_599);
not \U$7747 ( \9721 , RI9921e38_598);
not \U$7748 ( \9722 , RI9921eb0_597);
nor \U$7749 ( \9723 , \9719 , \9720 , \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7750 ( \9724 , RI9967078_223, \9723 );
nor \U$7751 ( \9725 , RI9921d48_600, \9720 , \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7752 ( \9726 , RI9967690_210, \9725 );
nor \U$7753 ( \9727 , \9719 , RI9921dc0_599, \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7754 ( \9728 , RI890fba0_197, \9727 );
nor \U$7755 ( \9729 , RI9921d48_600, RI9921dc0_599, \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7756 ( \9730 , RI8918b88_184, \9729 );
nor \U$7757 ( \9731 , \9719 , \9720 , RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7758 ( \9732 , RI89253b0_171, \9731 );
nor \U$7759 ( \9733 , RI9921d48_600, \9720 , RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7760 ( \9734 , RI8930dc8_158, \9733 );
nor \U$7761 ( \9735 , \9719 , RI9921dc0_599, RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7762 ( \9736 , RI8939db0_145, \9735 );
nor \U$7763 ( \9737 , RI9921d48_600, RI9921dc0_599, RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7764 ( \9738 , RI89465d8_132, \9737 );
nor \U$7765 ( \9739 , \9719 , \9720 , \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7766 ( \9740 , RI89ec640_119, \9739 );
nor \U$7767 ( \9741 , RI9921d48_600, \9720 , \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7768 ( \9742 , RI9776f80_106, \9741 );
nor \U$7769 ( \9743 , \9719 , RI9921dc0_599, \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7770 ( \9744 , RI9808480_93, \9743 );
nor \U$7771 ( \9745 , RI9921d48_600, RI9921dc0_599, \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7772 ( \9746 , RI9808a98_80, \9745 );
nor \U$7773 ( \9747 , \9719 , \9720 , RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7774 ( \9748 , RI9819730_67, \9747 );
nor \U$7775 ( \9749 , RI9921d48_600, \9720 , RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7776 ( \9750 , RI98abc38_54, \9749 );
nor \U$7777 ( \9751 , \9719 , RI9921dc0_599, RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7778 ( \9752 , RI98bc8d0_41, \9751 );
nor \U$7779 ( \9753 , RI9921d48_600, RI9921dc0_599, RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$7780 ( \9754 , RI994ddd0_28, \9753 );
or \U$7781 ( \9755 , \9718 , \9724 , \9726 , \9728 , \9730 , \9732 , \9734 , \9736 , \9738 , \9740 , \9742 , \9744 , \9746 , \9748 , \9750 , \9752 , \9754 );
buf \U$7782 ( \9756 , RI9921fa0_595);
buf \U$7783 ( \9757 , RI9922018_594);
buf \U$7784 ( \9758 , RI9922090_593);
buf \U$7785 ( \9759 , RI9922108_592);
buf \U$7786 ( \9760 , RI9922180_591);
buf \U$7787 ( \9761 , RI99221f8_590);
buf \U$7788 ( \9762 , RI9922270_589);
buf \U$7789 ( \9763 , RI99222e8_588);
buf \U$7790 ( \9764 , RI9921f28_596);
buf \U$7791 ( \9765 , RI9921d48_600);
buf \U$7792 ( \9766 , RI9921dc0_599);
buf \U$7793 ( \9767 , RI9921e38_598);
buf \U$7794 ( \9768 , RI9921eb0_597);
or \U$7795 ( \9769 , \9765 , \9766 , \9767 , \9768 );
and \U$7796 ( \9770 , \9764 , \9769 );
or \U$7797 ( \9771 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9770 );
buf \U$7798 ( \9772 , \9771 );
_DC g3a87 ( \9773_nG3a87 , \9755 , \9772 );
buf \U$7799 ( \9774 , \9773_nG3a87 );
not \U$7800 ( \9775 , \9774 );
xor \U$7801 ( \9776 , \9715 , \9775 );
xor \U$7802 ( \9777 , \9694 , \9711 );
buf \U$7803 ( \9778 , \9777 );
buf \U$7804 ( \9779 , \9778 );
and \U$7805 ( \9780 , RI995e3d8_237, \9717 );
and \U$7806 ( \9781 , RI99669e8_224, \9723 );
and \U$7807 ( \9782 , RI9967618_211, \9725 );
and \U$7808 ( \9783 , RI890fb28_198, \9727 );
and \U$7809 ( \9784 , RI8918b10_185, \9729 );
and \U$7810 ( \9785 , RI8925338_172, \9731 );
and \U$7811 ( \9786 , RI8930d50_159, \9733 );
and \U$7812 ( \9787 , RI8939d38_146, \9735 );
and \U$7813 ( \9788 , RI8946560_133, \9737 );
and \U$7814 ( \9789 , RI89ec5c8_120, \9739 );
and \U$7815 ( \9790 , RI9776f08_107, \9741 );
and \U$7816 ( \9791 , RI9808408_94, \9743 );
and \U$7817 ( \9792 , RI9808a20_81, \9745 );
and \U$7818 ( \9793 , RI98196b8_68, \9747 );
and \U$7819 ( \9794 , RI98abbc0_55, \9749 );
and \U$7820 ( \9795 , RI98bc858_42, \9751 );
and \U$7821 ( \9796 , RI994dd58_29, \9753 );
or \U$7822 ( \9797 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 );
_DC g3a63 ( \9798_nG3a63 , \9797 , \9772 );
buf \U$7823 ( \9799 , \9798_nG3a63 );
not \U$7824 ( \9800 , \9799 );
and \U$7825 ( \9801 , \9779 , \9800 );
xor \U$7826 ( \9802 , \9695 , \9710 );
buf \U$7827 ( \9803 , \9802 );
buf \U$7828 ( \9804 , \9803 );
and \U$7829 ( \9805 , RI9959fe0_238, \9717 );
and \U$7830 ( \9806 , RI995e978_225, \9723 );
and \U$7831 ( \9807 , RI99675a0_212, \9725 );
and \U$7832 ( \9808 , RI890fab0_199, \9727 );
and \U$7833 ( \9809 , RI8918a98_186, \9729 );
and \U$7834 ( \9810 , RI89252c0_173, \9731 );
and \U$7835 ( \9811 , RI8930cd8_160, \9733 );
and \U$7836 ( \9812 , RI8939cc0_147, \9735 );
and \U$7837 ( \9813 , RI89464e8_134, \9737 );
and \U$7838 ( \9814 , RI89ec550_121, \9739 );
and \U$7839 ( \9815 , RI9776e90_108, \9741 );
and \U$7840 ( \9816 , RI9808390_95, \9743 );
and \U$7841 ( \9817 , RI98089a8_82, \9745 );
and \U$7842 ( \9818 , RI9819640_69, \9747 );
and \U$7843 ( \9819 , RI98abb48_56, \9749 );
and \U$7844 ( \9820 , RI98bc7e0_43, \9751 );
and \U$7845 ( \9821 , RI994dce0_30, \9753 );
or \U$7846 ( \9822 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 );
_DC g38dc ( \9823_nG38dc , \9822 , \9772 );
buf \U$7847 ( \9824 , \9823_nG38dc );
not \U$7848 ( \9825 , \9824 );
and \U$7849 ( \9826 , \9804 , \9825 );
xor \U$7850 ( \9827 , \9696 , \9709 );
buf \U$7851 ( \9828 , \9827 );
buf \U$7852 ( \9829 , \9828 );
and \U$7853 ( \9830 , RI9959f68_239, \9717 );
and \U$7854 ( \9831 , RI995e900_226, \9723 );
and \U$7855 ( \9832 , RI9967528_213, \9725 );
and \U$7856 ( \9833 , RI890fa38_200, \9727 );
and \U$7857 ( \9834 , RI8918a20_187, \9729 );
and \U$7858 ( \9835 , RI8925248_174, \9731 );
and \U$7859 ( \9836 , RI8930c60_161, \9733 );
and \U$7860 ( \9837 , RI8939c48_148, \9735 );
and \U$7861 ( \9838 , RI8946470_135, \9737 );
and \U$7862 ( \9839 , RI89ec4d8_122, \9739 );
and \U$7863 ( \9840 , RI9776e18_109, \9741 );
and \U$7864 ( \9841 , RI9808318_96, \9743 );
and \U$7865 ( \9842 , RI9808930_83, \9745 );
and \U$7866 ( \9843 , RI98195c8_70, \9747 );
and \U$7867 ( \9844 , RI98abad0_57, \9749 );
and \U$7868 ( \9845 , RI98bc768_44, \9751 );
and \U$7869 ( \9846 , RI994dc68_31, \9753 );
or \U$7870 ( \9847 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 );
_DC g38b8 ( \9848_nG38b8 , \9847 , \9772 );
buf \U$7871 ( \9849 , \9848_nG38b8 );
not \U$7872 ( \9850 , \9849 );
and \U$7873 ( \9851 , \9829 , \9850 );
xor \U$7874 ( \9852 , \9697 , \9708 );
buf \U$7875 ( \9853 , \9852 );
buf \U$7876 ( \9854 , \9853 );
and \U$7877 ( \9855 , RI9959860_240, \9717 );
and \U$7878 ( \9856 , RI995e888_227, \9723 );
and \U$7879 ( \9857 , RI99674b0_214, \9725 );
and \U$7880 ( \9858 , RI890f9c0_201, \9727 );
and \U$7881 ( \9859 , RI89189a8_188, \9729 );
and \U$7882 ( \9860 , RI89251d0_175, \9731 );
and \U$7883 ( \9861 , RI8930be8_162, \9733 );
and \U$7884 ( \9862 , RI8939bd0_149, \9735 );
and \U$7885 ( \9863 , RI89463f8_136, \9737 );
and \U$7886 ( \9864 , RI89ec460_123, \9739 );
and \U$7887 ( \9865 , RI9776da0_110, \9741 );
and \U$7888 ( \9866 , RI98082a0_97, \9743 );
and \U$7889 ( \9867 , RI98088b8_84, \9745 );
and \U$7890 ( \9868 , RI9819550_71, \9747 );
and \U$7891 ( \9869 , RI98aba58_58, \9749 );
and \U$7892 ( \9870 , RI98bc6f0_45, \9751 );
and \U$7893 ( \9871 , RI994dbf0_32, \9753 );
or \U$7894 ( \9872 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 );
_DC g3743 ( \9873_nG3743 , \9872 , \9772 );
buf \U$7895 ( \9874 , \9873_nG3743 );
not \U$7896 ( \9875 , \9874 );
and \U$7897 ( \9876 , \9854 , \9875 );
xor \U$7898 ( \9877 , \9698 , \9707 );
buf \U$7899 ( \9878 , \9877 );
buf \U$7900 ( \9879 , \9878 );
and \U$7901 ( \9880 , RI994d998_241, \9717 );
and \U$7902 ( \9881 , RI995e810_228, \9723 );
and \U$7903 ( \9882 , RI9967438_215, \9725 );
and \U$7904 ( \9883 , RI890f948_202, \9727 );
and \U$7905 ( \9884 , RI8918930_189, \9729 );
and \U$7906 ( \9885 , RI8925158_176, \9731 );
and \U$7907 ( \9886 , RI8930b70_163, \9733 );
and \U$7908 ( \9887 , RI8939b58_150, \9735 );
and \U$7909 ( \9888 , RI8946380_137, \9737 );
and \U$7910 ( \9889 , RI89ec3e8_124, \9739 );
and \U$7911 ( \9890 , RI9776d28_111, \9741 );
and \U$7912 ( \9891 , RI9808228_98, \9743 );
and \U$7913 ( \9892 , RI9808840_85, \9745 );
and \U$7914 ( \9893 , RI98194d8_72, \9747 );
and \U$7915 ( \9894 , RI98ab9e0_59, \9749 );
and \U$7916 ( \9895 , RI98abff8_46, \9751 );
and \U$7917 ( \9896 , RI98bcc90_33, \9753 );
or \U$7918 ( \9897 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 );
_DC g371f ( \9898_nG371f , \9897 , \9772 );
buf \U$7919 ( \9899 , \9898_nG371f );
not \U$7920 ( \9900 , \9899 );
and \U$7921 ( \9901 , \9879 , \9900 );
xor \U$7922 ( \9902 , \9699 , \9706 );
buf \U$7923 ( \9903 , \9902 );
buf \U$7924 ( \9904 , \9903 );
and \U$7925 ( \9905 , RI994d920_242, \9717 );
and \U$7926 ( \9906 , RI995e798_229, \9723 );
and \U$7927 ( \9907 , RI99673c0_216, \9725 );
and \U$7928 ( \9908 , RI890f8d0_203, \9727 );
and \U$7929 ( \9909 , RI89188b8_190, \9729 );
and \U$7930 ( \9910 , RI89250e0_177, \9731 );
and \U$7931 ( \9911 , RI8930af8_164, \9733 );
and \U$7932 ( \9912 , RI8939ae0_151, \9735 );
and \U$7933 ( \9913 , RI8946308_138, \9737 );
and \U$7934 ( \9914 , RI89ec370_125, \9739 );
and \U$7935 ( \9915 , RI89ec988_112, \9741 );
and \U$7936 ( \9916 , RI97772c8_99, \9743 );
and \U$7937 ( \9917 , RI98087c8_86, \9745 );
and \U$7938 ( \9918 , RI9819460_73, \9747 );
and \U$7939 ( \9919 , RI98ab968_60, \9749 );
and \U$7940 ( \9920 , RI98abf80_47, \9751 );
and \U$7941 ( \9921 , RI98bcc18_34, \9753 );
or \U$7942 ( \9922 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 );
_DC g35e1 ( \9923_nG35e1 , \9922 , \9772 );
buf \U$7943 ( \9924 , \9923_nG35e1 );
not \U$7944 ( \9925 , \9924 );
and \U$7945 ( \9926 , \9904 , \9925 );
xor \U$7946 ( \9927 , \9700 , \9705 );
buf \U$7947 ( \9928 , \9927 );
buf \U$7948 ( \9929 , \9928 );
and \U$7949 ( \9930 , RI994d8a8_243, \9717 );
and \U$7950 ( \9931 , RI995e720_230, \9723 );
and \U$7951 ( \9932 , RI9967348_217, \9725 );
and \U$7952 ( \9933 , RI890f858_204, \9727 );
and \U$7953 ( \9934 , RI8918840_191, \9729 );
and \U$7954 ( \9935 , RI8925068_178, \9731 );
and \U$7955 ( \9936 , RI8930a80_165, \9733 );
and \U$7956 ( \9937 , RI8939a68_152, \9735 );
and \U$7957 ( \9938 , RI8946290_139, \9737 );
and \U$7958 ( \9939 , RI89ec2f8_126, \9739 );
and \U$7959 ( \9940 , RI89ec910_113, \9741 );
and \U$7960 ( \9941 , RI9777250_100, \9743 );
and \U$7961 ( \9942 , RI9808750_87, \9745 );
and \U$7962 ( \9943 , RI98193e8_74, \9747 );
and \U$7963 ( \9944 , RI98ab8f0_61, \9749 );
and \U$7964 ( \9945 , RI98abf08_48, \9751 );
and \U$7965 ( \9946 , RI98bcba0_35, \9753 );
or \U$7966 ( \9947 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 );
_DC g35bd ( \9948_nG35bd , \9947 , \9772 );
buf \U$7967 ( \9949 , \9948_nG35bd );
not \U$7968 ( \9950 , \9949 );
and \U$7969 ( \9951 , \9929 , \9950 );
xor \U$7970 ( \9952 , \9701 , \9704 );
buf \U$7971 ( \9953 , \9952 );
buf \U$7972 ( \9954 , \9953 );
and \U$7973 ( \9955 , RI994d830_244, \9717 );
and \U$7974 ( \9956 , RI995e6a8_231, \9723 );
and \U$7975 ( \9957 , RI99672d0_218, \9725 );
and \U$7976 ( \9958 , RI890f7e0_205, \9727 );
and \U$7977 ( \9959 , RI89187c8_192, \9729 );
and \U$7978 ( \9960 , RI8924ff0_179, \9731 );
and \U$7979 ( \9961 , RI8930a08_166, \9733 );
and \U$7980 ( \9962 , RI89399f0_153, \9735 );
and \U$7981 ( \9963 , RI8946218_140, \9737 );
and \U$7982 ( \9964 , RI89ec280_127, \9739 );
and \U$7983 ( \9965 , RI89ec898_114, \9741 );
and \U$7984 ( \9966 , RI97771d8_101, \9743 );
and \U$7985 ( \9967 , RI98086d8_88, \9745 );
and \U$7986 ( \9968 , RI9819370_75, \9747 );
and \U$7987 ( \9969 , RI98ab878_62, \9749 );
and \U$7988 ( \9970 , RI98abe90_49, \9751 );
and \U$7989 ( \9971 , RI98bcb28_36, \9753 );
or \U$7990 ( \9972 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 );
_DC g34b0 ( \9973_nG34b0 , \9972 , \9772 );
buf \U$7991 ( \9974 , \9973_nG34b0 );
not \U$7992 ( \9975 , \9974 );
and \U$7993 ( \9976 , \9954 , \9975 );
xor \U$7994 ( \9977 , \9702 , \9703 );
buf \U$7995 ( \9978 , \9977 );
buf \U$7996 ( \9979 , \9978 );
and \U$7997 ( \9980 , RI994d7b8_245, \9717 );
and \U$7998 ( \9981 , RI995e630_232, \9723 );
and \U$7999 ( \9982 , RI9967258_219, \9725 );
and \U$8000 ( \9983 , RI890f768_206, \9727 );
and \U$8001 ( \9984 , RI8918750_193, \9729 );
and \U$8002 ( \9985 , RI8924f78_180, \9731 );
and \U$8003 ( \9986 , RI8930990_167, \9733 );
and \U$8004 ( \9987 , RI8939978_154, \9735 );
and \U$8005 ( \9988 , RI89461a0_141, \9737 );
and \U$8006 ( \9989 , RI89ec208_128, \9739 );
and \U$8007 ( \9990 , RI89ec820_115, \9741 );
and \U$8008 ( \9991 , RI9777160_102, \9743 );
and \U$8009 ( \9992 , RI9808660_89, \9745 );
and \U$8010 ( \9993 , RI98192f8_76, \9747 );
and \U$8011 ( \9994 , RI98ab800_63, \9749 );
and \U$8012 ( \9995 , RI98abe18_50, \9751 );
and \U$8013 ( \9996 , RI98bcab0_37, \9753 );
or \U$8014 ( \9997 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 );
_DC g34c9 ( \9998_nG34c9 , \9997 , \9772 );
buf \U$8015 ( \9999 , \9998_nG34c9 );
not \U$8016 ( \10000 , \9999 );
and \U$8017 ( \10001 , \9979 , \10000 );
not \U$8018 ( \10002 , \9703 );
buf \U$8019 ( \10003 , \10002 );
buf \U$8020 ( \10004 , \10003 );
and \U$8021 ( \10005 , RI994d740_246, \9717 );
and \U$8022 ( \10006 , RI995e5b8_233, \9723 );
and \U$8023 ( \10007 , RI99671e0_220, \9725 );
and \U$8024 ( \10008 , RI890f6f0_207, \9727 );
and \U$8025 ( \10009 , RI89186d8_194, \9729 );
and \U$8026 ( \10010 , RI8924f00_181, \9731 );
and \U$8027 ( \10011 , RI8930918_168, \9733 );
and \U$8028 ( \10012 , RI8939900_155, \9735 );
and \U$8029 ( \10013 , RI8946128_142, \9737 );
and \U$8030 ( \10014 , RI89ec190_129, \9739 );
and \U$8031 ( \10015 , RI89ec7a8_116, \9741 );
and \U$8032 ( \10016 , RI97770e8_103, \9743 );
and \U$8033 ( \10017 , RI98085e8_90, \9745 );
and \U$8034 ( \10018 , RI9819280_77, \9747 );
and \U$8035 ( \10019 , RI98ab788_64, \9749 );
and \U$8036 ( \10020 , RI98abda0_51, \9751 );
and \U$8037 ( \10021 , RI98bca38_38, \9753 );
or \U$8038 ( \10022 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 );
_DC g3393 ( \10023_nG3393 , \10022 , \9772 );
buf \U$8039 ( \10024 , \10023_nG3393 );
not \U$8040 ( \10025 , \10024 );
and \U$8041 ( \10026 , \10004 , \10025 );
buf \U$8042 ( \10027 , RI994e4d8_13);
buf \U$8045 ( \10028 , \10027 );
and \U$8046 ( \10029 , RI994d6c8_247, \9717 );
and \U$8047 ( \10030 , RI995e540_234, \9723 );
and \U$8048 ( \10031 , RI9967168_221, \9725 );
and \U$8049 ( \10032 , RI890f678_208, \9727 );
and \U$8050 ( \10033 , RI8918660_195, \9729 );
and \U$8051 ( \10034 , RI8924e88_182, \9731 );
and \U$8052 ( \10035 , RI89308a0_169, \9733 );
and \U$8053 ( \10036 , RI8939888_156, \9735 );
and \U$8054 ( \10037 , RI89460b0_143, \9737 );
and \U$8055 ( \10038 , RI89ec118_130, \9739 );
and \U$8056 ( \10039 , RI89ec730_117, \9741 );
and \U$8057 ( \10040 , RI9777070_104, \9743 );
and \U$8058 ( \10041 , RI9808570_91, \9745 );
and \U$8059 ( \10042 , RI9819208_78, \9747 );
and \U$8060 ( \10043 , RI98ab710_65, \9749 );
and \U$8061 ( \10044 , RI98abd28_52, \9751 );
and \U$8062 ( \10045 , RI98bc9c0_39, \9753 );
or \U$8063 ( \10046 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 );
_DC g3377 ( \10047_nG3377 , \10046 , \9772 );
buf \U$8064 ( \10048 , \10047_nG3377 );
not \U$8065 ( \10049 , \10048 );
or \U$8066 ( \10050 , \10028 , \10049 );
and \U$8067 ( \10051 , \10025 , \10050 );
and \U$8068 ( \10052 , \10004 , \10050 );
or \U$8069 ( \10053 , \10026 , \10051 , \10052 );
and \U$8070 ( \10054 , \10000 , \10053 );
and \U$8071 ( \10055 , \9979 , \10053 );
or \U$8072 ( \10056 , \10001 , \10054 , \10055 );
and \U$8073 ( \10057 , \9975 , \10056 );
and \U$8074 ( \10058 , \9954 , \10056 );
or \U$8075 ( \10059 , \9976 , \10057 , \10058 );
and \U$8076 ( \10060 , \9950 , \10059 );
and \U$8077 ( \10061 , \9929 , \10059 );
or \U$8078 ( \10062 , \9951 , \10060 , \10061 );
and \U$8079 ( \10063 , \9925 , \10062 );
and \U$8080 ( \10064 , \9904 , \10062 );
or \U$8081 ( \10065 , \9926 , \10063 , \10064 );
and \U$8082 ( \10066 , \9900 , \10065 );
and \U$8083 ( \10067 , \9879 , \10065 );
or \U$8084 ( \10068 , \9901 , \10066 , \10067 );
and \U$8085 ( \10069 , \9875 , \10068 );
and \U$8086 ( \10070 , \9854 , \10068 );
or \U$8087 ( \10071 , \9876 , \10069 , \10070 );
and \U$8088 ( \10072 , \9850 , \10071 );
and \U$8089 ( \10073 , \9829 , \10071 );
or \U$8090 ( \10074 , \9851 , \10072 , \10073 );
and \U$8091 ( \10075 , \9825 , \10074 );
and \U$8092 ( \10076 , \9804 , \10074 );
or \U$8093 ( \10077 , \9826 , \10075 , \10076 );
and \U$8094 ( \10078 , \9800 , \10077 );
and \U$8095 ( \10079 , \9779 , \10077 );
or \U$8096 ( \10080 , \9801 , \10078 , \10079 );
xor \U$8097 ( \10081 , \9776 , \10080 );
buf g3a90_GF_PartitionCandidate( \10082_nG3a90 , \10081 );
buf \U$8098 ( \10083 , \10082_nG3a90 );
xor \U$8099 ( \10084 , \9779 , \9800 );
xor \U$8100 ( \10085 , \10084 , \10077 );
buf g3a6c_GF_PartitionCandidate( \10086_nG3a6c , \10085 );
buf \U$8101 ( \10087 , \10086_nG3a6c );
xor \U$8102 ( \10088 , \9804 , \9825 );
xor \U$8103 ( \10089 , \10088 , \10074 );
buf g38e5_GF_PartitionCandidate( \10090_nG38e5 , \10089 );
buf \U$8104 ( \10091 , \10090_nG38e5 );
and \U$8105 ( \10092 , \10087 , \10091 );
not \U$8106 ( \10093 , \10092 );
and \U$8107 ( \10094 , \10083 , \10093 );
not \U$8108 ( \10095 , \10094 );
buf \U$8109 ( \10096 , RI9921d48_600);
buf \U$8110 ( \10097 , RI9921fa0_595);
buf \U$8111 ( \10098 , RI9922018_594);
buf \U$8112 ( \10099 , RI9922090_593);
buf \U$8113 ( \10100 , RI9922108_592);
buf \U$8114 ( \10101 , RI9922180_591);
buf \U$8115 ( \10102 , RI99221f8_590);
buf \U$8116 ( \10103 , RI9922270_589);
buf \U$8117 ( \10104 , RI99222e8_588);
buf \U$8118 ( \10105 , RI9921f28_596);
nor \U$8119 ( \10106 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 );
buf \U$8120 ( \10107 , \10106 );
buf \U$8121 ( \10108 , \10107 );
xor \U$8122 ( \10109 , \10096 , \10108 );
buf \U$8123 ( \10110 , \10109 );
buf \U$8124 ( \10111 , RI9921dc0_599);
and \U$8125 ( \10112 , \10096 , \10108 );
xor \U$8126 ( \10113 , \10111 , \10112 );
buf \U$8127 ( \10114 , \10113 );
buf \U$8128 ( \10115 , RI9921e38_598);
and \U$8129 ( \10116 , \10111 , \10112 );
xor \U$8130 ( \10117 , \10115 , \10116 );
buf \U$8131 ( \10118 , \10117 );
buf \U$8132 ( \10119 , RI9921eb0_597);
and \U$8133 ( \10120 , \10115 , \10116 );
xor \U$8134 ( \10121 , \10119 , \10120 );
buf \U$8135 ( \10122 , \10121 );
buf \U$8136 ( \10123 , RI9921f28_596);
and \U$8137 ( \10124 , \10119 , \10120 );
xor \U$8138 ( \10125 , \10123 , \10124 );
buf \U$8139 ( \10126 , \10125 );
not \U$8140 ( \10127 , \10126 );
buf \U$8141 ( \10128 , RI9921fa0_595);
and \U$8142 ( \10129 , \10123 , \10124 );
xor \U$8143 ( \10130 , \10128 , \10129 );
buf \U$8144 ( \10131 , \10130 );
buf \U$8145 ( \10132 , RI9922018_594);
and \U$8146 ( \10133 , \10128 , \10129 );
xor \U$8147 ( \10134 , \10132 , \10133 );
buf \U$8148 ( \10135 , \10134 );
buf \U$8149 ( \10136 , RI9922090_593);
and \U$8150 ( \10137 , \10132 , \10133 );
xor \U$8151 ( \10138 , \10136 , \10137 );
buf \U$8152 ( \10139 , \10138 );
buf \U$8153 ( \10140 , RI9922108_592);
and \U$8154 ( \10141 , \10136 , \10137 );
xor \U$8155 ( \10142 , \10140 , \10141 );
buf \U$8156 ( \10143 , \10142 );
buf \U$8157 ( \10144 , RI9922180_591);
and \U$8158 ( \10145 , \10140 , \10141 );
xor \U$8159 ( \10146 , \10144 , \10145 );
buf \U$8160 ( \10147 , \10146 );
buf \U$8161 ( \10148 , RI99221f8_590);
and \U$8162 ( \10149 , \10144 , \10145 );
xor \U$8163 ( \10150 , \10148 , \10149 );
buf \U$8164 ( \10151 , \10150 );
buf \U$8165 ( \10152 , RI9922270_589);
and \U$8166 ( \10153 , \10148 , \10149 );
xor \U$8167 ( \10154 , \10152 , \10153 );
buf \U$8168 ( \10155 , \10154 );
buf \U$8169 ( \10156 , RI99222e8_588);
and \U$8170 ( \10157 , \10152 , \10153 );
xor \U$8171 ( \10158 , \10156 , \10157 );
buf \U$8172 ( \10159 , \10158 );
nor \U$8173 ( \10160 , \10110 , \10114 , \10118 , \10122 , \10127 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8174 ( \10161 , RI9922bd0_569, \10160 );
not \U$8175 ( \10162 , \10110 );
not \U$8176 ( \10163 , \10114 );
not \U$8177 ( \10164 , \10118 );
not \U$8178 ( \10165 , \10122 );
nor \U$8179 ( \10166 , \10162 , \10163 , \10164 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8180 ( \10167 , RI9923800_549, \10166 );
nor \U$8181 ( \10168 , \10110 , \10163 , \10164 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8182 ( \10169 , RI9924160_529, \10168 );
nor \U$8183 ( \10170 , \10162 , \10114 , \10164 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8184 ( \10171 , RI9924ac0_509, \10170 );
nor \U$8185 ( \10172 , \10110 , \10114 , \10164 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8186 ( \10173 , RI9925ab0_489, \10172 );
nor \U$8187 ( \10174 , \10162 , \10163 , \10118 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8188 ( \10175 , RI9926410_469, \10174 );
nor \U$8189 ( \10176 , \10110 , \10163 , \10118 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8190 ( \10177 , RI9926d70_449, \10176 );
nor \U$8191 ( \10178 , \10162 , \10114 , \10118 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8192 ( \10179 , RI9928120_429, \10178 );
nor \U$8193 ( \10180 , \10110 , \10114 , \10118 , \10165 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8194 ( \10181 , RI9928a80_409, \10180 );
nor \U$8195 ( \10182 , \10162 , \10163 , \10164 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8196 ( \10183 , RI992a1f0_389, \10182 );
nor \U$8197 ( \10184 , \10110 , \10163 , \10164 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8198 ( \10185 , RI992ab50_369, \10184 );
nor \U$8199 ( \10186 , \10162 , \10114 , \10164 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8200 ( \10187 , RI992b4b0_349, \10186 );
nor \U$8201 ( \10188 , \10110 , \10114 , \10164 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8202 ( \10189 , RI992cfe0_329, \10188 );
nor \U$8203 ( \10190 , \10162 , \10163 , \10118 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8204 ( \10191 , RI992eed0_309, \10190 );
nor \U$8205 ( \10192 , \10110 , \10163 , \10118 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8206 ( \10193 , RI992f830_289, \10192 );
nor \U$8207 ( \10194 , \10162 , \10114 , \10118 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8208 ( \10195 , RI9931ae0_269, \10194 );
nor \U$8209 ( \10196 , \10110 , \10114 , \10118 , \10122 , \10126 , \10131 , \10135 , \10139 , \10143 , \10147 , \10151 , \10155 , \10159 );
and \U$8210 ( \10197 , RI994d5d8_249, \10196 );
or \U$8211 ( \10198 , \10161 , \10167 , \10169 , \10171 , \10173 , \10175 , \10177 , \10179 , \10181 , \10183 , \10185 , \10187 , \10189 , \10191 , \10193 , \10195 , \10197 );
buf \U$8212 ( \10199 , \10131 );
buf \U$8213 ( \10200 , \10135 );
buf \U$8214 ( \10201 , \10139 );
buf \U$8215 ( \10202 , \10143 );
buf \U$8216 ( \10203 , \10147 );
buf \U$8217 ( \10204 , \10151 );
buf \U$8218 ( \10205 , \10155 );
buf \U$8219 ( \10206 , \10159 );
buf \U$8220 ( \10207 , \10126 );
buf \U$8221 ( \10208 , \10110 );
buf \U$8222 ( \10209 , \10114 );
buf \U$8223 ( \10210 , \10118 );
buf \U$8224 ( \10211 , \10122 );
or \U$8225 ( \10212 , \10208 , \10209 , \10210 , \10211 );
and \U$8226 ( \10213 , \10207 , \10212 );
or \U$8227 ( \10214 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10213 );
buf \U$8228 ( \10215 , \10214 );
_DC g4187 ( \10216_nG4187 , \10198 , \10215 );
buf \U$8229 ( \10217 , \10216_nG4187 );
buf \U$8230 ( \10218 , RI995f0f8_1);
and \U$8231 ( \10219 , \9693 , \9712 );
and \U$8232 ( \10220 , \10218 , \10219 );
buf \U$8233 ( \10221 , \10220 );
buf \U$8234 ( \10222 , \10221 );
xor \U$8235 ( \10223 , \10218 , \10219 );
buf \U$8236 ( \10224 , \10223 );
buf \U$8237 ( \10225 , \10224 );
and \U$8238 ( \10226 , RI995e4c8_235, \9717 );
and \U$8239 ( \10227 , RI99670f0_222, \9723 );
and \U$8240 ( \10228 , RI890f600_209, \9725 );
and \U$8241 ( \10229 , RI89185e8_196, \9727 );
and \U$8242 ( \10230 , RI8924e10_183, \9729 );
and \U$8243 ( \10231 , RI8930828_170, \9731 );
and \U$8244 ( \10232 , RI8939810_157, \9733 );
and \U$8245 ( \10233 , RI8946038_144, \9735 );
and \U$8246 ( \10234 , RI89ec0a0_131, \9737 );
and \U$8247 ( \10235 , RI89ec6b8_118, \9739 );
and \U$8248 ( \10236 , RI9776ff8_105, \9741 );
and \U$8249 ( \10237 , RI98084f8_92, \9743 );
and \U$8250 ( \10238 , RI9808b10_79, \9745 );
and \U$8251 ( \10239 , RI98197a8_66, \9747 );
and \U$8252 ( \10240 , RI98abcb0_53, \9749 );
and \U$8253 ( \10241 , RI98bc948_40, \9751 );
and \U$8254 ( \10242 , RI994de48_27, \9753 );
or \U$8255 ( \10243 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 );
_DC g3c4f ( \10244_nG3c4f , \10243 , \9772 );
buf \U$8256 ( \10245 , \10244_nG3c4f );
not \U$8257 ( \10246 , \10245 );
and \U$8258 ( \10247 , \10225 , \10246 );
and \U$8259 ( \10248 , \9715 , \9775 );
and \U$8260 ( \10249 , \9775 , \10080 );
and \U$8261 ( \10250 , \9715 , \10080 );
or \U$8262 ( \10251 , \10248 , \10249 , \10250 );
and \U$8263 ( \10252 , \10246 , \10251 );
and \U$8264 ( \10253 , \10225 , \10251 );
or \U$8265 ( \10254 , \10247 , \10252 , \10253 );
xnor \U$8266 ( \10255 , \10222 , \10254 );
buf g3c64_GF_PartitionCandidate( \10256_nG3c64 , \10255 );
buf \U$8267 ( \10257 , \10256_nG3c64 );
xor \U$8268 ( \10258 , \10225 , \10246 );
xor \U$8269 ( \10259 , \10258 , \10251 );
buf g3c58_GF_PartitionCandidate( \10260_nG3c58 , \10259 );
buf \U$8270 ( \10261 , \10260_nG3c58 );
xor \U$8271 ( \10262 , \10257 , \10261 );
xor \U$8272 ( \10263 , \10261 , \10083 );
not \U$8273 ( \10264 , \10263 );
and \U$8274 ( \10265 , \10262 , \10264 );
and \U$8275 ( \10266 , \10217 , \10265 );
and \U$8276 ( \10267 , RI9922f18_568, \10160 );
and \U$8277 ( \10268 , RI9923878_548, \10166 );
and \U$8278 ( \10269 , RI99241d8_528, \10168 );
and \U$8279 ( \10270 , RI9924b38_508, \10170 );
and \U$8280 ( \10271 , RI9925b28_488, \10172 );
and \U$8281 ( \10272 , RI9926488_468, \10174 );
and \U$8282 ( \10273 , RI9926de8_448, \10176 );
and \U$8283 ( \10274 , RI9928198_428, \10178 );
and \U$8284 ( \10275 , RI9928af8_408, \10180 );
and \U$8285 ( \10276 , RI992a268_388, \10182 );
and \U$8286 ( \10277 , RI992abc8_368, \10184 );
and \U$8287 ( \10278 , RI992c6f8_348, \10186 );
and \U$8288 ( \10279 , RI992d058_328, \10188 );
and \U$8289 ( \10280 , RI992ef48_308, \10190 );
and \U$8290 ( \10281 , RI992f8a8_288, \10192 );
and \U$8291 ( \10282 , RI9931b58_268, \10194 );
and \U$8292 ( \10283 , RI994d650_248, \10196 );
or \U$8293 ( \10284 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 );
_DC g427b ( \10285_nG427b , \10284 , \10215 );
buf \U$8294 ( \10286 , \10285_nG427b );
and \U$8295 ( \10287 , \10286 , \10263 );
nor \U$8296 ( \10288 , \10266 , \10287 );
and \U$8297 ( \10289 , \10261 , \10083 );
not \U$8298 ( \10290 , \10289 );
and \U$8299 ( \10291 , \10257 , \10290 );
xnor \U$8300 ( \10292 , \10288 , \10291 );
xor \U$8301 ( \10293 , \10095 , \10292 );
and \U$8303 ( \10294 , RI9922b58_570, \10160 );
and \U$8304 ( \10295 , RI9923788_550, \10166 );
and \U$8305 ( \10296 , RI99240e8_530, \10168 );
and \U$8306 ( \10297 , RI9924a48_510, \10170 );
and \U$8307 ( \10298 , RI9925a38_490, \10172 );
and \U$8308 ( \10299 , RI9926398_470, \10174 );
and \U$8309 ( \10300 , RI9926cf8_450, \10176 );
and \U$8310 ( \10301 , RI99280a8_430, \10178 );
and \U$8311 ( \10302 , RI9928a08_410, \10180 );
and \U$8312 ( \10303 , RI992a178_390, \10182 );
and \U$8313 ( \10304 , RI992aad8_370, \10184 );
and \U$8314 ( \10305 , RI992b438_350, \10186 );
and \U$8315 ( \10306 , RI992cf68_330, \10188 );
and \U$8316 ( \10307 , RI992ee58_310, \10190 );
and \U$8317 ( \10308 , RI992f7b8_290, \10192 );
and \U$8318 ( \10309 , RI9931a68_270, \10194 );
and \U$8319 ( \10310 , RI994d560_250, \10196 );
or \U$8320 ( \10311 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 );
_DC g40c5 ( \10312_nG40c5 , \10311 , \10215 );
buf \U$8321 ( \10313 , \10312_nG40c5 );
or \U$8322 ( \10314 , \10222 , \10254 );
not \U$8323 ( \10315 , \10314 );
buf g3e60_GF_PartitionCandidate( \10316_nG3e60 , \10315 );
buf \U$8324 ( \10317 , \10316_nG3e60 );
xor \U$8325 ( \10318 , \10317 , \10257 );
and \U$8326 ( \10319 , \10313 , \10318 );
nor \U$8327 ( \10320 , 1'b0 , \10319 );
xnor \U$8329 ( \10321 , \10320 , 1'b0 );
xor \U$8330 ( \10322 , \10293 , \10321 );
xor \U$8331 ( \10323 , 1'b0 , \10322 );
xor \U$8333 ( \10324 , \10083 , \10087 );
xor \U$8334 ( \10325 , \10087 , \10091 );
not \U$8335 ( \10326 , \10325 );
and \U$8336 ( \10327 , \10324 , \10326 );
and \U$8337 ( \10328 , \10286 , \10327 );
not \U$8338 ( \10329 , \10328 );
xnor \U$8339 ( \10330 , \10329 , \10094 );
and \U$8340 ( \10331 , \10313 , \10265 );
and \U$8341 ( \10332 , \10217 , \10263 );
nor \U$8342 ( \10333 , \10331 , \10332 );
xnor \U$8343 ( \10334 , \10333 , \10291 );
and \U$8344 ( \10335 , \10330 , \10334 );
or \U$8346 ( \10336 , 1'b0 , \10335 , 1'b0 );
xor \U$8348 ( \10337 , \10336 , 1'b0 );
xor \U$8350 ( \10338 , \10337 , 1'b0 );
and \U$8351 ( \10339 , \10323 , \10338 );
or \U$8352 ( \10340 , 1'b0 , 1'b0 , \10339 );
and \U$8355 ( \10341 , \10286 , \10265 );
not \U$8356 ( \10342 , \10341 );
xnor \U$8357 ( \10343 , \10342 , \10291 );
xor \U$8358 ( \10344 , 1'b0 , \10343 );
and \U$8360 ( \10345 , \10217 , \10318 );
nor \U$8361 ( \10346 , 1'b0 , \10345 );
xnor \U$8362 ( \10347 , \10346 , 1'b0 );
xor \U$8363 ( \10348 , \10344 , \10347 );
xor \U$8364 ( \10349 , 1'b0 , \10348 );
xor \U$8366 ( \10350 , \10349 , 1'b1 );
and \U$8367 ( \10351 , \10095 , \10292 );
and \U$8368 ( \10352 , \10292 , \10321 );
and \U$8369 ( \10353 , \10095 , \10321 );
or \U$8370 ( \10354 , \10351 , \10352 , \10353 );
xor \U$8372 ( \10355 , \10354 , 1'b0 );
xor \U$8374 ( \10356 , \10355 , 1'b0 );
xor \U$8375 ( \10357 , \10350 , \10356 );
and \U$8376 ( \10358 , \10340 , \10357 );
or \U$8378 ( \10359 , 1'b0 , \10358 , 1'b0 );
xor \U$8380 ( \10360 , \10359 , 1'b0 );
and \U$8382 ( \10361 , \10349 , 1'b1 );
and \U$8383 ( \10362 , 1'b1 , \10356 );
and \U$8384 ( \10363 , \10349 , \10356 );
or \U$8385 ( \10364 , \10361 , \10362 , \10363 );
xor \U$8386 ( \10365 , 1'b0 , \10364 );
not \U$8388 ( \10366 , \10291 );
and \U$8390 ( \10367 , \10286 , \10318 );
nor \U$8391 ( \10368 , 1'b0 , \10367 );
xnor \U$8392 ( \10369 , \10368 , 1'b0 );
xor \U$8393 ( \10370 , \10366 , \10369 );
xor \U$8395 ( \10371 , \10370 , 1'b0 );
xor \U$8396 ( \10372 , 1'b0 , \10371 );
xor \U$8398 ( \10373 , \10372 , 1'b0 );
and \U$8400 ( \10374 , \10343 , \10347 );
or \U$8402 ( \10375 , 1'b0 , \10374 , 1'b0 );
xor \U$8404 ( \10376 , \10375 , 1'b0 );
xor \U$8406 ( \10377 , \10376 , 1'b0 );
xor \U$8407 ( \10378 , \10373 , \10377 );
xor \U$8408 ( \10379 , \10365 , \10378 );
xor \U$8409 ( \10380 , \10360 , \10379 );
xor \U$8415 ( \10381 , \9829 , \9850 );
xor \U$8416 ( \10382 , \10381 , \10071 );
buf g38c1_GF_PartitionCandidate( \10383_nG38c1 , \10382 );
buf \U$8417 ( \10384 , \10383_nG38c1 );
xor \U$8418 ( \10385 , \10091 , \10384 );
xor \U$8419 ( \10386 , \9854 , \9875 );
xor \U$8420 ( \10387 , \10386 , \10068 );
buf g374c_GF_PartitionCandidate( \10388_nG374c , \10387 );
buf \U$8421 ( \10389 , \10388_nG374c );
xor \U$8422 ( \10390 , \10384 , \10389 );
not \U$8423 ( \10391 , \10390 );
and \U$8424 ( \10392 , \10385 , \10391 );
and \U$8425 ( \10393 , \10286 , \10392 );
not \U$8426 ( \10394 , \10393 );
and \U$8427 ( \10395 , \10384 , \10389 );
not \U$8428 ( \10396 , \10395 );
and \U$8429 ( \10397 , \10091 , \10396 );
xnor \U$8430 ( \10398 , \10394 , \10397 );
and \U$8431 ( \10399 , \10313 , \10327 );
and \U$8432 ( \10400 , \10217 , \10325 );
nor \U$8433 ( \10401 , \10399 , \10400 );
xnor \U$8434 ( \10402 , \10401 , \10094 );
and \U$8435 ( \10403 , \10398 , \10402 );
or \U$8437 ( \10404 , 1'b0 , \10403 , 1'b0 );
and \U$8438 ( \10405 , RI9922a68_572, \10160 );
and \U$8439 ( \10406 , RI9923698_552, \10166 );
and \U$8440 ( \10407 , RI9923ff8_532, \10168 );
and \U$8441 ( \10408 , RI9924958_512, \10170 );
and \U$8442 ( \10409 , RI9925948_492, \10172 );
and \U$8443 ( \10410 , RI99262a8_472, \10174 );
and \U$8444 ( \10411 , RI9926c08_452, \10176 );
and \U$8445 ( \10412 , RI9927fb8_432, \10178 );
and \U$8446 ( \10413 , RI9928918_412, \10180 );
and \U$8447 ( \10414 , RI9929278_392, \10182 );
and \U$8448 ( \10415 , RI992a9e8_372, \10184 );
and \U$8449 ( \10416 , RI992b348_352, \10186 );
and \U$8450 ( \10417 , RI992ce78_332, \10188 );
and \U$8451 ( \10418 , RI992ed68_312, \10190 );
and \U$8452 ( \10419 , RI992f6c8_292, \10192 );
and \U$8453 ( \10420 , RI9931978_272, \10194 );
and \U$8454 ( \10421 , RI994d470_252, \10196 );
or \U$8455 ( \10422 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 );
_DC g3f2a ( \10423_nG3f2a , \10422 , \10215 );
buf \U$8456 ( \10424 , \10423_nG3f2a );
and \U$8457 ( \10425 , \10424 , \10265 );
and \U$8458 ( \10426 , RI9922ae0_571, \10160 );
and \U$8459 ( \10427 , RI9923710_551, \10166 );
and \U$8460 ( \10428 , RI9924070_531, \10168 );
and \U$8461 ( \10429 , RI99249d0_511, \10170 );
and \U$8462 ( \10430 , RI99259c0_491, \10172 );
and \U$8463 ( \10431 , RI9926320_471, \10174 );
and \U$8464 ( \10432 , RI9926c80_451, \10176 );
and \U$8465 ( \10433 , RI9928030_431, \10178 );
and \U$8466 ( \10434 , RI9928990_411, \10180 );
and \U$8467 ( \10435 , RI992a100_391, \10182 );
and \U$8468 ( \10436 , RI992aa60_371, \10184 );
and \U$8469 ( \10437 , RI992b3c0_351, \10186 );
and \U$8470 ( \10438 , RI992cef0_331, \10188 );
and \U$8471 ( \10439 , RI992ede0_311, \10190 );
and \U$8472 ( \10440 , RI992f740_291, \10192 );
and \U$8473 ( \10441 , RI99319f0_271, \10194 );
and \U$8474 ( \10442 , RI994d4e8_251, \10196 );
or \U$8475 ( \10443 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 );
_DC g4004 ( \10444_nG4004 , \10443 , \10215 );
buf \U$8476 ( \10445 , \10444_nG4004 );
and \U$8477 ( \10446 , \10445 , \10263 );
nor \U$8478 ( \10447 , \10425 , \10446 );
xnor \U$8479 ( \10448 , \10447 , \10291 );
and \U$8481 ( \10449 , RI99229f0_573, \10160 );
and \U$8482 ( \10450 , RI9923620_553, \10166 );
and \U$8483 ( \10451 , RI9923f80_533, \10168 );
and \U$8484 ( \10452 , RI99248e0_513, \10170 );
and \U$8485 ( \10453 , RI99258d0_493, \10172 );
and \U$8486 ( \10454 , RI9926230_473, \10174 );
and \U$8487 ( \10455 , RI9926b90_453, \10176 );
and \U$8488 ( \10456 , RI9927f40_433, \10178 );
and \U$8489 ( \10457 , RI99288a0_413, \10180 );
and \U$8490 ( \10458 , RI9929200_393, \10182 );
and \U$8491 ( \10459 , RI992a970_373, \10184 );
and \U$8492 ( \10460 , RI992b2d0_353, \10186 );
and \U$8493 ( \10461 , RI992ce00_333, \10188 );
and \U$8494 ( \10462 , RI992ecf0_313, \10190 );
and \U$8495 ( \10463 , RI992f650_293, \10192 );
and \U$8496 ( \10464 , RI9931900_273, \10194 );
and \U$8497 ( \10465 , RI994d3f8_253, \10196 );
or \U$8498 ( \10466 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 );
_DC g3e3f ( \10467_nG3e3f , \10466 , \10215 );
buf \U$8499 ( \10468 , \10467_nG3e3f );
and \U$8500 ( \10469 , \10468 , \10318 );
nor \U$8501 ( \10470 , 1'b0 , \10469 );
xnor \U$8502 ( \10471 , \10470 , 1'b0 );
and \U$8503 ( \10472 , \10448 , \10471 );
or \U$8506 ( \10473 , \10472 , 1'b0 , 1'b0 );
and \U$8507 ( \10474 , \10404 , \10473 );
or \U$8510 ( \10475 , \10474 , 1'b0 , 1'b0 );
and \U$8513 ( \10476 , \10424 , \10318 );
nor \U$8514 ( \10477 , 1'b0 , \10476 );
xnor \U$8515 ( \10478 , \10477 , 1'b0 );
xor \U$8517 ( \10479 , \10478 , 1'b0 );
xor \U$8519 ( \10480 , \10479 , 1'b0 );
not \U$8520 ( \10481 , \10397 );
and \U$8521 ( \10482 , \10217 , \10327 );
and \U$8522 ( \10483 , \10286 , \10325 );
nor \U$8523 ( \10484 , \10482 , \10483 );
xnor \U$8524 ( \10485 , \10484 , \10094 );
xor \U$8525 ( \10486 , \10481 , \10485 );
and \U$8526 ( \10487 , \10445 , \10265 );
and \U$8527 ( \10488 , \10313 , \10263 );
nor \U$8528 ( \10489 , \10487 , \10488 );
xnor \U$8529 ( \10490 , \10489 , \10291 );
xor \U$8530 ( \10491 , \10486 , \10490 );
and \U$8531 ( \10492 , \10480 , \10491 );
or \U$8533 ( \10493 , 1'b0 , \10492 , 1'b0 );
and \U$8534 ( \10494 , \10475 , \10493 );
or \U$8535 ( \10495 , 1'b0 , 1'b0 , \10494 );
and \U$8537 ( \10496 , \10445 , \10318 );
nor \U$8538 ( \10497 , 1'b0 , \10496 );
xnor \U$8539 ( \10498 , \10497 , 1'b0 );
xor \U$8541 ( \10499 , \10498 , 1'b0 );
xor \U$8543 ( \10500 , \10499 , 1'b0 );
xor \U$8545 ( \10501 , 1'b0 , \10330 );
xor \U$8546 ( \10502 , \10501 , \10334 );
xor \U$8547 ( \10503 , \10500 , \10502 );
and \U$8549 ( \10504 , \10503 , 1'b1 );
and \U$8550 ( \10505 , \10481 , \10485 );
and \U$8551 ( \10506 , \10485 , \10490 );
and \U$8552 ( \10507 , \10481 , \10490 );
or \U$8553 ( \10508 , \10505 , \10506 , \10507 );
xor \U$8555 ( \10509 , \10508 , 1'b0 );
xor \U$8557 ( \10510 , \10509 , 1'b0 );
and \U$8558 ( \10511 , 1'b1 , \10510 );
and \U$8559 ( \10512 , \10503 , \10510 );
or \U$8560 ( \10513 , \10504 , \10511 , \10512 );
and \U$8561 ( \10514 , \10495 , \10513 );
xor \U$8563 ( \10515 , \10323 , 1'b0 );
xor \U$8564 ( \10516 , \10515 , \10338 );
and \U$8565 ( \10517 , \10513 , \10516 );
and \U$8566 ( \10518 , \10495 , \10516 );
or \U$8567 ( \10519 , \10514 , \10517 , \10518 );
xor \U$8569 ( \10520 , 1'b0 , \10340 );
xor \U$8570 ( \10521 , \10520 , \10357 );
and \U$8571 ( \10522 , \10519 , \10521 );
or \U$8572 ( \10523 , 1'b0 , 1'b0 , \10522 );
nand \U$8573 ( \10524 , \10380 , \10523 );
nor \U$8574 ( \10525 , \10380 , \10523 );
not \U$8575 ( \10526 , \10525 );
nand \U$8576 ( \10527 , \10524 , \10526 );
xor \U$8577 ( \10528 , \10004 , \10025 );
xor \U$8578 ( \10529 , \10528 , \10050 );
buf g339a_GF_PartitionCandidate( \10530_nG339a , \10529 );
buf \U$8579 ( \10531 , \10530_nG339a );
xor \U$8580 ( \10532 , \10028 , \10048 );
buf g337a_GF_PartitionCandidate( \10533_nG337a , \10532 );
buf \U$8581 ( \10534 , \10533_nG337a );
xor \U$8582 ( \10535 , \10531 , \10534 );
not \U$8583 ( \10536 , \10534 );
and \U$8584 ( \10537 , \10535 , \10536 );
and \U$8585 ( \10538 , \10468 , \10537 );
and \U$8586 ( \10539 , \10424 , \10534 );
nor \U$8587 ( \10540 , \10538 , \10539 );
xnor \U$8588 ( \10541 , \10540 , \10531 );
and \U$8589 ( \10542 , RI9922900_575, \10160 );
and \U$8590 ( \10543 , RI9923530_555, \10166 );
and \U$8591 ( \10544 , RI9923e90_535, \10168 );
and \U$8592 ( \10545 , RI99247f0_515, \10170 );
and \U$8593 ( \10546 , RI99257e0_495, \10172 );
and \U$8594 ( \10547 , RI9926140_475, \10174 );
and \U$8595 ( \10548 , RI9926aa0_455, \10176 );
and \U$8596 ( \10549 , RI9927e50_435, \10178 );
and \U$8597 ( \10550 , RI99287b0_415, \10180 );
and \U$8598 ( \10551 , RI9929110_395, \10182 );
and \U$8599 ( \10552 , RI992a880_375, \10184 );
and \U$8600 ( \10553 , RI992b1e0_355, \10186 );
and \U$8601 ( \10554 , RI992cd10_335, \10188 );
and \U$8602 ( \10555 , RI992d670_315, \10190 );
and \U$8603 ( \10556 , RI992f560_295, \10192 );
and \U$8604 ( \10557 , RI9931810_275, \10194 );
and \U$8605 ( \10558 , RI9935f50_255, \10196 );
or \U$8606 ( \10559 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 );
_DC g3c8c ( \10560_nG3c8c , \10559 , \10215 );
buf \U$8607 ( \10561 , \10560_nG3c8c );
xor \U$8608 ( \10562 , \9954 , \9975 );
xor \U$8609 ( \10563 , \10562 , \10056 );
buf g34d5_GF_PartitionCandidate( \10564_nG34d5 , \10563 );
buf \U$8610 ( \10565 , \10564_nG34d5 );
xor \U$8611 ( \10566 , \9979 , \10000 );
xor \U$8612 ( \10567 , \10566 , \10053 );
buf g34d9_GF_PartitionCandidate( \10568_nG34d9 , \10567 );
buf \U$8613 ( \10569 , \10568_nG34d9 );
xor \U$8614 ( \10570 , \10565 , \10569 );
xor \U$8615 ( \10571 , \10569 , \10531 );
not \U$8616 ( \10572 , \10571 );
and \U$8617 ( \10573 , \10570 , \10572 );
and \U$8618 ( \10574 , \10561 , \10573 );
and \U$8619 ( \10575 , RI9922978_574, \10160 );
and \U$8620 ( \10576 , RI99235a8_554, \10166 );
and \U$8621 ( \10577 , RI9923f08_534, \10168 );
and \U$8622 ( \10578 , RI9924868_514, \10170 );
and \U$8623 ( \10579 , RI9925858_494, \10172 );
and \U$8624 ( \10580 , RI99261b8_474, \10174 );
and \U$8625 ( \10581 , RI9926b18_454, \10176 );
and \U$8626 ( \10582 , RI9927ec8_434, \10178 );
and \U$8627 ( \10583 , RI9928828_414, \10180 );
and \U$8628 ( \10584 , RI9929188_394, \10182 );
and \U$8629 ( \10585 , RI992a8f8_374, \10184 );
and \U$8630 ( \10586 , RI992b258_354, \10186 );
and \U$8631 ( \10587 , RI992cd88_334, \10188 );
and \U$8632 ( \10588 , RI992d6e8_314, \10190 );
and \U$8633 ( \10589 , RI992f5d8_294, \10192 );
and \U$8634 ( \10590 , RI9931888_274, \10194 );
and \U$8635 ( \10591 , RI9935fc8_254, \10196 );
or \U$8636 ( \10592 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 );
_DC g3d60 ( \10593_nG3d60 , \10592 , \10215 );
buf \U$8637 ( \10594 , \10593_nG3d60 );
and \U$8638 ( \10595 , \10594 , \10571 );
nor \U$8639 ( \10596 , \10574 , \10595 );
and \U$8640 ( \10597 , \10569 , \10531 );
not \U$8641 ( \10598 , \10597 );
and \U$8642 ( \10599 , \10565 , \10598 );
xnor \U$8643 ( \10600 , \10596 , \10599 );
and \U$8644 ( \10601 , \10541 , \10600 );
and \U$8645 ( \10602 , RI9922810_577, \10160 );
and \U$8646 ( \10603 , RI9923440_557, \10166 );
and \U$8647 ( \10604 , RI9923da0_537, \10168 );
and \U$8648 ( \10605 , RI9924700_517, \10170 );
and \U$8649 ( \10606 , RI99256f0_497, \10172 );
and \U$8650 ( \10607 , RI9926050_477, \10174 );
and \U$8651 ( \10608 , RI99269b0_457, \10176 );
and \U$8652 ( \10609 , RI9927d60_437, \10178 );
and \U$8653 ( \10610 , RI99286c0_417, \10180 );
and \U$8654 ( \10611 , RI9929020_397, \10182 );
and \U$8655 ( \10612 , RI992a790_377, \10184 );
and \U$8656 ( \10613 , RI992b0f0_357, \10186 );
and \U$8657 ( \10614 , RI992cc20_337, \10188 );
and \U$8658 ( \10615 , RI992d580_317, \10190 );
and \U$8659 ( \10616 , RI992f470_297, \10192 );
and \U$8660 ( \10617 , RI9931720_277, \10194 );
and \U$8661 ( \10618 , RI9933d90_257, \10196 );
or \U$8662 ( \10619 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 );
_DC g3abf ( \10620_nG3abf , \10619 , \10215 );
buf \U$8663 ( \10621 , \10620_nG3abf );
xor \U$8664 ( \10622 , \9904 , \9925 );
xor \U$8665 ( \10623 , \10622 , \10062 );
buf g35ea_GF_PartitionCandidate( \10624_nG35ea , \10623 );
buf \U$8666 ( \10625 , \10624_nG35ea );
xor \U$8667 ( \10626 , \9929 , \9950 );
xor \U$8668 ( \10627 , \10626 , \10059 );
buf g35c6_GF_PartitionCandidate( \10628_nG35c6 , \10627 );
buf \U$8669 ( \10629 , \10628_nG35c6 );
xor \U$8670 ( \10630 , \10625 , \10629 );
xor \U$8671 ( \10631 , \10629 , \10565 );
not \U$8672 ( \10632 , \10631 );
and \U$8673 ( \10633 , \10630 , \10632 );
and \U$8674 ( \10634 , \10621 , \10633 );
and \U$8675 ( \10635 , RI9922888_576, \10160 );
and \U$8676 ( \10636 , RI99234b8_556, \10166 );
and \U$8677 ( \10637 , RI9923e18_536, \10168 );
and \U$8678 ( \10638 , RI9924778_516, \10170 );
and \U$8679 ( \10639 , RI9925768_496, \10172 );
and \U$8680 ( \10640 , RI99260c8_476, \10174 );
and \U$8681 ( \10641 , RI9926a28_456, \10176 );
and \U$8682 ( \10642 , RI9927dd8_436, \10178 );
and \U$8683 ( \10643 , RI9928738_416, \10180 );
and \U$8684 ( \10644 , RI9929098_396, \10182 );
and \U$8685 ( \10645 , RI992a808_376, \10184 );
and \U$8686 ( \10646 , RI992b168_356, \10186 );
and \U$8687 ( \10647 , RI992cc98_336, \10188 );
and \U$8688 ( \10648 , RI992d5f8_316, \10190 );
and \U$8689 ( \10649 , RI992f4e8_296, \10192 );
and \U$8690 ( \10650 , RI9931798_276, \10194 );
and \U$8691 ( \10651 , RI9935ed8_256, \10196 );
or \U$8692 ( \10652 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 );
_DC g3b96 ( \10653_nG3b96 , \10652 , \10215 );
buf \U$8693 ( \10654 , \10653_nG3b96 );
and \U$8694 ( \10655 , \10654 , \10631 );
nor \U$8695 ( \10656 , \10634 , \10655 );
and \U$8696 ( \10657 , \10629 , \10565 );
not \U$8697 ( \10658 , \10657 );
and \U$8698 ( \10659 , \10625 , \10658 );
xnor \U$8699 ( \10660 , \10656 , \10659 );
and \U$8700 ( \10661 , \10600 , \10660 );
and \U$8701 ( \10662 , \10541 , \10660 );
or \U$8702 ( \10663 , \10601 , \10661 , \10662 );
and \U$8703 ( \10664 , RI9922720_579, \10160 );
and \U$8704 ( \10665 , RI9923350_559, \10166 );
and \U$8705 ( \10666 , RI9923cb0_539, \10168 );
and \U$8706 ( \10667 , RI9924610_519, \10170 );
and \U$8707 ( \10668 , RI9925600_499, \10172 );
and \U$8708 ( \10669 , RI9925f60_479, \10174 );
and \U$8709 ( \10670 , RI99268c0_459, \10176 );
and \U$8710 ( \10671 , RI9927c70_439, \10178 );
and \U$8711 ( \10672 , RI99285d0_419, \10180 );
and \U$8712 ( \10673 , RI9928f30_399, \10182 );
and \U$8713 ( \10674 , RI992a6a0_379, \10184 );
and \U$8714 ( \10675 , RI992b000_359, \10186 );
and \U$8715 ( \10676 , RI992cb30_339, \10188 );
and \U$8716 ( \10677 , RI992d490_319, \10190 );
and \U$8717 ( \10678 , RI992f380_299, \10192 );
and \U$8718 ( \10679 , RI9931630_279, \10194 );
and \U$8719 ( \10680 , RI9933ca0_259, \10196 );
or \U$8720 ( \10681 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 );
_DC g3900 ( \10682_nG3900 , \10681 , \10215 );
buf \U$8721 ( \10683 , \10682_nG3900 );
xor \U$8722 ( \10684 , \9879 , \9900 );
xor \U$8723 ( \10685 , \10684 , \10065 );
buf g3728_GF_PartitionCandidate( \10686_nG3728 , \10685 );
buf \U$8724 ( \10687 , \10686_nG3728 );
xor \U$8725 ( \10688 , \10389 , \10687 );
xor \U$8726 ( \10689 , \10687 , \10625 );
not \U$8727 ( \10690 , \10689 );
and \U$8728 ( \10691 , \10688 , \10690 );
and \U$8729 ( \10692 , \10683 , \10691 );
and \U$8730 ( \10693 , RI9922798_578, \10160 );
and \U$8731 ( \10694 , RI99233c8_558, \10166 );
and \U$8732 ( \10695 , RI9923d28_538, \10168 );
and \U$8733 ( \10696 , RI9924688_518, \10170 );
and \U$8734 ( \10697 , RI9925678_498, \10172 );
and \U$8735 ( \10698 , RI9925fd8_478, \10174 );
and \U$8736 ( \10699 , RI9926938_458, \10176 );
and \U$8737 ( \10700 , RI9927ce8_438, \10178 );
and \U$8738 ( \10701 , RI9928648_418, \10180 );
and \U$8739 ( \10702 , RI9928fa8_398, \10182 );
and \U$8740 ( \10703 , RI992a718_378, \10184 );
and \U$8741 ( \10704 , RI992b078_358, \10186 );
and \U$8742 ( \10705 , RI992cba8_338, \10188 );
and \U$8743 ( \10706 , RI992d508_318, \10190 );
and \U$8744 ( \10707 , RI992f3f8_298, \10192 );
and \U$8745 ( \10708 , RI99316a8_278, \10194 );
and \U$8746 ( \10709 , RI9933d18_258, \10196 );
or \U$8747 ( \10710 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 );
_DC g39c9 ( \10711_nG39c9 , \10710 , \10215 );
buf \U$8748 ( \10712 , \10711_nG39c9 );
and \U$8749 ( \10713 , \10712 , \10689 );
nor \U$8750 ( \10714 , \10692 , \10713 );
and \U$8751 ( \10715 , \10687 , \10625 );
not \U$8752 ( \10716 , \10715 );
and \U$8753 ( \10717 , \10389 , \10716 );
xnor \U$8754 ( \10718 , \10714 , \10717 );
and \U$8755 ( \10719 , RI9922630_581, \10160 );
and \U$8756 ( \10720 , RI9923260_561, \10166 );
and \U$8757 ( \10721 , RI9923bc0_541, \10168 );
and \U$8758 ( \10722 , RI9924520_521, \10170 );
and \U$8759 ( \10723 , RI9925510_501, \10172 );
and \U$8760 ( \10724 , RI9925e70_481, \10174 );
and \U$8761 ( \10725 , RI99267d0_461, \10176 );
and \U$8762 ( \10726 , RI9927b80_441, \10178 );
and \U$8763 ( \10727 , RI99284e0_421, \10180 );
and \U$8764 ( \10728 , RI9928e40_401, \10182 );
and \U$8765 ( \10729 , RI992a5b0_381, \10184 );
and \U$8766 ( \10730 , RI992af10_361, \10186 );
and \U$8767 ( \10731 , RI992ca40_341, \10188 );
and \U$8768 ( \10732 , RI992d3a0_321, \10190 );
and \U$8769 ( \10733 , RI992f290_301, \10192 );
and \U$8770 ( \10734 , RI9931540_281, \10194 );
and \U$8771 ( \10735 , RI9933bb0_261, \10196 );
or \U$8772 ( \10736 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 );
_DC g3767 ( \10737_nG3767 , \10736 , \10215 );
buf \U$8773 ( \10738 , \10737_nG3767 );
and \U$8774 ( \10739 , \10738 , \10392 );
and \U$8775 ( \10740 , RI99226a8_580, \10160 );
and \U$8776 ( \10741 , RI99232d8_560, \10166 );
and \U$8777 ( \10742 , RI9923c38_540, \10168 );
and \U$8778 ( \10743 , RI9924598_520, \10170 );
and \U$8779 ( \10744 , RI9925588_500, \10172 );
and \U$8780 ( \10745 , RI9925ee8_480, \10174 );
and \U$8781 ( \10746 , RI9926848_460, \10176 );
and \U$8782 ( \10747 , RI9927bf8_440, \10178 );
and \U$8783 ( \10748 , RI9928558_420, \10180 );
and \U$8784 ( \10749 , RI9928eb8_400, \10182 );
and \U$8785 ( \10750 , RI992a628_380, \10184 );
and \U$8786 ( \10751 , RI992af88_360, \10186 );
and \U$8787 ( \10752 , RI992cab8_340, \10188 );
and \U$8788 ( \10753 , RI992d418_320, \10190 );
and \U$8789 ( \10754 , RI992f308_300, \10192 );
and \U$8790 ( \10755 , RI99315b8_280, \10194 );
and \U$8791 ( \10756 , RI9933c28_260, \10196 );
or \U$8792 ( \10757 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 );
_DC g381a ( \10758_nG381a , \10757 , \10215 );
buf \U$8793 ( \10759 , \10758_nG381a );
and \U$8794 ( \10760 , \10759 , \10390 );
nor \U$8795 ( \10761 , \10739 , \10760 );
xnor \U$8796 ( \10762 , \10761 , \10397 );
and \U$8797 ( \10763 , \10718 , \10762 );
and \U$8798 ( \10764 , RI9922540_583, \10160 );
and \U$8799 ( \10765 , RI9923170_563, \10166 );
and \U$8800 ( \10766 , RI9923ad0_543, \10168 );
and \U$8801 ( \10767 , RI9924430_523, \10170 );
and \U$8802 ( \10768 , RI9924d90_503, \10172 );
and \U$8803 ( \10769 , RI9925d80_483, \10174 );
and \U$8804 ( \10770 , RI99266e0_463, \10176 );
and \U$8805 ( \10771 , RI9927040_443, \10178 );
and \U$8806 ( \10772 , RI99283f0_423, \10180 );
and \U$8807 ( \10773 , RI9928d50_403, \10182 );
and \U$8808 ( \10774 , RI992a4c0_383, \10184 );
and \U$8809 ( \10775 , RI992ae20_363, \10186 );
and \U$8810 ( \10776 , RI992c950_343, \10188 );
and \U$8811 ( \10777 , RI992d2b0_323, \10190 );
and \U$8812 ( \10778 , RI992f1a0_303, \10192 );
and \U$8813 ( \10779 , RI9931450_283, \10194 );
and \U$8814 ( \10780 , RI9933ac0_263, \10196 );
or \U$8815 ( \10781 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 );
_DC g3603 ( \10782_nG3603 , \10781 , \10215 );
buf \U$8816 ( \10783 , \10782_nG3603 );
and \U$8817 ( \10784 , \10783 , \10327 );
and \U$8818 ( \10785 , RI99225b8_582, \10160 );
and \U$8819 ( \10786 , RI99231e8_562, \10166 );
and \U$8820 ( \10787 , RI9923b48_542, \10168 );
and \U$8821 ( \10788 , RI99244a8_522, \10170 );
and \U$8822 ( \10789 , RI9924e08_502, \10172 );
and \U$8823 ( \10790 , RI9925df8_482, \10174 );
and \U$8824 ( \10791 , RI9926758_462, \10176 );
and \U$8825 ( \10792 , RI9927b08_442, \10178 );
and \U$8826 ( \10793 , RI9928468_422, \10180 );
and \U$8827 ( \10794 , RI9928dc8_402, \10182 );
and \U$8828 ( \10795 , RI992a538_382, \10184 );
and \U$8829 ( \10796 , RI992ae98_362, \10186 );
and \U$8830 ( \10797 , RI992c9c8_342, \10188 );
and \U$8831 ( \10798 , RI992d328_322, \10190 );
and \U$8832 ( \10799 , RI992f218_302, \10192 );
and \U$8833 ( \10800 , RI99314c8_282, \10194 );
and \U$8834 ( \10801 , RI9933b38_262, \10196 );
or \U$8835 ( \10802 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 );
_DC g36aa ( \10803_nG36aa , \10802 , \10215 );
buf \U$8836 ( \10804 , \10803_nG36aa );
and \U$8837 ( \10805 , \10804 , \10325 );
nor \U$8838 ( \10806 , \10784 , \10805 );
xnor \U$8839 ( \10807 , \10806 , \10094 );
and \U$8840 ( \10808 , \10762 , \10807 );
and \U$8841 ( \10809 , \10718 , \10807 );
or \U$8842 ( \10810 , \10763 , \10808 , \10809 );
and \U$8843 ( \10811 , \10663 , \10810 );
and \U$8844 ( \10812 , RI9922450_585, \10160 );
and \U$8845 ( \10813 , RI9923080_565, \10166 );
and \U$8846 ( \10814 , RI99239e0_545, \10168 );
and \U$8847 ( \10815 , RI9924340_525, \10170 );
and \U$8848 ( \10816 , RI9924ca0_505, \10172 );
and \U$8849 ( \10817 , RI9925c90_485, \10174 );
and \U$8850 ( \10818 , RI99265f0_465, \10176 );
and \U$8851 ( \10819 , RI9926f50_445, \10178 );
and \U$8852 ( \10820 , RI9928300_425, \10180 );
and \U$8853 ( \10821 , RI9928c60_405, \10182 );
and \U$8854 ( \10822 , RI992a3d0_385, \10184 );
and \U$8855 ( \10823 , RI992ad30_365, \10186 );
and \U$8856 ( \10824 , RI992c860_345, \10188 );
and \U$8857 ( \10825 , RI992d1c0_325, \10190 );
and \U$8858 ( \10826 , RI992f0b0_305, \10192 );
and \U$8859 ( \10827 , RI9931360_285, \10194 );
and \U$8860 ( \10828 , RI99339d0_265, \10196 );
or \U$8861 ( \10829 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 );
_DC g3493 ( \10830_nG3493 , \10829 , \10215 );
buf \U$8862 ( \10831 , \10830_nG3493 );
and \U$8863 ( \10832 , \10831 , \10265 );
and \U$8864 ( \10833 , RI99224c8_584, \10160 );
and \U$8865 ( \10834 , RI99230f8_564, \10166 );
and \U$8866 ( \10835 , RI9923a58_544, \10168 );
and \U$8867 ( \10836 , RI99243b8_524, \10170 );
and \U$8868 ( \10837 , RI9924d18_504, \10172 );
and \U$8869 ( \10838 , RI9925d08_484, \10174 );
and \U$8870 ( \10839 , RI9926668_464, \10176 );
and \U$8871 ( \10840 , RI9926fc8_444, \10178 );
and \U$8872 ( \10841 , RI9928378_424, \10180 );
and \U$8873 ( \10842 , RI9928cd8_404, \10182 );
and \U$8874 ( \10843 , RI992a448_384, \10184 );
and \U$8875 ( \10844 , RI992ada8_364, \10186 );
and \U$8876 ( \10845 , RI992c8d8_344, \10188 );
and \U$8877 ( \10846 , RI992d238_324, \10190 );
and \U$8878 ( \10847 , RI992f128_304, \10192 );
and \U$8879 ( \10848 , RI99313d8_284, \10194 );
and \U$8880 ( \10849 , RI9933a48_264, \10196 );
or \U$8881 ( \10850 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 );
_DC g3564 ( \10851_nG3564 , \10850 , \10215 );
buf \U$8882 ( \10852 , \10851_nG3564 );
and \U$8883 ( \10853 , \10852 , \10263 );
nor \U$8884 ( \10854 , \10832 , \10853 );
xnor \U$8885 ( \10855 , \10854 , \10291 );
and \U$8887 ( \10856 , RI99223d8_586, \10160 );
and \U$8888 ( \10857 , RI9923008_566, \10166 );
and \U$8889 ( \10858 , RI9923968_546, \10168 );
and \U$8890 ( \10859 , RI99242c8_526, \10170 );
and \U$8891 ( \10860 , RI9924c28_506, \10172 );
and \U$8892 ( \10861 , RI9925c18_486, \10174 );
and \U$8893 ( \10862 , RI9926578_466, \10176 );
and \U$8894 ( \10863 , RI9926ed8_446, \10178 );
and \U$8895 ( \10864 , RI9928288_426, \10180 );
and \U$8896 ( \10865 , RI9928be8_406, \10182 );
and \U$8897 ( \10866 , RI992a358_386, \10184 );
and \U$8898 ( \10867 , RI992acb8_366, \10186 );
and \U$8899 ( \10868 , RI992c7e8_346, \10188 );
and \U$8900 ( \10869 , RI992d148_326, \10190 );
and \U$8901 ( \10870 , RI992f038_306, \10192 );
and \U$8902 ( \10871 , RI99312e8_286, \10194 );
and \U$8903 ( \10872 , RI9933958_266, \10196 );
or \U$8904 ( \10873 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 );
_DC g3451 ( \10874_nG3451 , \10873 , \10215 );
buf \U$8905 ( \10875 , \10874_nG3451 );
and \U$8906 ( \10876 , \10875 , \10318 );
nor \U$8907 ( \10877 , 1'b0 , \10876 );
xnor \U$8908 ( \10878 , \10877 , 1'b0 );
and \U$8909 ( \10879 , \10855 , \10878 );
and \U$8910 ( \10880 , \10810 , \10879 );
and \U$8911 ( \10881 , \10663 , \10879 );
or \U$8912 ( \10882 , \10811 , \10880 , \10881 );
and \U$8914 ( \10883 , \10804 , \10327 );
and \U$8915 ( \10884 , \10738 , \10325 );
nor \U$8916 ( \10885 , \10883 , \10884 );
xnor \U$8917 ( \10886 , \10885 , \10094 );
and \U$8918 ( \10887 , \10852 , \10265 );
and \U$8919 ( \10888 , \10783 , \10263 );
nor \U$8920 ( \10889 , \10887 , \10888 );
xnor \U$8921 ( \10890 , \10889 , \10291 );
xor \U$8922 ( \10891 , \10886 , \10890 );
and \U$8924 ( \10892 , \10831 , \10318 );
nor \U$8925 ( \10893 , 1'b0 , \10892 );
xnor \U$8926 ( \10894 , \10893 , 1'b0 );
xor \U$8927 ( \10895 , \10891 , \10894 );
and \U$8928 ( \10896 , \10654 , \10633 );
and \U$8929 ( \10897 , \10561 , \10631 );
nor \U$8930 ( \10898 , \10896 , \10897 );
xnor \U$8931 ( \10899 , \10898 , \10659 );
and \U$8932 ( \10900 , \10712 , \10691 );
and \U$8933 ( \10901 , \10621 , \10689 );
nor \U$8934 ( \10902 , \10900 , \10901 );
xnor \U$8935 ( \10903 , \10902 , \10717 );
xor \U$8936 ( \10904 , \10899 , \10903 );
and \U$8937 ( \10905 , \10759 , \10392 );
and \U$8938 ( \10906 , \10683 , \10390 );
nor \U$8939 ( \10907 , \10905 , \10906 );
xnor \U$8940 ( \10908 , \10907 , \10397 );
xor \U$8941 ( \10909 , \10904 , \10908 );
and \U$8942 ( \10910 , \10895 , \10909 );
or \U$8944 ( \10911 , 1'b0 , \10910 , 1'b0 );
xor \U$8945 ( \10912 , \10882 , \10911 );
and \U$8946 ( \10913 , \10783 , \10265 );
and \U$8947 ( \10914 , \10804 , \10263 );
nor \U$8948 ( \10915 , \10913 , \10914 );
xnor \U$8949 ( \10916 , \10915 , \10291 );
and \U$8951 ( \10917 , \10852 , \10318 );
nor \U$8952 ( \10918 , 1'b0 , \10917 );
xnor \U$8953 ( \10919 , \10918 , 1'b0 );
xor \U$8954 ( \10920 , \10916 , \10919 );
xor \U$8956 ( \10921 , \10920 , 1'b0 );
and \U$8957 ( \10922 , \10621 , \10691 );
and \U$8958 ( \10923 , \10654 , \10689 );
nor \U$8959 ( \10924 , \10922 , \10923 );
xnor \U$8960 ( \10925 , \10924 , \10717 );
and \U$8961 ( \10926 , \10683 , \10392 );
and \U$8962 ( \10927 , \10712 , \10390 );
nor \U$8963 ( \10928 , \10926 , \10927 );
xnor \U$8964 ( \10929 , \10928 , \10397 );
xor \U$8965 ( \10930 , \10925 , \10929 );
and \U$8966 ( \10931 , \10738 , \10327 );
and \U$8967 ( \10932 , \10759 , \10325 );
nor \U$8968 ( \10933 , \10931 , \10932 );
xnor \U$8969 ( \10934 , \10933 , \10094 );
xor \U$8970 ( \10935 , \10930 , \10934 );
xor \U$8971 ( \10936 , \10921 , \10935 );
and \U$8972 ( \10937 , \10445 , \10537 );
and \U$8973 ( \10938 , \10313 , \10534 );
nor \U$8974 ( \10939 , \10937 , \10938 );
xnor \U$8975 ( \10940 , \10939 , \10531 );
and \U$8976 ( \10941 , \10468 , \10573 );
and \U$8977 ( \10942 , \10424 , \10571 );
nor \U$8978 ( \10943 , \10941 , \10942 );
xnor \U$8979 ( \10944 , \10943 , \10599 );
xor \U$8980 ( \10945 , \10940 , \10944 );
and \U$8981 ( \10946 , \10561 , \10633 );
and \U$8982 ( \10947 , \10594 , \10631 );
nor \U$8983 ( \10948 , \10946 , \10947 );
xnor \U$8984 ( \10949 , \10948 , \10659 );
xor \U$8985 ( \10950 , \10945 , \10949 );
xor \U$8986 ( \10951 , \10936 , \10950 );
xor \U$8987 ( \10952 , \10912 , \10951 );
and \U$8989 ( \10953 , \10594 , \10537 );
and \U$8990 ( \10954 , \10468 , \10534 );
nor \U$8991 ( \10955 , \10953 , \10954 );
xnor \U$8992 ( \10956 , \10955 , \10531 );
and \U$8993 ( \10957 , \10654 , \10573 );
and \U$8994 ( \10958 , \10561 , \10571 );
nor \U$8995 ( \10959 , \10957 , \10958 );
xnor \U$8996 ( \10960 , \10959 , \10599 );
and \U$8997 ( \10961 , \10956 , \10960 );
or \U$8999 ( \10962 , 1'b0 , \10961 , 1'b0 );
and \U$9000 ( \10963 , \10712 , \10633 );
and \U$9001 ( \10964 , \10621 , \10631 );
nor \U$9002 ( \10965 , \10963 , \10964 );
xnor \U$9003 ( \10966 , \10965 , \10659 );
and \U$9004 ( \10967 , \10759 , \10691 );
and \U$9005 ( \10968 , \10683 , \10689 );
nor \U$9006 ( \10969 , \10967 , \10968 );
xnor \U$9007 ( \10970 , \10969 , \10717 );
and \U$9008 ( \10971 , \10966 , \10970 );
and \U$9009 ( \10972 , \10804 , \10392 );
and \U$9010 ( \10973 , \10738 , \10390 );
nor \U$9011 ( \10974 , \10972 , \10973 );
xnor \U$9012 ( \10975 , \10974 , \10397 );
and \U$9013 ( \10976 , \10970 , \10975 );
and \U$9014 ( \10977 , \10966 , \10975 );
or \U$9015 ( \10978 , \10971 , \10976 , \10977 );
and \U$9016 ( \10979 , \10962 , \10978 );
and \U$9017 ( \10980 , \10852 , \10327 );
and \U$9018 ( \10981 , \10783 , \10325 );
nor \U$9019 ( \10982 , \10980 , \10981 );
xnor \U$9020 ( \10983 , \10982 , \10094 );
and \U$9021 ( \10984 , \10875 , \10265 );
and \U$9022 ( \10985 , \10831 , \10263 );
nor \U$9023 ( \10986 , \10984 , \10985 );
xnor \U$9024 ( \10987 , \10986 , \10291 );
and \U$9025 ( \10988 , \10983 , \10987 );
and \U$9026 ( \10989 , RI9922360_587, \10160 );
and \U$9027 ( \10990 , RI9922f90_567, \10166 );
and \U$9028 ( \10991 , RI99238f0_547, \10168 );
and \U$9029 ( \10992 , RI9924250_527, \10170 );
and \U$9030 ( \10993 , RI9924bb0_507, \10172 );
and \U$9031 ( \10994 , RI9925ba0_487, \10174 );
and \U$9032 ( \10995 , RI9926500_467, \10176 );
and \U$9033 ( \10996 , RI9926e60_447, \10178 );
and \U$9034 ( \10997 , RI9928210_427, \10180 );
and \U$9035 ( \10998 , RI9928b70_407, \10182 );
and \U$9036 ( \10999 , RI992a2e0_387, \10184 );
and \U$9037 ( \11000 , RI992ac40_367, \10186 );
and \U$9038 ( \11001 , RI992c770_347, \10188 );
and \U$9039 ( \11002 , RI992d0d0_327, \10190 );
and \U$9040 ( \11003 , RI992efc0_307, \10192 );
and \U$9041 ( \11004 , RI992f920_287, \10194 );
and \U$9042 ( \11005 , RI99338e0_267, \10196 );
or \U$9043 ( \11006 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 );
_DC g333d ( \11007_nG333d , \11006 , \10215 );
buf \U$9044 ( \11008 , \11007_nG333d );
nand \U$9045 ( \11009 , \11008 , \10318 );
xnor \U$9046 ( \11010 , \11009 , 1'b0 );
and \U$9047 ( \11011 , \10987 , \11010 );
and \U$9048 ( \11012 , \10983 , \11010 );
or \U$9049 ( \11013 , \10988 , \11011 , \11012 );
and \U$9050 ( \11014 , \10978 , \11013 );
and \U$9051 ( \11015 , \10962 , \11013 );
or \U$9052 ( \11016 , \10979 , \11014 , \11015 );
xor \U$9053 ( \11017 , \10855 , \10878 );
xor \U$9054 ( \11018 , \10718 , \10762 );
xor \U$9055 ( \11019 , \11018 , \10807 );
and \U$9056 ( \11020 , \11017 , \11019 );
xor \U$9057 ( \11021 , \10541 , \10600 );
xor \U$9058 ( \11022 , \11021 , \10660 );
and \U$9059 ( \11023 , \11019 , \11022 );
and \U$9060 ( \11024 , \11017 , \11022 );
or \U$9061 ( \11025 , \11020 , \11023 , \11024 );
and \U$9062 ( \11026 , \11016 , \11025 );
and \U$9064 ( \11027 , \10424 , \10537 );
and \U$9065 ( \11028 , \10445 , \10534 );
nor \U$9066 ( \11029 , \11027 , \11028 );
xnor \U$9067 ( \11030 , \11029 , \10531 );
xor \U$9068 ( \11031 , 1'b0 , \11030 );
and \U$9069 ( \11032 , \10594 , \10573 );
and \U$9070 ( \11033 , \10468 , \10571 );
nor \U$9071 ( \11034 , \11032 , \11033 );
xnor \U$9072 ( \11035 , \11034 , \10599 );
xor \U$9073 ( \11036 , \11031 , \11035 );
and \U$9074 ( \11037 , \11025 , \11036 );
and \U$9075 ( \11038 , \11016 , \11036 );
or \U$9076 ( \11039 , \11026 , \11037 , \11038 );
xor \U$9078 ( \11040 , 1'b0 , \10895 );
xor \U$9079 ( \11041 , \11040 , \10909 );
xor \U$9080 ( \11042 , \10663 , \10810 );
xor \U$9081 ( \11043 , \11042 , \10879 );
and \U$9082 ( \11044 , \11041 , \11043 );
xor \U$9083 ( \11045 , \11039 , \11044 );
and \U$9085 ( \11046 , \11030 , \11035 );
or \U$9087 ( \11047 , 1'b0 , \11046 , 1'b0 );
and \U$9088 ( \11048 , \10899 , \10903 );
and \U$9089 ( \11049 , \10903 , \10908 );
and \U$9090 ( \11050 , \10899 , \10908 );
or \U$9091 ( \11051 , \11048 , \11049 , \11050 );
xor \U$9092 ( \11052 , \11047 , \11051 );
and \U$9093 ( \11053 , \10886 , \10890 );
and \U$9094 ( \11054 , \10890 , \10894 );
and \U$9095 ( \11055 , \10886 , \10894 );
or \U$9096 ( \11056 , \11053 , \11054 , \11055 );
xor \U$9097 ( \11057 , \11052 , \11056 );
xor \U$9098 ( \11058 , \11045 , \11057 );
xor \U$9099 ( \11059 , \10952 , \11058 );
and \U$9100 ( \11060 , \10561 , \10537 );
and \U$9101 ( \11061 , \10594 , \10534 );
nor \U$9102 ( \11062 , \11060 , \11061 );
xnor \U$9103 ( \11063 , \11062 , \10531 );
and \U$9104 ( \11064 , \10621 , \10573 );
and \U$9105 ( \11065 , \10654 , \10571 );
nor \U$9106 ( \11066 , \11064 , \11065 );
xnor \U$9107 ( \11067 , \11066 , \10599 );
and \U$9108 ( \11068 , \11063 , \11067 );
and \U$9109 ( \11069 , \10683 , \10633 );
and \U$9110 ( \11070 , \10712 , \10631 );
nor \U$9111 ( \11071 , \11069 , \11070 );
xnor \U$9112 ( \11072 , \11071 , \10659 );
and \U$9113 ( \11073 , \11067 , \11072 );
and \U$9114 ( \11074 , \11063 , \11072 );
or \U$9115 ( \11075 , \11068 , \11073 , \11074 );
and \U$9116 ( \11076 , \10738 , \10691 );
and \U$9117 ( \11077 , \10759 , \10689 );
nor \U$9118 ( \11078 , \11076 , \11077 );
xnor \U$9119 ( \11079 , \11078 , \10717 );
and \U$9120 ( \11080 , \10783 , \10392 );
and \U$9121 ( \11081 , \10804 , \10390 );
nor \U$9122 ( \11082 , \11080 , \11081 );
xnor \U$9123 ( \11083 , \11082 , \10397 );
and \U$9124 ( \11084 , \11079 , \11083 );
and \U$9125 ( \11085 , \10831 , \10327 );
and \U$9126 ( \11086 , \10852 , \10325 );
nor \U$9127 ( \11087 , \11085 , \11086 );
xnor \U$9128 ( \11088 , \11087 , \10094 );
and \U$9129 ( \11089 , \11083 , \11088 );
and \U$9130 ( \11090 , \11079 , \11088 );
or \U$9131 ( \11091 , \11084 , \11089 , \11090 );
and \U$9132 ( \11092 , \11075 , \11091 );
xor \U$9133 ( \11093 , \10983 , \10987 );
xor \U$9134 ( \11094 , \11093 , \11010 );
and \U$9135 ( \11095 , \11091 , \11094 );
and \U$9136 ( \11096 , \11075 , \11094 );
or \U$9137 ( \11097 , \11092 , \11095 , \11096 );
xor \U$9138 ( \11098 , \10966 , \10970 );
xor \U$9139 ( \11099 , \11098 , \10975 );
xor \U$9140 ( \11100 , 1'b0 , \10956 );
xor \U$9141 ( \11101 , \11100 , \10960 );
and \U$9142 ( \11102 , \11099 , \11101 );
and \U$9143 ( \11103 , \11097 , \11102 );
xor \U$9144 ( \11104 , \11017 , \11019 );
xor \U$9145 ( \11105 , \11104 , \11022 );
and \U$9146 ( \11106 , \11102 , \11105 );
and \U$9147 ( \11107 , \11097 , \11105 );
or \U$9148 ( \11108 , \11103 , \11106 , \11107 );
xor \U$9149 ( \11109 , \11041 , \11043 );
and \U$9150 ( \11110 , \11108 , \11109 );
xor \U$9151 ( \11111 , \11016 , \11025 );
xor \U$9152 ( \11112 , \11111 , \11036 );
and \U$9153 ( \11113 , \11109 , \11112 );
and \U$9154 ( \11114 , \11108 , \11112 );
or \U$9155 ( \11115 , \11110 , \11113 , \11114 );
nor \U$9156 ( \11116 , \11059 , \11115 );
and \U$9157 ( \11117 , \11039 , \11044 );
and \U$9158 ( \11118 , \11044 , \11057 );
and \U$9159 ( \11119 , \11039 , \11057 );
or \U$9160 ( \11120 , \11117 , \11118 , \11119 );
and \U$9161 ( \11121 , \10882 , \10911 );
and \U$9162 ( \11122 , \10911 , \10951 );
and \U$9163 ( \11123 , \10882 , \10951 );
or \U$9164 ( \11124 , \11121 , \11122 , \11123 );
and \U$9166 ( \11125 , \10313 , \10537 );
and \U$9167 ( \11126 , \10217 , \10534 );
nor \U$9168 ( \11127 , \11125 , \11126 );
xnor \U$9169 ( \11128 , \11127 , \10531 );
xor \U$9170 ( \11129 , 1'b0 , \11128 );
and \U$9171 ( \11130 , \10424 , \10573 );
and \U$9172 ( \11131 , \10445 , \10571 );
nor \U$9173 ( \11132 , \11130 , \11131 );
xnor \U$9174 ( \11133 , \11132 , \10599 );
xor \U$9175 ( \11134 , \11129 , \11133 );
and \U$9177 ( \11135 , \10759 , \10327 );
and \U$9178 ( \11136 , \10683 , \10325 );
nor \U$9179 ( \11137 , \11135 , \11136 );
xnor \U$9180 ( \11138 , \11137 , \10094 );
and \U$9181 ( \11139 , \10804 , \10265 );
and \U$9182 ( \11140 , \10738 , \10263 );
nor \U$9183 ( \11141 , \11139 , \11140 );
xnor \U$9184 ( \11142 , \11141 , \10291 );
xor \U$9185 ( \11143 , \11138 , \11142 );
and \U$9187 ( \11144 , \10783 , \10318 );
nor \U$9188 ( \11145 , 1'b0 , \11144 );
xnor \U$9189 ( \11146 , \11145 , 1'b0 );
xor \U$9190 ( \11147 , \11143 , \11146 );
xor \U$9191 ( \11148 , 1'b0 , \11147 );
xor \U$9192 ( \11149 , \11134 , \11148 );
and \U$9193 ( \11150 , \10940 , \10944 );
and \U$9194 ( \11151 , \10944 , \10949 );
and \U$9195 ( \11152 , \10940 , \10949 );
or \U$9196 ( \11153 , \11150 , \11151 , \11152 );
and \U$9197 ( \11154 , \10925 , \10929 );
and \U$9198 ( \11155 , \10929 , \10934 );
and \U$9199 ( \11156 , \10925 , \10934 );
or \U$9200 ( \11157 , \11154 , \11155 , \11156 );
xor \U$9201 ( \11158 , \11153 , \11157 );
and \U$9202 ( \11159 , \10916 , \10919 );
or \U$9205 ( \11160 , \11159 , 1'b0 , 1'b0 );
xor \U$9206 ( \11161 , \11158 , \11160 );
xor \U$9207 ( \11162 , \11149 , \11161 );
xor \U$9208 ( \11163 , \11124 , \11162 );
and \U$9209 ( \11164 , \11047 , \11051 );
and \U$9210 ( \11165 , \11051 , \11056 );
and \U$9211 ( \11166 , \11047 , \11056 );
or \U$9212 ( \11167 , \11164 , \11165 , \11166 );
and \U$9213 ( \11168 , \10921 , \10935 );
and \U$9214 ( \11169 , \10935 , \10950 );
and \U$9215 ( \11170 , \10921 , \10950 );
or \U$9216 ( \11171 , \11168 , \11169 , \11170 );
xor \U$9217 ( \11172 , \11167 , \11171 );
and \U$9218 ( \11173 , \10594 , \10633 );
and \U$9219 ( \11174 , \10468 , \10631 );
nor \U$9220 ( \11175 , \11173 , \11174 );
xnor \U$9221 ( \11176 , \11175 , \10659 );
and \U$9222 ( \11177 , \10654 , \10691 );
and \U$9223 ( \11178 , \10561 , \10689 );
nor \U$9224 ( \11179 , \11177 , \11178 );
xnor \U$9225 ( \11180 , \11179 , \10717 );
xor \U$9226 ( \11181 , \11176 , \11180 );
and \U$9227 ( \11182 , \10712 , \10392 );
and \U$9228 ( \11183 , \10621 , \10390 );
nor \U$9229 ( \11184 , \11182 , \11183 );
xnor \U$9230 ( \11185 , \11184 , \10397 );
xor \U$9231 ( \11186 , \11181 , \11185 );
xor \U$9232 ( \11187 , \11172 , \11186 );
xor \U$9233 ( \11188 , \11163 , \11187 );
xor \U$9234 ( \11189 , \11120 , \11188 );
and \U$9235 ( \11190 , \10952 , \11058 );
nor \U$9236 ( \11191 , \11189 , \11190 );
nor \U$9237 ( \11192 , \11116 , \11191 );
and \U$9238 ( \11193 , \11124 , \11162 );
and \U$9239 ( \11194 , \11162 , \11187 );
and \U$9240 ( \11195 , \11124 , \11187 );
or \U$9241 ( \11196 , \11193 , \11194 , \11195 );
and \U$9243 ( \11197 , \11128 , \11133 );
or \U$9245 ( \11198 , 1'b0 , \11197 , 1'b0 );
and \U$9246 ( \11199 , \11176 , \11180 );
and \U$9247 ( \11200 , \11180 , \11185 );
and \U$9248 ( \11201 , \11176 , \11185 );
or \U$9249 ( \11202 , \11199 , \11200 , \11201 );
xor \U$9250 ( \11203 , \11198 , \11202 );
and \U$9251 ( \11204 , \11138 , \11142 );
and \U$9252 ( \11205 , \11142 , \11146 );
and \U$9253 ( \11206 , \11138 , \11146 );
or \U$9254 ( \11207 , \11204 , \11205 , \11206 );
xor \U$9255 ( \11208 , \11203 , \11207 );
and \U$9256 ( \11209 , \11153 , \11157 );
and \U$9257 ( \11210 , \11157 , \11160 );
and \U$9258 ( \11211 , \11153 , \11160 );
or \U$9259 ( \11212 , \11209 , \11210 , \11211 );
xor \U$9261 ( \11213 , \11212 , 1'b0 );
and \U$9262 ( \11214 , \10217 , \10537 );
and \U$9263 ( \11215 , \10286 , \10534 );
nor \U$9264 ( \11216 , \11214 , \11215 );
xnor \U$9265 ( \11217 , \11216 , \10531 );
and \U$9266 ( \11218 , \10445 , \10573 );
and \U$9267 ( \11219 , \10313 , \10571 );
nor \U$9268 ( \11220 , \11218 , \11219 );
xnor \U$9269 ( \11221 , \11220 , \10599 );
xor \U$9270 ( \11222 , \11217 , \11221 );
and \U$9271 ( \11223 , \10468 , \10633 );
and \U$9272 ( \11224 , \10424 , \10631 );
nor \U$9273 ( \11225 , \11223 , \11224 );
xnor \U$9274 ( \11226 , \11225 , \10659 );
xor \U$9275 ( \11227 , \11222 , \11226 );
xor \U$9276 ( \11228 , \11213 , \11227 );
xor \U$9277 ( \11229 , \11208 , \11228 );
xor \U$9278 ( \11230 , \11196 , \11229 );
and \U$9279 ( \11231 , \11167 , \11171 );
and \U$9280 ( \11232 , \11171 , \11186 );
and \U$9281 ( \11233 , \11167 , \11186 );
or \U$9282 ( \11234 , \11231 , \11232 , \11233 );
and \U$9283 ( \11235 , \11134 , \11148 );
and \U$9284 ( \11236 , \11148 , \11161 );
and \U$9285 ( \11237 , \11134 , \11161 );
or \U$9286 ( \11238 , \11235 , \11236 , \11237 );
xor \U$9287 ( \11239 , \11234 , \11238 );
and \U$9289 ( \11240 , \10738 , \10265 );
and \U$9290 ( \11241 , \10759 , \10263 );
nor \U$9291 ( \11242 , \11240 , \11241 );
xnor \U$9292 ( \11243 , \11242 , \10291 );
and \U$9294 ( \11244 , \10804 , \10318 );
nor \U$9295 ( \11245 , 1'b0 , \11244 );
xnor \U$9296 ( \11246 , \11245 , 1'b0 );
xor \U$9297 ( \11247 , \11243 , \11246 );
xor \U$9299 ( \11248 , \11247 , 1'b0 );
xor \U$9300 ( \11249 , 1'b0 , \11248 );
and \U$9301 ( \11250 , \10561 , \10691 );
and \U$9302 ( \11251 , \10594 , \10689 );
nor \U$9303 ( \11252 , \11250 , \11251 );
xnor \U$9304 ( \11253 , \11252 , \10717 );
and \U$9305 ( \11254 , \10621 , \10392 );
and \U$9306 ( \11255 , \10654 , \10390 );
nor \U$9307 ( \11256 , \11254 , \11255 );
xnor \U$9308 ( \11257 , \11256 , \10397 );
xor \U$9309 ( \11258 , \11253 , \11257 );
and \U$9310 ( \11259 , \10683 , \10327 );
and \U$9311 ( \11260 , \10712 , \10325 );
nor \U$9312 ( \11261 , \11259 , \11260 );
xnor \U$9313 ( \11262 , \11261 , \10094 );
xor \U$9314 ( \11263 , \11258 , \11262 );
xor \U$9315 ( \11264 , \11249 , \11263 );
xor \U$9316 ( \11265 , \11239 , \11264 );
xor \U$9317 ( \11266 , \11230 , \11265 );
and \U$9318 ( \11267 , \11120 , \11188 );
nor \U$9319 ( \11268 , \11266 , \11267 );
and \U$9320 ( \11269 , \11234 , \11238 );
and \U$9321 ( \11270 , \11238 , \11264 );
and \U$9322 ( \11271 , \11234 , \11264 );
or \U$9323 ( \11272 , \11269 , \11270 , \11271 );
and \U$9324 ( \11273 , \11208 , \11228 );
xor \U$9325 ( \11274 , \11272 , \11273 );
and \U$9328 ( \11275 , \11212 , \11227 );
or \U$9329 ( \11276 , 1'b0 , 1'b0 , \11275 );
and \U$9331 ( \11277 , \10712 , \10327 );
and \U$9332 ( \11278 , \10621 , \10325 );
nor \U$9333 ( \11279 , \11277 , \11278 );
xnor \U$9334 ( \11280 , \11279 , \10094 );
and \U$9335 ( \11281 , \10759 , \10265 );
and \U$9336 ( \11282 , \10683 , \10263 );
nor \U$9337 ( \11283 , \11281 , \11282 );
xnor \U$9338 ( \11284 , \11283 , \10291 );
xor \U$9339 ( \11285 , \11280 , \11284 );
and \U$9341 ( \11286 , \10738 , \10318 );
nor \U$9342 ( \11287 , 1'b0 , \11286 );
xnor \U$9343 ( \11288 , \11287 , 1'b0 );
xor \U$9344 ( \11289 , \11285 , \11288 );
xor \U$9345 ( \11290 , 1'b0 , \11289 );
and \U$9346 ( \11291 , \10424 , \10633 );
and \U$9347 ( \11292 , \10445 , \10631 );
nor \U$9348 ( \11293 , \11291 , \11292 );
xnor \U$9349 ( \11294 , \11293 , \10659 );
and \U$9350 ( \11295 , \10594 , \10691 );
and \U$9351 ( \11296 , \10468 , \10689 );
nor \U$9352 ( \11297 , \11295 , \11296 );
xnor \U$9353 ( \11298 , \11297 , \10717 );
xor \U$9354 ( \11299 , \11294 , \11298 );
and \U$9355 ( \11300 , \10654 , \10392 );
and \U$9356 ( \11301 , \10561 , \10390 );
nor \U$9357 ( \11302 , \11300 , \11301 );
xnor \U$9358 ( \11303 , \11302 , \10397 );
xor \U$9359 ( \11304 , \11299 , \11303 );
xor \U$9360 ( \11305 , \11290 , \11304 );
and \U$9361 ( \11306 , \11217 , \11221 );
and \U$9362 ( \11307 , \11221 , \11226 );
and \U$9363 ( \11308 , \11217 , \11226 );
or \U$9364 ( \11309 , \11306 , \11307 , \11308 );
and \U$9365 ( \11310 , \11253 , \11257 );
and \U$9366 ( \11311 , \11257 , \11262 );
and \U$9367 ( \11312 , \11253 , \11262 );
or \U$9368 ( \11313 , \11310 , \11311 , \11312 );
xor \U$9369 ( \11314 , \11309 , \11313 );
and \U$9370 ( \11315 , \11243 , \11246 );
or \U$9373 ( \11316 , \11315 , 1'b0 , 1'b0 );
xor \U$9374 ( \11317 , \11314 , \11316 );
xor \U$9375 ( \11318 , \11305 , \11317 );
xor \U$9376 ( \11319 , \11276 , \11318 );
and \U$9377 ( \11320 , \11198 , \11202 );
and \U$9378 ( \11321 , \11202 , \11207 );
and \U$9379 ( \11322 , \11198 , \11207 );
or \U$9380 ( \11323 , \11320 , \11321 , \11322 );
and \U$9382 ( \11324 , \11248 , \11263 );
or \U$9384 ( \11325 , 1'b0 , \11324 , 1'b0 );
xor \U$9385 ( \11326 , \11323 , \11325 );
and \U$9387 ( \11327 , \10286 , \10537 );
not \U$9388 ( \11328 , \11327 );
xnor \U$9389 ( \11329 , \11328 , \10531 );
xor \U$9390 ( \11330 , 1'b0 , \11329 );
and \U$9391 ( \11331 , \10313 , \10573 );
and \U$9392 ( \11332 , \10217 , \10571 );
nor \U$9393 ( \11333 , \11331 , \11332 );
xnor \U$9394 ( \11334 , \11333 , \10599 );
xor \U$9395 ( \11335 , \11330 , \11334 );
xor \U$9396 ( \11336 , \11326 , \11335 );
xor \U$9397 ( \11337 , \11319 , \11336 );
xor \U$9398 ( \11338 , \11274 , \11337 );
and \U$9399 ( \11339 , \11196 , \11229 );
and \U$9400 ( \11340 , \11229 , \11265 );
and \U$9401 ( \11341 , \11196 , \11265 );
or \U$9402 ( \11342 , \11339 , \11340 , \11341 );
nor \U$9403 ( \11343 , \11338 , \11342 );
nor \U$9404 ( \11344 , \11268 , \11343 );
nand \U$9405 ( \11345 , \11192 , \11344 );
and \U$9406 ( \11346 , \11276 , \11318 );
and \U$9407 ( \11347 , \11318 , \11336 );
and \U$9408 ( \11348 , \11276 , \11336 );
or \U$9409 ( \11349 , \11346 , \11347 , \11348 );
and \U$9410 ( \11350 , \11309 , \11313 );
and \U$9411 ( \11351 , \11313 , \11316 );
and \U$9412 ( \11352 , \11309 , \11316 );
or \U$9413 ( \11353 , \11350 , \11351 , \11352 );
and \U$9415 ( \11354 , \11289 , \11304 );
or \U$9417 ( \11355 , 1'b0 , \11354 , 1'b0 );
xor \U$9418 ( \11356 , \11353 , \11355 );
and \U$9419 ( \11357 , \10468 , \10691 );
and \U$9420 ( \11358 , \10424 , \10689 );
nor \U$9421 ( \11359 , \11357 , \11358 );
xnor \U$9422 ( \11360 , \11359 , \10717 );
and \U$9423 ( \11361 , \10561 , \10392 );
and \U$9424 ( \11362 , \10594 , \10390 );
nor \U$9425 ( \11363 , \11361 , \11362 );
xnor \U$9426 ( \11364 , \11363 , \10397 );
xor \U$9427 ( \11365 , \11360 , \11364 );
and \U$9428 ( \11366 , \10621 , \10327 );
and \U$9429 ( \11367 , \10654 , \10325 );
nor \U$9430 ( \11368 , \11366 , \11367 );
xnor \U$9431 ( \11369 , \11368 , \10094 );
xor \U$9432 ( \11370 , \11365 , \11369 );
xor \U$9433 ( \11371 , \11356 , \11370 );
xor \U$9434 ( \11372 , \11349 , \11371 );
and \U$9435 ( \11373 , \11323 , \11325 );
and \U$9436 ( \11374 , \11325 , \11335 );
and \U$9437 ( \11375 , \11323 , \11335 );
or \U$9438 ( \11376 , \11373 , \11374 , \11375 );
and \U$9439 ( \11377 , \11305 , \11317 );
xor \U$9440 ( \11378 , \11376 , \11377 );
not \U$9441 ( \11379 , \10531 );
and \U$9442 ( \11380 , \10217 , \10573 );
and \U$9443 ( \11381 , \10286 , \10571 );
nor \U$9444 ( \11382 , \11380 , \11381 );
xnor \U$9445 ( \11383 , \11382 , \10599 );
xor \U$9446 ( \11384 , \11379 , \11383 );
and \U$9447 ( \11385 , \10445 , \10633 );
and \U$9448 ( \11386 , \10313 , \10631 );
nor \U$9449 ( \11387 , \11385 , \11386 );
xnor \U$9450 ( \11388 , \11387 , \10659 );
xor \U$9451 ( \11389 , \11384 , \11388 );
and \U$9453 ( \11390 , \10683 , \10265 );
and \U$9454 ( \11391 , \10712 , \10263 );
nor \U$9455 ( \11392 , \11390 , \11391 );
xnor \U$9456 ( \11393 , \11392 , \10291 );
and \U$9458 ( \11394 , \10759 , \10318 );
nor \U$9459 ( \11395 , 1'b0 , \11394 );
xnor \U$9460 ( \11396 , \11395 , 1'b0 );
xor \U$9461 ( \11397 , \11393 , \11396 );
xor \U$9463 ( \11398 , \11397 , 1'b0 );
xor \U$9464 ( \11399 , 1'b1 , \11398 );
xor \U$9465 ( \11400 , \11389 , \11399 );
and \U$9467 ( \11401 , \11329 , \11334 );
or \U$9469 ( \11402 , 1'b0 , \11401 , 1'b0 );
and \U$9470 ( \11403 , \11294 , \11298 );
and \U$9471 ( \11404 , \11298 , \11303 );
and \U$9472 ( \11405 , \11294 , \11303 );
or \U$9473 ( \11406 , \11403 , \11404 , \11405 );
xor \U$9474 ( \11407 , \11402 , \11406 );
and \U$9475 ( \11408 , \11280 , \11284 );
and \U$9476 ( \11409 , \11284 , \11288 );
and \U$9477 ( \11410 , \11280 , \11288 );
or \U$9478 ( \11411 , \11408 , \11409 , \11410 );
xor \U$9479 ( \11412 , \11407 , \11411 );
xor \U$9480 ( \11413 , \11400 , \11412 );
xor \U$9481 ( \11414 , \11378 , \11413 );
xor \U$9482 ( \11415 , \11372 , \11414 );
and \U$9483 ( \11416 , \11272 , \11273 );
and \U$9484 ( \11417 , \11273 , \11337 );
and \U$9485 ( \11418 , \11272 , \11337 );
or \U$9486 ( \11419 , \11416 , \11417 , \11418 );
nor \U$9487 ( \11420 , \11415 , \11419 );
and \U$9488 ( \11421 , \11376 , \11377 );
and \U$9489 ( \11422 , \11377 , \11413 );
and \U$9490 ( \11423 , \11376 , \11413 );
or \U$9491 ( \11424 , \11421 , \11422 , \11423 );
and \U$9492 ( \11425 , \11379 , \11383 );
and \U$9493 ( \11426 , \11383 , \11388 );
and \U$9494 ( \11427 , \11379 , \11388 );
or \U$9495 ( \11428 , \11425 , \11426 , \11427 );
and \U$9496 ( \11429 , \11360 , \11364 );
and \U$9497 ( \11430 , \11364 , \11369 );
and \U$9498 ( \11431 , \11360 , \11369 );
or \U$9499 ( \11432 , \11429 , \11430 , \11431 );
xor \U$9500 ( \11433 , \11428 , \11432 );
and \U$9501 ( \11434 , \11393 , \11396 );
or \U$9504 ( \11435 , \11434 , 1'b0 , 1'b0 );
xor \U$9505 ( \11436 , \11433 , \11435 );
and \U$9506 ( \11437 , \11402 , \11406 );
and \U$9507 ( \11438 , \11406 , \11411 );
and \U$9508 ( \11439 , \11402 , \11411 );
or \U$9509 ( \11440 , \11437 , \11438 , \11439 );
and \U$9512 ( \11441 , 1'b1 , \11398 );
or \U$9514 ( \11442 , 1'b0 , \11441 , 1'b0 );
xor \U$9515 ( \11443 , \11440 , \11442 );
and \U$9516 ( \11444 , \10712 , \10265 );
and \U$9517 ( \11445 , \10621 , \10263 );
nor \U$9518 ( \11446 , \11444 , \11445 );
xnor \U$9519 ( \11447 , \11446 , \10291 );
and \U$9521 ( \11448 , \10683 , \10318 );
nor \U$9522 ( \11449 , 1'b0 , \11448 );
xnor \U$9523 ( \11450 , \11449 , 1'b0 );
xor \U$9524 ( \11451 , \11447 , \11450 );
xor \U$9526 ( \11452 , \11451 , 1'b0 );
and \U$9527 ( \11453 , \10424 , \10691 );
and \U$9528 ( \11454 , \10445 , \10689 );
nor \U$9529 ( \11455 , \11453 , \11454 );
xnor \U$9530 ( \11456 , \11455 , \10717 );
and \U$9531 ( \11457 , \10594 , \10392 );
and \U$9532 ( \11458 , \10468 , \10390 );
nor \U$9533 ( \11459 , \11457 , \11458 );
xnor \U$9534 ( \11460 , \11459 , \10397 );
xor \U$9535 ( \11461 , \11456 , \11460 );
and \U$9536 ( \11462 , \10654 , \10327 );
and \U$9537 ( \11463 , \10561 , \10325 );
nor \U$9538 ( \11464 , \11462 , \11463 );
xnor \U$9539 ( \11465 , \11464 , \10094 );
xor \U$9540 ( \11466 , \11461 , \11465 );
xor \U$9541 ( \11467 , \11452 , \11466 );
and \U$9543 ( \11468 , \10286 , \10573 );
not \U$9544 ( \11469 , \11468 );
xnor \U$9545 ( \11470 , \11469 , \10599 );
xor \U$9546 ( \11471 , 1'b0 , \11470 );
and \U$9547 ( \11472 , \10313 , \10633 );
and \U$9548 ( \11473 , \10217 , \10631 );
nor \U$9549 ( \11474 , \11472 , \11473 );
xnor \U$9550 ( \11475 , \11474 , \10659 );
xor \U$9551 ( \11476 , \11471 , \11475 );
xor \U$9552 ( \11477 , \11467 , \11476 );
xor \U$9553 ( \11478 , \11443 , \11477 );
xor \U$9554 ( \11479 , \11436 , \11478 );
xor \U$9555 ( \11480 , \11424 , \11479 );
and \U$9556 ( \11481 , \11353 , \11355 );
and \U$9557 ( \11482 , \11355 , \11370 );
and \U$9558 ( \11483 , \11353 , \11370 );
or \U$9559 ( \11484 , \11481 , \11482 , \11483 );
and \U$9560 ( \11485 , \11389 , \11399 );
and \U$9561 ( \11486 , \11399 , \11412 );
and \U$9562 ( \11487 , \11389 , \11412 );
or \U$9563 ( \11488 , \11485 , \11486 , \11487 );
xor \U$9564 ( \11489 , \11484 , \11488 );
xor \U$9566 ( \11490 , \11489 , 1'b1 );
xor \U$9567 ( \11491 , \11480 , \11490 );
and \U$9568 ( \11492 , \11349 , \11371 );
and \U$9569 ( \11493 , \11371 , \11414 );
and \U$9570 ( \11494 , \11349 , \11414 );
or \U$9571 ( \11495 , \11492 , \11493 , \11494 );
nor \U$9572 ( \11496 , \11491 , \11495 );
nor \U$9573 ( \11497 , \11420 , \11496 );
and \U$9574 ( \11498 , \11484 , \11488 );
and \U$9575 ( \11499 , \11488 , 1'b1 );
and \U$9576 ( \11500 , \11484 , 1'b1 );
or \U$9577 ( \11501 , \11498 , \11499 , \11500 );
and \U$9578 ( \11502 , \11436 , \11478 );
xor \U$9579 ( \11503 , \11501 , \11502 );
and \U$9580 ( \11504 , \11440 , \11442 );
and \U$9581 ( \11505 , \11442 , \11477 );
and \U$9582 ( \11506 , \11440 , \11477 );
or \U$9583 ( \11507 , \11504 , \11505 , \11506 );
and \U$9585 ( \11508 , \10712 , \10318 );
nor \U$9586 ( \11509 , 1'b0 , \11508 );
xnor \U$9587 ( \11510 , \11509 , 1'b0 );
xor \U$9589 ( \11511 , \11510 , 1'b0 );
xor \U$9591 ( \11512 , \11511 , 1'b0 );
and \U$9592 ( \11513 , \10468 , \10392 );
and \U$9593 ( \11514 , \10424 , \10390 );
nor \U$9594 ( \11515 , \11513 , \11514 );
xnor \U$9595 ( \11516 , \11515 , \10397 );
and \U$9596 ( \11517 , \10561 , \10327 );
and \U$9597 ( \11518 , \10594 , \10325 );
nor \U$9598 ( \11519 , \11517 , \11518 );
xnor \U$9599 ( \11520 , \11519 , \10094 );
xor \U$9600 ( \11521 , \11516 , \11520 );
and \U$9601 ( \11522 , \10621 , \10265 );
and \U$9602 ( \11523 , \10654 , \10263 );
nor \U$9603 ( \11524 , \11522 , \11523 );
xnor \U$9604 ( \11525 , \11524 , \10291 );
xor \U$9605 ( \11526 , \11521 , \11525 );
xor \U$9606 ( \11527 , \11512 , \11526 );
not \U$9607 ( \11528 , \10599 );
and \U$9608 ( \11529 , \10217 , \10633 );
and \U$9609 ( \11530 , \10286 , \10631 );
nor \U$9610 ( \11531 , \11529 , \11530 );
xnor \U$9611 ( \11532 , \11531 , \10659 );
xor \U$9612 ( \11533 , \11528 , \11532 );
and \U$9613 ( \11534 , \10445 , \10691 );
and \U$9614 ( \11535 , \10313 , \10689 );
nor \U$9615 ( \11536 , \11534 , \11535 );
xnor \U$9616 ( \11537 , \11536 , \10717 );
xor \U$9617 ( \11538 , \11533 , \11537 );
xor \U$9618 ( \11539 , \11527 , \11538 );
xor \U$9620 ( \11540 , \11539 , 1'b0 );
and \U$9622 ( \11541 , \11470 , \11475 );
or \U$9624 ( \11542 , 1'b0 , \11541 , 1'b0 );
and \U$9625 ( \11543 , \11456 , \11460 );
and \U$9626 ( \11544 , \11460 , \11465 );
and \U$9627 ( \11545 , \11456 , \11465 );
or \U$9628 ( \11546 , \11543 , \11544 , \11545 );
xor \U$9629 ( \11547 , \11542 , \11546 );
and \U$9630 ( \11548 , \11447 , \11450 );
or \U$9633 ( \11549 , \11548 , 1'b0 , 1'b0 );
xor \U$9634 ( \11550 , \11547 , \11549 );
xor \U$9635 ( \11551 , \11540 , \11550 );
xor \U$9636 ( \11552 , \11507 , \11551 );
and \U$9637 ( \11553 , \11428 , \11432 );
and \U$9638 ( \11554 , \11432 , \11435 );
and \U$9639 ( \11555 , \11428 , \11435 );
or \U$9640 ( \11556 , \11553 , \11554 , \11555 );
xor \U$9642 ( \11557 , \11556 , 1'b0 );
and \U$9643 ( \11558 , \11452 , \11466 );
and \U$9644 ( \11559 , \11466 , \11476 );
and \U$9645 ( \11560 , \11452 , \11476 );
or \U$9646 ( \11561 , \11558 , \11559 , \11560 );
xor \U$9647 ( \11562 , \11557 , \11561 );
xor \U$9648 ( \11563 , \11552 , \11562 );
xor \U$9649 ( \11564 , \11503 , \11563 );
and \U$9650 ( \11565 , \11424 , \11479 );
and \U$9651 ( \11566 , \11479 , \11490 );
and \U$9652 ( \11567 , \11424 , \11490 );
or \U$9653 ( \11568 , \11565 , \11566 , \11567 );
nor \U$9654 ( \11569 , \11564 , \11568 );
and \U$9655 ( \11570 , \11507 , \11551 );
and \U$9656 ( \11571 , \11551 , \11562 );
and \U$9657 ( \11572 , \11507 , \11562 );
or \U$9658 ( \11573 , \11570 , \11571 , \11572 );
and \U$9659 ( \11574 , \11542 , \11546 );
and \U$9660 ( \11575 , \11546 , \11549 );
and \U$9661 ( \11576 , \11542 , \11549 );
or \U$9662 ( \11577 , \11574 , \11575 , \11576 );
xor \U$9664 ( \11578 , \11577 , 1'b0 );
and \U$9665 ( \11579 , \11512 , \11526 );
and \U$9666 ( \11580 , \11526 , \11538 );
and \U$9667 ( \11581 , \11512 , \11538 );
or \U$9668 ( \11582 , \11579 , \11580 , \11581 );
xor \U$9669 ( \11583 , \11578 , \11582 );
xor \U$9670 ( \11584 , \11573 , \11583 );
and \U$9673 ( \11585 , \11556 , \11561 );
or \U$9674 ( \11586 , 1'b0 , 1'b0 , \11585 );
and \U$9677 ( \11587 , \11539 , \11550 );
or \U$9678 ( \11588 , 1'b0 , 1'b0 , \11587 );
xor \U$9679 ( \11589 , \11586 , \11588 );
and \U$9680 ( \11590 , \10424 , \10392 );
and \U$9681 ( \11591 , \10445 , \10390 );
nor \U$9682 ( \11592 , \11590 , \11591 );
xnor \U$9683 ( \11593 , \11592 , \10397 );
and \U$9684 ( \11594 , \10594 , \10327 );
and \U$9685 ( \11595 , \10468 , \10325 );
nor \U$9686 ( \11596 , \11594 , \11595 );
xnor \U$9687 ( \11597 , \11596 , \10094 );
xor \U$9688 ( \11598 , \11593 , \11597 );
and \U$9689 ( \11599 , \10654 , \10265 );
and \U$9690 ( \11600 , \10561 , \10263 );
nor \U$9691 ( \11601 , \11599 , \11600 );
xnor \U$9692 ( \11602 , \11601 , \10291 );
xor \U$9693 ( \11603 , \11598 , \11602 );
and \U$9695 ( \11604 , \10286 , \10633 );
not \U$9696 ( \11605 , \11604 );
xnor \U$9697 ( \11606 , \11605 , \10659 );
xor \U$9698 ( \11607 , 1'b0 , \11606 );
and \U$9699 ( \11608 , \10313 , \10691 );
and \U$9700 ( \11609 , \10217 , \10689 );
nor \U$9701 ( \11610 , \11608 , \11609 );
xnor \U$9702 ( \11611 , \11610 , \10717 );
xor \U$9703 ( \11612 , \11607 , \11611 );
xor \U$9704 ( \11613 , \11603 , \11612 );
and \U$9707 ( \11614 , \10621 , \10318 );
nor \U$9708 ( \11615 , 1'b0 , \11614 );
xnor \U$9709 ( \11616 , \11615 , 1'b0 );
xor \U$9711 ( \11617 , \11616 , 1'b0 );
xor \U$9713 ( \11618 , \11617 , 1'b0 );
xnor \U$9714 ( \11619 , 1'b0 , \11618 );
xor \U$9715 ( \11620 , \11613 , \11619 );
and \U$9716 ( \11621 , \11528 , \11532 );
and \U$9717 ( \11622 , \11532 , \11537 );
and \U$9718 ( \11623 , \11528 , \11537 );
or \U$9719 ( \11624 , \11621 , \11622 , \11623 );
and \U$9720 ( \11625 , \11516 , \11520 );
and \U$9721 ( \11626 , \11520 , \11525 );
and \U$9722 ( \11627 , \11516 , \11525 );
or \U$9723 ( \11628 , \11625 , \11626 , \11627 );
xor \U$9724 ( \11629 , \11624 , \11628 );
xor \U$9726 ( \11630 , \11629 , 1'b0 );
xor \U$9727 ( \11631 , \11620 , \11630 );
xor \U$9728 ( \11632 , \11589 , \11631 );
xor \U$9729 ( \11633 , \11584 , \11632 );
and \U$9730 ( \11634 , \11501 , \11502 );
and \U$9731 ( \11635 , \11502 , \11563 );
and \U$9732 ( \11636 , \11501 , \11563 );
or \U$9733 ( \11637 , \11634 , \11635 , \11636 );
nor \U$9734 ( \11638 , \11633 , \11637 );
nor \U$9735 ( \11639 , \11569 , \11638 );
nand \U$9736 ( \11640 , \11497 , \11639 );
nor \U$9737 ( \11641 , \11345 , \11640 );
and \U$9738 ( \11642 , \11586 , \11588 );
and \U$9739 ( \11643 , \11588 , \11631 );
and \U$9740 ( \11644 , \11586 , \11631 );
or \U$9741 ( \11645 , \11642 , \11643 , \11644 );
and \U$9742 ( \11646 , \11624 , \11628 );
or \U$9745 ( \11647 , \11646 , 1'b0 , 1'b0 );
or \U$9746 ( \11648 , 1'b0 , \11618 );
xor \U$9747 ( \11649 , \11647 , \11648 );
and \U$9748 ( \11650 , \11603 , \11612 );
xor \U$9749 ( \11651 , \11649 , \11650 );
xor \U$9750 ( \11652 , \11645 , \11651 );
and \U$9753 ( \11653 , \11577 , \11582 );
or \U$9754 ( \11654 , 1'b0 , 1'b0 , \11653 );
and \U$9755 ( \11655 , \11613 , \11619 );
and \U$9756 ( \11656 , \11619 , \11630 );
and \U$9757 ( \11657 , \11613 , \11630 );
or \U$9758 ( \11658 , \11655 , \11656 , \11657 );
xor \U$9759 ( \11659 , \11654 , \11658 );
and \U$9761 ( \11660 , \10468 , \10327 );
and \U$9762 ( \11661 , \10424 , \10325 );
nor \U$9763 ( \11662 , \11660 , \11661 );
xnor \U$9764 ( \11663 , \11662 , \10094 );
and \U$9765 ( \11664 , \10561 , \10265 );
and \U$9766 ( \11665 , \10594 , \10263 );
nor \U$9767 ( \11666 , \11664 , \11665 );
xnor \U$9768 ( \11667 , \11666 , \10291 );
xor \U$9769 ( \11668 , \11663 , \11667 );
and \U$9771 ( \11669 , \10654 , \10318 );
nor \U$9772 ( \11670 , 1'b0 , \11669 );
xnor \U$9773 ( \11671 , \11670 , 1'b0 );
xor \U$9774 ( \11672 , \11668 , \11671 );
xor \U$9775 ( \11673 , 1'b0 , \11672 );
not \U$9776 ( \11674 , \10659 );
and \U$9777 ( \11675 , \10217 , \10691 );
and \U$9778 ( \11676 , \10286 , \10689 );
nor \U$9779 ( \11677 , \11675 , \11676 );
xnor \U$9780 ( \11678 , \11677 , \10717 );
xor \U$9781 ( \11679 , \11674 , \11678 );
and \U$9782 ( \11680 , \10445 , \10392 );
and \U$9783 ( \11681 , \10313 , \10390 );
nor \U$9784 ( \11682 , \11680 , \11681 );
xnor \U$9785 ( \11683 , \11682 , \10397 );
xor \U$9786 ( \11684 , \11679 , \11683 );
xor \U$9787 ( \11685 , \11673 , \11684 );
xor \U$9789 ( \11686 , \11685 , 1'b0 );
and \U$9791 ( \11687 , \11606 , \11611 );
or \U$9793 ( \11688 , 1'b0 , \11687 , 1'b0 );
and \U$9794 ( \11689 , \11593 , \11597 );
and \U$9795 ( \11690 , \11597 , \11602 );
and \U$9796 ( \11691 , \11593 , \11602 );
or \U$9797 ( \11692 , \11689 , \11690 , \11691 );
xor \U$9798 ( \11693 , \11688 , \11692 );
xor \U$9800 ( \11694 , \11693 , 1'b0 );
xor \U$9801 ( \11695 , \11686 , \11694 );
xor \U$9802 ( \11696 , \11659 , \11695 );
xor \U$9803 ( \11697 , \11652 , \11696 );
and \U$9804 ( \11698 , \11573 , \11583 );
and \U$9805 ( \11699 , \11583 , \11632 );
and \U$9806 ( \11700 , \11573 , \11632 );
or \U$9807 ( \11701 , \11698 , \11699 , \11700 );
nor \U$9808 ( \11702 , \11697 , \11701 );
and \U$9809 ( \11703 , \11654 , \11658 );
and \U$9810 ( \11704 , \11658 , \11695 );
and \U$9811 ( \11705 , \11654 , \11695 );
or \U$9812 ( \11706 , \11703 , \11704 , \11705 );
and \U$9813 ( \11707 , \11688 , \11692 );
or \U$9816 ( \11708 , \11707 , 1'b0 , 1'b0 );
xor \U$9818 ( \11709 , \11708 , 1'b0 );
and \U$9820 ( \11710 , \11672 , \11684 );
or \U$9822 ( \11711 , 1'b0 , \11710 , 1'b0 );
xor \U$9823 ( \11712 , \11709 , \11711 );
xor \U$9824 ( \11713 , \11706 , \11712 );
and \U$9825 ( \11714 , \11647 , \11648 );
and \U$9826 ( \11715 , \11648 , \11650 );
and \U$9827 ( \11716 , \11647 , \11650 );
or \U$9828 ( \11717 , \11714 , \11715 , \11716 );
and \U$9831 ( \11718 , \11685 , \11694 );
or \U$9832 ( \11719 , 1'b0 , 1'b0 , \11718 );
xor \U$9833 ( \11720 , \11717 , \11719 );
and \U$9834 ( \11721 , \10424 , \10327 );
and \U$9835 ( \11722 , \10445 , \10325 );
nor \U$9836 ( \11723 , \11721 , \11722 );
xnor \U$9837 ( \11724 , \11723 , \10094 );
and \U$9838 ( \11725 , \10594 , \10265 );
and \U$9839 ( \11726 , \10468 , \10263 );
nor \U$9840 ( \11727 , \11725 , \11726 );
xnor \U$9841 ( \11728 , \11727 , \10291 );
xor \U$9842 ( \11729 , \11724 , \11728 );
and \U$9844 ( \11730 , \10561 , \10318 );
nor \U$9845 ( \11731 , 1'b0 , \11730 );
xnor \U$9846 ( \11732 , \11731 , 1'b0 );
xor \U$9847 ( \11733 , \11729 , \11732 );
and \U$9849 ( \11734 , \10286 , \10691 );
not \U$9850 ( \11735 , \11734 );
xnor \U$9851 ( \11736 , \11735 , \10717 );
xor \U$9852 ( \11737 , 1'b0 , \11736 );
and \U$9853 ( \11738 , \10313 , \10392 );
and \U$9854 ( \11739 , \10217 , \10390 );
nor \U$9855 ( \11740 , \11738 , \11739 );
xnor \U$9856 ( \11741 , \11740 , \10397 );
xor \U$9857 ( \11742 , \11737 , \11741 );
xor \U$9858 ( \11743 , \11733 , \11742 );
xor \U$9860 ( \11744 , \11743 , 1'b1 );
and \U$9861 ( \11745 , \11674 , \11678 );
and \U$9862 ( \11746 , \11678 , \11683 );
and \U$9863 ( \11747 , \11674 , \11683 );
or \U$9864 ( \11748 , \11745 , \11746 , \11747 );
and \U$9865 ( \11749 , \11663 , \11667 );
and \U$9866 ( \11750 , \11667 , \11671 );
and \U$9867 ( \11751 , \11663 , \11671 );
or \U$9868 ( \11752 , \11749 , \11750 , \11751 );
xor \U$9869 ( \11753 , \11748 , \11752 );
xor \U$9871 ( \11754 , \11753 , 1'b0 );
xor \U$9872 ( \11755 , \11744 , \11754 );
xor \U$9873 ( \11756 , \11720 , \11755 );
xor \U$9874 ( \11757 , \11713 , \11756 );
and \U$9875 ( \11758 , \11645 , \11651 );
and \U$9876 ( \11759 , \11651 , \11696 );
and \U$9877 ( \11760 , \11645 , \11696 );
or \U$9878 ( \11761 , \11758 , \11759 , \11760 );
nor \U$9879 ( \11762 , \11757 , \11761 );
nor \U$9880 ( \11763 , \11702 , \11762 );
and \U$9881 ( \11764 , \11717 , \11719 );
and \U$9882 ( \11765 , \11719 , \11755 );
and \U$9883 ( \11766 , \11717 , \11755 );
or \U$9884 ( \11767 , \11764 , \11765 , \11766 );
and \U$9885 ( \11768 , \11748 , \11752 );
or \U$9888 ( \11769 , \11768 , 1'b0 , 1'b0 );
xor \U$9890 ( \11770 , \11769 , 1'b0 );
and \U$9891 ( \11771 , \11733 , \11742 );
xor \U$9892 ( \11772 , \11770 , \11771 );
xor \U$9893 ( \11773 , \11767 , \11772 );
and \U$9896 ( \11774 , \11708 , \11711 );
or \U$9897 ( \11775 , 1'b0 , 1'b0 , \11774 );
and \U$9898 ( \11776 , \11743 , 1'b1 );
and \U$9899 ( \11777 , 1'b1 , \11754 );
and \U$9900 ( \11778 , \11743 , \11754 );
or \U$9901 ( \11779 , \11776 , \11777 , \11778 );
xor \U$9902 ( \11780 , \11775 , \11779 );
and \U$9904 ( \11781 , \10468 , \10265 );
and \U$9905 ( \11782 , \10424 , \10263 );
nor \U$9906 ( \11783 , \11781 , \11782 );
xnor \U$9907 ( \11784 , \11783 , \10291 );
and \U$9909 ( \11785 , \10594 , \10318 );
nor \U$9910 ( \11786 , 1'b0 , \11785 );
xnor \U$9911 ( \11787 , \11786 , 1'b0 );
xor \U$9912 ( \11788 , \11784 , \11787 );
xor \U$9914 ( \11789 , \11788 , 1'b0 );
xor \U$9915 ( \11790 , 1'b0 , \11789 );
not \U$9916 ( \11791 , \10717 );
and \U$9917 ( \11792 , \10217 , \10392 );
and \U$9918 ( \11793 , \10286 , \10390 );
nor \U$9919 ( \11794 , \11792 , \11793 );
xnor \U$9920 ( \11795 , \11794 , \10397 );
xor \U$9921 ( \11796 , \11791 , \11795 );
and \U$9922 ( \11797 , \10445 , \10327 );
and \U$9923 ( \11798 , \10313 , \10325 );
nor \U$9924 ( \11799 , \11797 , \11798 );
xnor \U$9925 ( \11800 , \11799 , \10094 );
xor \U$9926 ( \11801 , \11796 , \11800 );
xor \U$9927 ( \11802 , \11790 , \11801 );
xor \U$9929 ( \11803 , \11802 , 1'b0 );
and \U$9931 ( \11804 , \11736 , \11741 );
or \U$9933 ( \11805 , 1'b0 , \11804 , 1'b0 );
and \U$9934 ( \11806 , \11724 , \11728 );
and \U$9935 ( \11807 , \11728 , \11732 );
and \U$9936 ( \11808 , \11724 , \11732 );
or \U$9937 ( \11809 , \11806 , \11807 , \11808 );
xor \U$9938 ( \11810 , \11805 , \11809 );
xor \U$9940 ( \11811 , \11810 , 1'b0 );
xor \U$9941 ( \11812 , \11803 , \11811 );
xor \U$9942 ( \11813 , \11780 , \11812 );
xor \U$9943 ( \11814 , \11773 , \11813 );
and \U$9944 ( \11815 , \11706 , \11712 );
and \U$9945 ( \11816 , \11712 , \11756 );
and \U$9946 ( \11817 , \11706 , \11756 );
or \U$9947 ( \11818 , \11815 , \11816 , \11817 );
nor \U$9948 ( \11819 , \11814 , \11818 );
and \U$9949 ( \11820 , \11775 , \11779 );
and \U$9950 ( \11821 , \11779 , \11812 );
and \U$9951 ( \11822 , \11775 , \11812 );
or \U$9952 ( \11823 , \11820 , \11821 , \11822 );
and \U$9953 ( \11824 , \11805 , \11809 );
or \U$9956 ( \11825 , \11824 , 1'b0 , 1'b0 );
xor \U$9958 ( \11826 , \11825 , 1'b0 );
and \U$9960 ( \11827 , \11789 , \11801 );
or \U$9962 ( \11828 , 1'b0 , \11827 , 1'b0 );
xor \U$9963 ( \11829 , \11826 , \11828 );
xor \U$9964 ( \11830 , \11823 , \11829 );
and \U$9967 ( \11831 , \11769 , \11771 );
or \U$9968 ( \11832 , 1'b0 , 1'b0 , \11831 );
and \U$9971 ( \11833 , \11802 , \11811 );
or \U$9972 ( \11834 , 1'b0 , 1'b0 , \11833 );
xor \U$9973 ( \11835 , \11832 , \11834 );
xor \U$9974 ( \11836 , \10448 , \10471 );
xor \U$9976 ( \11837 , \11836 , 1'b0 );
xor \U$9978 ( \11838 , 1'b0 , \10398 );
xor \U$9979 ( \11839 , \11838 , \10402 );
xor \U$9980 ( \11840 , \11837 , \11839 );
xor \U$9982 ( \11841 , \11840 , 1'b1 );
and \U$9983 ( \11842 , \11791 , \11795 );
and \U$9984 ( \11843 , \11795 , \11800 );
and \U$9985 ( \11844 , \11791 , \11800 );
or \U$9986 ( \11845 , \11842 , \11843 , \11844 );
and \U$9987 ( \11846 , \11784 , \11787 );
or \U$9990 ( \11847 , \11846 , 1'b0 , 1'b0 );
xor \U$9991 ( \11848 , \11845 , \11847 );
xor \U$9993 ( \11849 , \11848 , 1'b0 );
xor \U$9994 ( \11850 , \11841 , \11849 );
xor \U$9995 ( \11851 , \11835 , \11850 );
xor \U$9996 ( \11852 , \11830 , \11851 );
and \U$9997 ( \11853 , \11767 , \11772 );
and \U$9998 ( \11854 , \11772 , \11813 );
and \U$9999 ( \11855 , \11767 , \11813 );
or \U$10000 ( \11856 , \11853 , \11854 , \11855 );
nor \U$10001 ( \11857 , \11852 , \11856 );
nor \U$10002 ( \11858 , \11819 , \11857 );
nand \U$10003 ( \11859 , \11763 , \11858 );
and \U$10004 ( \11860 , \11832 , \11834 );
and \U$10005 ( \11861 , \11834 , \11850 );
and \U$10006 ( \11862 , \11832 , \11850 );
or \U$10007 ( \11863 , \11860 , \11861 , \11862 );
and \U$10008 ( \11864 , \11845 , \11847 );
or \U$10011 ( \11865 , \11864 , 1'b0 , 1'b0 );
xor \U$10013 ( \11866 , \11865 , 1'b0 );
and \U$10014 ( \11867 , \11837 , \11839 );
xor \U$10015 ( \11868 , \11866 , \11867 );
xor \U$10016 ( \11869 , \11863 , \11868 );
and \U$10019 ( \11870 , \11825 , \11828 );
or \U$10020 ( \11871 , 1'b0 , 1'b0 , \11870 );
and \U$10021 ( \11872 , \11840 , 1'b1 );
and \U$10022 ( \11873 , 1'b1 , \11849 );
and \U$10023 ( \11874 , \11840 , \11849 );
or \U$10024 ( \11875 , \11872 , \11873 , \11874 );
xor \U$10025 ( \11876 , \11871 , \11875 );
xor \U$10027 ( \11877 , 1'b0 , \10480 );
xor \U$10028 ( \11878 , \11877 , \10491 );
xor \U$10030 ( \11879 , \11878 , 1'b0 );
xor \U$10031 ( \11880 , \10404 , \10473 );
xor \U$10033 ( \11881 , \11880 , 1'b0 );
xor \U$10034 ( \11882 , \11879 , \11881 );
xor \U$10035 ( \11883 , \11876 , \11882 );
xor \U$10036 ( \11884 , \11869 , \11883 );
and \U$10037 ( \11885 , \11823 , \11829 );
and \U$10038 ( \11886 , \11829 , \11851 );
and \U$10039 ( \11887 , \11823 , \11851 );
or \U$10040 ( \11888 , \11885 , \11886 , \11887 );
nor \U$10041 ( \11889 , \11884 , \11888 );
and \U$10042 ( \11890 , \11871 , \11875 );
and \U$10043 ( \11891 , \11875 , \11882 );
and \U$10044 ( \11892 , \11871 , \11882 );
or \U$10045 ( \11893 , \11890 , \11891 , \11892 );
xor \U$10047 ( \11894 , \10475 , 1'b0 );
xor \U$10048 ( \11895 , \11894 , \10493 );
xor \U$10049 ( \11896 , \11893 , \11895 );
and \U$10052 ( \11897 , \11865 , \11867 );
or \U$10053 ( \11898 , 1'b0 , 1'b0 , \11897 );
and \U$10056 ( \11899 , \11878 , \11881 );
or \U$10057 ( \11900 , 1'b0 , 1'b0 , \11899 );
xor \U$10058 ( \11901 , \11898 , \11900 );
xor \U$10059 ( \11902 , \10503 , 1'b1 );
xor \U$10060 ( \11903 , \11902 , \10510 );
xor \U$10061 ( \11904 , \11901 , \11903 );
xor \U$10062 ( \11905 , \11896 , \11904 );
and \U$10063 ( \11906 , \11863 , \11868 );
and \U$10064 ( \11907 , \11868 , \11883 );
and \U$10065 ( \11908 , \11863 , \11883 );
or \U$10066 ( \11909 , \11906 , \11907 , \11908 );
nor \U$10067 ( \11910 , \11905 , \11909 );
nor \U$10068 ( \11911 , \11889 , \11910 );
and \U$10069 ( \11912 , \11898 , \11900 );
and \U$10070 ( \11913 , \11900 , \11903 );
and \U$10071 ( \11914 , \11898 , \11903 );
or \U$10072 ( \11915 , \11912 , \11913 , \11914 );
and \U$10074 ( \11916 , \10500 , \10502 );
xor \U$10075 ( \11917 , 1'b0 , \11916 );
xor \U$10076 ( \11918 , \11915 , \11917 );
xor \U$10077 ( \11919 , \10495 , \10513 );
xor \U$10078 ( \11920 , \11919 , \10516 );
xor \U$10079 ( \11921 , \11918 , \11920 );
and \U$10080 ( \11922 , \11893 , \11895 );
and \U$10081 ( \11923 , \11895 , \11904 );
and \U$10082 ( \11924 , \11893 , \11904 );
or \U$10083 ( \11925 , \11922 , \11923 , \11924 );
nor \U$10084 ( \11926 , \11921 , \11925 );
xor \U$10086 ( \11927 , \10519 , 1'b0 );
xor \U$10087 ( \11928 , \11927 , \10521 );
and \U$10088 ( \11929 , \11915 , \11917 );
and \U$10089 ( \11930 , \11917 , \11920 );
and \U$10090 ( \11931 , \11915 , \11920 );
or \U$10091 ( \11932 , \11929 , \11930 , \11931 );
nor \U$10092 ( \11933 , \11928 , \11932 );
nor \U$10093 ( \11934 , \11926 , \11933 );
nand \U$10094 ( \11935 , \11911 , \11934 );
nor \U$10095 ( \11936 , \11859 , \11935 );
nand \U$10096 ( \11937 , \11641 , \11936 );
and \U$10097 ( \11938 , \10738 , \10537 );
and \U$10098 ( \11939 , \10759 , \10534 );
nor \U$10099 ( \11940 , \11938 , \11939 );
xnor \U$10100 ( \11941 , \11940 , \10531 );
and \U$10101 ( \11942 , \10783 , \10573 );
and \U$10102 ( \11943 , \10804 , \10571 );
nor \U$10103 ( \11944 , \11942 , \11943 );
xnor \U$10104 ( \11945 , \11944 , \10599 );
and \U$10105 ( \11946 , \11941 , \11945 );
and \U$10106 ( \11947 , \10831 , \10633 );
and \U$10107 ( \11948 , \10852 , \10631 );
nor \U$10108 ( \11949 , \11947 , \11948 );
xnor \U$10109 ( \11950 , \11949 , \10659 );
and \U$10110 ( \11951 , \11945 , \11950 );
and \U$10111 ( \11952 , \11941 , \11950 );
or \U$10112 ( \11953 , \11946 , \11951 , \11952 );
and \U$10113 ( \11954 , \10852 , \10633 );
and \U$10114 ( \11955 , \10783 , \10631 );
nor \U$10115 ( \11956 , \11954 , \11955 );
xnor \U$10116 ( \11957 , \11956 , \10659 );
and \U$10117 ( \11958 , \10875 , \10691 );
and \U$10118 ( \11959 , \10831 , \10689 );
nor \U$10119 ( \11960 , \11958 , \11959 );
xnor \U$10120 ( \11961 , \11960 , \10717 );
xor \U$10121 ( \11962 , \11957 , \11961 );
nand \U$10122 ( \11963 , \11008 , \10390 );
xnor \U$10123 ( \11964 , \11963 , \10397 );
xor \U$10124 ( \11965 , \11962 , \11964 );
and \U$10125 ( \11966 , \11953 , \11965 );
and \U$10126 ( \11967 , \10759 , \10537 );
and \U$10127 ( \11968 , \10683 , \10534 );
nor \U$10128 ( \11969 , \11967 , \11968 );
xnor \U$10129 ( \11970 , \11969 , \10531 );
xor \U$10130 ( \11971 , \10397 , \11970 );
and \U$10131 ( \11972 , \10804 , \10573 );
and \U$10132 ( \11973 , \10738 , \10571 );
nor \U$10133 ( \11974 , \11972 , \11973 );
xnor \U$10134 ( \11975 , \11974 , \10599 );
xor \U$10135 ( \11976 , \11971 , \11975 );
and \U$10136 ( \11977 , \11965 , \11976 );
and \U$10137 ( \11978 , \11953 , \11976 );
or \U$10138 ( \11979 , \11966 , \11977 , \11978 );
and \U$10139 ( \11980 , \11008 , \10392 );
and \U$10140 ( \11981 , \10875 , \10390 );
nor \U$10141 ( \11982 , \11980 , \11981 );
xnor \U$10142 ( \11983 , \11982 , \10397 );
and \U$10143 ( \11984 , \10683 , \10537 );
and \U$10144 ( \11985 , \10712 , \10534 );
nor \U$10145 ( \11986 , \11984 , \11985 );
xnor \U$10146 ( \11987 , \11986 , \10531 );
and \U$10147 ( \11988 , \10738 , \10573 );
and \U$10148 ( \11989 , \10759 , \10571 );
nor \U$10149 ( \11990 , \11988 , \11989 );
xnor \U$10150 ( \11991 , \11990 , \10599 );
xor \U$10151 ( \11992 , \11987 , \11991 );
and \U$10152 ( \11993 , \10783 , \10633 );
and \U$10153 ( \11994 , \10804 , \10631 );
nor \U$10154 ( \11995 , \11993 , \11994 );
xnor \U$10155 ( \11996 , \11995 , \10659 );
xor \U$10156 ( \11997 , \11992 , \11996 );
xor \U$10157 ( \11998 , \11983 , \11997 );
xor \U$10158 ( \11999 , \11979 , \11998 );
and \U$10159 ( \12000 , \10397 , \11970 );
and \U$10160 ( \12001 , \11970 , \11975 );
and \U$10161 ( \12002 , \10397 , \11975 );
or \U$10162 ( \12003 , \12000 , \12001 , \12002 );
and \U$10163 ( \12004 , \11957 , \11961 );
and \U$10164 ( \12005 , \11961 , \11964 );
and \U$10165 ( \12006 , \11957 , \11964 );
or \U$10166 ( \12007 , \12004 , \12005 , \12006 );
xor \U$10167 ( \12008 , \12003 , \12007 );
and \U$10168 ( \12009 , \10831 , \10691 );
and \U$10169 ( \12010 , \10852 , \10689 );
nor \U$10170 ( \12011 , \12009 , \12010 );
xnor \U$10171 ( \12012 , \12011 , \10717 );
xor \U$10172 ( \12013 , \12008 , \12012 );
xor \U$10173 ( \12014 , \11999 , \12013 );
and \U$10174 ( \12015 , \10804 , \10537 );
and \U$10175 ( \12016 , \10738 , \10534 );
nor \U$10176 ( \12017 , \12015 , \12016 );
xnor \U$10177 ( \12018 , \12017 , \10531 );
and \U$10178 ( \12019 , \10717 , \12018 );
and \U$10179 ( \12020 , \10852 , \10573 );
and \U$10180 ( \12021 , \10783 , \10571 );
nor \U$10181 ( \12022 , \12020 , \12021 );
xnor \U$10182 ( \12023 , \12022 , \10599 );
and \U$10183 ( \12024 , \12018 , \12023 );
and \U$10184 ( \12025 , \10717 , \12023 );
or \U$10185 ( \12026 , \12019 , \12024 , \12025 );
and \U$10186 ( \12027 , \10875 , \10633 );
and \U$10187 ( \12028 , \10831 , \10631 );
nor \U$10188 ( \12029 , \12027 , \12028 );
xnor \U$10189 ( \12030 , \12029 , \10659 );
nand \U$10190 ( \12031 , \11008 , \10689 );
xnor \U$10191 ( \12032 , \12031 , \10717 );
and \U$10192 ( \12033 , \12030 , \12032 );
and \U$10193 ( \12034 , \12026 , \12033 );
and \U$10194 ( \12035 , \11008 , \10691 );
and \U$10195 ( \12036 , \10875 , \10689 );
nor \U$10196 ( \12037 , \12035 , \12036 );
xnor \U$10197 ( \12038 , \12037 , \10717 );
and \U$10198 ( \12039 , \12033 , \12038 );
and \U$10199 ( \12040 , \12026 , \12038 );
or \U$10200 ( \12041 , \12034 , \12039 , \12040 );
xor \U$10201 ( \12042 , \11953 , \11965 );
xor \U$10202 ( \12043 , \12042 , \11976 );
and \U$10203 ( \12044 , \12041 , \12043 );
nor \U$10204 ( \12045 , \12014 , \12044 );
and \U$10205 ( \12046 , \11987 , \11991 );
and \U$10206 ( \12047 , \11991 , \11996 );
and \U$10207 ( \12048 , \11987 , \11996 );
or \U$10208 ( \12049 , \12046 , \12047 , \12048 );
nand \U$10209 ( \12050 , \11008 , \10325 );
xnor \U$10210 ( \12051 , \12050 , \10094 );
xor \U$10211 ( \12052 , \12049 , \12051 );
and \U$10212 ( \12053 , \10804 , \10633 );
and \U$10213 ( \12054 , \10738 , \10631 );
nor \U$10214 ( \12055 , \12053 , \12054 );
xnor \U$10215 ( \12056 , \12055 , \10659 );
and \U$10216 ( \12057 , \10852 , \10691 );
and \U$10217 ( \12058 , \10783 , \10689 );
nor \U$10218 ( \12059 , \12057 , \12058 );
xnor \U$10219 ( \12060 , \12059 , \10717 );
xor \U$10220 ( \12061 , \12056 , \12060 );
and \U$10221 ( \12062 , \10875 , \10392 );
and \U$10222 ( \12063 , \10831 , \10390 );
nor \U$10223 ( \12064 , \12062 , \12063 );
xnor \U$10224 ( \12065 , \12064 , \10397 );
xor \U$10225 ( \12066 , \12061 , \12065 );
xor \U$10226 ( \12067 , \12052 , \12066 );
and \U$10227 ( \12068 , \12003 , \12007 );
and \U$10228 ( \12069 , \12007 , \12012 );
and \U$10229 ( \12070 , \12003 , \12012 );
or \U$10230 ( \12071 , \12068 , \12069 , \12070 );
and \U$10231 ( \12072 , \11983 , \11997 );
xor \U$10232 ( \12073 , \12071 , \12072 );
and \U$10233 ( \12074 , \10712 , \10537 );
and \U$10234 ( \12075 , \10621 , \10534 );
nor \U$10235 ( \12076 , \12074 , \12075 );
xnor \U$10236 ( \12077 , \12076 , \10531 );
xor \U$10237 ( \12078 , \10094 , \12077 );
and \U$10238 ( \12079 , \10759 , \10573 );
and \U$10239 ( \12080 , \10683 , \10571 );
nor \U$10240 ( \12081 , \12079 , \12080 );
xnor \U$10241 ( \12082 , \12081 , \10599 );
xor \U$10242 ( \12083 , \12078 , \12082 );
xor \U$10243 ( \12084 , \12073 , \12083 );
xor \U$10244 ( \12085 , \12067 , \12084 );
and \U$10245 ( \12086 , \11979 , \11998 );
and \U$10246 ( \12087 , \11998 , \12013 );
and \U$10247 ( \12088 , \11979 , \12013 );
or \U$10248 ( \12089 , \12086 , \12087 , \12088 );
nor \U$10249 ( \12090 , \12085 , \12089 );
nor \U$10250 ( \12091 , \12045 , \12090 );
and \U$10251 ( \12092 , \12071 , \12072 );
and \U$10252 ( \12093 , \12072 , \12083 );
and \U$10253 ( \12094 , \12071 , \12083 );
or \U$10254 ( \12095 , \12092 , \12093 , \12094 );
and \U$10255 ( \12096 , \12049 , \12051 );
and \U$10256 ( \12097 , \12051 , \12066 );
and \U$10257 ( \12098 , \12049 , \12066 );
or \U$10258 ( \12099 , \12096 , \12097 , \12098 );
and \U$10259 ( \12100 , \10621 , \10537 );
and \U$10260 ( \12101 , \10654 , \10534 );
nor \U$10261 ( \12102 , \12100 , \12101 );
xnor \U$10262 ( \12103 , \12102 , \10531 );
and \U$10263 ( \12104 , \10683 , \10573 );
and \U$10264 ( \12105 , \10712 , \10571 );
nor \U$10265 ( \12106 , \12104 , \12105 );
xnor \U$10266 ( \12107 , \12106 , \10599 );
xor \U$10267 ( \12108 , \12103 , \12107 );
and \U$10268 ( \12109 , \10738 , \10633 );
and \U$10269 ( \12110 , \10759 , \10631 );
nor \U$10270 ( \12111 , \12109 , \12110 );
xnor \U$10271 ( \12112 , \12111 , \10659 );
xor \U$10272 ( \12113 , \12108 , \12112 );
xor \U$10273 ( \12114 , \12099 , \12113 );
and \U$10274 ( \12115 , \10094 , \12077 );
and \U$10275 ( \12116 , \12077 , \12082 );
and \U$10276 ( \12117 , \10094 , \12082 );
or \U$10277 ( \12118 , \12115 , \12116 , \12117 );
and \U$10278 ( \12119 , \12056 , \12060 );
and \U$10279 ( \12120 , \12060 , \12065 );
and \U$10280 ( \12121 , \12056 , \12065 );
or \U$10281 ( \12122 , \12119 , \12120 , \12121 );
xor \U$10282 ( \12123 , \12118 , \12122 );
and \U$10283 ( \12124 , \10783 , \10691 );
and \U$10284 ( \12125 , \10804 , \10689 );
nor \U$10285 ( \12126 , \12124 , \12125 );
xnor \U$10286 ( \12127 , \12126 , \10717 );
and \U$10287 ( \12128 , \10831 , \10392 );
and \U$10288 ( \12129 , \10852 , \10390 );
nor \U$10289 ( \12130 , \12128 , \12129 );
xnor \U$10290 ( \12131 , \12130 , \10397 );
xor \U$10291 ( \12132 , \12127 , \12131 );
and \U$10292 ( \12133 , \11008 , \10327 );
and \U$10293 ( \12134 , \10875 , \10325 );
nor \U$10294 ( \12135 , \12133 , \12134 );
xnor \U$10295 ( \12136 , \12135 , \10094 );
xor \U$10296 ( \12137 , \12132 , \12136 );
xor \U$10297 ( \12138 , \12123 , \12137 );
xor \U$10298 ( \12139 , \12114 , \12138 );
xor \U$10299 ( \12140 , \12095 , \12139 );
and \U$10300 ( \12141 , \12067 , \12084 );
nor \U$10301 ( \12142 , \12140 , \12141 );
and \U$10302 ( \12143 , \12099 , \12113 );
and \U$10303 ( \12144 , \12113 , \12138 );
and \U$10304 ( \12145 , \12099 , \12138 );
or \U$10305 ( \12146 , \12143 , \12144 , \12145 );
and \U$10306 ( \12147 , \12118 , \12122 );
and \U$10307 ( \12148 , \12122 , \12137 );
and \U$10308 ( \12149 , \12118 , \12137 );
or \U$10309 ( \12150 , \12147 , \12148 , \12149 );
nand \U$10310 ( \12151 , \11008 , \10263 );
xnor \U$10311 ( \12152 , \12151 , \10291 );
and \U$10312 ( \12153 , \10759 , \10633 );
and \U$10313 ( \12154 , \10683 , \10631 );
nor \U$10314 ( \12155 , \12153 , \12154 );
xnor \U$10315 ( \12156 , \12155 , \10659 );
and \U$10316 ( \12157 , \10804 , \10691 );
and \U$10317 ( \12158 , \10738 , \10689 );
nor \U$10318 ( \12159 , \12157 , \12158 );
xnor \U$10319 ( \12160 , \12159 , \10717 );
xor \U$10320 ( \12161 , \12156 , \12160 );
and \U$10321 ( \12162 , \10852 , \10392 );
and \U$10322 ( \12163 , \10783 , \10390 );
nor \U$10323 ( \12164 , \12162 , \12163 );
xnor \U$10324 ( \12165 , \12164 , \10397 );
xor \U$10325 ( \12166 , \12161 , \12165 );
xor \U$10326 ( \12167 , \12152 , \12166 );
and \U$10327 ( \12168 , \10654 , \10537 );
and \U$10328 ( \12169 , \10561 , \10534 );
nor \U$10329 ( \12170 , \12168 , \12169 );
xnor \U$10330 ( \12171 , \12170 , \10531 );
xor \U$10331 ( \12172 , \10291 , \12171 );
and \U$10332 ( \12173 , \10712 , \10573 );
and \U$10333 ( \12174 , \10621 , \10571 );
nor \U$10334 ( \12175 , \12173 , \12174 );
xnor \U$10335 ( \12176 , \12175 , \10599 );
xor \U$10336 ( \12177 , \12172 , \12176 );
xor \U$10337 ( \12178 , \12167 , \12177 );
xor \U$10338 ( \12179 , \12150 , \12178 );
and \U$10339 ( \12180 , \12103 , \12107 );
and \U$10340 ( \12181 , \12107 , \12112 );
and \U$10341 ( \12182 , \12103 , \12112 );
or \U$10342 ( \12183 , \12180 , \12181 , \12182 );
and \U$10343 ( \12184 , \12127 , \12131 );
and \U$10344 ( \12185 , \12131 , \12136 );
and \U$10345 ( \12186 , \12127 , \12136 );
or \U$10346 ( \12187 , \12184 , \12185 , \12186 );
xor \U$10347 ( \12188 , \12183 , \12187 );
and \U$10348 ( \12189 , \10875 , \10327 );
and \U$10349 ( \12190 , \10831 , \10325 );
nor \U$10350 ( \12191 , \12189 , \12190 );
xnor \U$10351 ( \12192 , \12191 , \10094 );
xor \U$10352 ( \12193 , \12188 , \12192 );
xor \U$10353 ( \12194 , \12179 , \12193 );
xor \U$10354 ( \12195 , \12146 , \12194 );
and \U$10355 ( \12196 , \12095 , \12139 );
nor \U$10356 ( \12197 , \12195 , \12196 );
nor \U$10357 ( \12198 , \12142 , \12197 );
nand \U$10358 ( \12199 , \12091 , \12198 );
and \U$10359 ( \12200 , \12150 , \12178 );
and \U$10360 ( \12201 , \12178 , \12193 );
and \U$10361 ( \12202 , \12150 , \12193 );
or \U$10362 ( \12203 , \12200 , \12201 , \12202 );
xor \U$10363 ( \12204 , \11063 , \11067 );
xor \U$10364 ( \12205 , \12204 , \11072 );
and \U$10365 ( \12206 , \10291 , \12171 );
and \U$10366 ( \12207 , \12171 , \12176 );
and \U$10367 ( \12208 , \10291 , \12176 );
or \U$10368 ( \12209 , \12206 , \12207 , \12208 );
and \U$10369 ( \12210 , \12156 , \12160 );
and \U$10370 ( \12211 , \12160 , \12165 );
and \U$10371 ( \12212 , \12156 , \12165 );
or \U$10372 ( \12213 , \12210 , \12211 , \12212 );
xor \U$10373 ( \12214 , \12209 , \12213 );
and \U$10374 ( \12215 , \11008 , \10265 );
and \U$10375 ( \12216 , \10875 , \10263 );
nor \U$10376 ( \12217 , \12215 , \12216 );
xnor \U$10377 ( \12218 , \12217 , \10291 );
xor \U$10378 ( \12219 , \12214 , \12218 );
xor \U$10379 ( \12220 , \12205 , \12219 );
xor \U$10380 ( \12221 , \12203 , \12220 );
and \U$10381 ( \12222 , \12183 , \12187 );
and \U$10382 ( \12223 , \12187 , \12192 );
and \U$10383 ( \12224 , \12183 , \12192 );
or \U$10384 ( \12225 , \12222 , \12223 , \12224 );
and \U$10385 ( \12226 , \12152 , \12166 );
and \U$10386 ( \12227 , \12166 , \12177 );
and \U$10387 ( \12228 , \12152 , \12177 );
or \U$10388 ( \12229 , \12226 , \12227 , \12228 );
xor \U$10389 ( \12230 , \12225 , \12229 );
xor \U$10390 ( \12231 , \11079 , \11083 );
xor \U$10391 ( \12232 , \12231 , \11088 );
xor \U$10392 ( \12233 , \12230 , \12232 );
xor \U$10393 ( \12234 , \12221 , \12233 );
and \U$10394 ( \12235 , \12146 , \12194 );
nor \U$10395 ( \12236 , \12234 , \12235 );
and \U$10396 ( \12237 , \12225 , \12229 );
and \U$10397 ( \12238 , \12229 , \12232 );
and \U$10398 ( \12239 , \12225 , \12232 );
or \U$10399 ( \12240 , \12237 , \12238 , \12239 );
and \U$10400 ( \12241 , \12205 , \12219 );
xor \U$10401 ( \12242 , \12240 , \12241 );
and \U$10402 ( \12243 , \12209 , \12213 );
and \U$10403 ( \12244 , \12213 , \12218 );
and \U$10404 ( \12245 , \12209 , \12218 );
or \U$10405 ( \12246 , \12243 , \12244 , \12245 );
xor \U$10406 ( \12247 , \11099 , \11101 );
xor \U$10407 ( \12248 , \12246 , \12247 );
xor \U$10408 ( \12249 , \11075 , \11091 );
xor \U$10409 ( \12250 , \12249 , \11094 );
xor \U$10410 ( \12251 , \12248 , \12250 );
xor \U$10411 ( \12252 , \12242 , \12251 );
and \U$10412 ( \12253 , \12203 , \12220 );
and \U$10413 ( \12254 , \12220 , \12233 );
and \U$10414 ( \12255 , \12203 , \12233 );
or \U$10415 ( \12256 , \12253 , \12254 , \12255 );
nor \U$10416 ( \12257 , \12252 , \12256 );
nor \U$10417 ( \12258 , \12236 , \12257 );
and \U$10418 ( \12259 , \12246 , \12247 );
and \U$10419 ( \12260 , \12247 , \12250 );
and \U$10420 ( \12261 , \12246 , \12250 );
or \U$10421 ( \12262 , \12259 , \12260 , \12261 );
xor \U$10422 ( \12263 , \10962 , \10978 );
xor \U$10423 ( \12264 , \12263 , \11013 );
xor \U$10424 ( \12265 , \12262 , \12264 );
xor \U$10425 ( \12266 , \11097 , \11102 );
xor \U$10426 ( \12267 , \12266 , \11105 );
xor \U$10427 ( \12268 , \12265 , \12267 );
and \U$10428 ( \12269 , \12240 , \12241 );
and \U$10429 ( \12270 , \12241 , \12251 );
and \U$10430 ( \12271 , \12240 , \12251 );
or \U$10431 ( \12272 , \12269 , \12270 , \12271 );
nor \U$10432 ( \12273 , \12268 , \12272 );
xor \U$10433 ( \12274 , \11108 , \11109 );
xor \U$10434 ( \12275 , \12274 , \11112 );
and \U$10435 ( \12276 , \12262 , \12264 );
and \U$10436 ( \12277 , \12264 , \12267 );
and \U$10437 ( \12278 , \12262 , \12267 );
or \U$10438 ( \12279 , \12276 , \12277 , \12278 );
nor \U$10439 ( \12280 , \12275 , \12279 );
nor \U$10440 ( \12281 , \12273 , \12280 );
nand \U$10441 ( \12282 , \12258 , \12281 );
nor \U$10442 ( \12283 , \12199 , \12282 );
and \U$10443 ( \12284 , \10852 , \10537 );
and \U$10444 ( \12285 , \10783 , \10534 );
nor \U$10445 ( \12286 , \12284 , \12285 );
xnor \U$10446 ( \12287 , \12286 , \10531 );
and \U$10447 ( \12288 , \10659 , \12287 );
and \U$10448 ( \12289 , \10875 , \10573 );
and \U$10449 ( \12290 , \10831 , \10571 );
nor \U$10450 ( \12291 , \12289 , \12290 );
xnor \U$10451 ( \12292 , \12291 , \10599 );
and \U$10452 ( \12293 , \12287 , \12292 );
and \U$10453 ( \12294 , \10659 , \12292 );
or \U$10454 ( \12295 , \12288 , \12293 , \12294 );
and \U$10455 ( \12296 , \10783 , \10537 );
and \U$10456 ( \12297 , \10804 , \10534 );
nor \U$10457 ( \12298 , \12296 , \12297 );
xnor \U$10458 ( \12299 , \12298 , \10531 );
and \U$10459 ( \12300 , \10831 , \10573 );
and \U$10460 ( \12301 , \10852 , \10571 );
nor \U$10461 ( \12302 , \12300 , \12301 );
xnor \U$10462 ( \12303 , \12302 , \10599 );
xor \U$10463 ( \12304 , \12299 , \12303 );
and \U$10464 ( \12305 , \11008 , \10633 );
and \U$10465 ( \12306 , \10875 , \10631 );
nor \U$10466 ( \12307 , \12305 , \12306 );
xnor \U$10467 ( \12308 , \12307 , \10659 );
xor \U$10468 ( \12309 , \12304 , \12308 );
xor \U$10469 ( \12310 , \12295 , \12309 );
nand \U$10470 ( \12311 , \11008 , \10631 );
xnor \U$10471 ( \12312 , \12311 , \10659 );
xor \U$10472 ( \12313 , \10659 , \12287 );
xor \U$10473 ( \12314 , \12313 , \12292 );
and \U$10474 ( \12315 , \12312 , \12314 );
nor \U$10475 ( \12316 , \12310 , \12315 );
and \U$10476 ( \12317 , \12299 , \12303 );
and \U$10477 ( \12318 , \12303 , \12308 );
and \U$10478 ( \12319 , \12299 , \12308 );
or \U$10479 ( \12320 , \12317 , \12318 , \12319 );
xor \U$10480 ( \12321 , \12030 , \12032 );
xor \U$10481 ( \12322 , \12320 , \12321 );
xor \U$10482 ( \12323 , \10717 , \12018 );
xor \U$10483 ( \12324 , \12323 , \12023 );
xor \U$10484 ( \12325 , \12322 , \12324 );
and \U$10485 ( \12326 , \12295 , \12309 );
nor \U$10486 ( \12327 , \12325 , \12326 );
nor \U$10487 ( \12328 , \12316 , \12327 );
xor \U$10488 ( \12329 , \11941 , \11945 );
xor \U$10489 ( \12330 , \12329 , \11950 );
xor \U$10490 ( \12331 , \12026 , \12033 );
xor \U$10491 ( \12332 , \12331 , \12038 );
xor \U$10492 ( \12333 , \12330 , \12332 );
and \U$10493 ( \12334 , \12320 , \12321 );
and \U$10494 ( \12335 , \12321 , \12324 );
and \U$10495 ( \12336 , \12320 , \12324 );
or \U$10496 ( \12337 , \12334 , \12335 , \12336 );
nor \U$10497 ( \12338 , \12333 , \12337 );
xor \U$10498 ( \12339 , \12041 , \12043 );
and \U$10499 ( \12340 , \12330 , \12332 );
nor \U$10500 ( \12341 , \12339 , \12340 );
nor \U$10501 ( \12342 , \12338 , \12341 );
nand \U$10502 ( \12343 , \12328 , \12342 );
and \U$10503 ( \12344 , \10831 , \10537 );
and \U$10504 ( \12345 , \10852 , \10534 );
nor \U$10505 ( \12346 , \12344 , \12345 );
xnor \U$10506 ( \12347 , \12346 , \10531 );
and \U$10507 ( \12348 , \11008 , \10573 );
and \U$10508 ( \12349 , \10875 , \10571 );
nor \U$10509 ( \12350 , \12348 , \12349 );
xnor \U$10510 ( \12351 , \12350 , \10599 );
xor \U$10511 ( \12352 , \12347 , \12351 );
and \U$10512 ( \12353 , \10875 , \10537 );
and \U$10513 ( \12354 , \10831 , \10534 );
nor \U$10514 ( \12355 , \12353 , \12354 );
xnor \U$10515 ( \12356 , \12355 , \10531 );
and \U$10516 ( \12357 , \12356 , \10599 );
nor \U$10517 ( \12358 , \12352 , \12357 );
xor \U$10518 ( \12359 , \12312 , \12314 );
and \U$10519 ( \12360 , \12347 , \12351 );
nor \U$10520 ( \12361 , \12359 , \12360 );
nor \U$10521 ( \12362 , \12358 , \12361 );
xor \U$10522 ( \12363 , \12356 , \10599 );
nand \U$10523 ( \12364 , \11008 , \10571 );
xnor \U$10524 ( \12365 , \12364 , \10599 );
nor \U$10525 ( \12366 , \12363 , \12365 );
and \U$10526 ( \12367 , \11008 , \10537 );
and \U$10527 ( \12368 , \10875 , \10534 );
nor \U$10528 ( \12369 , \12367 , \12368 );
xnor \U$10529 ( \12370 , \12369 , \10531 );
nand \U$10530 ( \12371 , \11008 , \10534 );
xnor \U$10531 ( \12372 , \12371 , \10531 );
and \U$10532 ( \12373 , \12372 , \10531 );
nand \U$10533 ( \12374 , \12370 , \12373 );
or \U$10534 ( \12375 , \12366 , \12374 );
nand \U$10535 ( \12376 , \12363 , \12365 );
nand \U$10536 ( \12377 , \12375 , \12376 );
and \U$10537 ( \12378 , \12362 , \12377 );
nand \U$10538 ( \12379 , \12352 , \12357 );
or \U$10539 ( \12380 , \12361 , \12379 );
nand \U$10540 ( \12381 , \12359 , \12360 );
nand \U$10541 ( \12382 , \12380 , \12381 );
nor \U$10542 ( \12383 , \12378 , \12382 );
or \U$10543 ( \12384 , \12343 , \12383 );
nand \U$10544 ( \12385 , \12310 , \12315 );
or \U$10545 ( \12386 , \12327 , \12385 );
nand \U$10546 ( \12387 , \12325 , \12326 );
nand \U$10547 ( \12388 , \12386 , \12387 );
and \U$10548 ( \12389 , \12342 , \12388 );
nand \U$10549 ( \12390 , \12333 , \12337 );
or \U$10550 ( \12391 , \12341 , \12390 );
nand \U$10551 ( \12392 , \12339 , \12340 );
nand \U$10552 ( \12393 , \12391 , \12392 );
nor \U$10553 ( \12394 , \12389 , \12393 );
nand \U$10554 ( \12395 , \12384 , \12394 );
and \U$10555 ( \12396 , \12283 , \12395 );
nand \U$10556 ( \12397 , \12014 , \12044 );
or \U$10557 ( \12398 , \12090 , \12397 );
nand \U$10558 ( \12399 , \12085 , \12089 );
nand \U$10559 ( \12400 , \12398 , \12399 );
and \U$10560 ( \12401 , \12198 , \12400 );
nand \U$10561 ( \12402 , \12140 , \12141 );
or \U$10562 ( \12403 , \12197 , \12402 );
nand \U$10563 ( \12404 , \12195 , \12196 );
nand \U$10564 ( \12405 , \12403 , \12404 );
nor \U$10565 ( \12406 , \12401 , \12405 );
or \U$10566 ( \12407 , \12282 , \12406 );
nand \U$10567 ( \12408 , \12234 , \12235 );
or \U$10568 ( \12409 , \12257 , \12408 );
nand \U$10569 ( \12410 , \12252 , \12256 );
nand \U$10570 ( \12411 , \12409 , \12410 );
and \U$10571 ( \12412 , \12281 , \12411 );
nand \U$10572 ( \12413 , \12268 , \12272 );
or \U$10573 ( \12414 , \12280 , \12413 );
nand \U$10574 ( \12415 , \12275 , \12279 );
nand \U$10575 ( \12416 , \12414 , \12415 );
nor \U$10576 ( \12417 , \12412 , \12416 );
nand \U$10577 ( \12418 , \12407 , \12417 );
nor \U$10578 ( \12419 , \12396 , \12418 );
or \U$10579 ( \12420 , \11937 , \12419 );
nand \U$10580 ( \12421 , \11059 , \11115 );
or \U$10581 ( \12422 , \11191 , \12421 );
nand \U$10582 ( \12423 , \11189 , \11190 );
nand \U$10583 ( \12424 , \12422 , \12423 );
and \U$10584 ( \12425 , \11344 , \12424 );
nand \U$10585 ( \12426 , \11266 , \11267 );
or \U$10586 ( \12427 , \11343 , \12426 );
nand \U$10587 ( \12428 , \11338 , \11342 );
nand \U$10588 ( \12429 , \12427 , \12428 );
nor \U$10589 ( \12430 , \12425 , \12429 );
or \U$10590 ( \12431 , \11640 , \12430 );
nand \U$10591 ( \12432 , \11415 , \11419 );
or \U$10592 ( \12433 , \11496 , \12432 );
nand \U$10593 ( \12434 , \11491 , \11495 );
nand \U$10594 ( \12435 , \12433 , \12434 );
and \U$10595 ( \12436 , \11639 , \12435 );
nand \U$10596 ( \12437 , \11564 , \11568 );
or \U$10597 ( \12438 , \11638 , \12437 );
nand \U$10598 ( \12439 , \11633 , \11637 );
nand \U$10599 ( \12440 , \12438 , \12439 );
nor \U$10600 ( \12441 , \12436 , \12440 );
nand \U$10601 ( \12442 , \12431 , \12441 );
and \U$10602 ( \12443 , \11936 , \12442 );
nand \U$10603 ( \12444 , \11697 , \11701 );
or \U$10604 ( \12445 , \11762 , \12444 );
nand \U$10605 ( \12446 , \11757 , \11761 );
nand \U$10606 ( \12447 , \12445 , \12446 );
and \U$10607 ( \12448 , \11858 , \12447 );
nand \U$10608 ( \12449 , \11814 , \11818 );
or \U$10609 ( \12450 , \11857 , \12449 );
nand \U$10610 ( \12451 , \11852 , \11856 );
nand \U$10611 ( \12452 , \12450 , \12451 );
nor \U$10612 ( \12453 , \12448 , \12452 );
or \U$10613 ( \12454 , \11935 , \12453 );
nand \U$10614 ( \12455 , \11884 , \11888 );
or \U$10615 ( \12456 , \11910 , \12455 );
nand \U$10616 ( \12457 , \11905 , \11909 );
nand \U$10617 ( \12458 , \12456 , \12457 );
and \U$10618 ( \12459 , \11934 , \12458 );
nand \U$10619 ( \12460 , \11921 , \11925 );
or \U$10620 ( \12461 , \11933 , \12460 );
nand \U$10621 ( \12462 , \11928 , \11932 );
nand \U$10622 ( \12463 , \12461 , \12462 );
nor \U$10623 ( \12464 , \12459 , \12463 );
nand \U$10624 ( \12465 , \12454 , \12464 );
nor \U$10625 ( \12466 , \12443 , \12465 );
nand \U$10626 ( \12467 , \12420 , \12466 );
not \U$10627 ( \12468 , \12467 );
xor \U$10628 ( \12469 , \10527 , \12468 );
buf g4b72_GF_PartitionCandidate( \12470_nG4b72 , \12469 );
buf \U$10633 ( \12471 , RI995f080_2);
buf \U$10634 ( \12472 , RI995f008_3);
buf \U$10635 ( \12473 , RI995ef90_4);
buf \U$10636 ( \12474 , RI995ef18_5);
buf \U$10637 ( \12475 , RI995eea0_6);
buf \U$10638 ( \12476 , RI995ee28_7);
buf \U$10639 ( \12477 , RI995edb0_8);
buf \U$10640 ( \12478 , RI995ed38_9);
buf \U$10641 ( \12479 , RI995ecc0_10);
buf \U$10642 ( \12480 , RI995ec48_11);
buf \U$10643 ( \12481 , RI995ebd0_12);
and \U$10644 ( \12482 , \12480 , \12481 );
and \U$10645 ( \12483 , \12479 , \12482 );
and \U$10646 ( \12484 , \12478 , \12483 );
and \U$10647 ( \12485 , \12477 , \12484 );
and \U$10648 ( \12486 , \12476 , \12485 );
and \U$10649 ( \12487 , \12475 , \12486 );
and \U$10650 ( \12488 , \12474 , \12487 );
and \U$10651 ( \12489 , \12473 , \12488 );
and \U$10652 ( \12490 , \12472 , \12489 );
xor \U$10653 ( \12491 , \12471 , \12490 );
buf \U$10654 ( \12492 , \12491 );
buf \U$10655 ( \12493 , \12492 );
buf \U$10656 ( \12494 , RI9921d48_600);
buf \U$10657 ( \12495 , RI9921f28_596);
buf \U$10658 ( \12496 , RI9921fa0_595);
buf \U$10659 ( \12497 , RI9922018_594);
buf \U$10660 ( \12498 , RI9922090_593);
buf \U$10661 ( \12499 , RI9922108_592);
buf \U$10662 ( \12500 , RI9922180_591);
buf \U$10663 ( \12501 , RI99221f8_590);
buf \U$10664 ( \12502 , RI9922270_589);
buf \U$10665 ( \12503 , RI99222e8_588);
buf \U$10666 ( \12504 , RI9921d48_600);
buf \U$10667 ( \12505 , RI9921dc0_599);
buf \U$10668 ( \12506 , RI9921e38_598);
buf \U$10669 ( \12507 , RI9921eb0_597);
and \U$10670 ( \12508 , \12504 , \12505 , \12506 , \12507 );
nor \U$10671 ( \12509 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12508 );
buf \U$10672 ( \12510 , \12509 );
buf \U$10673 ( \12511 , \12510 );
xor \U$10674 ( \12512 , \12494 , \12511 );
buf \U$10675 ( \12513 , \12512 );
buf \U$10676 ( \12514 , RI9921dc0_599);
and \U$10677 ( \12515 , \12494 , \12511 );
xor \U$10678 ( \12516 , \12514 , \12515 );
buf \U$10679 ( \12517 , \12516 );
buf \U$10680 ( \12518 , RI9921e38_598);
and \U$10681 ( \12519 , \12514 , \12515 );
xor \U$10682 ( \12520 , \12518 , \12519 );
buf \U$10683 ( \12521 , \12520 );
buf \U$10684 ( \12522 , RI9921eb0_597);
and \U$10685 ( \12523 , \12518 , \12519 );
xor \U$10686 ( \12524 , \12522 , \12523 );
buf \U$10687 ( \12525 , \12524 );
buf \U$10688 ( \12526 , RI9921f28_596);
and \U$10689 ( \12527 , \12522 , \12523 );
xor \U$10690 ( \12528 , \12526 , \12527 );
buf \U$10691 ( \12529 , \12528 );
not \U$10692 ( \12530 , \12529 );
buf \U$10693 ( \12531 , RI9921fa0_595);
and \U$10694 ( \12532 , \12526 , \12527 );
xor \U$10695 ( \12533 , \12531 , \12532 );
buf \U$10696 ( \12534 , \12533 );
buf \U$10697 ( \12535 , RI9922018_594);
and \U$10698 ( \12536 , \12531 , \12532 );
xor \U$10699 ( \12537 , \12535 , \12536 );
buf \U$10700 ( \12538 , \12537 );
buf \U$10701 ( \12539 , RI9922090_593);
and \U$10702 ( \12540 , \12535 , \12536 );
xor \U$10703 ( \12541 , \12539 , \12540 );
buf \U$10704 ( \12542 , \12541 );
buf \U$10705 ( \12543 , RI9922108_592);
and \U$10706 ( \12544 , \12539 , \12540 );
xor \U$10707 ( \12545 , \12543 , \12544 );
buf \U$10708 ( \12546 , \12545 );
buf \U$10709 ( \12547 , RI9922180_591);
and \U$10710 ( \12548 , \12543 , \12544 );
xor \U$10711 ( \12549 , \12547 , \12548 );
buf \U$10712 ( \12550 , \12549 );
buf \U$10713 ( \12551 , RI99221f8_590);
and \U$10714 ( \12552 , \12547 , \12548 );
xor \U$10715 ( \12553 , \12551 , \12552 );
buf \U$10716 ( \12554 , \12553 );
buf \U$10717 ( \12555 , RI9922270_589);
and \U$10718 ( \12556 , \12551 , \12552 );
xor \U$10719 ( \12557 , \12555 , \12556 );
buf \U$10720 ( \12558 , \12557 );
buf \U$10721 ( \12559 , RI99222e8_588);
and \U$10722 ( \12560 , \12555 , \12556 );
xor \U$10723 ( \12561 , \12559 , \12560 );
buf \U$10724 ( \12562 , \12561 );
nor \U$10725 ( \12563 , \12513 , \12517 , \12521 , \12525 , \12530 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10726 ( \12564 , RI995e450_236, \12563 );
not \U$10727 ( \12565 , \12513 );
not \U$10728 ( \12566 , \12517 );
not \U$10729 ( \12567 , \12521 );
not \U$10730 ( \12568 , \12525 );
nor \U$10731 ( \12569 , \12565 , \12566 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10732 ( \12570 , RI9967078_223, \12569 );
nor \U$10733 ( \12571 , \12513 , \12566 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10734 ( \12572 , RI9967690_210, \12571 );
nor \U$10735 ( \12573 , \12565 , \12517 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10736 ( \12574 , RI890fba0_197, \12573 );
nor \U$10737 ( \12575 , \12513 , \12517 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10738 ( \12576 , RI8918b88_184, \12575 );
nor \U$10739 ( \12577 , \12565 , \12566 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10740 ( \12578 , RI89253b0_171, \12577 );
nor \U$10741 ( \12579 , \12513 , \12566 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10742 ( \12580 , RI8930dc8_158, \12579 );
nor \U$10743 ( \12581 , \12565 , \12517 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10744 ( \12582 , RI8939db0_145, \12581 );
nor \U$10745 ( \12583 , \12513 , \12517 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10746 ( \12584 , RI89465d8_132, \12583 );
nor \U$10747 ( \12585 , \12565 , \12566 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10748 ( \12586 , RI89ec640_119, \12585 );
nor \U$10749 ( \12587 , \12513 , \12566 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10750 ( \12588 , RI9776f80_106, \12587 );
nor \U$10751 ( \12589 , \12565 , \12517 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10752 ( \12590 , RI9808480_93, \12589 );
nor \U$10753 ( \12591 , \12513 , \12517 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10754 ( \12592 , RI9808a98_80, \12591 );
nor \U$10755 ( \12593 , \12565 , \12566 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10756 ( \12594 , RI9819730_67, \12593 );
nor \U$10757 ( \12595 , \12513 , \12566 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10758 ( \12596 , RI98abc38_54, \12595 );
nor \U$10759 ( \12597 , \12565 , \12517 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10760 ( \12598 , RI98bc8d0_41, \12597 );
nor \U$10761 ( \12599 , \12513 , \12517 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$10762 ( \12600 , RI994ddd0_28, \12599 );
or \U$10763 ( \12601 , \12564 , \12570 , \12572 , \12574 , \12576 , \12578 , \12580 , \12582 , \12584 , \12586 , \12588 , \12590 , \12592 , \12594 , \12596 , \12598 , \12600 );
buf \U$10764 ( \12602 , \12534 );
buf \U$10765 ( \12603 , \12538 );
buf \U$10766 ( \12604 , \12542 );
buf \U$10767 ( \12605 , \12546 );
buf \U$10768 ( \12606 , \12550 );
buf \U$10769 ( \12607 , \12554 );
buf \U$10770 ( \12608 , \12558 );
buf \U$10771 ( \12609 , \12562 );
buf \U$10772 ( \12610 , \12529 );
buf \U$10773 ( \12611 , \12513 );
buf \U$10774 ( \12612 , \12517 );
buf \U$10775 ( \12613 , \12521 );
buf \U$10776 ( \12614 , \12525 );
or \U$10777 ( \12615 , \12611 , \12612 , \12613 , \12614 );
and \U$10778 ( \12616 , \12610 , \12615 );
or \U$10779 ( \12617 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12616 );
buf \U$10780 ( \12618 , \12617 );
_DC g3b20 ( \12619_nG3b20 , \12601 , \12618 );
buf \U$10781 ( \12620 , \12619_nG3b20 );
not \U$10782 ( \12621 , \12620 );
xor \U$10783 ( \12622 , \12493 , \12621 );
xor \U$10784 ( \12623 , \12472 , \12489 );
buf \U$10785 ( \12624 , \12623 );
buf \U$10786 ( \12625 , \12624 );
and \U$10787 ( \12626 , RI995e3d8_237, \12563 );
and \U$10788 ( \12627 , RI99669e8_224, \12569 );
and \U$10789 ( \12628 , RI9967618_211, \12571 );
and \U$10790 ( \12629 , RI890fb28_198, \12573 );
and \U$10791 ( \12630 , RI8918b10_185, \12575 );
and \U$10792 ( \12631 , RI8925338_172, \12577 );
and \U$10793 ( \12632 , RI8930d50_159, \12579 );
and \U$10794 ( \12633 , RI8939d38_146, \12581 );
and \U$10795 ( \12634 , RI8946560_133, \12583 );
and \U$10796 ( \12635 , RI89ec5c8_120, \12585 );
and \U$10797 ( \12636 , RI9776f08_107, \12587 );
and \U$10798 ( \12637 , RI9808408_94, \12589 );
and \U$10799 ( \12638 , RI9808a20_81, \12591 );
and \U$10800 ( \12639 , RI98196b8_68, \12593 );
and \U$10801 ( \12640 , RI98abbc0_55, \12595 );
and \U$10802 ( \12641 , RI98bc858_42, \12597 );
and \U$10803 ( \12642 , RI994dd58_29, \12599 );
or \U$10804 ( \12643 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 );
_DC g3afc ( \12644_nG3afc , \12643 , \12618 );
buf \U$10805 ( \12645 , \12644_nG3afc );
not \U$10806 ( \12646 , \12645 );
and \U$10807 ( \12647 , \12625 , \12646 );
xor \U$10808 ( \12648 , \12473 , \12488 );
buf \U$10809 ( \12649 , \12648 );
buf \U$10810 ( \12650 , \12649 );
and \U$10811 ( \12651 , RI9959fe0_238, \12563 );
and \U$10812 ( \12652 , RI995e978_225, \12569 );
and \U$10813 ( \12653 , RI99675a0_212, \12571 );
and \U$10814 ( \12654 , RI890fab0_199, \12573 );
and \U$10815 ( \12655 , RI8918a98_186, \12575 );
and \U$10816 ( \12656 , RI89252c0_173, \12577 );
and \U$10817 ( \12657 , RI8930cd8_160, \12579 );
and \U$10818 ( \12658 , RI8939cc0_147, \12581 );
and \U$10819 ( \12659 , RI89464e8_134, \12583 );
and \U$10820 ( \12660 , RI89ec550_121, \12585 );
and \U$10821 ( \12661 , RI9776e90_108, \12587 );
and \U$10822 ( \12662 , RI9808390_95, \12589 );
and \U$10823 ( \12663 , RI98089a8_82, \12591 );
and \U$10824 ( \12664 , RI9819640_69, \12593 );
and \U$10825 ( \12665 , RI98abb48_56, \12595 );
and \U$10826 ( \12666 , RI98bc7e0_43, \12597 );
and \U$10827 ( \12667 , RI994dce0_30, \12599 );
or \U$10828 ( \12668 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 );
_DC g3969 ( \12669_nG3969 , \12668 , \12618 );
buf \U$10829 ( \12670 , \12669_nG3969 );
not \U$10830 ( \12671 , \12670 );
and \U$10831 ( \12672 , \12650 , \12671 );
xor \U$10832 ( \12673 , \12474 , \12487 );
buf \U$10833 ( \12674 , \12673 );
buf \U$10834 ( \12675 , \12674 );
and \U$10835 ( \12676 , RI9959f68_239, \12563 );
and \U$10836 ( \12677 , RI995e900_226, \12569 );
and \U$10837 ( \12678 , RI9967528_213, \12571 );
and \U$10838 ( \12679 , RI890fa38_200, \12573 );
and \U$10839 ( \12680 , RI8918a20_187, \12575 );
and \U$10840 ( \12681 , RI8925248_174, \12577 );
and \U$10841 ( \12682 , RI8930c60_161, \12579 );
and \U$10842 ( \12683 , RI8939c48_148, \12581 );
and \U$10843 ( \12684 , RI8946470_135, \12583 );
and \U$10844 ( \12685 , RI89ec4d8_122, \12585 );
and \U$10845 ( \12686 , RI9776e18_109, \12587 );
and \U$10846 ( \12687 , RI9808318_96, \12589 );
and \U$10847 ( \12688 , RI9808930_83, \12591 );
and \U$10848 ( \12689 , RI98195c8_70, \12593 );
and \U$10849 ( \12690 , RI98abad0_57, \12595 );
and \U$10850 ( \12691 , RI98bc768_44, \12597 );
and \U$10851 ( \12692 , RI994dc68_31, \12599 );
or \U$10852 ( \12693 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 );
_DC g3945 ( \12694_nG3945 , \12693 , \12618 );
buf \U$10853 ( \12695 , \12694_nG3945 );
not \U$10854 ( \12696 , \12695 );
and \U$10855 ( \12697 , \12675 , \12696 );
xor \U$10856 ( \12698 , \12475 , \12486 );
buf \U$10857 ( \12699 , \12698 );
buf \U$10858 ( \12700 , \12699 );
and \U$10859 ( \12701 , RI9959860_240, \12563 );
and \U$10860 ( \12702 , RI995e888_227, \12569 );
and \U$10861 ( \12703 , RI99674b0_214, \12571 );
and \U$10862 ( \12704 , RI890f9c0_201, \12573 );
and \U$10863 ( \12705 , RI89189a8_188, \12575 );
and \U$10864 ( \12706 , RI89251d0_175, \12577 );
and \U$10865 ( \12707 , RI8930be8_162, \12579 );
and \U$10866 ( \12708 , RI8939bd0_149, \12581 );
and \U$10867 ( \12709 , RI89463f8_136, \12583 );
and \U$10868 ( \12710 , RI89ec460_123, \12585 );
and \U$10869 ( \12711 , RI9776da0_110, \12587 );
and \U$10870 ( \12712 , RI98082a0_97, \12589 );
and \U$10871 ( \12713 , RI98088b8_84, \12591 );
and \U$10872 ( \12714 , RI9819550_71, \12593 );
and \U$10873 ( \12715 , RI98aba58_58, \12595 );
and \U$10874 ( \12716 , RI98bc6f0_45, \12597 );
and \U$10875 ( \12717 , RI994dbf0_32, \12599 );
or \U$10876 ( \12718 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 );
_DC g37c6 ( \12719_nG37c6 , \12718 , \12618 );
buf \U$10877 ( \12720 , \12719_nG37c6 );
not \U$10878 ( \12721 , \12720 );
and \U$10879 ( \12722 , \12700 , \12721 );
xor \U$10880 ( \12723 , \12476 , \12485 );
buf \U$10881 ( \12724 , \12723 );
buf \U$10882 ( \12725 , \12724 );
and \U$10883 ( \12726 , RI994d998_241, \12563 );
and \U$10884 ( \12727 , RI995e810_228, \12569 );
and \U$10885 ( \12728 , RI9967438_215, \12571 );
and \U$10886 ( \12729 , RI890f948_202, \12573 );
and \U$10887 ( \12730 , RI8918930_189, \12575 );
and \U$10888 ( \12731 , RI8925158_176, \12577 );
and \U$10889 ( \12732 , RI8930b70_163, \12579 );
and \U$10890 ( \12733 , RI8939b58_150, \12581 );
and \U$10891 ( \12734 , RI8946380_137, \12583 );
and \U$10892 ( \12735 , RI89ec3e8_124, \12585 );
and \U$10893 ( \12736 , RI9776d28_111, \12587 );
and \U$10894 ( \12737 , RI9808228_98, \12589 );
and \U$10895 ( \12738 , RI9808840_85, \12591 );
and \U$10896 ( \12739 , RI98194d8_72, \12593 );
and \U$10897 ( \12740 , RI98ab9e0_59, \12595 );
and \U$10898 ( \12741 , RI98abff8_46, \12597 );
and \U$10899 ( \12742 , RI98bcc90_33, \12599 );
or \U$10900 ( \12743 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 );
_DC g37a2 ( \12744_nG37a2 , \12743 , \12618 );
buf \U$10901 ( \12745 , \12744_nG37a2 );
not \U$10902 ( \12746 , \12745 );
and \U$10903 ( \12747 , \12725 , \12746 );
xor \U$10904 ( \12748 , \12477 , \12484 );
buf \U$10905 ( \12749 , \12748 );
buf \U$10906 ( \12750 , \12749 );
and \U$10907 ( \12751 , RI994d920_242, \12563 );
and \U$10908 ( \12752 , RI995e798_229, \12569 );
and \U$10909 ( \12753 , RI99673c0_216, \12571 );
and \U$10910 ( \12754 , RI890f8d0_203, \12573 );
and \U$10911 ( \12755 , RI89188b8_190, \12575 );
and \U$10912 ( \12756 , RI89250e0_177, \12577 );
and \U$10913 ( \12757 , RI8930af8_164, \12579 );
and \U$10914 ( \12758 , RI8939ae0_151, \12581 );
and \U$10915 ( \12759 , RI8946308_138, \12583 );
and \U$10916 ( \12760 , RI89ec370_125, \12585 );
and \U$10917 ( \12761 , RI89ec988_112, \12587 );
and \U$10918 ( \12762 , RI97772c8_99, \12589 );
and \U$10919 ( \12763 , RI98087c8_86, \12591 );
and \U$10920 ( \12764 , RI9819460_73, \12593 );
and \U$10921 ( \12765 , RI98ab968_60, \12595 );
and \U$10922 ( \12766 , RI98abf80_47, \12597 );
and \U$10923 ( \12767 , RI98bcc18_34, \12599 );
or \U$10924 ( \12768 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 );
_DC g3657 ( \12769_nG3657 , \12768 , \12618 );
buf \U$10925 ( \12770 , \12769_nG3657 );
not \U$10926 ( \12771 , \12770 );
and \U$10927 ( \12772 , \12750 , \12771 );
xor \U$10928 ( \12773 , \12478 , \12483 );
buf \U$10929 ( \12774 , \12773 );
buf \U$10930 ( \12775 , \12774 );
and \U$10931 ( \12776 , RI994d8a8_243, \12563 );
and \U$10932 ( \12777 , RI995e720_230, \12569 );
and \U$10933 ( \12778 , RI9967348_217, \12571 );
and \U$10934 ( \12779 , RI890f858_204, \12573 );
and \U$10935 ( \12780 , RI8918840_191, \12575 );
and \U$10936 ( \12781 , RI8925068_178, \12577 );
and \U$10937 ( \12782 , RI8930a80_165, \12579 );
and \U$10938 ( \12783 , RI8939a68_152, \12581 );
and \U$10939 ( \12784 , RI8946290_139, \12583 );
and \U$10940 ( \12785 , RI89ec2f8_126, \12585 );
and \U$10941 ( \12786 , RI89ec910_113, \12587 );
and \U$10942 ( \12787 , RI9777250_100, \12589 );
and \U$10943 ( \12788 , RI9808750_87, \12591 );
and \U$10944 ( \12789 , RI98193e8_74, \12593 );
and \U$10945 ( \12790 , RI98ab8f0_61, \12595 );
and \U$10946 ( \12791 , RI98abf08_48, \12597 );
and \U$10947 ( \12792 , RI98bcba0_35, \12599 );
or \U$10948 ( \12793 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 );
_DC g3633 ( \12794_nG3633 , \12793 , \12618 );
buf \U$10949 ( \12795 , \12794_nG3633 );
not \U$10950 ( \12796 , \12795 );
and \U$10951 ( \12797 , \12775 , \12796 );
xor \U$10952 ( \12798 , \12479 , \12482 );
buf \U$10953 ( \12799 , \12798 );
buf \U$10954 ( \12800 , \12799 );
and \U$10955 ( \12801 , RI994d830_244, \12563 );
and \U$10956 ( \12802 , RI995e6a8_231, \12569 );
and \U$10957 ( \12803 , RI99672d0_218, \12571 );
and \U$10958 ( \12804 , RI890f7e0_205, \12573 );
and \U$10959 ( \12805 , RI89187c8_192, \12575 );
and \U$10960 ( \12806 , RI8924ff0_179, \12577 );
and \U$10961 ( \12807 , RI8930a08_166, \12579 );
and \U$10962 ( \12808 , RI89399f0_153, \12581 );
and \U$10963 ( \12809 , RI8946218_140, \12583 );
and \U$10964 ( \12810 , RI89ec280_127, \12585 );
and \U$10965 ( \12811 , RI89ec898_114, \12587 );
and \U$10966 ( \12812 , RI97771d8_101, \12589 );
and \U$10967 ( \12813 , RI98086d8_88, \12591 );
and \U$10968 ( \12814 , RI9819370_75, \12593 );
and \U$10969 ( \12815 , RI98ab878_62, \12595 );
and \U$10970 ( \12816 , RI98abe90_49, \12597 );
and \U$10971 ( \12817 , RI98bcb28_36, \12599 );
or \U$10972 ( \12818 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 );
_DC g3518 ( \12819_nG3518 , \12818 , \12618 );
buf \U$10973 ( \12820 , \12819_nG3518 );
not \U$10974 ( \12821 , \12820 );
and \U$10975 ( \12822 , \12800 , \12821 );
xor \U$10976 ( \12823 , \12480 , \12481 );
buf \U$10977 ( \12824 , \12823 );
buf \U$10978 ( \12825 , \12824 );
and \U$10979 ( \12826 , RI994d7b8_245, \12563 );
and \U$10980 ( \12827 , RI995e630_232, \12569 );
and \U$10981 ( \12828 , RI9967258_219, \12571 );
and \U$10982 ( \12829 , RI890f768_206, \12573 );
and \U$10983 ( \12830 , RI8918750_193, \12575 );
and \U$10984 ( \12831 , RI8924f78_180, \12577 );
and \U$10985 ( \12832 , RI8930990_167, \12579 );
and \U$10986 ( \12833 , RI8939978_154, \12581 );
and \U$10987 ( \12834 , RI89461a0_141, \12583 );
and \U$10988 ( \12835 , RI89ec208_128, \12585 );
and \U$10989 ( \12836 , RI89ec820_115, \12587 );
and \U$10990 ( \12837 , RI9777160_102, \12589 );
and \U$10991 ( \12838 , RI9808660_89, \12591 );
and \U$10992 ( \12839 , RI98192f8_76, \12593 );
and \U$10993 ( \12840 , RI98ab800_63, \12595 );
and \U$10994 ( \12841 , RI98abe18_50, \12597 );
and \U$10995 ( \12842 , RI98bcab0_37, \12599 );
or \U$10996 ( \12843 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 );
_DC g3531 ( \12844_nG3531 , \12843 , \12618 );
buf \U$10997 ( \12845 , \12844_nG3531 );
not \U$10998 ( \12846 , \12845 );
and \U$10999 ( \12847 , \12825 , \12846 );
not \U$11000 ( \12848 , \12481 );
buf \U$11001 ( \12849 , \12848 );
buf \U$11002 ( \12850 , \12849 );
and \U$11003 ( \12851 , RI994d740_246, \12563 );
and \U$11004 ( \12852 , RI995e5b8_233, \12569 );
and \U$11005 ( \12853 , RI99671e0_220, \12571 );
and \U$11006 ( \12854 , RI890f6f0_207, \12573 );
and \U$11007 ( \12855 , RI89186d8_194, \12575 );
and \U$11008 ( \12856 , RI8924f00_181, \12577 );
and \U$11009 ( \12857 , RI8930918_168, \12579 );
and \U$11010 ( \12858 , RI8939900_155, \12581 );
and \U$11011 ( \12859 , RI8946128_142, \12583 );
and \U$11012 ( \12860 , RI89ec190_129, \12585 );
and \U$11013 ( \12861 , RI89ec7a8_116, \12587 );
and \U$11014 ( \12862 , RI97770e8_103, \12589 );
and \U$11015 ( \12863 , RI98085e8_90, \12591 );
and \U$11016 ( \12864 , RI9819280_77, \12593 );
and \U$11017 ( \12865 , RI98ab788_64, \12595 );
and \U$11018 ( \12866 , RI98abda0_51, \12597 );
and \U$11019 ( \12867 , RI98bca38_38, \12599 );
or \U$11020 ( \12868 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 );
_DC g342e ( \12869_nG342e , \12868 , \12618 );
buf \U$11021 ( \12870 , \12869_nG342e );
not \U$11022 ( \12871 , \12870 );
and \U$11023 ( \12872 , \12850 , \12871 );
buf \U$11024 ( \12873 , RI994e4d8_13);
buf \U$11027 ( \12874 , \12873 );
and \U$11028 ( \12875 , RI994d6c8_247, \12563 );
and \U$11029 ( \12876 , RI995e540_234, \12569 );
and \U$11030 ( \12877 , RI9967168_221, \12571 );
and \U$11031 ( \12878 , RI890f678_208, \12573 );
and \U$11032 ( \12879 , RI8918660_195, \12575 );
and \U$11033 ( \12880 , RI8924e88_182, \12577 );
and \U$11034 ( \12881 , RI89308a0_169, \12579 );
and \U$11035 ( \12882 , RI8939888_156, \12581 );
and \U$11036 ( \12883 , RI89460b0_143, \12583 );
and \U$11037 ( \12884 , RI89ec118_130, \12585 );
and \U$11038 ( \12885 , RI89ec730_117, \12587 );
and \U$11039 ( \12886 , RI9777070_104, \12589 );
and \U$11040 ( \12887 , RI9808570_91, \12591 );
and \U$11041 ( \12888 , RI9819208_78, \12593 );
and \U$11042 ( \12889 , RI98ab710_65, \12595 );
and \U$11043 ( \12890 , RI98abd28_52, \12597 );
and \U$11044 ( \12891 , RI98bc9c0_39, \12599 );
or \U$11045 ( \12892 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 );
_DC g3412 ( \12893_nG3412 , \12892 , \12618 );
buf \U$11046 ( \12894 , \12893_nG3412 );
not \U$11047 ( \12895 , \12894 );
or \U$11048 ( \12896 , \12874 , \12895 );
and \U$11049 ( \12897 , \12871 , \12896 );
and \U$11050 ( \12898 , \12850 , \12896 );
or \U$11051 ( \12899 , \12872 , \12897 , \12898 );
and \U$11052 ( \12900 , \12846 , \12899 );
and \U$11053 ( \12901 , \12825 , \12899 );
or \U$11054 ( \12902 , \12847 , \12900 , \12901 );
and \U$11055 ( \12903 , \12821 , \12902 );
and \U$11056 ( \12904 , \12800 , \12902 );
or \U$11057 ( \12905 , \12822 , \12903 , \12904 );
and \U$11058 ( \12906 , \12796 , \12905 );
and \U$11059 ( \12907 , \12775 , \12905 );
or \U$11060 ( \12908 , \12797 , \12906 , \12907 );
and \U$11061 ( \12909 , \12771 , \12908 );
and \U$11062 ( \12910 , \12750 , \12908 );
or \U$11063 ( \12911 , \12772 , \12909 , \12910 );
and \U$11064 ( \12912 , \12746 , \12911 );
and \U$11065 ( \12913 , \12725 , \12911 );
or \U$11066 ( \12914 , \12747 , \12912 , \12913 );
and \U$11067 ( \12915 , \12721 , \12914 );
and \U$11068 ( \12916 , \12700 , \12914 );
or \U$11069 ( \12917 , \12722 , \12915 , \12916 );
and \U$11070 ( \12918 , \12696 , \12917 );
and \U$11071 ( \12919 , \12675 , \12917 );
or \U$11072 ( \12920 , \12697 , \12918 , \12919 );
and \U$11073 ( \12921 , \12671 , \12920 );
and \U$11074 ( \12922 , \12650 , \12920 );
or \U$11075 ( \12923 , \12672 , \12921 , \12922 );
and \U$11076 ( \12924 , \12646 , \12923 );
and \U$11077 ( \12925 , \12625 , \12923 );
or \U$11078 ( \12926 , \12647 , \12924 , \12925 );
xor \U$11079 ( \12927 , \12622 , \12926 );
buf g3b29_GF_PartitionCandidate( \12928_nG3b29 , \12927 );
buf \U$11080 ( \12929 , \12928_nG3b29 );
xor \U$11081 ( \12930 , \12625 , \12646 );
xor \U$11082 ( \12931 , \12930 , \12923 );
buf g3b05_GF_PartitionCandidate( \12932_nG3b05 , \12931 );
buf \U$11083 ( \12933 , \12932_nG3b05 );
xor \U$11084 ( \12934 , \12650 , \12671 );
xor \U$11085 ( \12935 , \12934 , \12920 );
buf g3972_GF_PartitionCandidate( \12936_nG3972 , \12935 );
buf \U$11086 ( \12937 , \12936_nG3972 );
and \U$11087 ( \12938 , \12933 , \12937 );
not \U$11088 ( \12939 , \12938 );
and \U$11089 ( \12940 , \12929 , \12939 );
not \U$11090 ( \12941 , \12940 );
buf \U$11091 ( \12942 , \12513 );
buf \U$11092 ( \12943 , \12534 );
buf \U$11093 ( \12944 , \12538 );
buf \U$11094 ( \12945 , \12542 );
buf \U$11095 ( \12946 , \12546 );
buf \U$11096 ( \12947 , \12550 );
buf \U$11097 ( \12948 , \12554 );
buf \U$11098 ( \12949 , \12558 );
buf \U$11099 ( \12950 , \12562 );
buf \U$11100 ( \12951 , \12529 );
nor \U$11101 ( \12952 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 );
buf \U$11102 ( \12953 , \12952 );
buf \U$11103 ( \12954 , \12953 );
xor \U$11104 ( \12955 , \12942 , \12954 );
buf \U$11105 ( \12956 , \12955 );
buf \U$11106 ( \12957 , \12517 );
and \U$11107 ( \12958 , \12942 , \12954 );
xor \U$11108 ( \12959 , \12957 , \12958 );
buf \U$11109 ( \12960 , \12959 );
buf \U$11110 ( \12961 , \12521 );
and \U$11111 ( \12962 , \12957 , \12958 );
xor \U$11112 ( \12963 , \12961 , \12962 );
buf \U$11113 ( \12964 , \12963 );
buf \U$11114 ( \12965 , \12525 );
and \U$11115 ( \12966 , \12961 , \12962 );
xor \U$11116 ( \12967 , \12965 , \12966 );
buf \U$11117 ( \12968 , \12967 );
buf \U$11118 ( \12969 , \12529 );
and \U$11119 ( \12970 , \12965 , \12966 );
xor \U$11120 ( \12971 , \12969 , \12970 );
buf \U$11121 ( \12972 , \12971 );
not \U$11122 ( \12973 , \12972 );
buf \U$11123 ( \12974 , \12534 );
and \U$11124 ( \12975 , \12969 , \12970 );
xor \U$11125 ( \12976 , \12974 , \12975 );
buf \U$11126 ( \12977 , \12976 );
buf \U$11127 ( \12978 , \12538 );
and \U$11128 ( \12979 , \12974 , \12975 );
xor \U$11129 ( \12980 , \12978 , \12979 );
buf \U$11130 ( \12981 , \12980 );
buf \U$11131 ( \12982 , \12542 );
and \U$11132 ( \12983 , \12978 , \12979 );
xor \U$11133 ( \12984 , \12982 , \12983 );
buf \U$11134 ( \12985 , \12984 );
buf \U$11135 ( \12986 , \12546 );
and \U$11136 ( \12987 , \12982 , \12983 );
xor \U$11137 ( \12988 , \12986 , \12987 );
buf \U$11138 ( \12989 , \12988 );
buf \U$11139 ( \12990 , \12550 );
and \U$11140 ( \12991 , \12986 , \12987 );
xor \U$11141 ( \12992 , \12990 , \12991 );
buf \U$11142 ( \12993 , \12992 );
buf \U$11143 ( \12994 , \12554 );
and \U$11144 ( \12995 , \12990 , \12991 );
xor \U$11145 ( \12996 , \12994 , \12995 );
buf \U$11146 ( \12997 , \12996 );
buf \U$11147 ( \12998 , \12558 );
and \U$11148 ( \12999 , \12994 , \12995 );
xor \U$11149 ( \13000 , \12998 , \12999 );
buf \U$11150 ( \13001 , \13000 );
buf \U$11151 ( \13002 , \12562 );
and \U$11152 ( \13003 , \12998 , \12999 );
xor \U$11153 ( \13004 , \13002 , \13003 );
buf \U$11154 ( \13005 , \13004 );
nor \U$11155 ( \13006 , \12956 , \12960 , \12964 , \12968 , \12973 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11156 ( \13007 , RI9922bd0_569, \13006 );
not \U$11157 ( \13008 , \12956 );
not \U$11158 ( \13009 , \12960 );
not \U$11159 ( \13010 , \12964 );
not \U$11160 ( \13011 , \12968 );
nor \U$11161 ( \13012 , \13008 , \13009 , \13010 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11162 ( \13013 , RI9923800_549, \13012 );
nor \U$11163 ( \13014 , \12956 , \13009 , \13010 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11164 ( \13015 , RI9924160_529, \13014 );
nor \U$11165 ( \13016 , \13008 , \12960 , \13010 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11166 ( \13017 , RI9924ac0_509, \13016 );
nor \U$11167 ( \13018 , \12956 , \12960 , \13010 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11168 ( \13019 , RI9925ab0_489, \13018 );
nor \U$11169 ( \13020 , \13008 , \13009 , \12964 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11170 ( \13021 , RI9926410_469, \13020 );
nor \U$11171 ( \13022 , \12956 , \13009 , \12964 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11172 ( \13023 , RI9926d70_449, \13022 );
nor \U$11173 ( \13024 , \13008 , \12960 , \12964 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11174 ( \13025 , RI9928120_429, \13024 );
nor \U$11175 ( \13026 , \12956 , \12960 , \12964 , \13011 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11176 ( \13027 , RI9928a80_409, \13026 );
nor \U$11177 ( \13028 , \13008 , \13009 , \13010 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11178 ( \13029 , RI992a1f0_389, \13028 );
nor \U$11179 ( \13030 , \12956 , \13009 , \13010 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11180 ( \13031 , RI992ab50_369, \13030 );
nor \U$11181 ( \13032 , \13008 , \12960 , \13010 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11182 ( \13033 , RI992b4b0_349, \13032 );
nor \U$11183 ( \13034 , \12956 , \12960 , \13010 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11184 ( \13035 , RI992cfe0_329, \13034 );
nor \U$11185 ( \13036 , \13008 , \13009 , \12964 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11186 ( \13037 , RI992eed0_309, \13036 );
nor \U$11187 ( \13038 , \12956 , \13009 , \12964 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11188 ( \13039 , RI992f830_289, \13038 );
nor \U$11189 ( \13040 , \13008 , \12960 , \12964 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11190 ( \13041 , RI9931ae0_269, \13040 );
nor \U$11191 ( \13042 , \12956 , \12960 , \12964 , \12968 , \12972 , \12977 , \12981 , \12985 , \12989 , \12993 , \12997 , \13001 , \13005 );
and \U$11192 ( \13043 , RI994d5d8_249, \13042 );
or \U$11193 ( \13044 , \13007 , \13013 , \13015 , \13017 , \13019 , \13021 , \13023 , \13025 , \13027 , \13029 , \13031 , \13033 , \13035 , \13037 , \13039 , \13041 , \13043 );
buf \U$11194 ( \13045 , \12977 );
buf \U$11195 ( \13046 , \12981 );
buf \U$11196 ( \13047 , \12985 );
buf \U$11197 ( \13048 , \12989 );
buf \U$11198 ( \13049 , \12993 );
buf \U$11199 ( \13050 , \12997 );
buf \U$11200 ( \13051 , \13001 );
buf \U$11201 ( \13052 , \13005 );
buf \U$11202 ( \13053 , \12972 );
buf \U$11203 ( \13054 , \12956 );
buf \U$11204 ( \13055 , \12960 );
buf \U$11205 ( \13056 , \12964 );
buf \U$11206 ( \13057 , \12968 );
or \U$11207 ( \13058 , \13054 , \13055 , \13056 , \13057 );
and \U$11208 ( \13059 , \13053 , \13058 );
or \U$11209 ( \13060 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13059 );
buf \U$11210 ( \13061 , \13060 );
_DC g41fa ( \13062_nG41fa , \13044 , \13061 );
buf \U$11211 ( \13063 , \13062_nG41fa );
buf \U$11212 ( \13064 , RI995f0f8_1);
and \U$11213 ( \13065 , \12471 , \12490 );
and \U$11214 ( \13066 , \13064 , \13065 );
buf \U$11215 ( \13067 , \13066 );
buf \U$11216 ( \13068 , \13067 );
xor \U$11217 ( \13069 , \13064 , \13065 );
buf \U$11218 ( \13070 , \13069 );
buf \U$11219 ( \13071 , \13070 );
and \U$11220 ( \13072 , RI995e4c8_235, \12563 );
and \U$11221 ( \13073 , RI99670f0_222, \12569 );
and \U$11222 ( \13074 , RI890f600_209, \12571 );
and \U$11223 ( \13075 , RI89185e8_196, \12573 );
and \U$11224 ( \13076 , RI8924e10_183, \12575 );
and \U$11225 ( \13077 , RI8930828_170, \12577 );
and \U$11226 ( \13078 , RI8939810_157, \12579 );
and \U$11227 ( \13079 , RI8946038_144, \12581 );
and \U$11228 ( \13080 , RI89ec0a0_131, \12583 );
and \U$11229 ( \13081 , RI89ec6b8_118, \12585 );
and \U$11230 ( \13082 , RI9776ff8_105, \12587 );
and \U$11231 ( \13083 , RI98084f8_92, \12589 );
and \U$11232 ( \13084 , RI9808b10_79, \12591 );
and \U$11233 ( \13085 , RI98197a8_66, \12593 );
and \U$11234 ( \13086 , RI98abcb0_53, \12595 );
and \U$11235 ( \13087 , RI98bc948_40, \12597 );
and \U$11236 ( \13088 , RI994de48_27, \12599 );
or \U$11237 ( \13089 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 );
_DC g3cdb ( \13090_nG3cdb , \13089 , \12618 );
buf \U$11238 ( \13091 , \13090_nG3cdb );
not \U$11239 ( \13092 , \13091 );
and \U$11240 ( \13093 , \13071 , \13092 );
and \U$11241 ( \13094 , \12493 , \12621 );
and \U$11242 ( \13095 , \12621 , \12926 );
and \U$11243 ( \13096 , \12493 , \12926 );
or \U$11244 ( \13097 , \13094 , \13095 , \13096 );
and \U$11245 ( \13098 , \13092 , \13097 );
and \U$11246 ( \13099 , \13071 , \13097 );
or \U$11247 ( \13100 , \13093 , \13098 , \13099 );
xnor \U$11248 ( \13101 , \13068 , \13100 );
buf g3cf0_GF_PartitionCandidate( \13102_nG3cf0 , \13101 );
buf \U$11249 ( \13103 , \13102_nG3cf0 );
xor \U$11250 ( \13104 , \13071 , \13092 );
xor \U$11251 ( \13105 , \13104 , \13097 );
buf g3ce4_GF_PartitionCandidate( \13106_nG3ce4 , \13105 );
buf \U$11252 ( \13107 , \13106_nG3ce4 );
xor \U$11253 ( \13108 , \13103 , \13107 );
xor \U$11254 ( \13109 , \13107 , \12929 );
not \U$11255 ( \13110 , \13109 );
and \U$11256 ( \13111 , \13108 , \13110 );
and \U$11257 ( \13112 , \13063 , \13111 );
and \U$11258 ( \13113 , RI9922f18_568, \13006 );
and \U$11259 ( \13114 , RI9923878_548, \13012 );
and \U$11260 ( \13115 , RI99241d8_528, \13014 );
and \U$11261 ( \13116 , RI9924b38_508, \13016 );
and \U$11262 ( \13117 , RI9925b28_488, \13018 );
and \U$11263 ( \13118 , RI9926488_468, \13020 );
and \U$11264 ( \13119 , RI9926de8_448, \13022 );
and \U$11265 ( \13120 , RI9928198_428, \13024 );
and \U$11266 ( \13121 , RI9928af8_408, \13026 );
and \U$11267 ( \13122 , RI992a268_388, \13028 );
and \U$11268 ( \13123 , RI992abc8_368, \13030 );
and \U$11269 ( \13124 , RI992c6f8_348, \13032 );
and \U$11270 ( \13125 , RI992d058_328, \13034 );
and \U$11271 ( \13126 , RI992ef48_308, \13036 );
and \U$11272 ( \13127 , RI992f8a8_288, \13038 );
and \U$11273 ( \13128 , RI9931b58_268, \13040 );
and \U$11274 ( \13129 , RI994d650_248, \13042 );
or \U$11275 ( \13130 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 );
_DC g42ef ( \13131_nG42ef , \13130 , \13061 );
buf \U$11276 ( \13132 , \13131_nG42ef );
and \U$11277 ( \13133 , \13132 , \13109 );
nor \U$11278 ( \13134 , \13112 , \13133 );
and \U$11279 ( \13135 , \13107 , \12929 );
not \U$11280 ( \13136 , \13135 );
and \U$11281 ( \13137 , \13103 , \13136 );
xnor \U$11282 ( \13138 , \13134 , \13137 );
xor \U$11283 ( \13139 , \12941 , \13138 );
and \U$11285 ( \13140 , RI9922b58_570, \13006 );
and \U$11286 ( \13141 , RI9923788_550, \13012 );
and \U$11287 ( \13142 , RI99240e8_530, \13014 );
and \U$11288 ( \13143 , RI9924a48_510, \13016 );
and \U$11289 ( \13144 , RI9925a38_490, \13018 );
and \U$11290 ( \13145 , RI9926398_470, \13020 );
and \U$11291 ( \13146 , RI9926cf8_450, \13022 );
and \U$11292 ( \13147 , RI99280a8_430, \13024 );
and \U$11293 ( \13148 , RI9928a08_410, \13026 );
and \U$11294 ( \13149 , RI992a178_390, \13028 );
and \U$11295 ( \13150 , RI992aad8_370, \13030 );
and \U$11296 ( \13151 , RI992b438_350, \13032 );
and \U$11297 ( \13152 , RI992cf68_330, \13034 );
and \U$11298 ( \13153 , RI992ee58_310, \13036 );
and \U$11299 ( \13154 , RI992f7b8_290, \13038 );
and \U$11300 ( \13155 , RI9931a68_270, \13040 );
and \U$11301 ( \13156 , RI994d560_250, \13042 );
or \U$11302 ( \13157 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 );
_DC g4131 ( \13158_nG4131 , \13157 , \13061 );
buf \U$11303 ( \13159 , \13158_nG4131 );
or \U$11304 ( \13160 , \13068 , \13100 );
not \U$11305 ( \13161 , \13160 );
buf g3eca_GF_PartitionCandidate( \13162_nG3eca , \13161 );
buf \U$11306 ( \13163 , \13162_nG3eca );
xor \U$11307 ( \13164 , \13163 , \13103 );
and \U$11308 ( \13165 , \13159 , \13164 );
nor \U$11309 ( \13166 , 1'b0 , \13165 );
xnor \U$11311 ( \13167 , \13166 , 1'b0 );
xor \U$11312 ( \13168 , \13139 , \13167 );
xor \U$11313 ( \13169 , 1'b0 , \13168 );
xor \U$11315 ( \13170 , \12929 , \12933 );
xor \U$11316 ( \13171 , \12933 , \12937 );
not \U$11317 ( \13172 , \13171 );
and \U$11318 ( \13173 , \13170 , \13172 );
and \U$11319 ( \13174 , \13132 , \13173 );
not \U$11320 ( \13175 , \13174 );
xnor \U$11321 ( \13176 , \13175 , \12940 );
and \U$11322 ( \13177 , \13159 , \13111 );
and \U$11323 ( \13178 , \13063 , \13109 );
nor \U$11324 ( \13179 , \13177 , \13178 );
xnor \U$11325 ( \13180 , \13179 , \13137 );
and \U$11326 ( \13181 , \13176 , \13180 );
or \U$11328 ( \13182 , 1'b0 , \13181 , 1'b0 );
xor \U$11330 ( \13183 , \13182 , 1'b0 );
xor \U$11332 ( \13184 , \13183 , 1'b0 );
and \U$11333 ( \13185 , \13169 , \13184 );
or \U$11334 ( \13186 , 1'b0 , 1'b0 , \13185 );
and \U$11337 ( \13187 , \13132 , \13111 );
not \U$11338 ( \13188 , \13187 );
xnor \U$11339 ( \13189 , \13188 , \13137 );
xor \U$11340 ( \13190 , 1'b0 , \13189 );
and \U$11342 ( \13191 , \13063 , \13164 );
nor \U$11343 ( \13192 , 1'b0 , \13191 );
xnor \U$11344 ( \13193 , \13192 , 1'b0 );
xor \U$11345 ( \13194 , \13190 , \13193 );
xor \U$11346 ( \13195 , 1'b0 , \13194 );
xor \U$11348 ( \13196 , \13195 , 1'b1 );
and \U$11349 ( \13197 , \12941 , \13138 );
and \U$11350 ( \13198 , \13138 , \13167 );
and \U$11351 ( \13199 , \12941 , \13167 );
or \U$11352 ( \13200 , \13197 , \13198 , \13199 );
xor \U$11354 ( \13201 , \13200 , 1'b0 );
xor \U$11356 ( \13202 , \13201 , 1'b0 );
xor \U$11357 ( \13203 , \13196 , \13202 );
and \U$11358 ( \13204 , \13186 , \13203 );
or \U$11360 ( \13205 , 1'b0 , \13204 , 1'b0 );
xor \U$11362 ( \13206 , \13205 , 1'b0 );
and \U$11364 ( \13207 , \13195 , 1'b1 );
and \U$11365 ( \13208 , 1'b1 , \13202 );
and \U$11366 ( \13209 , \13195 , \13202 );
or \U$11367 ( \13210 , \13207 , \13208 , \13209 );
xor \U$11368 ( \13211 , 1'b0 , \13210 );
not \U$11370 ( \13212 , \13137 );
and \U$11372 ( \13213 , \13132 , \13164 );
nor \U$11373 ( \13214 , 1'b0 , \13213 );
xnor \U$11374 ( \13215 , \13214 , 1'b0 );
xor \U$11375 ( \13216 , \13212 , \13215 );
xor \U$11377 ( \13217 , \13216 , 1'b0 );
xor \U$11378 ( \13218 , 1'b0 , \13217 );
xor \U$11380 ( \13219 , \13218 , 1'b0 );
and \U$11382 ( \13220 , \13189 , \13193 );
or \U$11384 ( \13221 , 1'b0 , \13220 , 1'b0 );
xor \U$11386 ( \13222 , \13221 , 1'b0 );
xor \U$11388 ( \13223 , \13222 , 1'b0 );
xor \U$11389 ( \13224 , \13219 , \13223 );
xor \U$11390 ( \13225 , \13211 , \13224 );
xor \U$11391 ( \13226 , \13206 , \13225 );
xor \U$11397 ( \13227 , \12675 , \12696 );
xor \U$11398 ( \13228 , \13227 , \12917 );
buf g394e_GF_PartitionCandidate( \13229_nG394e , \13228 );
buf \U$11399 ( \13230 , \13229_nG394e );
xor \U$11400 ( \13231 , \12937 , \13230 );
xor \U$11401 ( \13232 , \12700 , \12721 );
xor \U$11402 ( \13233 , \13232 , \12914 );
buf g37cf_GF_PartitionCandidate( \13234_nG37cf , \13233 );
buf \U$11403 ( \13235 , \13234_nG37cf );
xor \U$11404 ( \13236 , \13230 , \13235 );
not \U$11405 ( \13237 , \13236 );
and \U$11406 ( \13238 , \13231 , \13237 );
and \U$11407 ( \13239 , \13132 , \13238 );
not \U$11408 ( \13240 , \13239 );
and \U$11409 ( \13241 , \13230 , \13235 );
not \U$11410 ( \13242 , \13241 );
and \U$11411 ( \13243 , \12937 , \13242 );
xnor \U$11412 ( \13244 , \13240 , \13243 );
and \U$11413 ( \13245 , \13159 , \13173 );
and \U$11414 ( \13246 , \13063 , \13171 );
nor \U$11415 ( \13247 , \13245 , \13246 );
xnor \U$11416 ( \13248 , \13247 , \12940 );
and \U$11417 ( \13249 , \13244 , \13248 );
or \U$11419 ( \13250 , 1'b0 , \13249 , 1'b0 );
and \U$11420 ( \13251 , RI9922a68_572, \13006 );
and \U$11421 ( \13252 , RI9923698_552, \13012 );
and \U$11422 ( \13253 , RI9923ff8_532, \13014 );
and \U$11423 ( \13254 , RI9924958_512, \13016 );
and \U$11424 ( \13255 , RI9925948_492, \13018 );
and \U$11425 ( \13256 , RI99262a8_472, \13020 );
and \U$11426 ( \13257 , RI9926c08_452, \13022 );
and \U$11427 ( \13258 , RI9927fb8_432, \13024 );
and \U$11428 ( \13259 , RI9928918_412, \13026 );
and \U$11429 ( \13260 , RI9929278_392, \13028 );
and \U$11430 ( \13261 , RI992a9e8_372, \13030 );
and \U$11431 ( \13262 , RI992b348_352, \13032 );
and \U$11432 ( \13263 , RI992ce78_332, \13034 );
and \U$11433 ( \13264 , RI992ed68_312, \13036 );
and \U$11434 ( \13265 , RI992f6c8_292, \13038 );
and \U$11435 ( \13266 , RI9931978_272, \13040 );
and \U$11436 ( \13267 , RI994d470_252, \13042 );
or \U$11437 ( \13268 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 );
_DC g3f92 ( \13269_nG3f92 , \13268 , \13061 );
buf \U$11438 ( \13270 , \13269_nG3f92 );
and \U$11439 ( \13271 , \13270 , \13111 );
and \U$11440 ( \13272 , RI9922ae0_571, \13006 );
and \U$11441 ( \13273 , RI9923710_551, \13012 );
and \U$11442 ( \13274 , RI9924070_531, \13014 );
and \U$11443 ( \13275 , RI99249d0_511, \13016 );
and \U$11444 ( \13276 , RI99259c0_491, \13018 );
and \U$11445 ( \13277 , RI9926320_471, \13020 );
and \U$11446 ( \13278 , RI9926c80_451, \13022 );
and \U$11447 ( \13279 , RI9928030_431, \13024 );
and \U$11448 ( \13280 , RI9928990_411, \13026 );
and \U$11449 ( \13281 , RI992a100_391, \13028 );
and \U$11450 ( \13282 , RI992aa60_371, \13030 );
and \U$11451 ( \13283 , RI992b3c0_351, \13032 );
and \U$11452 ( \13284 , RI992cef0_331, \13034 );
and \U$11453 ( \13285 , RI992ede0_311, \13036 );
and \U$11454 ( \13286 , RI992f740_291, \13038 );
and \U$11455 ( \13287 , RI99319f0_271, \13040 );
and \U$11456 ( \13288 , RI994d4e8_251, \13042 );
or \U$11457 ( \13289 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 );
_DC g4070 ( \13290_nG4070 , \13289 , \13061 );
buf \U$11458 ( \13291 , \13290_nG4070 );
and \U$11459 ( \13292 , \13291 , \13109 );
nor \U$11460 ( \13293 , \13271 , \13292 );
xnor \U$11461 ( \13294 , \13293 , \13137 );
and \U$11463 ( \13295 , RI99229f0_573, \13006 );
and \U$11464 ( \13296 , RI9923620_553, \13012 );
and \U$11465 ( \13297 , RI9923f80_533, \13014 );
and \U$11466 ( \13298 , RI99248e0_513, \13016 );
and \U$11467 ( \13299 , RI99258d0_493, \13018 );
and \U$11468 ( \13300 , RI9926230_473, \13020 );
and \U$11469 ( \13301 , RI9926b90_453, \13022 );
and \U$11470 ( \13302 , RI9927f40_433, \13024 );
and \U$11471 ( \13303 , RI99288a0_413, \13026 );
and \U$11472 ( \13304 , RI9929200_393, \13028 );
and \U$11473 ( \13305 , RI992a970_373, \13030 );
and \U$11474 ( \13306 , RI992b2d0_353, \13032 );
and \U$11475 ( \13307 , RI992ce00_333, \13034 );
and \U$11476 ( \13308 , RI992ecf0_313, \13036 );
and \U$11477 ( \13309 , RI992f650_293, \13038 );
and \U$11478 ( \13310 , RI9931900_273, \13040 );
and \U$11479 ( \13311 , RI994d3f8_253, \13042 );
or \U$11480 ( \13312 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 );
_DC g3ea9 ( \13313_nG3ea9 , \13312 , \13061 );
buf \U$11481 ( \13314 , \13313_nG3ea9 );
and \U$11482 ( \13315 , \13314 , \13164 );
nor \U$11483 ( \13316 , 1'b0 , \13315 );
xnor \U$11484 ( \13317 , \13316 , 1'b0 );
and \U$11485 ( \13318 , \13294 , \13317 );
or \U$11488 ( \13319 , \13318 , 1'b0 , 1'b0 );
and \U$11489 ( \13320 , \13250 , \13319 );
or \U$11492 ( \13321 , \13320 , 1'b0 , 1'b0 );
and \U$11495 ( \13322 , \13270 , \13164 );
nor \U$11496 ( \13323 , 1'b0 , \13322 );
xnor \U$11497 ( \13324 , \13323 , 1'b0 );
xor \U$11499 ( \13325 , \13324 , 1'b0 );
xor \U$11501 ( \13326 , \13325 , 1'b0 );
not \U$11502 ( \13327 , \13243 );
and \U$11503 ( \13328 , \13063 , \13173 );
and \U$11504 ( \13329 , \13132 , \13171 );
nor \U$11505 ( \13330 , \13328 , \13329 );
xnor \U$11506 ( \13331 , \13330 , \12940 );
xor \U$11507 ( \13332 , \13327 , \13331 );
and \U$11508 ( \13333 , \13291 , \13111 );
and \U$11509 ( \13334 , \13159 , \13109 );
nor \U$11510 ( \13335 , \13333 , \13334 );
xnor \U$11511 ( \13336 , \13335 , \13137 );
xor \U$11512 ( \13337 , \13332 , \13336 );
and \U$11513 ( \13338 , \13326 , \13337 );
or \U$11515 ( \13339 , 1'b0 , \13338 , 1'b0 );
and \U$11516 ( \13340 , \13321 , \13339 );
or \U$11517 ( \13341 , 1'b0 , 1'b0 , \13340 );
and \U$11519 ( \13342 , \13291 , \13164 );
nor \U$11520 ( \13343 , 1'b0 , \13342 );
xnor \U$11521 ( \13344 , \13343 , 1'b0 );
xor \U$11523 ( \13345 , \13344 , 1'b0 );
xor \U$11525 ( \13346 , \13345 , 1'b0 );
xor \U$11527 ( \13347 , 1'b0 , \13176 );
xor \U$11528 ( \13348 , \13347 , \13180 );
xor \U$11529 ( \13349 , \13346 , \13348 );
and \U$11531 ( \13350 , \13349 , 1'b1 );
and \U$11532 ( \13351 , \13327 , \13331 );
and \U$11533 ( \13352 , \13331 , \13336 );
and \U$11534 ( \13353 , \13327 , \13336 );
or \U$11535 ( \13354 , \13351 , \13352 , \13353 );
xor \U$11537 ( \13355 , \13354 , 1'b0 );
xor \U$11539 ( \13356 , \13355 , 1'b0 );
and \U$11540 ( \13357 , 1'b1 , \13356 );
and \U$11541 ( \13358 , \13349 , \13356 );
or \U$11542 ( \13359 , \13350 , \13357 , \13358 );
and \U$11543 ( \13360 , \13341 , \13359 );
xor \U$11545 ( \13361 , \13169 , 1'b0 );
xor \U$11546 ( \13362 , \13361 , \13184 );
and \U$11547 ( \13363 , \13359 , \13362 );
and \U$11548 ( \13364 , \13341 , \13362 );
or \U$11549 ( \13365 , \13360 , \13363 , \13364 );
xor \U$11551 ( \13366 , 1'b0 , \13186 );
xor \U$11552 ( \13367 , \13366 , \13203 );
and \U$11553 ( \13368 , \13365 , \13367 );
or \U$11554 ( \13369 , 1'b0 , 1'b0 , \13368 );
nand \U$11555 ( \13370 , \13226 , \13369 );
nor \U$11556 ( \13371 , \13226 , \13369 );
not \U$11557 ( \13372 , \13371 );
nand \U$11558 ( \13373 , \13370 , \13372 );
xor \U$11559 ( \13374 , \12850 , \12871 );
xor \U$11560 ( \13375 , \13374 , \12896 );
buf g3435_GF_PartitionCandidate( \13376_nG3435 , \13375 );
buf \U$11561 ( \13377 , \13376_nG3435 );
xor \U$11562 ( \13378 , \12874 , \12894 );
buf g3415_GF_PartitionCandidate( \13379_nG3415 , \13378 );
buf \U$11563 ( \13380 , \13379_nG3415 );
xor \U$11564 ( \13381 , \13377 , \13380 );
not \U$11565 ( \13382 , \13380 );
and \U$11566 ( \13383 , \13381 , \13382 );
and \U$11567 ( \13384 , \13314 , \13383 );
and \U$11568 ( \13385 , \13270 , \13380 );
nor \U$11569 ( \13386 , \13384 , \13385 );
xnor \U$11570 ( \13387 , \13386 , \13377 );
and \U$11571 ( \13388 , RI9922900_575, \13006 );
and \U$11572 ( \13389 , RI9923530_555, \13012 );
and \U$11573 ( \13390 , RI9923e90_535, \13014 );
and \U$11574 ( \13391 , RI99247f0_515, \13016 );
and \U$11575 ( \13392 , RI99257e0_495, \13018 );
and \U$11576 ( \13393 , RI9926140_475, \13020 );
and \U$11577 ( \13394 , RI9926aa0_455, \13022 );
and \U$11578 ( \13395 , RI9927e50_435, \13024 );
and \U$11579 ( \13396 , RI99287b0_415, \13026 );
and \U$11580 ( \13397 , RI9929110_395, \13028 );
and \U$11581 ( \13398 , RI992a880_375, \13030 );
and \U$11582 ( \13399 , RI992b1e0_355, \13032 );
and \U$11583 ( \13400 , RI992cd10_335, \13034 );
and \U$11584 ( \13401 , RI992d670_315, \13036 );
and \U$11585 ( \13402 , RI992f560_295, \13038 );
and \U$11586 ( \13403 , RI9931810_275, \13040 );
and \U$11587 ( \13404 , RI9935f50_255, \13042 );
or \U$11588 ( \13405 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 );
_DC g3d18 ( \13406_nG3d18 , \13405 , \13061 );
buf \U$11589 ( \13407 , \13406_nG3d18 );
xor \U$11590 ( \13408 , \12800 , \12821 );
xor \U$11591 ( \13409 , \13408 , \12902 );
buf g353d_GF_PartitionCandidate( \13410_nG353d , \13409 );
buf \U$11592 ( \13411 , \13410_nG353d );
xor \U$11593 ( \13412 , \12825 , \12846 );
xor \U$11594 ( \13413 , \13412 , \12899 );
buf g3541_GF_PartitionCandidate( \13414_nG3541 , \13413 );
buf \U$11595 ( \13415 , \13414_nG3541 );
xor \U$11596 ( \13416 , \13411 , \13415 );
xor \U$11597 ( \13417 , \13415 , \13377 );
not \U$11598 ( \13418 , \13417 );
and \U$11599 ( \13419 , \13416 , \13418 );
and \U$11600 ( \13420 , \13407 , \13419 );
and \U$11601 ( \13421 , RI9922978_574, \13006 );
and \U$11602 ( \13422 , RI99235a8_554, \13012 );
and \U$11603 ( \13423 , RI9923f08_534, \13014 );
and \U$11604 ( \13424 , RI9924868_514, \13016 );
and \U$11605 ( \13425 , RI9925858_494, \13018 );
and \U$11606 ( \13426 , RI99261b8_474, \13020 );
and \U$11607 ( \13427 , RI9926b18_454, \13022 );
and \U$11608 ( \13428 , RI9927ec8_434, \13024 );
and \U$11609 ( \13429 , RI9928828_414, \13026 );
and \U$11610 ( \13430 , RI9929188_394, \13028 );
and \U$11611 ( \13431 , RI992a8f8_374, \13030 );
and \U$11612 ( \13432 , RI992b258_354, \13032 );
and \U$11613 ( \13433 , RI992cd88_334, \13034 );
and \U$11614 ( \13434 , RI992d6e8_314, \13036 );
and \U$11615 ( \13435 , RI992f5d8_294, \13038 );
and \U$11616 ( \13436 , RI9931888_274, \13040 );
and \U$11617 ( \13437 , RI9935fc8_254, \13042 );
or \U$11618 ( \13438 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 );
_DC g3dc5 ( \13439_nG3dc5 , \13438 , \13061 );
buf \U$11619 ( \13440 , \13439_nG3dc5 );
and \U$11620 ( \13441 , \13440 , \13417 );
nor \U$11621 ( \13442 , \13420 , \13441 );
and \U$11622 ( \13443 , \13415 , \13377 );
not \U$11623 ( \13444 , \13443 );
and \U$11624 ( \13445 , \13411 , \13444 );
xnor \U$11625 ( \13446 , \13442 , \13445 );
and \U$11626 ( \13447 , \13387 , \13446 );
and \U$11627 ( \13448 , RI9922810_577, \13006 );
and \U$11628 ( \13449 , RI9923440_557, \13012 );
and \U$11629 ( \13450 , RI9923da0_537, \13014 );
and \U$11630 ( \13451 , RI9924700_517, \13016 );
and \U$11631 ( \13452 , RI99256f0_497, \13018 );
and \U$11632 ( \13453 , RI9926050_477, \13020 );
and \U$11633 ( \13454 , RI99269b0_457, \13022 );
and \U$11634 ( \13455 , RI9927d60_437, \13024 );
and \U$11635 ( \13456 , RI99286c0_417, \13026 );
and \U$11636 ( \13457 , RI9929020_397, \13028 );
and \U$11637 ( \13458 , RI992a790_377, \13030 );
and \U$11638 ( \13459 , RI992b0f0_357, \13032 );
and \U$11639 ( \13460 , RI992cc20_337, \13034 );
and \U$11640 ( \13461 , RI992d580_317, \13036 );
and \U$11641 ( \13462 , RI992f470_297, \13038 );
and \U$11642 ( \13463 , RI9931720_277, \13040 );
and \U$11643 ( \13464 , RI9933d90_257, \13042 );
or \U$11644 ( \13465 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 );
_DC g3b58 ( \13466_nG3b58 , \13465 , \13061 );
buf \U$11645 ( \13467 , \13466_nG3b58 );
xor \U$11646 ( \13468 , \12750 , \12771 );
xor \U$11647 ( \13469 , \13468 , \12908 );
buf g3660_GF_PartitionCandidate( \13470_nG3660 , \13469 );
buf \U$11648 ( \13471 , \13470_nG3660 );
xor \U$11649 ( \13472 , \12775 , \12796 );
xor \U$11650 ( \13473 , \13472 , \12905 );
buf g363c_GF_PartitionCandidate( \13474_nG363c , \13473 );
buf \U$11651 ( \13475 , \13474_nG363c );
xor \U$11652 ( \13476 , \13471 , \13475 );
xor \U$11653 ( \13477 , \13475 , \13411 );
not \U$11654 ( \13478 , \13477 );
and \U$11655 ( \13479 , \13476 , \13478 );
and \U$11656 ( \13480 , \13467 , \13479 );
and \U$11657 ( \13481 , RI9922888_576, \13006 );
and \U$11658 ( \13482 , RI99234b8_556, \13012 );
and \U$11659 ( \13483 , RI9923e18_536, \13014 );
and \U$11660 ( \13484 , RI9924778_516, \13016 );
and \U$11661 ( \13485 , RI9925768_496, \13018 );
and \U$11662 ( \13486 , RI99260c8_476, \13020 );
and \U$11663 ( \13487 , RI9926a28_456, \13022 );
and \U$11664 ( \13488 , RI9927dd8_436, \13024 );
and \U$11665 ( \13489 , RI9928738_416, \13026 );
and \U$11666 ( \13490 , RI9929098_396, \13028 );
and \U$11667 ( \13491 , RI992a808_376, \13030 );
and \U$11668 ( \13492 , RI992b168_356, \13032 );
and \U$11669 ( \13493 , RI992cc98_336, \13034 );
and \U$11670 ( \13494 , RI992d5f8_316, \13036 );
and \U$11671 ( \13495 , RI992f4e8_296, \13038 );
and \U$11672 ( \13496 , RI9931798_276, \13040 );
and \U$11673 ( \13497 , RI9935ed8_256, \13042 );
or \U$11674 ( \13498 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 );
_DC g3bf0 ( \13499_nG3bf0 , \13498 , \13061 );
buf \U$11675 ( \13500 , \13499_nG3bf0 );
and \U$11676 ( \13501 , \13500 , \13477 );
nor \U$11677 ( \13502 , \13480 , \13501 );
and \U$11678 ( \13503 , \13475 , \13411 );
not \U$11679 ( \13504 , \13503 );
and \U$11680 ( \13505 , \13471 , \13504 );
xnor \U$11681 ( \13506 , \13502 , \13505 );
and \U$11682 ( \13507 , \13446 , \13506 );
and \U$11683 ( \13508 , \13387 , \13506 );
or \U$11684 ( \13509 , \13447 , \13507 , \13508 );
and \U$11685 ( \13510 , RI9922720_579, \13006 );
and \U$11686 ( \13511 , RI9923350_559, \13012 );
and \U$11687 ( \13512 , RI9923cb0_539, \13014 );
and \U$11688 ( \13513 , RI9924610_519, \13016 );
and \U$11689 ( \13514 , RI9925600_499, \13018 );
and \U$11690 ( \13515 , RI9925f60_479, \13020 );
and \U$11691 ( \13516 , RI99268c0_459, \13022 );
and \U$11692 ( \13517 , RI9927c70_439, \13024 );
and \U$11693 ( \13518 , RI99285d0_419, \13026 );
and \U$11694 ( \13519 , RI9928f30_399, \13028 );
and \U$11695 ( \13520 , RI992a6a0_379, \13030 );
and \U$11696 ( \13521 , RI992b000_359, \13032 );
and \U$11697 ( \13522 , RI992cb30_339, \13034 );
and \U$11698 ( \13523 , RI992d490_319, \13036 );
and \U$11699 ( \13524 , RI992f380_299, \13038 );
and \U$11700 ( \13525 , RI9931630_279, \13040 );
and \U$11701 ( \13526 , RI9933ca0_259, \13042 );
or \U$11702 ( \13527 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 );
_DC g398d ( \13528_nG398d , \13527 , \13061 );
buf \U$11703 ( \13529 , \13528_nG398d );
xor \U$11704 ( \13530 , \12725 , \12746 );
xor \U$11705 ( \13531 , \13530 , \12911 );
buf g37ab_GF_PartitionCandidate( \13532_nG37ab , \13531 );
buf \U$11706 ( \13533 , \13532_nG37ab );
xor \U$11707 ( \13534 , \13235 , \13533 );
xor \U$11708 ( \13535 , \13533 , \13471 );
not \U$11709 ( \13536 , \13535 );
and \U$11710 ( \13537 , \13534 , \13536 );
and \U$11711 ( \13538 , \13529 , \13537 );
and \U$11712 ( \13539 , RI9922798_578, \13006 );
and \U$11713 ( \13540 , RI99233c8_558, \13012 );
and \U$11714 ( \13541 , RI9923d28_538, \13014 );
and \U$11715 ( \13542 , RI9924688_518, \13016 );
and \U$11716 ( \13543 , RI9925678_498, \13018 );
and \U$11717 ( \13544 , RI9925fd8_478, \13020 );
and \U$11718 ( \13545 , RI9926938_458, \13022 );
and \U$11719 ( \13546 , RI9927ce8_438, \13024 );
and \U$11720 ( \13547 , RI9928648_418, \13026 );
and \U$11721 ( \13548 , RI9928fa8_398, \13028 );
and \U$11722 ( \13549 , RI992a718_378, \13030 );
and \U$11723 ( \13550 , RI992b078_358, \13032 );
and \U$11724 ( \13551 , RI992cba8_338, \13034 );
and \U$11725 ( \13552 , RI992d508_318, \13036 );
and \U$11726 ( \13553 , RI992f3f8_298, \13038 );
and \U$11727 ( \13554 , RI99316a8_278, \13040 );
and \U$11728 ( \13555 , RI9933d18_258, \13042 );
or \U$11729 ( \13556 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 );
_DC g3a17 ( \13557_nG3a17 , \13556 , \13061 );
buf \U$11730 ( \13558 , \13557_nG3a17 );
and \U$11731 ( \13559 , \13558 , \13535 );
nor \U$11732 ( \13560 , \13538 , \13559 );
and \U$11733 ( \13561 , \13533 , \13471 );
not \U$11734 ( \13562 , \13561 );
and \U$11735 ( \13563 , \13235 , \13562 );
xnor \U$11736 ( \13564 , \13560 , \13563 );
and \U$11737 ( \13565 , RI9922630_581, \13006 );
and \U$11738 ( \13566 , RI9923260_561, \13012 );
and \U$11739 ( \13567 , RI9923bc0_541, \13014 );
and \U$11740 ( \13568 , RI9924520_521, \13016 );
and \U$11741 ( \13569 , RI9925510_501, \13018 );
and \U$11742 ( \13570 , RI9925e70_481, \13020 );
and \U$11743 ( \13571 , RI99267d0_461, \13022 );
and \U$11744 ( \13572 , RI9927b80_441, \13024 );
and \U$11745 ( \13573 , RI99284e0_421, \13026 );
and \U$11746 ( \13574 , RI9928e40_401, \13028 );
and \U$11747 ( \13575 , RI992a5b0_381, \13030 );
and \U$11748 ( \13576 , RI992af10_361, \13032 );
and \U$11749 ( \13577 , RI992ca40_341, \13034 );
and \U$11750 ( \13578 , RI992d3a0_321, \13036 );
and \U$11751 ( \13579 , RI992f290_301, \13038 );
and \U$11752 ( \13580 , RI9931540_281, \13040 );
and \U$11753 ( \13581 , RI9933bb0_261, \13042 );
or \U$11754 ( \13582 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 );
_DC g37ea ( \13583_nG37ea , \13582 , \13061 );
buf \U$11755 ( \13584 , \13583_nG37ea );
and \U$11756 ( \13585 , \13584 , \13238 );
and \U$11757 ( \13586 , RI99226a8_580, \13006 );
and \U$11758 ( \13587 , RI99232d8_560, \13012 );
and \U$11759 ( \13588 , RI9923c38_540, \13014 );
and \U$11760 ( \13589 , RI9924598_520, \13016 );
and \U$11761 ( \13590 , RI9925588_500, \13018 );
and \U$11762 ( \13591 , RI9925ee8_480, \13020 );
and \U$11763 ( \13592 , RI9926848_460, \13022 );
and \U$11764 ( \13593 , RI9927bf8_440, \13024 );
and \U$11765 ( \13594 , RI9928558_420, \13026 );
and \U$11766 ( \13595 , RI9928eb8_400, \13028 );
and \U$11767 ( \13596 , RI992a628_380, \13030 );
and \U$11768 ( \13597 , RI992af88_360, \13032 );
and \U$11769 ( \13598 , RI992cab8_340, \13034 );
and \U$11770 ( \13599 , RI992d418_320, \13036 );
and \U$11771 ( \13600 , RI992f308_300, \13038 );
and \U$11772 ( \13601 , RI99315b8_280, \13040 );
and \U$11773 ( \13602 , RI9933c28_260, \13042 );
or \U$11774 ( \13603 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 );
_DC g385e ( \13604_nG385e , \13603 , \13061 );
buf \U$11775 ( \13605 , \13604_nG385e );
and \U$11776 ( \13606 , \13605 , \13236 );
nor \U$11777 ( \13607 , \13585 , \13606 );
xnor \U$11778 ( \13608 , \13607 , \13243 );
and \U$11779 ( \13609 , \13564 , \13608 );
and \U$11780 ( \13610 , RI9922540_583, \13006 );
and \U$11781 ( \13611 , RI9923170_563, \13012 );
and \U$11782 ( \13612 , RI9923ad0_543, \13014 );
and \U$11783 ( \13613 , RI9924430_523, \13016 );
and \U$11784 ( \13614 , RI9924d90_503, \13018 );
and \U$11785 ( \13615 , RI9925d80_483, \13020 );
and \U$11786 ( \13616 , RI99266e0_463, \13022 );
and \U$11787 ( \13617 , RI9927040_443, \13024 );
and \U$11788 ( \13618 , RI99283f0_423, \13026 );
and \U$11789 ( \13619 , RI9928d50_403, \13028 );
and \U$11790 ( \13620 , RI992a4c0_383, \13030 );
and \U$11791 ( \13621 , RI992ae20_363, \13032 );
and \U$11792 ( \13622 , RI992c950_343, \13034 );
and \U$11793 ( \13623 , RI992d2b0_323, \13036 );
and \U$11794 ( \13624 , RI992f1a0_303, \13038 );
and \U$11795 ( \13625 , RI9931450_283, \13040 );
and \U$11796 ( \13626 , RI9933ac0_263, \13042 );
or \U$11797 ( \13627 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 );
_DC g3679 ( \13628_nG3679 , \13627 , \13061 );
buf \U$11798 ( \13629 , \13628_nG3679 );
and \U$11799 ( \13630 , \13629 , \13173 );
and \U$11800 ( \13631 , RI99225b8_582, \13006 );
and \U$11801 ( \13632 , RI99231e8_562, \13012 );
and \U$11802 ( \13633 , RI9923b48_542, \13014 );
and \U$11803 ( \13634 , RI99244a8_522, \13016 );
and \U$11804 ( \13635 , RI9924e08_502, \13018 );
and \U$11805 ( \13636 , RI9925df8_482, \13020 );
and \U$11806 ( \13637 , RI9926758_462, \13022 );
and \U$11807 ( \13638 , RI9927b08_442, \13024 );
and \U$11808 ( \13639 , RI9928468_422, \13026 );
and \U$11809 ( \13640 , RI9928dc8_402, \13028 );
and \U$11810 ( \13641 , RI992a538_382, \13030 );
and \U$11811 ( \13642 , RI992ae98_362, \13032 );
and \U$11812 ( \13643 , RI992c9c8_342, \13034 );
and \U$11813 ( \13644 , RI992d328_322, \13036 );
and \U$11814 ( \13645 , RI992f218_302, \13038 );
and \U$11815 ( \13646 , RI99314c8_282, \13040 );
and \U$11816 ( \13647 , RI9933b38_262, \13042 );
or \U$11817 ( \13648 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 );
_DC g36e0 ( \13649_nG36e0 , \13648 , \13061 );
buf \U$11818 ( \13650 , \13649_nG36e0 );
and \U$11819 ( \13651 , \13650 , \13171 );
nor \U$11820 ( \13652 , \13630 , \13651 );
xnor \U$11821 ( \13653 , \13652 , \12940 );
and \U$11822 ( \13654 , \13608 , \13653 );
and \U$11823 ( \13655 , \13564 , \13653 );
or \U$11824 ( \13656 , \13609 , \13654 , \13655 );
and \U$11825 ( \13657 , \13509 , \13656 );
and \U$11826 ( \13658 , RI9922450_585, \13006 );
and \U$11827 ( \13659 , RI9923080_565, \13012 );
and \U$11828 ( \13660 , RI99239e0_545, \13014 );
and \U$11829 ( \13661 , RI9924340_525, \13016 );
and \U$11830 ( \13662 , RI9924ca0_505, \13018 );
and \U$11831 ( \13663 , RI9925c90_485, \13020 );
and \U$11832 ( \13664 , RI99265f0_465, \13022 );
and \U$11833 ( \13665 , RI9926f50_445, \13024 );
and \U$11834 ( \13666 , RI9928300_425, \13026 );
and \U$11835 ( \13667 , RI9928c60_405, \13028 );
and \U$11836 ( \13668 , RI992a3d0_385, \13030 );
and \U$11837 ( \13669 , RI992ad30_365, \13032 );
and \U$11838 ( \13670 , RI992c860_345, \13034 );
and \U$11839 ( \13671 , RI992d1c0_325, \13036 );
and \U$11840 ( \13672 , RI992f0b0_305, \13038 );
and \U$11841 ( \13673 , RI9931360_285, \13040 );
and \U$11842 ( \13674 , RI99339d0_265, \13042 );
or \U$11843 ( \13675 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 );
_DC g34fb ( \13676_nG34fb , \13675 , \13061 );
buf \U$11844 ( \13677 , \13676_nG34fb );
and \U$11845 ( \13678 , \13677 , \13111 );
and \U$11846 ( \13679 , RI99224c8_584, \13006 );
and \U$11847 ( \13680 , RI99230f8_564, \13012 );
and \U$11848 ( \13681 , RI9923a58_544, \13014 );
and \U$11849 ( \13682 , RI99243b8_524, \13016 );
and \U$11850 ( \13683 , RI9924d18_504, \13018 );
and \U$11851 ( \13684 , RI9925d08_484, \13020 );
and \U$11852 ( \13685 , RI9926668_464, \13022 );
and \U$11853 ( \13686 , RI9926fc8_444, \13024 );
and \U$11854 ( \13687 , RI9928378_424, \13026 );
and \U$11855 ( \13688 , RI9928cd8_404, \13028 );
and \U$11856 ( \13689 , RI992a448_384, \13030 );
and \U$11857 ( \13690 , RI992ada8_364, \13032 );
and \U$11858 ( \13691 , RI992c8d8_344, \13034 );
and \U$11859 ( \13692 , RI992d238_324, \13036 );
and \U$11860 ( \13693 , RI992f128_304, \13038 );
and \U$11861 ( \13694 , RI99313d8_284, \13040 );
and \U$11862 ( \13695 , RI9933a48_264, \13042 );
or \U$11863 ( \13696 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 );
_DC g358e ( \13697_nG358e , \13696 , \13061 );
buf \U$11864 ( \13698 , \13697_nG358e );
and \U$11865 ( \13699 , \13698 , \13109 );
nor \U$11866 ( \13700 , \13678 , \13699 );
xnor \U$11867 ( \13701 , \13700 , \13137 );
and \U$11869 ( \13702 , RI99223d8_586, \13006 );
and \U$11870 ( \13703 , RI9923008_566, \13012 );
and \U$11871 ( \13704 , RI9923968_546, \13014 );
and \U$11872 ( \13705 , RI99242c8_526, \13016 );
and \U$11873 ( \13706 , RI9924c28_506, \13018 );
and \U$11874 ( \13707 , RI9925c18_486, \13020 );
and \U$11875 ( \13708 , RI9926578_466, \13022 );
and \U$11876 ( \13709 , RI9926ed8_446, \13024 );
and \U$11877 ( \13710 , RI9928288_426, \13026 );
and \U$11878 ( \13711 , RI9928be8_406, \13028 );
and \U$11879 ( \13712 , RI992a358_386, \13030 );
and \U$11880 ( \13713 , RI992acb8_366, \13032 );
and \U$11881 ( \13714 , RI992c7e8_346, \13034 );
and \U$11882 ( \13715 , RI992d148_326, \13036 );
and \U$11883 ( \13716 , RI992f038_306, \13038 );
and \U$11884 ( \13717 , RI99312e8_286, \13040 );
and \U$11885 ( \13718 , RI9933958_266, \13042 );
or \U$11886 ( \13719 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 );
_DC g3473 ( \13720_nG3473 , \13719 , \13061 );
buf \U$11887 ( \13721 , \13720_nG3473 );
and \U$11888 ( \13722 , \13721 , \13164 );
nor \U$11889 ( \13723 , 1'b0 , \13722 );
xnor \U$11890 ( \13724 , \13723 , 1'b0 );
and \U$11891 ( \13725 , \13701 , \13724 );
and \U$11892 ( \13726 , \13656 , \13725 );
and \U$11893 ( \13727 , \13509 , \13725 );
or \U$11894 ( \13728 , \13657 , \13726 , \13727 );
and \U$11896 ( \13729 , \13650 , \13173 );
and \U$11897 ( \13730 , \13584 , \13171 );
nor \U$11898 ( \13731 , \13729 , \13730 );
xnor \U$11899 ( \13732 , \13731 , \12940 );
and \U$11900 ( \13733 , \13698 , \13111 );
and \U$11901 ( \13734 , \13629 , \13109 );
nor \U$11902 ( \13735 , \13733 , \13734 );
xnor \U$11903 ( \13736 , \13735 , \13137 );
xor \U$11904 ( \13737 , \13732 , \13736 );
and \U$11906 ( \13738 , \13677 , \13164 );
nor \U$11907 ( \13739 , 1'b0 , \13738 );
xnor \U$11908 ( \13740 , \13739 , 1'b0 );
xor \U$11909 ( \13741 , \13737 , \13740 );
and \U$11910 ( \13742 , \13500 , \13479 );
and \U$11911 ( \13743 , \13407 , \13477 );
nor \U$11912 ( \13744 , \13742 , \13743 );
xnor \U$11913 ( \13745 , \13744 , \13505 );
and \U$11914 ( \13746 , \13558 , \13537 );
and \U$11915 ( \13747 , \13467 , \13535 );
nor \U$11916 ( \13748 , \13746 , \13747 );
xnor \U$11917 ( \13749 , \13748 , \13563 );
xor \U$11918 ( \13750 , \13745 , \13749 );
and \U$11919 ( \13751 , \13605 , \13238 );
and \U$11920 ( \13752 , \13529 , \13236 );
nor \U$11921 ( \13753 , \13751 , \13752 );
xnor \U$11922 ( \13754 , \13753 , \13243 );
xor \U$11923 ( \13755 , \13750 , \13754 );
and \U$11924 ( \13756 , \13741 , \13755 );
or \U$11926 ( \13757 , 1'b0 , \13756 , 1'b0 );
xor \U$11927 ( \13758 , \13728 , \13757 );
and \U$11928 ( \13759 , \13629 , \13111 );
and \U$11929 ( \13760 , \13650 , \13109 );
nor \U$11930 ( \13761 , \13759 , \13760 );
xnor \U$11931 ( \13762 , \13761 , \13137 );
and \U$11933 ( \13763 , \13698 , \13164 );
nor \U$11934 ( \13764 , 1'b0 , \13763 );
xnor \U$11935 ( \13765 , \13764 , 1'b0 );
xor \U$11936 ( \13766 , \13762 , \13765 );
xor \U$11938 ( \13767 , \13766 , 1'b0 );
and \U$11939 ( \13768 , \13467 , \13537 );
and \U$11940 ( \13769 , \13500 , \13535 );
nor \U$11941 ( \13770 , \13768 , \13769 );
xnor \U$11942 ( \13771 , \13770 , \13563 );
and \U$11943 ( \13772 , \13529 , \13238 );
and \U$11944 ( \13773 , \13558 , \13236 );
nor \U$11945 ( \13774 , \13772 , \13773 );
xnor \U$11946 ( \13775 , \13774 , \13243 );
xor \U$11947 ( \13776 , \13771 , \13775 );
and \U$11948 ( \13777 , \13584 , \13173 );
and \U$11949 ( \13778 , \13605 , \13171 );
nor \U$11950 ( \13779 , \13777 , \13778 );
xnor \U$11951 ( \13780 , \13779 , \12940 );
xor \U$11952 ( \13781 , \13776 , \13780 );
xor \U$11953 ( \13782 , \13767 , \13781 );
and \U$11954 ( \13783 , \13291 , \13383 );
and \U$11955 ( \13784 , \13159 , \13380 );
nor \U$11956 ( \13785 , \13783 , \13784 );
xnor \U$11957 ( \13786 , \13785 , \13377 );
and \U$11958 ( \13787 , \13314 , \13419 );
and \U$11959 ( \13788 , \13270 , \13417 );
nor \U$11960 ( \13789 , \13787 , \13788 );
xnor \U$11961 ( \13790 , \13789 , \13445 );
xor \U$11962 ( \13791 , \13786 , \13790 );
and \U$11963 ( \13792 , \13407 , \13479 );
and \U$11964 ( \13793 , \13440 , \13477 );
nor \U$11965 ( \13794 , \13792 , \13793 );
xnor \U$11966 ( \13795 , \13794 , \13505 );
xor \U$11967 ( \13796 , \13791 , \13795 );
xor \U$11968 ( \13797 , \13782 , \13796 );
xor \U$11969 ( \13798 , \13758 , \13797 );
and \U$11971 ( \13799 , \13440 , \13383 );
and \U$11972 ( \13800 , \13314 , \13380 );
nor \U$11973 ( \13801 , \13799 , \13800 );
xnor \U$11974 ( \13802 , \13801 , \13377 );
and \U$11975 ( \13803 , \13500 , \13419 );
and \U$11976 ( \13804 , \13407 , \13417 );
nor \U$11977 ( \13805 , \13803 , \13804 );
xnor \U$11978 ( \13806 , \13805 , \13445 );
and \U$11979 ( \13807 , \13802 , \13806 );
or \U$11981 ( \13808 , 1'b0 , \13807 , 1'b0 );
and \U$11982 ( \13809 , \13558 , \13479 );
and \U$11983 ( \13810 , \13467 , \13477 );
nor \U$11984 ( \13811 , \13809 , \13810 );
xnor \U$11985 ( \13812 , \13811 , \13505 );
and \U$11986 ( \13813 , \13605 , \13537 );
and \U$11987 ( \13814 , \13529 , \13535 );
nor \U$11988 ( \13815 , \13813 , \13814 );
xnor \U$11989 ( \13816 , \13815 , \13563 );
and \U$11990 ( \13817 , \13812 , \13816 );
and \U$11991 ( \13818 , \13650 , \13238 );
and \U$11992 ( \13819 , \13584 , \13236 );
nor \U$11993 ( \13820 , \13818 , \13819 );
xnor \U$11994 ( \13821 , \13820 , \13243 );
and \U$11995 ( \13822 , \13816 , \13821 );
and \U$11996 ( \13823 , \13812 , \13821 );
or \U$11997 ( \13824 , \13817 , \13822 , \13823 );
and \U$11998 ( \13825 , \13808 , \13824 );
and \U$11999 ( \13826 , \13698 , \13173 );
and \U$12000 ( \13827 , \13629 , \13171 );
nor \U$12001 ( \13828 , \13826 , \13827 );
xnor \U$12002 ( \13829 , \13828 , \12940 );
and \U$12003 ( \13830 , \13721 , \13111 );
and \U$12004 ( \13831 , \13677 , \13109 );
nor \U$12005 ( \13832 , \13830 , \13831 );
xnor \U$12006 ( \13833 , \13832 , \13137 );
and \U$12007 ( \13834 , \13829 , \13833 );
and \U$12008 ( \13835 , RI9922360_587, \13006 );
and \U$12009 ( \13836 , RI9922f90_567, \13012 );
and \U$12010 ( \13837 , RI99238f0_547, \13014 );
and \U$12011 ( \13838 , RI9924250_527, \13016 );
and \U$12012 ( \13839 , RI9924bb0_507, \13018 );
and \U$12013 ( \13840 , RI9925ba0_487, \13020 );
and \U$12014 ( \13841 , RI9926500_467, \13022 );
and \U$12015 ( \13842 , RI9926e60_447, \13024 );
and \U$12016 ( \13843 , RI9928210_427, \13026 );
and \U$12017 ( \13844 , RI9928b70_407, \13028 );
and \U$12018 ( \13845 , RI992a2e0_387, \13030 );
and \U$12019 ( \13846 , RI992ac40_367, \13032 );
and \U$12020 ( \13847 , RI992c770_347, \13034 );
and \U$12021 ( \13848 , RI992d0d0_327, \13036 );
and \U$12022 ( \13849 , RI992efc0_307, \13038 );
and \U$12023 ( \13850 , RI992f920_287, \13040 );
and \U$12024 ( \13851 , RI99338e0_267, \13042 );
or \U$12025 ( \13852 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 );
_DC g33d8 ( \13853_nG33d8 , \13852 , \13061 );
buf \U$12026 ( \13854 , \13853_nG33d8 );
nand \U$12027 ( \13855 , \13854 , \13164 );
xnor \U$12028 ( \13856 , \13855 , 1'b0 );
and \U$12029 ( \13857 , \13833 , \13856 );
and \U$12030 ( \13858 , \13829 , \13856 );
or \U$12031 ( \13859 , \13834 , \13857 , \13858 );
and \U$12032 ( \13860 , \13824 , \13859 );
and \U$12033 ( \13861 , \13808 , \13859 );
or \U$12034 ( \13862 , \13825 , \13860 , \13861 );
xor \U$12035 ( \13863 , \13701 , \13724 );
xor \U$12036 ( \13864 , \13564 , \13608 );
xor \U$12037 ( \13865 , \13864 , \13653 );
and \U$12038 ( \13866 , \13863 , \13865 );
xor \U$12039 ( \13867 , \13387 , \13446 );
xor \U$12040 ( \13868 , \13867 , \13506 );
and \U$12041 ( \13869 , \13865 , \13868 );
and \U$12042 ( \13870 , \13863 , \13868 );
or \U$12043 ( \13871 , \13866 , \13869 , \13870 );
and \U$12044 ( \13872 , \13862 , \13871 );
and \U$12046 ( \13873 , \13270 , \13383 );
and \U$12047 ( \13874 , \13291 , \13380 );
nor \U$12048 ( \13875 , \13873 , \13874 );
xnor \U$12049 ( \13876 , \13875 , \13377 );
xor \U$12050 ( \13877 , 1'b0 , \13876 );
and \U$12051 ( \13878 , \13440 , \13419 );
and \U$12052 ( \13879 , \13314 , \13417 );
nor \U$12053 ( \13880 , \13878 , \13879 );
xnor \U$12054 ( \13881 , \13880 , \13445 );
xor \U$12055 ( \13882 , \13877 , \13881 );
and \U$12056 ( \13883 , \13871 , \13882 );
and \U$12057 ( \13884 , \13862 , \13882 );
or \U$12058 ( \13885 , \13872 , \13883 , \13884 );
xor \U$12060 ( \13886 , 1'b0 , \13741 );
xor \U$12061 ( \13887 , \13886 , \13755 );
xor \U$12062 ( \13888 , \13509 , \13656 );
xor \U$12063 ( \13889 , \13888 , \13725 );
and \U$12064 ( \13890 , \13887 , \13889 );
xor \U$12065 ( \13891 , \13885 , \13890 );
and \U$12067 ( \13892 , \13876 , \13881 );
or \U$12069 ( \13893 , 1'b0 , \13892 , 1'b0 );
and \U$12070 ( \13894 , \13745 , \13749 );
and \U$12071 ( \13895 , \13749 , \13754 );
and \U$12072 ( \13896 , \13745 , \13754 );
or \U$12073 ( \13897 , \13894 , \13895 , \13896 );
xor \U$12074 ( \13898 , \13893 , \13897 );
and \U$12075 ( \13899 , \13732 , \13736 );
and \U$12076 ( \13900 , \13736 , \13740 );
and \U$12077 ( \13901 , \13732 , \13740 );
or \U$12078 ( \13902 , \13899 , \13900 , \13901 );
xor \U$12079 ( \13903 , \13898 , \13902 );
xor \U$12080 ( \13904 , \13891 , \13903 );
xor \U$12081 ( \13905 , \13798 , \13904 );
and \U$12082 ( \13906 , \13407 , \13383 );
and \U$12083 ( \13907 , \13440 , \13380 );
nor \U$12084 ( \13908 , \13906 , \13907 );
xnor \U$12085 ( \13909 , \13908 , \13377 );
and \U$12086 ( \13910 , \13467 , \13419 );
and \U$12087 ( \13911 , \13500 , \13417 );
nor \U$12088 ( \13912 , \13910 , \13911 );
xnor \U$12089 ( \13913 , \13912 , \13445 );
and \U$12090 ( \13914 , \13909 , \13913 );
and \U$12091 ( \13915 , \13529 , \13479 );
and \U$12092 ( \13916 , \13558 , \13477 );
nor \U$12093 ( \13917 , \13915 , \13916 );
xnor \U$12094 ( \13918 , \13917 , \13505 );
and \U$12095 ( \13919 , \13913 , \13918 );
and \U$12096 ( \13920 , \13909 , \13918 );
or \U$12097 ( \13921 , \13914 , \13919 , \13920 );
and \U$12098 ( \13922 , \13584 , \13537 );
and \U$12099 ( \13923 , \13605 , \13535 );
nor \U$12100 ( \13924 , \13922 , \13923 );
xnor \U$12101 ( \13925 , \13924 , \13563 );
and \U$12102 ( \13926 , \13629 , \13238 );
and \U$12103 ( \13927 , \13650 , \13236 );
nor \U$12104 ( \13928 , \13926 , \13927 );
xnor \U$12105 ( \13929 , \13928 , \13243 );
and \U$12106 ( \13930 , \13925 , \13929 );
and \U$12107 ( \13931 , \13677 , \13173 );
and \U$12108 ( \13932 , \13698 , \13171 );
nor \U$12109 ( \13933 , \13931 , \13932 );
xnor \U$12110 ( \13934 , \13933 , \12940 );
and \U$12111 ( \13935 , \13929 , \13934 );
and \U$12112 ( \13936 , \13925 , \13934 );
or \U$12113 ( \13937 , \13930 , \13935 , \13936 );
and \U$12114 ( \13938 , \13921 , \13937 );
xor \U$12115 ( \13939 , \13829 , \13833 );
xor \U$12116 ( \13940 , \13939 , \13856 );
and \U$12117 ( \13941 , \13937 , \13940 );
and \U$12118 ( \13942 , \13921 , \13940 );
or \U$12119 ( \13943 , \13938 , \13941 , \13942 );
xor \U$12120 ( \13944 , \13812 , \13816 );
xor \U$12121 ( \13945 , \13944 , \13821 );
xor \U$12122 ( \13946 , 1'b0 , \13802 );
xor \U$12123 ( \13947 , \13946 , \13806 );
and \U$12124 ( \13948 , \13945 , \13947 );
and \U$12125 ( \13949 , \13943 , \13948 );
xor \U$12126 ( \13950 , \13863 , \13865 );
xor \U$12127 ( \13951 , \13950 , \13868 );
and \U$12128 ( \13952 , \13948 , \13951 );
and \U$12129 ( \13953 , \13943 , \13951 );
or \U$12130 ( \13954 , \13949 , \13952 , \13953 );
xor \U$12131 ( \13955 , \13887 , \13889 );
and \U$12132 ( \13956 , \13954 , \13955 );
xor \U$12133 ( \13957 , \13862 , \13871 );
xor \U$12134 ( \13958 , \13957 , \13882 );
and \U$12135 ( \13959 , \13955 , \13958 );
and \U$12136 ( \13960 , \13954 , \13958 );
or \U$12137 ( \13961 , \13956 , \13959 , \13960 );
nor \U$12138 ( \13962 , \13905 , \13961 );
and \U$12139 ( \13963 , \13885 , \13890 );
and \U$12140 ( \13964 , \13890 , \13903 );
and \U$12141 ( \13965 , \13885 , \13903 );
or \U$12142 ( \13966 , \13963 , \13964 , \13965 );
and \U$12143 ( \13967 , \13728 , \13757 );
and \U$12144 ( \13968 , \13757 , \13797 );
and \U$12145 ( \13969 , \13728 , \13797 );
or \U$12146 ( \13970 , \13967 , \13968 , \13969 );
and \U$12148 ( \13971 , \13159 , \13383 );
and \U$12149 ( \13972 , \13063 , \13380 );
nor \U$12150 ( \13973 , \13971 , \13972 );
xnor \U$12151 ( \13974 , \13973 , \13377 );
xor \U$12152 ( \13975 , 1'b0 , \13974 );
and \U$12153 ( \13976 , \13270 , \13419 );
and \U$12154 ( \13977 , \13291 , \13417 );
nor \U$12155 ( \13978 , \13976 , \13977 );
xnor \U$12156 ( \13979 , \13978 , \13445 );
xor \U$12157 ( \13980 , \13975 , \13979 );
and \U$12159 ( \13981 , \13605 , \13173 );
and \U$12160 ( \13982 , \13529 , \13171 );
nor \U$12161 ( \13983 , \13981 , \13982 );
xnor \U$12162 ( \13984 , \13983 , \12940 );
and \U$12163 ( \13985 , \13650 , \13111 );
and \U$12164 ( \13986 , \13584 , \13109 );
nor \U$12165 ( \13987 , \13985 , \13986 );
xnor \U$12166 ( \13988 , \13987 , \13137 );
xor \U$12167 ( \13989 , \13984 , \13988 );
and \U$12169 ( \13990 , \13629 , \13164 );
nor \U$12170 ( \13991 , 1'b0 , \13990 );
xnor \U$12171 ( \13992 , \13991 , 1'b0 );
xor \U$12172 ( \13993 , \13989 , \13992 );
xor \U$12173 ( \13994 , 1'b0 , \13993 );
xor \U$12174 ( \13995 , \13980 , \13994 );
and \U$12175 ( \13996 , \13786 , \13790 );
and \U$12176 ( \13997 , \13790 , \13795 );
and \U$12177 ( \13998 , \13786 , \13795 );
or \U$12178 ( \13999 , \13996 , \13997 , \13998 );
and \U$12179 ( \14000 , \13771 , \13775 );
and \U$12180 ( \14001 , \13775 , \13780 );
and \U$12181 ( \14002 , \13771 , \13780 );
or \U$12182 ( \14003 , \14000 , \14001 , \14002 );
xor \U$12183 ( \14004 , \13999 , \14003 );
and \U$12184 ( \14005 , \13762 , \13765 );
or \U$12187 ( \14006 , \14005 , 1'b0 , 1'b0 );
xor \U$12188 ( \14007 , \14004 , \14006 );
xor \U$12189 ( \14008 , \13995 , \14007 );
xor \U$12190 ( \14009 , \13970 , \14008 );
and \U$12191 ( \14010 , \13893 , \13897 );
and \U$12192 ( \14011 , \13897 , \13902 );
and \U$12193 ( \14012 , \13893 , \13902 );
or \U$12194 ( \14013 , \14010 , \14011 , \14012 );
and \U$12195 ( \14014 , \13767 , \13781 );
and \U$12196 ( \14015 , \13781 , \13796 );
and \U$12197 ( \14016 , \13767 , \13796 );
or \U$12198 ( \14017 , \14014 , \14015 , \14016 );
xor \U$12199 ( \14018 , \14013 , \14017 );
and \U$12200 ( \14019 , \13440 , \13479 );
and \U$12201 ( \14020 , \13314 , \13477 );
nor \U$12202 ( \14021 , \14019 , \14020 );
xnor \U$12203 ( \14022 , \14021 , \13505 );
and \U$12204 ( \14023 , \13500 , \13537 );
and \U$12205 ( \14024 , \13407 , \13535 );
nor \U$12206 ( \14025 , \14023 , \14024 );
xnor \U$12207 ( \14026 , \14025 , \13563 );
xor \U$12208 ( \14027 , \14022 , \14026 );
and \U$12209 ( \14028 , \13558 , \13238 );
and \U$12210 ( \14029 , \13467 , \13236 );
nor \U$12211 ( \14030 , \14028 , \14029 );
xnor \U$12212 ( \14031 , \14030 , \13243 );
xor \U$12213 ( \14032 , \14027 , \14031 );
xor \U$12214 ( \14033 , \14018 , \14032 );
xor \U$12215 ( \14034 , \14009 , \14033 );
xor \U$12216 ( \14035 , \13966 , \14034 );
and \U$12217 ( \14036 , \13798 , \13904 );
nor \U$12218 ( \14037 , \14035 , \14036 );
nor \U$12219 ( \14038 , \13962 , \14037 );
and \U$12220 ( \14039 , \13970 , \14008 );
and \U$12221 ( \14040 , \14008 , \14033 );
and \U$12222 ( \14041 , \13970 , \14033 );
or \U$12223 ( \14042 , \14039 , \14040 , \14041 );
and \U$12225 ( \14043 , \13974 , \13979 );
or \U$12227 ( \14044 , 1'b0 , \14043 , 1'b0 );
and \U$12228 ( \14045 , \14022 , \14026 );
and \U$12229 ( \14046 , \14026 , \14031 );
and \U$12230 ( \14047 , \14022 , \14031 );
or \U$12231 ( \14048 , \14045 , \14046 , \14047 );
xor \U$12232 ( \14049 , \14044 , \14048 );
and \U$12233 ( \14050 , \13984 , \13988 );
and \U$12234 ( \14051 , \13988 , \13992 );
and \U$12235 ( \14052 , \13984 , \13992 );
or \U$12236 ( \14053 , \14050 , \14051 , \14052 );
xor \U$12237 ( \14054 , \14049 , \14053 );
and \U$12238 ( \14055 , \13999 , \14003 );
and \U$12239 ( \14056 , \14003 , \14006 );
and \U$12240 ( \14057 , \13999 , \14006 );
or \U$12241 ( \14058 , \14055 , \14056 , \14057 );
xor \U$12243 ( \14059 , \14058 , 1'b0 );
and \U$12244 ( \14060 , \13063 , \13383 );
and \U$12245 ( \14061 , \13132 , \13380 );
nor \U$12246 ( \14062 , \14060 , \14061 );
xnor \U$12247 ( \14063 , \14062 , \13377 );
and \U$12248 ( \14064 , \13291 , \13419 );
and \U$12249 ( \14065 , \13159 , \13417 );
nor \U$12250 ( \14066 , \14064 , \14065 );
xnor \U$12251 ( \14067 , \14066 , \13445 );
xor \U$12252 ( \14068 , \14063 , \14067 );
and \U$12253 ( \14069 , \13314 , \13479 );
and \U$12254 ( \14070 , \13270 , \13477 );
nor \U$12255 ( \14071 , \14069 , \14070 );
xnor \U$12256 ( \14072 , \14071 , \13505 );
xor \U$12257 ( \14073 , \14068 , \14072 );
xor \U$12258 ( \14074 , \14059 , \14073 );
xor \U$12259 ( \14075 , \14054 , \14074 );
xor \U$12260 ( \14076 , \14042 , \14075 );
and \U$12261 ( \14077 , \14013 , \14017 );
and \U$12262 ( \14078 , \14017 , \14032 );
and \U$12263 ( \14079 , \14013 , \14032 );
or \U$12264 ( \14080 , \14077 , \14078 , \14079 );
and \U$12265 ( \14081 , \13980 , \13994 );
and \U$12266 ( \14082 , \13994 , \14007 );
and \U$12267 ( \14083 , \13980 , \14007 );
or \U$12268 ( \14084 , \14081 , \14082 , \14083 );
xor \U$12269 ( \14085 , \14080 , \14084 );
and \U$12271 ( \14086 , \13584 , \13111 );
and \U$12272 ( \14087 , \13605 , \13109 );
nor \U$12273 ( \14088 , \14086 , \14087 );
xnor \U$12274 ( \14089 , \14088 , \13137 );
and \U$12276 ( \14090 , \13650 , \13164 );
nor \U$12277 ( \14091 , 1'b0 , \14090 );
xnor \U$12278 ( \14092 , \14091 , 1'b0 );
xor \U$12279 ( \14093 , \14089 , \14092 );
xor \U$12281 ( \14094 , \14093 , 1'b0 );
xor \U$12282 ( \14095 , 1'b0 , \14094 );
and \U$12283 ( \14096 , \13407 , \13537 );
and \U$12284 ( \14097 , \13440 , \13535 );
nor \U$12285 ( \14098 , \14096 , \14097 );
xnor \U$12286 ( \14099 , \14098 , \13563 );
and \U$12287 ( \14100 , \13467 , \13238 );
and \U$12288 ( \14101 , \13500 , \13236 );
nor \U$12289 ( \14102 , \14100 , \14101 );
xnor \U$12290 ( \14103 , \14102 , \13243 );
xor \U$12291 ( \14104 , \14099 , \14103 );
and \U$12292 ( \14105 , \13529 , \13173 );
and \U$12293 ( \14106 , \13558 , \13171 );
nor \U$12294 ( \14107 , \14105 , \14106 );
xnor \U$12295 ( \14108 , \14107 , \12940 );
xor \U$12296 ( \14109 , \14104 , \14108 );
xor \U$12297 ( \14110 , \14095 , \14109 );
xor \U$12298 ( \14111 , \14085 , \14110 );
xor \U$12299 ( \14112 , \14076 , \14111 );
and \U$12300 ( \14113 , \13966 , \14034 );
nor \U$12301 ( \14114 , \14112 , \14113 );
and \U$12302 ( \14115 , \14080 , \14084 );
and \U$12303 ( \14116 , \14084 , \14110 );
and \U$12304 ( \14117 , \14080 , \14110 );
or \U$12305 ( \14118 , \14115 , \14116 , \14117 );
and \U$12306 ( \14119 , \14054 , \14074 );
xor \U$12307 ( \14120 , \14118 , \14119 );
and \U$12310 ( \14121 , \14058 , \14073 );
or \U$12311 ( \14122 , 1'b0 , 1'b0 , \14121 );
and \U$12313 ( \14123 , \13558 , \13173 );
and \U$12314 ( \14124 , \13467 , \13171 );
nor \U$12315 ( \14125 , \14123 , \14124 );
xnor \U$12316 ( \14126 , \14125 , \12940 );
and \U$12317 ( \14127 , \13605 , \13111 );
and \U$12318 ( \14128 , \13529 , \13109 );
nor \U$12319 ( \14129 , \14127 , \14128 );
xnor \U$12320 ( \14130 , \14129 , \13137 );
xor \U$12321 ( \14131 , \14126 , \14130 );
and \U$12323 ( \14132 , \13584 , \13164 );
nor \U$12324 ( \14133 , 1'b0 , \14132 );
xnor \U$12325 ( \14134 , \14133 , 1'b0 );
xor \U$12326 ( \14135 , \14131 , \14134 );
xor \U$12327 ( \14136 , 1'b0 , \14135 );
and \U$12328 ( \14137 , \13270 , \13479 );
and \U$12329 ( \14138 , \13291 , \13477 );
nor \U$12330 ( \14139 , \14137 , \14138 );
xnor \U$12331 ( \14140 , \14139 , \13505 );
and \U$12332 ( \14141 , \13440 , \13537 );
and \U$12333 ( \14142 , \13314 , \13535 );
nor \U$12334 ( \14143 , \14141 , \14142 );
xnor \U$12335 ( \14144 , \14143 , \13563 );
xor \U$12336 ( \14145 , \14140 , \14144 );
and \U$12337 ( \14146 , \13500 , \13238 );
and \U$12338 ( \14147 , \13407 , \13236 );
nor \U$12339 ( \14148 , \14146 , \14147 );
xnor \U$12340 ( \14149 , \14148 , \13243 );
xor \U$12341 ( \14150 , \14145 , \14149 );
xor \U$12342 ( \14151 , \14136 , \14150 );
and \U$12343 ( \14152 , \14063 , \14067 );
and \U$12344 ( \14153 , \14067 , \14072 );
and \U$12345 ( \14154 , \14063 , \14072 );
or \U$12346 ( \14155 , \14152 , \14153 , \14154 );
and \U$12347 ( \14156 , \14099 , \14103 );
and \U$12348 ( \14157 , \14103 , \14108 );
and \U$12349 ( \14158 , \14099 , \14108 );
or \U$12350 ( \14159 , \14156 , \14157 , \14158 );
xor \U$12351 ( \14160 , \14155 , \14159 );
and \U$12352 ( \14161 , \14089 , \14092 );
or \U$12355 ( \14162 , \14161 , 1'b0 , 1'b0 );
xor \U$12356 ( \14163 , \14160 , \14162 );
xor \U$12357 ( \14164 , \14151 , \14163 );
xor \U$12358 ( \14165 , \14122 , \14164 );
and \U$12359 ( \14166 , \14044 , \14048 );
and \U$12360 ( \14167 , \14048 , \14053 );
and \U$12361 ( \14168 , \14044 , \14053 );
or \U$12362 ( \14169 , \14166 , \14167 , \14168 );
and \U$12364 ( \14170 , \14094 , \14109 );
or \U$12366 ( \14171 , 1'b0 , \14170 , 1'b0 );
xor \U$12367 ( \14172 , \14169 , \14171 );
and \U$12369 ( \14173 , \13132 , \13383 );
not \U$12370 ( \14174 , \14173 );
xnor \U$12371 ( \14175 , \14174 , \13377 );
xor \U$12372 ( \14176 , 1'b0 , \14175 );
and \U$12373 ( \14177 , \13159 , \13419 );
and \U$12374 ( \14178 , \13063 , \13417 );
nor \U$12375 ( \14179 , \14177 , \14178 );
xnor \U$12376 ( \14180 , \14179 , \13445 );
xor \U$12377 ( \14181 , \14176 , \14180 );
xor \U$12378 ( \14182 , \14172 , \14181 );
xor \U$12379 ( \14183 , \14165 , \14182 );
xor \U$12380 ( \14184 , \14120 , \14183 );
and \U$12381 ( \14185 , \14042 , \14075 );
and \U$12382 ( \14186 , \14075 , \14111 );
and \U$12383 ( \14187 , \14042 , \14111 );
or \U$12384 ( \14188 , \14185 , \14186 , \14187 );
nor \U$12385 ( \14189 , \14184 , \14188 );
nor \U$12386 ( \14190 , \14114 , \14189 );
nand \U$12387 ( \14191 , \14038 , \14190 );
and \U$12388 ( \14192 , \14122 , \14164 );
and \U$12389 ( \14193 , \14164 , \14182 );
and \U$12390 ( \14194 , \14122 , \14182 );
or \U$12391 ( \14195 , \14192 , \14193 , \14194 );
and \U$12392 ( \14196 , \14155 , \14159 );
and \U$12393 ( \14197 , \14159 , \14162 );
and \U$12394 ( \14198 , \14155 , \14162 );
or \U$12395 ( \14199 , \14196 , \14197 , \14198 );
and \U$12397 ( \14200 , \14135 , \14150 );
or \U$12399 ( \14201 , 1'b0 , \14200 , 1'b0 );
xor \U$12400 ( \14202 , \14199 , \14201 );
and \U$12401 ( \14203 , \13314 , \13537 );
and \U$12402 ( \14204 , \13270 , \13535 );
nor \U$12403 ( \14205 , \14203 , \14204 );
xnor \U$12404 ( \14206 , \14205 , \13563 );
and \U$12405 ( \14207 , \13407 , \13238 );
and \U$12406 ( \14208 , \13440 , \13236 );
nor \U$12407 ( \14209 , \14207 , \14208 );
xnor \U$12408 ( \14210 , \14209 , \13243 );
xor \U$12409 ( \14211 , \14206 , \14210 );
and \U$12410 ( \14212 , \13467 , \13173 );
and \U$12411 ( \14213 , \13500 , \13171 );
nor \U$12412 ( \14214 , \14212 , \14213 );
xnor \U$12413 ( \14215 , \14214 , \12940 );
xor \U$12414 ( \14216 , \14211 , \14215 );
xor \U$12415 ( \14217 , \14202 , \14216 );
xor \U$12416 ( \14218 , \14195 , \14217 );
and \U$12417 ( \14219 , \14169 , \14171 );
and \U$12418 ( \14220 , \14171 , \14181 );
and \U$12419 ( \14221 , \14169 , \14181 );
or \U$12420 ( \14222 , \14219 , \14220 , \14221 );
and \U$12421 ( \14223 , \14151 , \14163 );
xor \U$12422 ( \14224 , \14222 , \14223 );
not \U$12423 ( \14225 , \13377 );
and \U$12424 ( \14226 , \13063 , \13419 );
and \U$12425 ( \14227 , \13132 , \13417 );
nor \U$12426 ( \14228 , \14226 , \14227 );
xnor \U$12427 ( \14229 , \14228 , \13445 );
xor \U$12428 ( \14230 , \14225 , \14229 );
and \U$12429 ( \14231 , \13291 , \13479 );
and \U$12430 ( \14232 , \13159 , \13477 );
nor \U$12431 ( \14233 , \14231 , \14232 );
xnor \U$12432 ( \14234 , \14233 , \13505 );
xor \U$12433 ( \14235 , \14230 , \14234 );
and \U$12435 ( \14236 , \13529 , \13111 );
and \U$12436 ( \14237 , \13558 , \13109 );
nor \U$12437 ( \14238 , \14236 , \14237 );
xnor \U$12438 ( \14239 , \14238 , \13137 );
and \U$12440 ( \14240 , \13605 , \13164 );
nor \U$12441 ( \14241 , 1'b0 , \14240 );
xnor \U$12442 ( \14242 , \14241 , 1'b0 );
xor \U$12443 ( \14243 , \14239 , \14242 );
xor \U$12445 ( \14244 , \14243 , 1'b0 );
xor \U$12446 ( \14245 , 1'b1 , \14244 );
xor \U$12447 ( \14246 , \14235 , \14245 );
and \U$12449 ( \14247 , \14175 , \14180 );
or \U$12451 ( \14248 , 1'b0 , \14247 , 1'b0 );
and \U$12452 ( \14249 , \14140 , \14144 );
and \U$12453 ( \14250 , \14144 , \14149 );
and \U$12454 ( \14251 , \14140 , \14149 );
or \U$12455 ( \14252 , \14249 , \14250 , \14251 );
xor \U$12456 ( \14253 , \14248 , \14252 );
and \U$12457 ( \14254 , \14126 , \14130 );
and \U$12458 ( \14255 , \14130 , \14134 );
and \U$12459 ( \14256 , \14126 , \14134 );
or \U$12460 ( \14257 , \14254 , \14255 , \14256 );
xor \U$12461 ( \14258 , \14253 , \14257 );
xor \U$12462 ( \14259 , \14246 , \14258 );
xor \U$12463 ( \14260 , \14224 , \14259 );
xor \U$12464 ( \14261 , \14218 , \14260 );
and \U$12465 ( \14262 , \14118 , \14119 );
and \U$12466 ( \14263 , \14119 , \14183 );
and \U$12467 ( \14264 , \14118 , \14183 );
or \U$12468 ( \14265 , \14262 , \14263 , \14264 );
nor \U$12469 ( \14266 , \14261 , \14265 );
and \U$12470 ( \14267 , \14222 , \14223 );
and \U$12471 ( \14268 , \14223 , \14259 );
and \U$12472 ( \14269 , \14222 , \14259 );
or \U$12473 ( \14270 , \14267 , \14268 , \14269 );
and \U$12474 ( \14271 , \14225 , \14229 );
and \U$12475 ( \14272 , \14229 , \14234 );
and \U$12476 ( \14273 , \14225 , \14234 );
or \U$12477 ( \14274 , \14271 , \14272 , \14273 );
and \U$12478 ( \14275 , \14206 , \14210 );
and \U$12479 ( \14276 , \14210 , \14215 );
and \U$12480 ( \14277 , \14206 , \14215 );
or \U$12481 ( \14278 , \14275 , \14276 , \14277 );
xor \U$12482 ( \14279 , \14274 , \14278 );
and \U$12483 ( \14280 , \14239 , \14242 );
or \U$12486 ( \14281 , \14280 , 1'b0 , 1'b0 );
xor \U$12487 ( \14282 , \14279 , \14281 );
and \U$12488 ( \14283 , \14248 , \14252 );
and \U$12489 ( \14284 , \14252 , \14257 );
and \U$12490 ( \14285 , \14248 , \14257 );
or \U$12491 ( \14286 , \14283 , \14284 , \14285 );
and \U$12494 ( \14287 , 1'b1 , \14244 );
or \U$12496 ( \14288 , 1'b0 , \14287 , 1'b0 );
xor \U$12497 ( \14289 , \14286 , \14288 );
and \U$12498 ( \14290 , \13558 , \13111 );
and \U$12499 ( \14291 , \13467 , \13109 );
nor \U$12500 ( \14292 , \14290 , \14291 );
xnor \U$12501 ( \14293 , \14292 , \13137 );
and \U$12503 ( \14294 , \13529 , \13164 );
nor \U$12504 ( \14295 , 1'b0 , \14294 );
xnor \U$12505 ( \14296 , \14295 , 1'b0 );
xor \U$12506 ( \14297 , \14293 , \14296 );
xor \U$12508 ( \14298 , \14297 , 1'b0 );
and \U$12509 ( \14299 , \13270 , \13537 );
and \U$12510 ( \14300 , \13291 , \13535 );
nor \U$12511 ( \14301 , \14299 , \14300 );
xnor \U$12512 ( \14302 , \14301 , \13563 );
and \U$12513 ( \14303 , \13440 , \13238 );
and \U$12514 ( \14304 , \13314 , \13236 );
nor \U$12515 ( \14305 , \14303 , \14304 );
xnor \U$12516 ( \14306 , \14305 , \13243 );
xor \U$12517 ( \14307 , \14302 , \14306 );
and \U$12518 ( \14308 , \13500 , \13173 );
and \U$12519 ( \14309 , \13407 , \13171 );
nor \U$12520 ( \14310 , \14308 , \14309 );
xnor \U$12521 ( \14311 , \14310 , \12940 );
xor \U$12522 ( \14312 , \14307 , \14311 );
xor \U$12523 ( \14313 , \14298 , \14312 );
and \U$12525 ( \14314 , \13132 , \13419 );
not \U$12526 ( \14315 , \14314 );
xnor \U$12527 ( \14316 , \14315 , \13445 );
xor \U$12528 ( \14317 , 1'b0 , \14316 );
and \U$12529 ( \14318 , \13159 , \13479 );
and \U$12530 ( \14319 , \13063 , \13477 );
nor \U$12531 ( \14320 , \14318 , \14319 );
xnor \U$12532 ( \14321 , \14320 , \13505 );
xor \U$12533 ( \14322 , \14317 , \14321 );
xor \U$12534 ( \14323 , \14313 , \14322 );
xor \U$12535 ( \14324 , \14289 , \14323 );
xor \U$12536 ( \14325 , \14282 , \14324 );
xor \U$12537 ( \14326 , \14270 , \14325 );
and \U$12538 ( \14327 , \14199 , \14201 );
and \U$12539 ( \14328 , \14201 , \14216 );
and \U$12540 ( \14329 , \14199 , \14216 );
or \U$12541 ( \14330 , \14327 , \14328 , \14329 );
and \U$12542 ( \14331 , \14235 , \14245 );
and \U$12543 ( \14332 , \14245 , \14258 );
and \U$12544 ( \14333 , \14235 , \14258 );
or \U$12545 ( \14334 , \14331 , \14332 , \14333 );
xor \U$12546 ( \14335 , \14330 , \14334 );
xor \U$12548 ( \14336 , \14335 , 1'b1 );
xor \U$12549 ( \14337 , \14326 , \14336 );
and \U$12550 ( \14338 , \14195 , \14217 );
and \U$12551 ( \14339 , \14217 , \14260 );
and \U$12552 ( \14340 , \14195 , \14260 );
or \U$12553 ( \14341 , \14338 , \14339 , \14340 );
nor \U$12554 ( \14342 , \14337 , \14341 );
nor \U$12555 ( \14343 , \14266 , \14342 );
and \U$12556 ( \14344 , \14330 , \14334 );
and \U$12557 ( \14345 , \14334 , 1'b1 );
and \U$12558 ( \14346 , \14330 , 1'b1 );
or \U$12559 ( \14347 , \14344 , \14345 , \14346 );
and \U$12560 ( \14348 , \14282 , \14324 );
xor \U$12561 ( \14349 , \14347 , \14348 );
and \U$12562 ( \14350 , \14286 , \14288 );
and \U$12563 ( \14351 , \14288 , \14323 );
and \U$12564 ( \14352 , \14286 , \14323 );
or \U$12565 ( \14353 , \14350 , \14351 , \14352 );
and \U$12567 ( \14354 , \13558 , \13164 );
nor \U$12568 ( \14355 , 1'b0 , \14354 );
xnor \U$12569 ( \14356 , \14355 , 1'b0 );
xor \U$12571 ( \14357 , \14356 , 1'b0 );
xor \U$12573 ( \14358 , \14357 , 1'b0 );
and \U$12574 ( \14359 , \13314 , \13238 );
and \U$12575 ( \14360 , \13270 , \13236 );
nor \U$12576 ( \14361 , \14359 , \14360 );
xnor \U$12577 ( \14362 , \14361 , \13243 );
and \U$12578 ( \14363 , \13407 , \13173 );
and \U$12579 ( \14364 , \13440 , \13171 );
nor \U$12580 ( \14365 , \14363 , \14364 );
xnor \U$12581 ( \14366 , \14365 , \12940 );
xor \U$12582 ( \14367 , \14362 , \14366 );
and \U$12583 ( \14368 , \13467 , \13111 );
and \U$12584 ( \14369 , \13500 , \13109 );
nor \U$12585 ( \14370 , \14368 , \14369 );
xnor \U$12586 ( \14371 , \14370 , \13137 );
xor \U$12587 ( \14372 , \14367 , \14371 );
xor \U$12588 ( \14373 , \14358 , \14372 );
not \U$12589 ( \14374 , \13445 );
and \U$12590 ( \14375 , \13063 , \13479 );
and \U$12591 ( \14376 , \13132 , \13477 );
nor \U$12592 ( \14377 , \14375 , \14376 );
xnor \U$12593 ( \14378 , \14377 , \13505 );
xor \U$12594 ( \14379 , \14374 , \14378 );
and \U$12595 ( \14380 , \13291 , \13537 );
and \U$12596 ( \14381 , \13159 , \13535 );
nor \U$12597 ( \14382 , \14380 , \14381 );
xnor \U$12598 ( \14383 , \14382 , \13563 );
xor \U$12599 ( \14384 , \14379 , \14383 );
xor \U$12600 ( \14385 , \14373 , \14384 );
xor \U$12602 ( \14386 , \14385 , 1'b0 );
and \U$12604 ( \14387 , \14316 , \14321 );
or \U$12606 ( \14388 , 1'b0 , \14387 , 1'b0 );
and \U$12607 ( \14389 , \14302 , \14306 );
and \U$12608 ( \14390 , \14306 , \14311 );
and \U$12609 ( \14391 , \14302 , \14311 );
or \U$12610 ( \14392 , \14389 , \14390 , \14391 );
xor \U$12611 ( \14393 , \14388 , \14392 );
and \U$12612 ( \14394 , \14293 , \14296 );
or \U$12615 ( \14395 , \14394 , 1'b0 , 1'b0 );
xor \U$12616 ( \14396 , \14393 , \14395 );
xor \U$12617 ( \14397 , \14386 , \14396 );
xor \U$12618 ( \14398 , \14353 , \14397 );
and \U$12619 ( \14399 , \14274 , \14278 );
and \U$12620 ( \14400 , \14278 , \14281 );
and \U$12621 ( \14401 , \14274 , \14281 );
or \U$12622 ( \14402 , \14399 , \14400 , \14401 );
xor \U$12624 ( \14403 , \14402 , 1'b0 );
and \U$12625 ( \14404 , \14298 , \14312 );
and \U$12626 ( \14405 , \14312 , \14322 );
and \U$12627 ( \14406 , \14298 , \14322 );
or \U$12628 ( \14407 , \14404 , \14405 , \14406 );
xor \U$12629 ( \14408 , \14403 , \14407 );
xor \U$12630 ( \14409 , \14398 , \14408 );
xor \U$12631 ( \14410 , \14349 , \14409 );
and \U$12632 ( \14411 , \14270 , \14325 );
and \U$12633 ( \14412 , \14325 , \14336 );
and \U$12634 ( \14413 , \14270 , \14336 );
or \U$12635 ( \14414 , \14411 , \14412 , \14413 );
nor \U$12636 ( \14415 , \14410 , \14414 );
and \U$12637 ( \14416 , \14353 , \14397 );
and \U$12638 ( \14417 , \14397 , \14408 );
and \U$12639 ( \14418 , \14353 , \14408 );
or \U$12640 ( \14419 , \14416 , \14417 , \14418 );
and \U$12641 ( \14420 , \14388 , \14392 );
and \U$12642 ( \14421 , \14392 , \14395 );
and \U$12643 ( \14422 , \14388 , \14395 );
or \U$12644 ( \14423 , \14420 , \14421 , \14422 );
xor \U$12646 ( \14424 , \14423 , 1'b0 );
and \U$12647 ( \14425 , \14358 , \14372 );
and \U$12648 ( \14426 , \14372 , \14384 );
and \U$12649 ( \14427 , \14358 , \14384 );
or \U$12650 ( \14428 , \14425 , \14426 , \14427 );
xor \U$12651 ( \14429 , \14424 , \14428 );
xor \U$12652 ( \14430 , \14419 , \14429 );
and \U$12655 ( \14431 , \14402 , \14407 );
or \U$12656 ( \14432 , 1'b0 , 1'b0 , \14431 );
and \U$12659 ( \14433 , \14385 , \14396 );
or \U$12660 ( \14434 , 1'b0 , 1'b0 , \14433 );
xor \U$12661 ( \14435 , \14432 , \14434 );
and \U$12662 ( \14436 , \13270 , \13238 );
and \U$12663 ( \14437 , \13291 , \13236 );
nor \U$12664 ( \14438 , \14436 , \14437 );
xnor \U$12665 ( \14439 , \14438 , \13243 );
and \U$12666 ( \14440 , \13440 , \13173 );
and \U$12667 ( \14441 , \13314 , \13171 );
nor \U$12668 ( \14442 , \14440 , \14441 );
xnor \U$12669 ( \14443 , \14442 , \12940 );
xor \U$12670 ( \14444 , \14439 , \14443 );
and \U$12671 ( \14445 , \13500 , \13111 );
and \U$12672 ( \14446 , \13407 , \13109 );
nor \U$12673 ( \14447 , \14445 , \14446 );
xnor \U$12674 ( \14448 , \14447 , \13137 );
xor \U$12675 ( \14449 , \14444 , \14448 );
and \U$12677 ( \14450 , \13132 , \13479 );
not \U$12678 ( \14451 , \14450 );
xnor \U$12679 ( \14452 , \14451 , \13505 );
xor \U$12680 ( \14453 , 1'b0 , \14452 );
and \U$12681 ( \14454 , \13159 , \13537 );
and \U$12682 ( \14455 , \13063 , \13535 );
nor \U$12683 ( \14456 , \14454 , \14455 );
xnor \U$12684 ( \14457 , \14456 , \13563 );
xor \U$12685 ( \14458 , \14453 , \14457 );
xor \U$12686 ( \14459 , \14449 , \14458 );
and \U$12689 ( \14460 , \13467 , \13164 );
nor \U$12690 ( \14461 , 1'b0 , \14460 );
xnor \U$12691 ( \14462 , \14461 , 1'b0 );
xor \U$12693 ( \14463 , \14462 , 1'b0 );
xor \U$12695 ( \14464 , \14463 , 1'b0 );
xnor \U$12696 ( \14465 , 1'b0 , \14464 );
xor \U$12697 ( \14466 , \14459 , \14465 );
and \U$12698 ( \14467 , \14374 , \14378 );
and \U$12699 ( \14468 , \14378 , \14383 );
and \U$12700 ( \14469 , \14374 , \14383 );
or \U$12701 ( \14470 , \14467 , \14468 , \14469 );
and \U$12702 ( \14471 , \14362 , \14366 );
and \U$12703 ( \14472 , \14366 , \14371 );
and \U$12704 ( \14473 , \14362 , \14371 );
or \U$12705 ( \14474 , \14471 , \14472 , \14473 );
xor \U$12706 ( \14475 , \14470 , \14474 );
xor \U$12708 ( \14476 , \14475 , 1'b0 );
xor \U$12709 ( \14477 , \14466 , \14476 );
xor \U$12710 ( \14478 , \14435 , \14477 );
xor \U$12711 ( \14479 , \14430 , \14478 );
and \U$12712 ( \14480 , \14347 , \14348 );
and \U$12713 ( \14481 , \14348 , \14409 );
and \U$12714 ( \14482 , \14347 , \14409 );
or \U$12715 ( \14483 , \14480 , \14481 , \14482 );
nor \U$12716 ( \14484 , \14479 , \14483 );
nor \U$12717 ( \14485 , \14415 , \14484 );
nand \U$12718 ( \14486 , \14343 , \14485 );
nor \U$12719 ( \14487 , \14191 , \14486 );
and \U$12720 ( \14488 , \14432 , \14434 );
and \U$12721 ( \14489 , \14434 , \14477 );
and \U$12722 ( \14490 , \14432 , \14477 );
or \U$12723 ( \14491 , \14488 , \14489 , \14490 );
and \U$12724 ( \14492 , \14470 , \14474 );
or \U$12727 ( \14493 , \14492 , 1'b0 , 1'b0 );
or \U$12728 ( \14494 , 1'b0 , \14464 );
xor \U$12729 ( \14495 , \14493 , \14494 );
and \U$12730 ( \14496 , \14449 , \14458 );
xor \U$12731 ( \14497 , \14495 , \14496 );
xor \U$12732 ( \14498 , \14491 , \14497 );
and \U$12735 ( \14499 , \14423 , \14428 );
or \U$12736 ( \14500 , 1'b0 , 1'b0 , \14499 );
and \U$12737 ( \14501 , \14459 , \14465 );
and \U$12738 ( \14502 , \14465 , \14476 );
and \U$12739 ( \14503 , \14459 , \14476 );
or \U$12740 ( \14504 , \14501 , \14502 , \14503 );
xor \U$12741 ( \14505 , \14500 , \14504 );
and \U$12743 ( \14506 , \13314 , \13173 );
and \U$12744 ( \14507 , \13270 , \13171 );
nor \U$12745 ( \14508 , \14506 , \14507 );
xnor \U$12746 ( \14509 , \14508 , \12940 );
and \U$12747 ( \14510 , \13407 , \13111 );
and \U$12748 ( \14511 , \13440 , \13109 );
nor \U$12749 ( \14512 , \14510 , \14511 );
xnor \U$12750 ( \14513 , \14512 , \13137 );
xor \U$12751 ( \14514 , \14509 , \14513 );
and \U$12753 ( \14515 , \13500 , \13164 );
nor \U$12754 ( \14516 , 1'b0 , \14515 );
xnor \U$12755 ( \14517 , \14516 , 1'b0 );
xor \U$12756 ( \14518 , \14514 , \14517 );
xor \U$12757 ( \14519 , 1'b0 , \14518 );
not \U$12758 ( \14520 , \13505 );
and \U$12759 ( \14521 , \13063 , \13537 );
and \U$12760 ( \14522 , \13132 , \13535 );
nor \U$12761 ( \14523 , \14521 , \14522 );
xnor \U$12762 ( \14524 , \14523 , \13563 );
xor \U$12763 ( \14525 , \14520 , \14524 );
and \U$12764 ( \14526 , \13291 , \13238 );
and \U$12765 ( \14527 , \13159 , \13236 );
nor \U$12766 ( \14528 , \14526 , \14527 );
xnor \U$12767 ( \14529 , \14528 , \13243 );
xor \U$12768 ( \14530 , \14525 , \14529 );
xor \U$12769 ( \14531 , \14519 , \14530 );
xor \U$12771 ( \14532 , \14531 , 1'b0 );
and \U$12773 ( \14533 , \14452 , \14457 );
or \U$12775 ( \14534 , 1'b0 , \14533 , 1'b0 );
and \U$12776 ( \14535 , \14439 , \14443 );
and \U$12777 ( \14536 , \14443 , \14448 );
and \U$12778 ( \14537 , \14439 , \14448 );
or \U$12779 ( \14538 , \14535 , \14536 , \14537 );
xor \U$12780 ( \14539 , \14534 , \14538 );
xor \U$12782 ( \14540 , \14539 , 1'b0 );
xor \U$12783 ( \14541 , \14532 , \14540 );
xor \U$12784 ( \14542 , \14505 , \14541 );
xor \U$12785 ( \14543 , \14498 , \14542 );
and \U$12786 ( \14544 , \14419 , \14429 );
and \U$12787 ( \14545 , \14429 , \14478 );
and \U$12788 ( \14546 , \14419 , \14478 );
or \U$12789 ( \14547 , \14544 , \14545 , \14546 );
nor \U$12790 ( \14548 , \14543 , \14547 );
and \U$12791 ( \14549 , \14500 , \14504 );
and \U$12792 ( \14550 , \14504 , \14541 );
and \U$12793 ( \14551 , \14500 , \14541 );
or \U$12794 ( \14552 , \14549 , \14550 , \14551 );
and \U$12795 ( \14553 , \14534 , \14538 );
or \U$12798 ( \14554 , \14553 , 1'b0 , 1'b0 );
xor \U$12800 ( \14555 , \14554 , 1'b0 );
and \U$12802 ( \14556 , \14518 , \14530 );
or \U$12804 ( \14557 , 1'b0 , \14556 , 1'b0 );
xor \U$12805 ( \14558 , \14555 , \14557 );
xor \U$12806 ( \14559 , \14552 , \14558 );
and \U$12807 ( \14560 , \14493 , \14494 );
and \U$12808 ( \14561 , \14494 , \14496 );
and \U$12809 ( \14562 , \14493 , \14496 );
or \U$12810 ( \14563 , \14560 , \14561 , \14562 );
and \U$12813 ( \14564 , \14531 , \14540 );
or \U$12814 ( \14565 , 1'b0 , 1'b0 , \14564 );
xor \U$12815 ( \14566 , \14563 , \14565 );
and \U$12816 ( \14567 , \13270 , \13173 );
and \U$12817 ( \14568 , \13291 , \13171 );
nor \U$12818 ( \14569 , \14567 , \14568 );
xnor \U$12819 ( \14570 , \14569 , \12940 );
and \U$12820 ( \14571 , \13440 , \13111 );
and \U$12821 ( \14572 , \13314 , \13109 );
nor \U$12822 ( \14573 , \14571 , \14572 );
xnor \U$12823 ( \14574 , \14573 , \13137 );
xor \U$12824 ( \14575 , \14570 , \14574 );
and \U$12826 ( \14576 , \13407 , \13164 );
nor \U$12827 ( \14577 , 1'b0 , \14576 );
xnor \U$12828 ( \14578 , \14577 , 1'b0 );
xor \U$12829 ( \14579 , \14575 , \14578 );
and \U$12831 ( \14580 , \13132 , \13537 );
not \U$12832 ( \14581 , \14580 );
xnor \U$12833 ( \14582 , \14581 , \13563 );
xor \U$12834 ( \14583 , 1'b0 , \14582 );
and \U$12835 ( \14584 , \13159 , \13238 );
and \U$12836 ( \14585 , \13063 , \13236 );
nor \U$12837 ( \14586 , \14584 , \14585 );
xnor \U$12838 ( \14587 , \14586 , \13243 );
xor \U$12839 ( \14588 , \14583 , \14587 );
xor \U$12840 ( \14589 , \14579 , \14588 );
xor \U$12842 ( \14590 , \14589 , 1'b1 );
and \U$12843 ( \14591 , \14520 , \14524 );
and \U$12844 ( \14592 , \14524 , \14529 );
and \U$12845 ( \14593 , \14520 , \14529 );
or \U$12846 ( \14594 , \14591 , \14592 , \14593 );
and \U$12847 ( \14595 , \14509 , \14513 );
and \U$12848 ( \14596 , \14513 , \14517 );
and \U$12849 ( \14597 , \14509 , \14517 );
or \U$12850 ( \14598 , \14595 , \14596 , \14597 );
xor \U$12851 ( \14599 , \14594 , \14598 );
xor \U$12853 ( \14600 , \14599 , 1'b0 );
xor \U$12854 ( \14601 , \14590 , \14600 );
xor \U$12855 ( \14602 , \14566 , \14601 );
xor \U$12856 ( \14603 , \14559 , \14602 );
and \U$12857 ( \14604 , \14491 , \14497 );
and \U$12858 ( \14605 , \14497 , \14542 );
and \U$12859 ( \14606 , \14491 , \14542 );
or \U$12860 ( \14607 , \14604 , \14605 , \14606 );
nor \U$12861 ( \14608 , \14603 , \14607 );
nor \U$12862 ( \14609 , \14548 , \14608 );
and \U$12863 ( \14610 , \14563 , \14565 );
and \U$12864 ( \14611 , \14565 , \14601 );
and \U$12865 ( \14612 , \14563 , \14601 );
or \U$12866 ( \14613 , \14610 , \14611 , \14612 );
and \U$12867 ( \14614 , \14594 , \14598 );
or \U$12870 ( \14615 , \14614 , 1'b0 , 1'b0 );
xor \U$12872 ( \14616 , \14615 , 1'b0 );
and \U$12873 ( \14617 , \14579 , \14588 );
xor \U$12874 ( \14618 , \14616 , \14617 );
xor \U$12875 ( \14619 , \14613 , \14618 );
and \U$12878 ( \14620 , \14554 , \14557 );
or \U$12879 ( \14621 , 1'b0 , 1'b0 , \14620 );
and \U$12880 ( \14622 , \14589 , 1'b1 );
and \U$12881 ( \14623 , 1'b1 , \14600 );
and \U$12882 ( \14624 , \14589 , \14600 );
or \U$12883 ( \14625 , \14622 , \14623 , \14624 );
xor \U$12884 ( \14626 , \14621 , \14625 );
and \U$12886 ( \14627 , \13314 , \13111 );
and \U$12887 ( \14628 , \13270 , \13109 );
nor \U$12888 ( \14629 , \14627 , \14628 );
xnor \U$12889 ( \14630 , \14629 , \13137 );
and \U$12891 ( \14631 , \13440 , \13164 );
nor \U$12892 ( \14632 , 1'b0 , \14631 );
xnor \U$12893 ( \14633 , \14632 , 1'b0 );
xor \U$12894 ( \14634 , \14630 , \14633 );
xor \U$12896 ( \14635 , \14634 , 1'b0 );
xor \U$12897 ( \14636 , 1'b0 , \14635 );
not \U$12898 ( \14637 , \13563 );
and \U$12899 ( \14638 , \13063 , \13238 );
and \U$12900 ( \14639 , \13132 , \13236 );
nor \U$12901 ( \14640 , \14638 , \14639 );
xnor \U$12902 ( \14641 , \14640 , \13243 );
xor \U$12903 ( \14642 , \14637 , \14641 );
and \U$12904 ( \14643 , \13291 , \13173 );
and \U$12905 ( \14644 , \13159 , \13171 );
nor \U$12906 ( \14645 , \14643 , \14644 );
xnor \U$12907 ( \14646 , \14645 , \12940 );
xor \U$12908 ( \14647 , \14642 , \14646 );
xor \U$12909 ( \14648 , \14636 , \14647 );
xor \U$12911 ( \14649 , \14648 , 1'b0 );
and \U$12913 ( \14650 , \14582 , \14587 );
or \U$12915 ( \14651 , 1'b0 , \14650 , 1'b0 );
and \U$12916 ( \14652 , \14570 , \14574 );
and \U$12917 ( \14653 , \14574 , \14578 );
and \U$12918 ( \14654 , \14570 , \14578 );
or \U$12919 ( \14655 , \14652 , \14653 , \14654 );
xor \U$12920 ( \14656 , \14651 , \14655 );
xor \U$12922 ( \14657 , \14656 , 1'b0 );
xor \U$12923 ( \14658 , \14649 , \14657 );
xor \U$12924 ( \14659 , \14626 , \14658 );
xor \U$12925 ( \14660 , \14619 , \14659 );
and \U$12926 ( \14661 , \14552 , \14558 );
and \U$12927 ( \14662 , \14558 , \14602 );
and \U$12928 ( \14663 , \14552 , \14602 );
or \U$12929 ( \14664 , \14661 , \14662 , \14663 );
nor \U$12930 ( \14665 , \14660 , \14664 );
and \U$12931 ( \14666 , \14621 , \14625 );
and \U$12932 ( \14667 , \14625 , \14658 );
and \U$12933 ( \14668 , \14621 , \14658 );
or \U$12934 ( \14669 , \14666 , \14667 , \14668 );
and \U$12935 ( \14670 , \14651 , \14655 );
or \U$12938 ( \14671 , \14670 , 1'b0 , 1'b0 );
xor \U$12940 ( \14672 , \14671 , 1'b0 );
and \U$12942 ( \14673 , \14635 , \14647 );
or \U$12944 ( \14674 , 1'b0 , \14673 , 1'b0 );
xor \U$12945 ( \14675 , \14672 , \14674 );
xor \U$12946 ( \14676 , \14669 , \14675 );
and \U$12949 ( \14677 , \14615 , \14617 );
or \U$12950 ( \14678 , 1'b0 , 1'b0 , \14677 );
and \U$12953 ( \14679 , \14648 , \14657 );
or \U$12954 ( \14680 , 1'b0 , 1'b0 , \14679 );
xor \U$12955 ( \14681 , \14678 , \14680 );
xor \U$12956 ( \14682 , \13294 , \13317 );
xor \U$12958 ( \14683 , \14682 , 1'b0 );
xor \U$12960 ( \14684 , 1'b0 , \13244 );
xor \U$12961 ( \14685 , \14684 , \13248 );
xor \U$12962 ( \14686 , \14683 , \14685 );
xor \U$12964 ( \14687 , \14686 , 1'b1 );
and \U$12965 ( \14688 , \14637 , \14641 );
and \U$12966 ( \14689 , \14641 , \14646 );
and \U$12967 ( \14690 , \14637 , \14646 );
or \U$12968 ( \14691 , \14688 , \14689 , \14690 );
and \U$12969 ( \14692 , \14630 , \14633 );
or \U$12972 ( \14693 , \14692 , 1'b0 , 1'b0 );
xor \U$12973 ( \14694 , \14691 , \14693 );
xor \U$12975 ( \14695 , \14694 , 1'b0 );
xor \U$12976 ( \14696 , \14687 , \14695 );
xor \U$12977 ( \14697 , \14681 , \14696 );
xor \U$12978 ( \14698 , \14676 , \14697 );
and \U$12979 ( \14699 , \14613 , \14618 );
and \U$12980 ( \14700 , \14618 , \14659 );
and \U$12981 ( \14701 , \14613 , \14659 );
or \U$12982 ( \14702 , \14699 , \14700 , \14701 );
nor \U$12983 ( \14703 , \14698 , \14702 );
nor \U$12984 ( \14704 , \14665 , \14703 );
nand \U$12985 ( \14705 , \14609 , \14704 );
and \U$12986 ( \14706 , \14678 , \14680 );
and \U$12987 ( \14707 , \14680 , \14696 );
and \U$12988 ( \14708 , \14678 , \14696 );
or \U$12989 ( \14709 , \14706 , \14707 , \14708 );
and \U$12990 ( \14710 , \14691 , \14693 );
or \U$12993 ( \14711 , \14710 , 1'b0 , 1'b0 );
xor \U$12995 ( \14712 , \14711 , 1'b0 );
and \U$12996 ( \14713 , \14683 , \14685 );
xor \U$12997 ( \14714 , \14712 , \14713 );
xor \U$12998 ( \14715 , \14709 , \14714 );
and \U$13001 ( \14716 , \14671 , \14674 );
or \U$13002 ( \14717 , 1'b0 , 1'b0 , \14716 );
and \U$13003 ( \14718 , \14686 , 1'b1 );
and \U$13004 ( \14719 , 1'b1 , \14695 );
and \U$13005 ( \14720 , \14686 , \14695 );
or \U$13006 ( \14721 , \14718 , \14719 , \14720 );
xor \U$13007 ( \14722 , \14717 , \14721 );
xor \U$13009 ( \14723 , 1'b0 , \13326 );
xor \U$13010 ( \14724 , \14723 , \13337 );
xor \U$13012 ( \14725 , \14724 , 1'b0 );
xor \U$13013 ( \14726 , \13250 , \13319 );
xor \U$13015 ( \14727 , \14726 , 1'b0 );
xor \U$13016 ( \14728 , \14725 , \14727 );
xor \U$13017 ( \14729 , \14722 , \14728 );
xor \U$13018 ( \14730 , \14715 , \14729 );
and \U$13019 ( \14731 , \14669 , \14675 );
and \U$13020 ( \14732 , \14675 , \14697 );
and \U$13021 ( \14733 , \14669 , \14697 );
or \U$13022 ( \14734 , \14731 , \14732 , \14733 );
nor \U$13023 ( \14735 , \14730 , \14734 );
and \U$13024 ( \14736 , \14717 , \14721 );
and \U$13025 ( \14737 , \14721 , \14728 );
and \U$13026 ( \14738 , \14717 , \14728 );
or \U$13027 ( \14739 , \14736 , \14737 , \14738 );
xor \U$13029 ( \14740 , \13321 , 1'b0 );
xor \U$13030 ( \14741 , \14740 , \13339 );
xor \U$13031 ( \14742 , \14739 , \14741 );
and \U$13034 ( \14743 , \14711 , \14713 );
or \U$13035 ( \14744 , 1'b0 , 1'b0 , \14743 );
and \U$13038 ( \14745 , \14724 , \14727 );
or \U$13039 ( \14746 , 1'b0 , 1'b0 , \14745 );
xor \U$13040 ( \14747 , \14744 , \14746 );
xor \U$13041 ( \14748 , \13349 , 1'b1 );
xor \U$13042 ( \14749 , \14748 , \13356 );
xor \U$13043 ( \14750 , \14747 , \14749 );
xor \U$13044 ( \14751 , \14742 , \14750 );
and \U$13045 ( \14752 , \14709 , \14714 );
and \U$13046 ( \14753 , \14714 , \14729 );
and \U$13047 ( \14754 , \14709 , \14729 );
or \U$13048 ( \14755 , \14752 , \14753 , \14754 );
nor \U$13049 ( \14756 , \14751 , \14755 );
nor \U$13050 ( \14757 , \14735 , \14756 );
and \U$13051 ( \14758 , \14744 , \14746 );
and \U$13052 ( \14759 , \14746 , \14749 );
and \U$13053 ( \14760 , \14744 , \14749 );
or \U$13054 ( \14761 , \14758 , \14759 , \14760 );
and \U$13056 ( \14762 , \13346 , \13348 );
xor \U$13057 ( \14763 , 1'b0 , \14762 );
xor \U$13058 ( \14764 , \14761 , \14763 );
xor \U$13059 ( \14765 , \13341 , \13359 );
xor \U$13060 ( \14766 , \14765 , \13362 );
xor \U$13061 ( \14767 , \14764 , \14766 );
and \U$13062 ( \14768 , \14739 , \14741 );
and \U$13063 ( \14769 , \14741 , \14750 );
and \U$13064 ( \14770 , \14739 , \14750 );
or \U$13065 ( \14771 , \14768 , \14769 , \14770 );
nor \U$13066 ( \14772 , \14767 , \14771 );
xor \U$13068 ( \14773 , \13365 , 1'b0 );
xor \U$13069 ( \14774 , \14773 , \13367 );
and \U$13070 ( \14775 , \14761 , \14763 );
and \U$13071 ( \14776 , \14763 , \14766 );
and \U$13072 ( \14777 , \14761 , \14766 );
or \U$13073 ( \14778 , \14775 , \14776 , \14777 );
nor \U$13074 ( \14779 , \14774 , \14778 );
nor \U$13075 ( \14780 , \14772 , \14779 );
nand \U$13076 ( \14781 , \14757 , \14780 );
nor \U$13077 ( \14782 , \14705 , \14781 );
nand \U$13078 ( \14783 , \14487 , \14782 );
and \U$13079 ( \14784 , \13584 , \13383 );
and \U$13080 ( \14785 , \13605 , \13380 );
nor \U$13081 ( \14786 , \14784 , \14785 );
xnor \U$13082 ( \14787 , \14786 , \13377 );
and \U$13083 ( \14788 , \13629 , \13419 );
and \U$13084 ( \14789 , \13650 , \13417 );
nor \U$13085 ( \14790 , \14788 , \14789 );
xnor \U$13086 ( \14791 , \14790 , \13445 );
and \U$13087 ( \14792 , \14787 , \14791 );
and \U$13088 ( \14793 , \13677 , \13479 );
and \U$13089 ( \14794 , \13698 , \13477 );
nor \U$13090 ( \14795 , \14793 , \14794 );
xnor \U$13091 ( \14796 , \14795 , \13505 );
and \U$13092 ( \14797 , \14791 , \14796 );
and \U$13093 ( \14798 , \14787 , \14796 );
or \U$13094 ( \14799 , \14792 , \14797 , \14798 );
and \U$13095 ( \14800 , \13698 , \13479 );
and \U$13096 ( \14801 , \13629 , \13477 );
nor \U$13097 ( \14802 , \14800 , \14801 );
xnor \U$13098 ( \14803 , \14802 , \13505 );
and \U$13099 ( \14804 , \13721 , \13537 );
and \U$13100 ( \14805 , \13677 , \13535 );
nor \U$13101 ( \14806 , \14804 , \14805 );
xnor \U$13102 ( \14807 , \14806 , \13563 );
xor \U$13103 ( \14808 , \14803 , \14807 );
nand \U$13104 ( \14809 , \13854 , \13236 );
xnor \U$13105 ( \14810 , \14809 , \13243 );
xor \U$13106 ( \14811 , \14808 , \14810 );
and \U$13107 ( \14812 , \14799 , \14811 );
and \U$13108 ( \14813 , \13605 , \13383 );
and \U$13109 ( \14814 , \13529 , \13380 );
nor \U$13110 ( \14815 , \14813 , \14814 );
xnor \U$13111 ( \14816 , \14815 , \13377 );
xor \U$13112 ( \14817 , \13243 , \14816 );
and \U$13113 ( \14818 , \13650 , \13419 );
and \U$13114 ( \14819 , \13584 , \13417 );
nor \U$13115 ( \14820 , \14818 , \14819 );
xnor \U$13116 ( \14821 , \14820 , \13445 );
xor \U$13117 ( \14822 , \14817 , \14821 );
and \U$13118 ( \14823 , \14811 , \14822 );
and \U$13119 ( \14824 , \14799 , \14822 );
or \U$13120 ( \14825 , \14812 , \14823 , \14824 );
and \U$13121 ( \14826 , \13854 , \13238 );
and \U$13122 ( \14827 , \13721 , \13236 );
nor \U$13123 ( \14828 , \14826 , \14827 );
xnor \U$13124 ( \14829 , \14828 , \13243 );
and \U$13125 ( \14830 , \13529 , \13383 );
and \U$13126 ( \14831 , \13558 , \13380 );
nor \U$13127 ( \14832 , \14830 , \14831 );
xnor \U$13128 ( \14833 , \14832 , \13377 );
and \U$13129 ( \14834 , \13584 , \13419 );
and \U$13130 ( \14835 , \13605 , \13417 );
nor \U$13131 ( \14836 , \14834 , \14835 );
xnor \U$13132 ( \14837 , \14836 , \13445 );
xor \U$13133 ( \14838 , \14833 , \14837 );
and \U$13134 ( \14839 , \13629 , \13479 );
and \U$13135 ( \14840 , \13650 , \13477 );
nor \U$13136 ( \14841 , \14839 , \14840 );
xnor \U$13137 ( \14842 , \14841 , \13505 );
xor \U$13138 ( \14843 , \14838 , \14842 );
xor \U$13139 ( \14844 , \14829 , \14843 );
xor \U$13140 ( \14845 , \14825 , \14844 );
and \U$13141 ( \14846 , \13243 , \14816 );
and \U$13142 ( \14847 , \14816 , \14821 );
and \U$13143 ( \14848 , \13243 , \14821 );
or \U$13144 ( \14849 , \14846 , \14847 , \14848 );
and \U$13145 ( \14850 , \14803 , \14807 );
and \U$13146 ( \14851 , \14807 , \14810 );
and \U$13147 ( \14852 , \14803 , \14810 );
or \U$13148 ( \14853 , \14850 , \14851 , \14852 );
xor \U$13149 ( \14854 , \14849 , \14853 );
and \U$13150 ( \14855 , \13677 , \13537 );
and \U$13151 ( \14856 , \13698 , \13535 );
nor \U$13152 ( \14857 , \14855 , \14856 );
xnor \U$13153 ( \14858 , \14857 , \13563 );
xor \U$13154 ( \14859 , \14854 , \14858 );
xor \U$13155 ( \14860 , \14845 , \14859 );
and \U$13156 ( \14861 , \13650 , \13383 );
and \U$13157 ( \14862 , \13584 , \13380 );
nor \U$13158 ( \14863 , \14861 , \14862 );
xnor \U$13159 ( \14864 , \14863 , \13377 );
and \U$13160 ( \14865 , \13563 , \14864 );
and \U$13161 ( \14866 , \13698 , \13419 );
and \U$13162 ( \14867 , \13629 , \13417 );
nor \U$13163 ( \14868 , \14866 , \14867 );
xnor \U$13164 ( \14869 , \14868 , \13445 );
and \U$13165 ( \14870 , \14864 , \14869 );
and \U$13166 ( \14871 , \13563 , \14869 );
or \U$13167 ( \14872 , \14865 , \14870 , \14871 );
and \U$13168 ( \14873 , \13721 , \13479 );
and \U$13169 ( \14874 , \13677 , \13477 );
nor \U$13170 ( \14875 , \14873 , \14874 );
xnor \U$13171 ( \14876 , \14875 , \13505 );
nand \U$13172 ( \14877 , \13854 , \13535 );
xnor \U$13173 ( \14878 , \14877 , \13563 );
and \U$13174 ( \14879 , \14876 , \14878 );
and \U$13175 ( \14880 , \14872 , \14879 );
and \U$13176 ( \14881 , \13854 , \13537 );
and \U$13177 ( \14882 , \13721 , \13535 );
nor \U$13178 ( \14883 , \14881 , \14882 );
xnor \U$13179 ( \14884 , \14883 , \13563 );
and \U$13180 ( \14885 , \14879 , \14884 );
and \U$13181 ( \14886 , \14872 , \14884 );
or \U$13182 ( \14887 , \14880 , \14885 , \14886 );
xor \U$13183 ( \14888 , \14799 , \14811 );
xor \U$13184 ( \14889 , \14888 , \14822 );
and \U$13185 ( \14890 , \14887 , \14889 );
nor \U$13186 ( \14891 , \14860 , \14890 );
and \U$13187 ( \14892 , \14833 , \14837 );
and \U$13188 ( \14893 , \14837 , \14842 );
and \U$13189 ( \14894 , \14833 , \14842 );
or \U$13190 ( \14895 , \14892 , \14893 , \14894 );
nand \U$13191 ( \14896 , \13854 , \13171 );
xnor \U$13192 ( \14897 , \14896 , \12940 );
xor \U$13193 ( \14898 , \14895 , \14897 );
and \U$13194 ( \14899 , \13650 , \13479 );
and \U$13195 ( \14900 , \13584 , \13477 );
nor \U$13196 ( \14901 , \14899 , \14900 );
xnor \U$13197 ( \14902 , \14901 , \13505 );
and \U$13198 ( \14903 , \13698 , \13537 );
and \U$13199 ( \14904 , \13629 , \13535 );
nor \U$13200 ( \14905 , \14903 , \14904 );
xnor \U$13201 ( \14906 , \14905 , \13563 );
xor \U$13202 ( \14907 , \14902 , \14906 );
and \U$13203 ( \14908 , \13721 , \13238 );
and \U$13204 ( \14909 , \13677 , \13236 );
nor \U$13205 ( \14910 , \14908 , \14909 );
xnor \U$13206 ( \14911 , \14910 , \13243 );
xor \U$13207 ( \14912 , \14907 , \14911 );
xor \U$13208 ( \14913 , \14898 , \14912 );
and \U$13209 ( \14914 , \14849 , \14853 );
and \U$13210 ( \14915 , \14853 , \14858 );
and \U$13211 ( \14916 , \14849 , \14858 );
or \U$13212 ( \14917 , \14914 , \14915 , \14916 );
and \U$13213 ( \14918 , \14829 , \14843 );
xor \U$13214 ( \14919 , \14917 , \14918 );
and \U$13215 ( \14920 , \13558 , \13383 );
and \U$13216 ( \14921 , \13467 , \13380 );
nor \U$13217 ( \14922 , \14920 , \14921 );
xnor \U$13218 ( \14923 , \14922 , \13377 );
xor \U$13219 ( \14924 , \12940 , \14923 );
and \U$13220 ( \14925 , \13605 , \13419 );
and \U$13221 ( \14926 , \13529 , \13417 );
nor \U$13222 ( \14927 , \14925 , \14926 );
xnor \U$13223 ( \14928 , \14927 , \13445 );
xor \U$13224 ( \14929 , \14924 , \14928 );
xor \U$13225 ( \14930 , \14919 , \14929 );
xor \U$13226 ( \14931 , \14913 , \14930 );
and \U$13227 ( \14932 , \14825 , \14844 );
and \U$13228 ( \14933 , \14844 , \14859 );
and \U$13229 ( \14934 , \14825 , \14859 );
or \U$13230 ( \14935 , \14932 , \14933 , \14934 );
nor \U$13231 ( \14936 , \14931 , \14935 );
nor \U$13232 ( \14937 , \14891 , \14936 );
and \U$13233 ( \14938 , \14917 , \14918 );
and \U$13234 ( \14939 , \14918 , \14929 );
and \U$13235 ( \14940 , \14917 , \14929 );
or \U$13236 ( \14941 , \14938 , \14939 , \14940 );
and \U$13237 ( \14942 , \14895 , \14897 );
and \U$13238 ( \14943 , \14897 , \14912 );
and \U$13239 ( \14944 , \14895 , \14912 );
or \U$13240 ( \14945 , \14942 , \14943 , \14944 );
and \U$13241 ( \14946 , \13467 , \13383 );
and \U$13242 ( \14947 , \13500 , \13380 );
nor \U$13243 ( \14948 , \14946 , \14947 );
xnor \U$13244 ( \14949 , \14948 , \13377 );
and \U$13245 ( \14950 , \13529 , \13419 );
and \U$13246 ( \14951 , \13558 , \13417 );
nor \U$13247 ( \14952 , \14950 , \14951 );
xnor \U$13248 ( \14953 , \14952 , \13445 );
xor \U$13249 ( \14954 , \14949 , \14953 );
and \U$13250 ( \14955 , \13584 , \13479 );
and \U$13251 ( \14956 , \13605 , \13477 );
nor \U$13252 ( \14957 , \14955 , \14956 );
xnor \U$13253 ( \14958 , \14957 , \13505 );
xor \U$13254 ( \14959 , \14954 , \14958 );
xor \U$13255 ( \14960 , \14945 , \14959 );
and \U$13256 ( \14961 , \12940 , \14923 );
and \U$13257 ( \14962 , \14923 , \14928 );
and \U$13258 ( \14963 , \12940 , \14928 );
or \U$13259 ( \14964 , \14961 , \14962 , \14963 );
and \U$13260 ( \14965 , \14902 , \14906 );
and \U$13261 ( \14966 , \14906 , \14911 );
and \U$13262 ( \14967 , \14902 , \14911 );
or \U$13263 ( \14968 , \14965 , \14966 , \14967 );
xor \U$13264 ( \14969 , \14964 , \14968 );
and \U$13265 ( \14970 , \13629 , \13537 );
and \U$13266 ( \14971 , \13650 , \13535 );
nor \U$13267 ( \14972 , \14970 , \14971 );
xnor \U$13268 ( \14973 , \14972 , \13563 );
and \U$13269 ( \14974 , \13677 , \13238 );
and \U$13270 ( \14975 , \13698 , \13236 );
nor \U$13271 ( \14976 , \14974 , \14975 );
xnor \U$13272 ( \14977 , \14976 , \13243 );
xor \U$13273 ( \14978 , \14973 , \14977 );
and \U$13274 ( \14979 , \13854 , \13173 );
and \U$13275 ( \14980 , \13721 , \13171 );
nor \U$13276 ( \14981 , \14979 , \14980 );
xnor \U$13277 ( \14982 , \14981 , \12940 );
xor \U$13278 ( \14983 , \14978 , \14982 );
xor \U$13279 ( \14984 , \14969 , \14983 );
xor \U$13280 ( \14985 , \14960 , \14984 );
xor \U$13281 ( \14986 , \14941 , \14985 );
and \U$13282 ( \14987 , \14913 , \14930 );
nor \U$13283 ( \14988 , \14986 , \14987 );
and \U$13284 ( \14989 , \14945 , \14959 );
and \U$13285 ( \14990 , \14959 , \14984 );
and \U$13286 ( \14991 , \14945 , \14984 );
or \U$13287 ( \14992 , \14989 , \14990 , \14991 );
and \U$13288 ( \14993 , \14964 , \14968 );
and \U$13289 ( \14994 , \14968 , \14983 );
and \U$13290 ( \14995 , \14964 , \14983 );
or \U$13291 ( \14996 , \14993 , \14994 , \14995 );
nand \U$13292 ( \14997 , \13854 , \13109 );
xnor \U$13293 ( \14998 , \14997 , \13137 );
and \U$13294 ( \14999 , \13605 , \13479 );
and \U$13295 ( \15000 , \13529 , \13477 );
nor \U$13296 ( \15001 , \14999 , \15000 );
xnor \U$13297 ( \15002 , \15001 , \13505 );
and \U$13298 ( \15003 , \13650 , \13537 );
and \U$13299 ( \15004 , \13584 , \13535 );
nor \U$13300 ( \15005 , \15003 , \15004 );
xnor \U$13301 ( \15006 , \15005 , \13563 );
xor \U$13302 ( \15007 , \15002 , \15006 );
and \U$13303 ( \15008 , \13698 , \13238 );
and \U$13304 ( \15009 , \13629 , \13236 );
nor \U$13305 ( \15010 , \15008 , \15009 );
xnor \U$13306 ( \15011 , \15010 , \13243 );
xor \U$13307 ( \15012 , \15007 , \15011 );
xor \U$13308 ( \15013 , \14998 , \15012 );
and \U$13309 ( \15014 , \13500 , \13383 );
and \U$13310 ( \15015 , \13407 , \13380 );
nor \U$13311 ( \15016 , \15014 , \15015 );
xnor \U$13312 ( \15017 , \15016 , \13377 );
xor \U$13313 ( \15018 , \13137 , \15017 );
and \U$13314 ( \15019 , \13558 , \13419 );
and \U$13315 ( \15020 , \13467 , \13417 );
nor \U$13316 ( \15021 , \15019 , \15020 );
xnor \U$13317 ( \15022 , \15021 , \13445 );
xor \U$13318 ( \15023 , \15018 , \15022 );
xor \U$13319 ( \15024 , \15013 , \15023 );
xor \U$13320 ( \15025 , \14996 , \15024 );
and \U$13321 ( \15026 , \14949 , \14953 );
and \U$13322 ( \15027 , \14953 , \14958 );
and \U$13323 ( \15028 , \14949 , \14958 );
or \U$13324 ( \15029 , \15026 , \15027 , \15028 );
and \U$13325 ( \15030 , \14973 , \14977 );
and \U$13326 ( \15031 , \14977 , \14982 );
and \U$13327 ( \15032 , \14973 , \14982 );
or \U$13328 ( \15033 , \15030 , \15031 , \15032 );
xor \U$13329 ( \15034 , \15029 , \15033 );
and \U$13330 ( \15035 , \13721 , \13173 );
and \U$13331 ( \15036 , \13677 , \13171 );
nor \U$13332 ( \15037 , \15035 , \15036 );
xnor \U$13333 ( \15038 , \15037 , \12940 );
xor \U$13334 ( \15039 , \15034 , \15038 );
xor \U$13335 ( \15040 , \15025 , \15039 );
xor \U$13336 ( \15041 , \14992 , \15040 );
and \U$13337 ( \15042 , \14941 , \14985 );
nor \U$13338 ( \15043 , \15041 , \15042 );
nor \U$13339 ( \15044 , \14988 , \15043 );
nand \U$13340 ( \15045 , \14937 , \15044 );
and \U$13341 ( \15046 , \14996 , \15024 );
and \U$13342 ( \15047 , \15024 , \15039 );
and \U$13343 ( \15048 , \14996 , \15039 );
or \U$13344 ( \15049 , \15046 , \15047 , \15048 );
xor \U$13345 ( \15050 , \13909 , \13913 );
xor \U$13346 ( \15051 , \15050 , \13918 );
and \U$13347 ( \15052 , \13137 , \15017 );
and \U$13348 ( \15053 , \15017 , \15022 );
and \U$13349 ( \15054 , \13137 , \15022 );
or \U$13350 ( \15055 , \15052 , \15053 , \15054 );
and \U$13351 ( \15056 , \15002 , \15006 );
and \U$13352 ( \15057 , \15006 , \15011 );
and \U$13353 ( \15058 , \15002 , \15011 );
or \U$13354 ( \15059 , \15056 , \15057 , \15058 );
xor \U$13355 ( \15060 , \15055 , \15059 );
and \U$13356 ( \15061 , \13854 , \13111 );
and \U$13357 ( \15062 , \13721 , \13109 );
nor \U$13358 ( \15063 , \15061 , \15062 );
xnor \U$13359 ( \15064 , \15063 , \13137 );
xor \U$13360 ( \15065 , \15060 , \15064 );
xor \U$13361 ( \15066 , \15051 , \15065 );
xor \U$13362 ( \15067 , \15049 , \15066 );
and \U$13363 ( \15068 , \15029 , \15033 );
and \U$13364 ( \15069 , \15033 , \15038 );
and \U$13365 ( \15070 , \15029 , \15038 );
or \U$13366 ( \15071 , \15068 , \15069 , \15070 );
and \U$13367 ( \15072 , \14998 , \15012 );
and \U$13368 ( \15073 , \15012 , \15023 );
and \U$13369 ( \15074 , \14998 , \15023 );
or \U$13370 ( \15075 , \15072 , \15073 , \15074 );
xor \U$13371 ( \15076 , \15071 , \15075 );
xor \U$13372 ( \15077 , \13925 , \13929 );
xor \U$13373 ( \15078 , \15077 , \13934 );
xor \U$13374 ( \15079 , \15076 , \15078 );
xor \U$13375 ( \15080 , \15067 , \15079 );
and \U$13376 ( \15081 , \14992 , \15040 );
nor \U$13377 ( \15082 , \15080 , \15081 );
and \U$13378 ( \15083 , \15071 , \15075 );
and \U$13379 ( \15084 , \15075 , \15078 );
and \U$13380 ( \15085 , \15071 , \15078 );
or \U$13381 ( \15086 , \15083 , \15084 , \15085 );
and \U$13382 ( \15087 , \15051 , \15065 );
xor \U$13383 ( \15088 , \15086 , \15087 );
and \U$13384 ( \15089 , \15055 , \15059 );
and \U$13385 ( \15090 , \15059 , \15064 );
and \U$13386 ( \15091 , \15055 , \15064 );
or \U$13387 ( \15092 , \15089 , \15090 , \15091 );
xor \U$13388 ( \15093 , \13945 , \13947 );
xor \U$13389 ( \15094 , \15092 , \15093 );
xor \U$13390 ( \15095 , \13921 , \13937 );
xor \U$13391 ( \15096 , \15095 , \13940 );
xor \U$13392 ( \15097 , \15094 , \15096 );
xor \U$13393 ( \15098 , \15088 , \15097 );
and \U$13394 ( \15099 , \15049 , \15066 );
and \U$13395 ( \15100 , \15066 , \15079 );
and \U$13396 ( \15101 , \15049 , \15079 );
or \U$13397 ( \15102 , \15099 , \15100 , \15101 );
nor \U$13398 ( \15103 , \15098 , \15102 );
nor \U$13399 ( \15104 , \15082 , \15103 );
and \U$13400 ( \15105 , \15092 , \15093 );
and \U$13401 ( \15106 , \15093 , \15096 );
and \U$13402 ( \15107 , \15092 , \15096 );
or \U$13403 ( \15108 , \15105 , \15106 , \15107 );
xor \U$13404 ( \15109 , \13808 , \13824 );
xor \U$13405 ( \15110 , \15109 , \13859 );
xor \U$13406 ( \15111 , \15108 , \15110 );
xor \U$13407 ( \15112 , \13943 , \13948 );
xor \U$13408 ( \15113 , \15112 , \13951 );
xor \U$13409 ( \15114 , \15111 , \15113 );
and \U$13410 ( \15115 , \15086 , \15087 );
and \U$13411 ( \15116 , \15087 , \15097 );
and \U$13412 ( \15117 , \15086 , \15097 );
or \U$13413 ( \15118 , \15115 , \15116 , \15117 );
nor \U$13414 ( \15119 , \15114 , \15118 );
xor \U$13415 ( \15120 , \13954 , \13955 );
xor \U$13416 ( \15121 , \15120 , \13958 );
and \U$13417 ( \15122 , \15108 , \15110 );
and \U$13418 ( \15123 , \15110 , \15113 );
and \U$13419 ( \15124 , \15108 , \15113 );
or \U$13420 ( \15125 , \15122 , \15123 , \15124 );
nor \U$13421 ( \15126 , \15121 , \15125 );
nor \U$13422 ( \15127 , \15119 , \15126 );
nand \U$13423 ( \15128 , \15104 , \15127 );
nor \U$13424 ( \15129 , \15045 , \15128 );
and \U$13425 ( \15130 , \13698 , \13383 );
and \U$13426 ( \15131 , \13629 , \13380 );
nor \U$13427 ( \15132 , \15130 , \15131 );
xnor \U$13428 ( \15133 , \15132 , \13377 );
and \U$13429 ( \15134 , \13505 , \15133 );
and \U$13430 ( \15135 , \13721 , \13419 );
and \U$13431 ( \15136 , \13677 , \13417 );
nor \U$13432 ( \15137 , \15135 , \15136 );
xnor \U$13433 ( \15138 , \15137 , \13445 );
and \U$13434 ( \15139 , \15133 , \15138 );
and \U$13435 ( \15140 , \13505 , \15138 );
or \U$13436 ( \15141 , \15134 , \15139 , \15140 );
and \U$13437 ( \15142 , \13629 , \13383 );
and \U$13438 ( \15143 , \13650 , \13380 );
nor \U$13439 ( \15144 , \15142 , \15143 );
xnor \U$13440 ( \15145 , \15144 , \13377 );
and \U$13441 ( \15146 , \13677 , \13419 );
and \U$13442 ( \15147 , \13698 , \13417 );
nor \U$13443 ( \15148 , \15146 , \15147 );
xnor \U$13444 ( \15149 , \15148 , \13445 );
xor \U$13445 ( \15150 , \15145 , \15149 );
and \U$13446 ( \15151 , \13854 , \13479 );
and \U$13447 ( \15152 , \13721 , \13477 );
nor \U$13448 ( \15153 , \15151 , \15152 );
xnor \U$13449 ( \15154 , \15153 , \13505 );
xor \U$13450 ( \15155 , \15150 , \15154 );
xor \U$13451 ( \15156 , \15141 , \15155 );
nand \U$13452 ( \15157 , \13854 , \13477 );
xnor \U$13453 ( \15158 , \15157 , \13505 );
xor \U$13454 ( \15159 , \13505 , \15133 );
xor \U$13455 ( \15160 , \15159 , \15138 );
and \U$13456 ( \15161 , \15158 , \15160 );
nor \U$13457 ( \15162 , \15156 , \15161 );
and \U$13458 ( \15163 , \15145 , \15149 );
and \U$13459 ( \15164 , \15149 , \15154 );
and \U$13460 ( \15165 , \15145 , \15154 );
or \U$13461 ( \15166 , \15163 , \15164 , \15165 );
xor \U$13462 ( \15167 , \14876 , \14878 );
xor \U$13463 ( \15168 , \15166 , \15167 );
xor \U$13464 ( \15169 , \13563 , \14864 );
xor \U$13465 ( \15170 , \15169 , \14869 );
xor \U$13466 ( \15171 , \15168 , \15170 );
and \U$13467 ( \15172 , \15141 , \15155 );
nor \U$13468 ( \15173 , \15171 , \15172 );
nor \U$13469 ( \15174 , \15162 , \15173 );
xor \U$13470 ( \15175 , \14787 , \14791 );
xor \U$13471 ( \15176 , \15175 , \14796 );
xor \U$13472 ( \15177 , \14872 , \14879 );
xor \U$13473 ( \15178 , \15177 , \14884 );
xor \U$13474 ( \15179 , \15176 , \15178 );
and \U$13475 ( \15180 , \15166 , \15167 );
and \U$13476 ( \15181 , \15167 , \15170 );
and \U$13477 ( \15182 , \15166 , \15170 );
or \U$13478 ( \15183 , \15180 , \15181 , \15182 );
nor \U$13479 ( \15184 , \15179 , \15183 );
xor \U$13480 ( \15185 , \14887 , \14889 );
and \U$13481 ( \15186 , \15176 , \15178 );
nor \U$13482 ( \15187 , \15185 , \15186 );
nor \U$13483 ( \15188 , \15184 , \15187 );
nand \U$13484 ( \15189 , \15174 , \15188 );
and \U$13485 ( \15190 , \13677 , \13383 );
and \U$13486 ( \15191 , \13698 , \13380 );
nor \U$13487 ( \15192 , \15190 , \15191 );
xnor \U$13488 ( \15193 , \15192 , \13377 );
and \U$13489 ( \15194 , \13854 , \13419 );
and \U$13490 ( \15195 , \13721 , \13417 );
nor \U$13491 ( \15196 , \15194 , \15195 );
xnor \U$13492 ( \15197 , \15196 , \13445 );
xor \U$13493 ( \15198 , \15193 , \15197 );
and \U$13494 ( \15199 , \13721 , \13383 );
and \U$13495 ( \15200 , \13677 , \13380 );
nor \U$13496 ( \15201 , \15199 , \15200 );
xnor \U$13497 ( \15202 , \15201 , \13377 );
and \U$13498 ( \15203 , \15202 , \13445 );
nor \U$13499 ( \15204 , \15198 , \15203 );
xor \U$13500 ( \15205 , \15158 , \15160 );
and \U$13501 ( \15206 , \15193 , \15197 );
nor \U$13502 ( \15207 , \15205 , \15206 );
nor \U$13503 ( \15208 , \15204 , \15207 );
xor \U$13504 ( \15209 , \15202 , \13445 );
nand \U$13505 ( \15210 , \13854 , \13417 );
xnor \U$13506 ( \15211 , \15210 , \13445 );
nor \U$13507 ( \15212 , \15209 , \15211 );
and \U$13508 ( \15213 , \13854 , \13383 );
and \U$13509 ( \15214 , \13721 , \13380 );
nor \U$13510 ( \15215 , \15213 , \15214 );
xnor \U$13511 ( \15216 , \15215 , \13377 );
nand \U$13512 ( \15217 , \13854 , \13380 );
xnor \U$13513 ( \15218 , \15217 , \13377 );
and \U$13514 ( \15219 , \15218 , \13377 );
nand \U$13515 ( \15220 , \15216 , \15219 );
or \U$13516 ( \15221 , \15212 , \15220 );
nand \U$13517 ( \15222 , \15209 , \15211 );
nand \U$13518 ( \15223 , \15221 , \15222 );
and \U$13519 ( \15224 , \15208 , \15223 );
nand \U$13520 ( \15225 , \15198 , \15203 );
or \U$13521 ( \15226 , \15207 , \15225 );
nand \U$13522 ( \15227 , \15205 , \15206 );
nand \U$13523 ( \15228 , \15226 , \15227 );
nor \U$13524 ( \15229 , \15224 , \15228 );
or \U$13525 ( \15230 , \15189 , \15229 );
nand \U$13526 ( \15231 , \15156 , \15161 );
or \U$13527 ( \15232 , \15173 , \15231 );
nand \U$13528 ( \15233 , \15171 , \15172 );
nand \U$13529 ( \15234 , \15232 , \15233 );
and \U$13530 ( \15235 , \15188 , \15234 );
nand \U$13531 ( \15236 , \15179 , \15183 );
or \U$13532 ( \15237 , \15187 , \15236 );
nand \U$13533 ( \15238 , \15185 , \15186 );
nand \U$13534 ( \15239 , \15237 , \15238 );
nor \U$13535 ( \15240 , \15235 , \15239 );
nand \U$13536 ( \15241 , \15230 , \15240 );
and \U$13537 ( \15242 , \15129 , \15241 );
nand \U$13538 ( \15243 , \14860 , \14890 );
or \U$13539 ( \15244 , \14936 , \15243 );
nand \U$13540 ( \15245 , \14931 , \14935 );
nand \U$13541 ( \15246 , \15244 , \15245 );
and \U$13542 ( \15247 , \15044 , \15246 );
nand \U$13543 ( \15248 , \14986 , \14987 );
or \U$13544 ( \15249 , \15043 , \15248 );
nand \U$13545 ( \15250 , \15041 , \15042 );
nand \U$13546 ( \15251 , \15249 , \15250 );
nor \U$13547 ( \15252 , \15247 , \15251 );
or \U$13548 ( \15253 , \15128 , \15252 );
nand \U$13549 ( \15254 , \15080 , \15081 );
or \U$13550 ( \15255 , \15103 , \15254 );
nand \U$13551 ( \15256 , \15098 , \15102 );
nand \U$13552 ( \15257 , \15255 , \15256 );
and \U$13553 ( \15258 , \15127 , \15257 );
nand \U$13554 ( \15259 , \15114 , \15118 );
or \U$13555 ( \15260 , \15126 , \15259 );
nand \U$13556 ( \15261 , \15121 , \15125 );
nand \U$13557 ( \15262 , \15260 , \15261 );
nor \U$13558 ( \15263 , \15258 , \15262 );
nand \U$13559 ( \15264 , \15253 , \15263 );
nor \U$13560 ( \15265 , \15242 , \15264 );
or \U$13561 ( \15266 , \14783 , \15265 );
nand \U$13562 ( \15267 , \13905 , \13961 );
or \U$13563 ( \15268 , \14037 , \15267 );
nand \U$13564 ( \15269 , \14035 , \14036 );
nand \U$13565 ( \15270 , \15268 , \15269 );
and \U$13566 ( \15271 , \14190 , \15270 );
nand \U$13567 ( \15272 , \14112 , \14113 );
or \U$13568 ( \15273 , \14189 , \15272 );
nand \U$13569 ( \15274 , \14184 , \14188 );
nand \U$13570 ( \15275 , \15273 , \15274 );
nor \U$13571 ( \15276 , \15271 , \15275 );
or \U$13572 ( \15277 , \14486 , \15276 );
nand \U$13573 ( \15278 , \14261 , \14265 );
or \U$13574 ( \15279 , \14342 , \15278 );
nand \U$13575 ( \15280 , \14337 , \14341 );
nand \U$13576 ( \15281 , \15279 , \15280 );
and \U$13577 ( \15282 , \14485 , \15281 );
nand \U$13578 ( \15283 , \14410 , \14414 );
or \U$13579 ( \15284 , \14484 , \15283 );
nand \U$13580 ( \15285 , \14479 , \14483 );
nand \U$13581 ( \15286 , \15284 , \15285 );
nor \U$13582 ( \15287 , \15282 , \15286 );
nand \U$13583 ( \15288 , \15277 , \15287 );
and \U$13584 ( \15289 , \14782 , \15288 );
nand \U$13585 ( \15290 , \14543 , \14547 );
or \U$13586 ( \15291 , \14608 , \15290 );
nand \U$13587 ( \15292 , \14603 , \14607 );
nand \U$13588 ( \15293 , \15291 , \15292 );
and \U$13589 ( \15294 , \14704 , \15293 );
nand \U$13590 ( \15295 , \14660 , \14664 );
or \U$13591 ( \15296 , \14703 , \15295 );
nand \U$13592 ( \15297 , \14698 , \14702 );
nand \U$13593 ( \15298 , \15296 , \15297 );
nor \U$13594 ( \15299 , \15294 , \15298 );
or \U$13595 ( \15300 , \14781 , \15299 );
nand \U$13596 ( \15301 , \14730 , \14734 );
or \U$13597 ( \15302 , \14756 , \15301 );
nand \U$13598 ( \15303 , \14751 , \14755 );
nand \U$13599 ( \15304 , \15302 , \15303 );
and \U$13600 ( \15305 , \14780 , \15304 );
nand \U$13601 ( \15306 , \14767 , \14771 );
or \U$13602 ( \15307 , \14779 , \15306 );
nand \U$13603 ( \15308 , \14774 , \14778 );
nand \U$13604 ( \15309 , \15307 , \15308 );
nor \U$13605 ( \15310 , \15305 , \15309 );
nand \U$13606 ( \15311 , \15300 , \15310 );
nor \U$13607 ( \15312 , \15289 , \15311 );
nand \U$13608 ( \15313 , \15266 , \15312 );
not \U$13609 ( \15314 , \15313 );
xor \U$13610 ( \15315 , \13373 , \15314 );
buf g4ba0_GF_PartitionCandidate( \15316_nG4ba0 , \15315 );
buf \U$13611 ( \15317 , RI995f0f8_1);
buf \U$13612 ( \15318 , RI995f080_2);
buf \U$13613 ( \15319 , RI995f008_3);
buf \U$13614 ( \15320 , RI995ef90_4);
buf \U$13615 ( \15321 , RI995ef18_5);
buf \U$13616 ( \15322 , RI995eea0_6);
buf \U$13617 ( \15323 , RI995ee28_7);
buf \U$13618 ( \15324 , RI995edb0_8);
buf \U$13619 ( \15325 , RI995ed38_9);
buf \U$13620 ( \15326 , RI995ecc0_10);
buf \U$13621 ( \15327 , RI995ec48_11);
buf \U$13622 ( \15328 , RI995ebd0_12);
not \U$13623 ( \15329 , RI99216b8_614);
buf \U$13624 ( \15330 , \15329 );
and \U$13625 ( \15331 , \15328 , \15330 );
and \U$13626 ( \15332 , \15327 , \15331 );
and \U$13627 ( \15333 , \15326 , \15332 );
and \U$13628 ( \15334 , \15325 , \15333 );
and \U$13629 ( \15335 , \15324 , \15334 );
and \U$13630 ( \15336 , \15323 , \15335 );
and \U$13631 ( \15337 , \15322 , \15336 );
and \U$13632 ( \15338 , \15321 , \15337 );
and \U$13633 ( \15339 , \15320 , \15338 );
and \U$13634 ( \15340 , \15319 , \15339 );
and \U$13635 ( \15341 , \15318 , \15340 );
xor \U$13636 ( \15342 , \15317 , \15341 );
buf \U$13637 ( \15343 , \15342 );
buf \U$13638 ( \15344 , \15343 );
not \U$13639 ( \15345 , \15344 );
nor \U$13640 ( \15346 , \12513 , \12517 , \12521 , \12525 , \12530 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13641 ( \15347 , RI995e4c8_235, \15346 );
nor \U$13642 ( \15348 , \12565 , \12566 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13643 ( \15349 , RI99670f0_222, \15348 );
nor \U$13644 ( \15350 , \12513 , \12566 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13645 ( \15351 , RI890f600_209, \15350 );
nor \U$13646 ( \15352 , \12565 , \12517 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13647 ( \15353 , RI89185e8_196, \15352 );
nor \U$13648 ( \15354 , \12513 , \12517 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13649 ( \15355 , RI8924e10_183, \15354 );
nor \U$13650 ( \15356 , \12565 , \12566 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13651 ( \15357 , RI8930828_170, \15356 );
nor \U$13652 ( \15358 , \12513 , \12566 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13653 ( \15359 , RI8939810_157, \15358 );
nor \U$13654 ( \15360 , \12565 , \12517 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13655 ( \15361 , RI8946038_144, \15360 );
nor \U$13656 ( \15362 , \12513 , \12517 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13657 ( \15363 , RI89ec0a0_131, \15362 );
nor \U$13658 ( \15364 , \12565 , \12566 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13659 ( \15365 , RI89ec6b8_118, \15364 );
nor \U$13660 ( \15366 , \12513 , \12566 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13661 ( \15367 , RI9776ff8_105, \15366 );
nor \U$13662 ( \15368 , \12565 , \12517 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13663 ( \15369 , RI98084f8_92, \15368 );
nor \U$13664 ( \15370 , \12513 , \12517 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13665 ( \15371 , RI9808b10_79, \15370 );
nor \U$13666 ( \15372 , \12565 , \12566 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13667 ( \15373 , RI98197a8_66, \15372 );
nor \U$13668 ( \15374 , \12513 , \12566 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13669 ( \15375 , RI98abcb0_53, \15374 );
nor \U$13670 ( \15376 , \12565 , \12517 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13671 ( \15377 , RI98bc948_40, \15376 );
nor \U$13672 ( \15378 , \12513 , \12517 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$13673 ( \15379 , RI994de48_27, \15378 );
or \U$13674 ( \15380 , \15347 , \15349 , \15351 , \15353 , \15355 , \15357 , \15359 , \15361 , \15363 , \15365 , \15367 , \15369 , \15371 , \15373 , \15375 , \15377 , \15379 );
buf \U$13675 ( \15381 , \12534 );
buf \U$13676 ( \15382 , \12538 );
buf \U$13677 ( \15383 , \12542 );
buf \U$13678 ( \15384 , \12546 );
buf \U$13679 ( \15385 , \12550 );
buf \U$13680 ( \15386 , \12554 );
buf \U$13681 ( \15387 , \12558 );
buf \U$13682 ( \15388 , \12562 );
buf \U$13683 ( \15389 , \12529 );
buf \U$13684 ( \15390 , \12513 );
buf \U$13685 ( \15391 , \12517 );
buf \U$13686 ( \15392 , \12521 );
buf \U$13687 ( \15393 , \12525 );
or \U$13688 ( \15394 , \15390 , \15391 , \15392 , \15393 );
and \U$13689 ( \15395 , \15389 , \15394 );
or \U$13690 ( \15396 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15395 );
buf \U$13691 ( \15397 , \15396 );
_DC g1512 ( \15398_nG1512 , \15380 , \15397 );
buf \U$13692 ( \15399 , \15398_nG1512 );
and \U$13693 ( \15400 , \15345 , \15399 );
xor \U$13694 ( \15401 , \15318 , \15340 );
buf \U$13695 ( \15402 , \15401 );
buf \U$13696 ( \15403 , \15402 );
not \U$13697 ( \15404 , \15403 );
and \U$13698 ( \15405 , RI995e450_236, \15346 );
and \U$13699 ( \15406 , RI9967078_223, \15348 );
and \U$13700 ( \15407 , RI9967690_210, \15350 );
and \U$13701 ( \15408 , RI890fba0_197, \15352 );
and \U$13702 ( \15409 , RI8918b88_184, \15354 );
and \U$13703 ( \15410 , RI89253b0_171, \15356 );
and \U$13704 ( \15411 , RI8930dc8_158, \15358 );
and \U$13705 ( \15412 , RI8939db0_145, \15360 );
and \U$13706 ( \15413 , RI89465d8_132, \15362 );
and \U$13707 ( \15414 , RI89ec640_119, \15364 );
and \U$13708 ( \15415 , RI9776f80_106, \15366 );
and \U$13709 ( \15416 , RI9808480_93, \15368 );
and \U$13710 ( \15417 , RI9808a98_80, \15370 );
and \U$13711 ( \15418 , RI9819730_67, \15372 );
and \U$13712 ( \15419 , RI98abc38_54, \15374 );
and \U$13713 ( \15420 , RI98bc8d0_41, \15376 );
and \U$13714 ( \15421 , RI994ddd0_28, \15378 );
or \U$13715 ( \15422 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 );
_DC g152b ( \15423_nG152b , \15422 , \15397 );
buf \U$13716 ( \15424 , \15423_nG152b );
and \U$13717 ( \15425 , \15404 , \15424 );
xor \U$13718 ( \15426 , \15319 , \15339 );
buf \U$13719 ( \15427 , \15426 );
buf \U$13720 ( \15428 , \15427 );
not \U$13721 ( \15429 , \15428 );
and \U$13722 ( \15430 , RI995e3d8_237, \15346 );
and \U$13723 ( \15431 , RI99669e8_224, \15348 );
and \U$13724 ( \15432 , RI9967618_211, \15350 );
and \U$13725 ( \15433 , RI890fb28_198, \15352 );
and \U$13726 ( \15434 , RI8918b10_185, \15354 );
and \U$13727 ( \15435 , RI8925338_172, \15356 );
and \U$13728 ( \15436 , RI8930d50_159, \15358 );
and \U$13729 ( \15437 , RI8939d38_146, \15360 );
and \U$13730 ( \15438 , RI8946560_133, \15362 );
and \U$13731 ( \15439 , RI89ec5c8_120, \15364 );
and \U$13732 ( \15440 , RI9776f08_107, \15366 );
and \U$13733 ( \15441 , RI9808408_94, \15368 );
and \U$13734 ( \15442 , RI9808a20_81, \15370 );
and \U$13735 ( \15443 , RI98196b8_68, \15372 );
and \U$13736 ( \15444 , RI98abbc0_55, \15374 );
and \U$13737 ( \15445 , RI98bc858_42, \15376 );
and \U$13738 ( \15446 , RI994dd58_29, \15378 );
or \U$13739 ( \15447 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 );
_DC g1544 ( \15448_nG1544 , \15447 , \15397 );
buf \U$13740 ( \15449 , \15448_nG1544 );
and \U$13741 ( \15450 , \15429 , \15449 );
xor \U$13742 ( \15451 , \15320 , \15338 );
buf \U$13743 ( \15452 , \15451 );
buf \U$13744 ( \15453 , \15452 );
not \U$13745 ( \15454 , \15453 );
and \U$13746 ( \15455 , RI9959fe0_238, \15346 );
and \U$13747 ( \15456 , RI995e978_225, \15348 );
and \U$13748 ( \15457 , RI99675a0_212, \15350 );
and \U$13749 ( \15458 , RI890fab0_199, \15352 );
and \U$13750 ( \15459 , RI8918a98_186, \15354 );
and \U$13751 ( \15460 , RI89252c0_173, \15356 );
and \U$13752 ( \15461 , RI8930cd8_160, \15358 );
and \U$13753 ( \15462 , RI8939cc0_147, \15360 );
and \U$13754 ( \15463 , RI89464e8_134, \15362 );
and \U$13755 ( \15464 , RI89ec550_121, \15364 );
and \U$13756 ( \15465 , RI9776e90_108, \15366 );
and \U$13757 ( \15466 , RI9808390_95, \15368 );
and \U$13758 ( \15467 , RI98089a8_82, \15370 );
and \U$13759 ( \15468 , RI9819640_69, \15372 );
and \U$13760 ( \15469 , RI98abb48_56, \15374 );
and \U$13761 ( \15470 , RI98bc7e0_43, \15376 );
and \U$13762 ( \15471 , RI994dce0_30, \15378 );
or \U$13763 ( \15472 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 );
_DC g155d ( \15473_nG155d , \15472 , \15397 );
buf \U$13764 ( \15474 , \15473_nG155d );
and \U$13765 ( \15475 , \15454 , \15474 );
xor \U$13766 ( \15476 , \15321 , \15337 );
buf \U$13767 ( \15477 , \15476 );
buf \U$13768 ( \15478 , \15477 );
not \U$13769 ( \15479 , \15478 );
and \U$13770 ( \15480 , RI9959f68_239, \15346 );
and \U$13771 ( \15481 , RI995e900_226, \15348 );
and \U$13772 ( \15482 , RI9967528_213, \15350 );
and \U$13773 ( \15483 , RI890fa38_200, \15352 );
and \U$13774 ( \15484 , RI8918a20_187, \15354 );
and \U$13775 ( \15485 , RI8925248_174, \15356 );
and \U$13776 ( \15486 , RI8930c60_161, \15358 );
and \U$13777 ( \15487 , RI8939c48_148, \15360 );
and \U$13778 ( \15488 , RI8946470_135, \15362 );
and \U$13779 ( \15489 , RI89ec4d8_122, \15364 );
and \U$13780 ( \15490 , RI9776e18_109, \15366 );
and \U$13781 ( \15491 , RI9808318_96, \15368 );
and \U$13782 ( \15492 , RI9808930_83, \15370 );
and \U$13783 ( \15493 , RI98195c8_70, \15372 );
and \U$13784 ( \15494 , RI98abad0_57, \15374 );
and \U$13785 ( \15495 , RI98bc768_44, \15376 );
and \U$13786 ( \15496 , RI994dc68_31, \15378 );
or \U$13787 ( \15497 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 );
_DC g1576 ( \15498_nG1576 , \15497 , \15397 );
buf \U$13788 ( \15499 , \15498_nG1576 );
and \U$13789 ( \15500 , \15479 , \15499 );
xor \U$13790 ( \15501 , \15322 , \15336 );
buf \U$13791 ( \15502 , \15501 );
buf \U$13792 ( \15503 , \15502 );
not \U$13793 ( \15504 , \15503 );
and \U$13794 ( \15505 , RI9959860_240, \15346 );
and \U$13795 ( \15506 , RI995e888_227, \15348 );
and \U$13796 ( \15507 , RI99674b0_214, \15350 );
and \U$13797 ( \15508 , RI890f9c0_201, \15352 );
and \U$13798 ( \15509 , RI89189a8_188, \15354 );
and \U$13799 ( \15510 , RI89251d0_175, \15356 );
and \U$13800 ( \15511 , RI8930be8_162, \15358 );
and \U$13801 ( \15512 , RI8939bd0_149, \15360 );
and \U$13802 ( \15513 , RI89463f8_136, \15362 );
and \U$13803 ( \15514 , RI89ec460_123, \15364 );
and \U$13804 ( \15515 , RI9776da0_110, \15366 );
and \U$13805 ( \15516 , RI98082a0_97, \15368 );
and \U$13806 ( \15517 , RI98088b8_84, \15370 );
and \U$13807 ( \15518 , RI9819550_71, \15372 );
and \U$13808 ( \15519 , RI98aba58_58, \15374 );
and \U$13809 ( \15520 , RI98bc6f0_45, \15376 );
and \U$13810 ( \15521 , RI994dbf0_32, \15378 );
or \U$13811 ( \15522 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 );
_DC g158f ( \15523_nG158f , \15522 , \15397 );
buf \U$13812 ( \15524 , \15523_nG158f );
and \U$13813 ( \15525 , \15504 , \15524 );
xor \U$13814 ( \15526 , \15323 , \15335 );
buf \U$13815 ( \15527 , \15526 );
buf \U$13816 ( \15528 , \15527 );
not \U$13817 ( \15529 , \15528 );
and \U$13818 ( \15530 , RI994d998_241, \15346 );
and \U$13819 ( \15531 , RI995e810_228, \15348 );
and \U$13820 ( \15532 , RI9967438_215, \15350 );
and \U$13821 ( \15533 , RI890f948_202, \15352 );
and \U$13822 ( \15534 , RI8918930_189, \15354 );
and \U$13823 ( \15535 , RI8925158_176, \15356 );
and \U$13824 ( \15536 , RI8930b70_163, \15358 );
and \U$13825 ( \15537 , RI8939b58_150, \15360 );
and \U$13826 ( \15538 , RI8946380_137, \15362 );
and \U$13827 ( \15539 , RI89ec3e8_124, \15364 );
and \U$13828 ( \15540 , RI9776d28_111, \15366 );
and \U$13829 ( \15541 , RI9808228_98, \15368 );
and \U$13830 ( \15542 , RI9808840_85, \15370 );
and \U$13831 ( \15543 , RI98194d8_72, \15372 );
and \U$13832 ( \15544 , RI98ab9e0_59, \15374 );
and \U$13833 ( \15545 , RI98abff8_46, \15376 );
and \U$13834 ( \15546 , RI98bcc90_33, \15378 );
or \U$13835 ( \15547 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 );
_DC g15a8 ( \15548_nG15a8 , \15547 , \15397 );
buf \U$13836 ( \15549 , \15548_nG15a8 );
and \U$13837 ( \15550 , \15529 , \15549 );
xor \U$13838 ( \15551 , \15324 , \15334 );
buf \U$13839 ( \15552 , \15551 );
buf \U$13840 ( \15553 , \15552 );
not \U$13841 ( \15554 , \15553 );
and \U$13842 ( \15555 , RI994d920_242, \15346 );
and \U$13843 ( \15556 , RI995e798_229, \15348 );
and \U$13844 ( \15557 , RI99673c0_216, \15350 );
and \U$13845 ( \15558 , RI890f8d0_203, \15352 );
and \U$13846 ( \15559 , RI89188b8_190, \15354 );
and \U$13847 ( \15560 , RI89250e0_177, \15356 );
and \U$13848 ( \15561 , RI8930af8_164, \15358 );
and \U$13849 ( \15562 , RI8939ae0_151, \15360 );
and \U$13850 ( \15563 , RI8946308_138, \15362 );
and \U$13851 ( \15564 , RI89ec370_125, \15364 );
and \U$13852 ( \15565 , RI89ec988_112, \15366 );
and \U$13853 ( \15566 , RI97772c8_99, \15368 );
and \U$13854 ( \15567 , RI98087c8_86, \15370 );
and \U$13855 ( \15568 , RI9819460_73, \15372 );
and \U$13856 ( \15569 , RI98ab968_60, \15374 );
and \U$13857 ( \15570 , RI98abf80_47, \15376 );
and \U$13858 ( \15571 , RI98bcc18_34, \15378 );
or \U$13859 ( \15572 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 );
_DC g15c1 ( \15573_nG15c1 , \15572 , \15397 );
buf \U$13860 ( \15574 , \15573_nG15c1 );
and \U$13861 ( \15575 , \15554 , \15574 );
xor \U$13862 ( \15576 , \15325 , \15333 );
buf \U$13863 ( \15577 , \15576 );
buf \U$13864 ( \15578 , \15577 );
not \U$13865 ( \15579 , \15578 );
and \U$13866 ( \15580 , RI994d8a8_243, \15346 );
and \U$13867 ( \15581 , RI995e720_230, \15348 );
and \U$13868 ( \15582 , RI9967348_217, \15350 );
and \U$13869 ( \15583 , RI890f858_204, \15352 );
and \U$13870 ( \15584 , RI8918840_191, \15354 );
and \U$13871 ( \15585 , RI8925068_178, \15356 );
and \U$13872 ( \15586 , RI8930a80_165, \15358 );
and \U$13873 ( \15587 , RI8939a68_152, \15360 );
and \U$13874 ( \15588 , RI8946290_139, \15362 );
and \U$13875 ( \15589 , RI89ec2f8_126, \15364 );
and \U$13876 ( \15590 , RI89ec910_113, \15366 );
and \U$13877 ( \15591 , RI9777250_100, \15368 );
and \U$13878 ( \15592 , RI9808750_87, \15370 );
and \U$13879 ( \15593 , RI98193e8_74, \15372 );
and \U$13880 ( \15594 , RI98ab8f0_61, \15374 );
and \U$13881 ( \15595 , RI98abf08_48, \15376 );
and \U$13882 ( \15596 , RI98bcba0_35, \15378 );
or \U$13883 ( \15597 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 );
_DC g15da ( \15598_nG15da , \15597 , \15397 );
buf \U$13884 ( \15599 , \15598_nG15da );
and \U$13885 ( \15600 , \15579 , \15599 );
xor \U$13886 ( \15601 , \15326 , \15332 );
buf \U$13887 ( \15602 , \15601 );
buf \U$13888 ( \15603 , \15602 );
not \U$13889 ( \15604 , \15603 );
and \U$13890 ( \15605 , RI994d830_244, \15346 );
and \U$13891 ( \15606 , RI995e6a8_231, \15348 );
and \U$13892 ( \15607 , RI99672d0_218, \15350 );
and \U$13893 ( \15608 , RI890f7e0_205, \15352 );
and \U$13894 ( \15609 , RI89187c8_192, \15354 );
and \U$13895 ( \15610 , RI8924ff0_179, \15356 );
and \U$13896 ( \15611 , RI8930a08_166, \15358 );
and \U$13897 ( \15612 , RI89399f0_153, \15360 );
and \U$13898 ( \15613 , RI8946218_140, \15362 );
and \U$13899 ( \15614 , RI89ec280_127, \15364 );
and \U$13900 ( \15615 , RI89ec898_114, \15366 );
and \U$13901 ( \15616 , RI97771d8_101, \15368 );
and \U$13902 ( \15617 , RI98086d8_88, \15370 );
and \U$13903 ( \15618 , RI9819370_75, \15372 );
and \U$13904 ( \15619 , RI98ab878_62, \15374 );
and \U$13905 ( \15620 , RI98abe90_49, \15376 );
and \U$13906 ( \15621 , RI98bcb28_36, \15378 );
or \U$13907 ( \15622 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 );
_DC g15f3 ( \15623_nG15f3 , \15622 , \15397 );
buf \U$13908 ( \15624 , \15623_nG15f3 );
and \U$13909 ( \15625 , \15604 , \15624 );
xor \U$13910 ( \15626 , \15327 , \15331 );
buf \U$13911 ( \15627 , \15626 );
buf \U$13912 ( \15628 , \15627 );
not \U$13913 ( \15629 , \15628 );
and \U$13914 ( \15630 , RI994d7b8_245, \15346 );
and \U$13915 ( \15631 , RI995e630_232, \15348 );
and \U$13916 ( \15632 , RI9967258_219, \15350 );
and \U$13917 ( \15633 , RI890f768_206, \15352 );
and \U$13918 ( \15634 , RI8918750_193, \15354 );
and \U$13919 ( \15635 , RI8924f78_180, \15356 );
and \U$13920 ( \15636 , RI8930990_167, \15358 );
and \U$13921 ( \15637 , RI8939978_154, \15360 );
and \U$13922 ( \15638 , RI89461a0_141, \15362 );
and \U$13923 ( \15639 , RI89ec208_128, \15364 );
and \U$13924 ( \15640 , RI89ec820_115, \15366 );
and \U$13925 ( \15641 , RI9777160_102, \15368 );
and \U$13926 ( \15642 , RI9808660_89, \15370 );
and \U$13927 ( \15643 , RI98192f8_76, \15372 );
and \U$13928 ( \15644 , RI98ab800_63, \15374 );
and \U$13929 ( \15645 , RI98abe18_50, \15376 );
and \U$13930 ( \15646 , RI98bcab0_37, \15378 );
or \U$13931 ( \15647 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 );
_DC g160c ( \15648_nG160c , \15647 , \15397 );
buf \U$13932 ( \15649 , \15648_nG160c );
and \U$13933 ( \15650 , \15629 , \15649 );
xor \U$13934 ( \15651 , \15328 , \15330 );
buf \U$13935 ( \15652 , \15651 );
buf \U$13936 ( \15653 , \15652 );
not \U$13937 ( \15654 , \15653 );
and \U$13938 ( \15655 , RI994d740_246, \15346 );
and \U$13939 ( \15656 , RI995e5b8_233, \15348 );
and \U$13940 ( \15657 , RI99671e0_220, \15350 );
and \U$13941 ( \15658 , RI890f6f0_207, \15352 );
and \U$13942 ( \15659 , RI89186d8_194, \15354 );
and \U$13943 ( \15660 , RI8924f00_181, \15356 );
and \U$13944 ( \15661 , RI8930918_168, \15358 );
and \U$13945 ( \15662 , RI8939900_155, \15360 );
and \U$13946 ( \15663 , RI8946128_142, \15362 );
and \U$13947 ( \15664 , RI89ec190_129, \15364 );
and \U$13948 ( \15665 , RI89ec7a8_116, \15366 );
and \U$13949 ( \15666 , RI97770e8_103, \15368 );
and \U$13950 ( \15667 , RI98085e8_90, \15370 );
and \U$13951 ( \15668 , RI9819280_77, \15372 );
and \U$13952 ( \15669 , RI98ab788_64, \15374 );
and \U$13953 ( \15670 , RI98abda0_51, \15376 );
and \U$13954 ( \15671 , RI98bca38_38, \15378 );
or \U$13955 ( \15672 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 );
_DC g1625 ( \15673_nG1625 , \15672 , \15397 );
buf \U$13956 ( \15674 , \15673_nG1625 );
and \U$13957 ( \15675 , \15654 , \15674 );
buf \U$13958 ( \15676 , RI994e4d8_13);
buf \U$13961 ( \15677 , \15676 );
not \U$13962 ( \15678 , \15677 );
and \U$13963 ( \15679 , RI994d6c8_247, \15346 );
and \U$13964 ( \15680 , RI995e540_234, \15348 );
and \U$13965 ( \15681 , RI9967168_221, \15350 );
and \U$13966 ( \15682 , RI890f678_208, \15352 );
and \U$13967 ( \15683 , RI8918660_195, \15354 );
and \U$13968 ( \15684 , RI8924e88_182, \15356 );
and \U$13969 ( \15685 , RI89308a0_169, \15358 );
and \U$13970 ( \15686 , RI8939888_156, \15360 );
and \U$13971 ( \15687 , RI89460b0_143, \15362 );
and \U$13972 ( \15688 , RI89ec118_130, \15364 );
and \U$13973 ( \15689 , RI89ec730_117, \15366 );
and \U$13974 ( \15690 , RI9777070_104, \15368 );
and \U$13975 ( \15691 , RI9808570_91, \15370 );
and \U$13976 ( \15692 , RI9819208_78, \15372 );
and \U$13977 ( \15693 , RI98ab710_65, \15374 );
and \U$13978 ( \15694 , RI98abd28_52, \15376 );
and \U$13979 ( \15695 , RI98bc9c0_39, \15378 );
or \U$13980 ( \15696 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 );
_DC g163f ( \15697_nG163f , \15696 , \15397 );
buf \U$13981 ( \15698 , \15697_nG163f );
and \U$13982 ( \15699 , \15678 , \15698 );
xnor \U$13983 ( \15700 , \15653 , \15674 );
and \U$13984 ( \15701 , \15699 , \15700 );
or \U$13985 ( \15702 , \15675 , \15701 );
xnor \U$13986 ( \15703 , \15628 , \15649 );
and \U$13987 ( \15704 , \15702 , \15703 );
or \U$13988 ( \15705 , \15650 , \15704 );
xnor \U$13989 ( \15706 , \15603 , \15624 );
and \U$13990 ( \15707 , \15705 , \15706 );
or \U$13991 ( \15708 , \15625 , \15707 );
xnor \U$13992 ( \15709 , \15578 , \15599 );
and \U$13993 ( \15710 , \15708 , \15709 );
or \U$13994 ( \15711 , \15600 , \15710 );
xnor \U$13995 ( \15712 , \15553 , \15574 );
and \U$13996 ( \15713 , \15711 , \15712 );
or \U$13997 ( \15714 , \15575 , \15713 );
xnor \U$13998 ( \15715 , \15528 , \15549 );
and \U$13999 ( \15716 , \15714 , \15715 );
or \U$14000 ( \15717 , \15550 , \15716 );
xnor \U$14001 ( \15718 , \15503 , \15524 );
and \U$14002 ( \15719 , \15717 , \15718 );
or \U$14003 ( \15720 , \15525 , \15719 );
xnor \U$14004 ( \15721 , \15478 , \15499 );
and \U$14005 ( \15722 , \15720 , \15721 );
or \U$14006 ( \15723 , \15500 , \15722 );
xnor \U$14007 ( \15724 , \15453 , \15474 );
and \U$14008 ( \15725 , \15723 , \15724 );
or \U$14009 ( \15726 , \15475 , \15725 );
xnor \U$14010 ( \15727 , \15428 , \15449 );
and \U$14011 ( \15728 , \15726 , \15727 );
or \U$14012 ( \15729 , \15450 , \15728 );
xnor \U$14013 ( \15730 , \15403 , \15424 );
and \U$14014 ( \15731 , \15729 , \15730 );
or \U$14015 ( \15732 , \15425 , \15731 );
xnor \U$14016 ( \15733 , \15344 , \15399 );
and \U$14017 ( \15734 , \15732 , \15733 );
or \U$14018 ( \15735 , \15400 , \15734 );
not \U$14019 ( \15736 , \15735 );
buf \U$14020 ( \15737 , \15736 );
buf \U$14021 ( \15738 , RI9921f28_596);
buf \U$14022 ( \15739 , RI9921fa0_595);
buf \U$14023 ( \15740 , RI9922018_594);
buf \U$14024 ( \15741 , RI9922090_593);
buf \U$14025 ( \15742 , RI9922108_592);
buf \U$14026 ( \15743 , RI9922180_591);
buf \U$14027 ( \15744 , RI99221f8_590);
buf \U$14028 ( \15745 , RI9922270_589);
buf \U$14029 ( \15746 , RI99222e8_588);
buf \U$14030 ( \15747 , RI9921d48_600);
buf \U$14031 ( \15748 , RI9921dc0_599);
buf \U$14032 ( \15749 , RI9921e38_598);
buf \U$14033 ( \15750 , RI9921eb0_597);
and \U$14034 ( \15751 , \15747 , \15748 , \15749 , \15750 );
nor \U$14035 ( \15752 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15751 );
buf \U$14036 ( \15753 , \15752 );
and \U$14037 ( \15754 , \15737 , \15753 );
nor \U$14038 ( \15755 , RI9921d48_600, RI9921dc0_599, RI9921e38_598, RI9921eb0_597, \9716 , RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14039 ( \15756 , RI995e4c8_235, \15755 );
nor \U$14040 ( \15757 , \9719 , \9720 , \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14041 ( \15758 , RI99670f0_222, \15757 );
nor \U$14042 ( \15759 , RI9921d48_600, \9720 , \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14043 ( \15760 , RI890f600_209, \15759 );
nor \U$14044 ( \15761 , \9719 , RI9921dc0_599, \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14045 ( \15762 , RI89185e8_196, \15761 );
nor \U$14046 ( \15763 , RI9921d48_600, RI9921dc0_599, \9721 , \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14047 ( \15764 , RI8924e10_183, \15763 );
nor \U$14048 ( \15765 , \9719 , \9720 , RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14049 ( \15766 , RI8930828_170, \15765 );
nor \U$14050 ( \15767 , RI9921d48_600, \9720 , RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14051 ( \15768 , RI8939810_157, \15767 );
nor \U$14052 ( \15769 , \9719 , RI9921dc0_599, RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14053 ( \15770 , RI8946038_144, \15769 );
nor \U$14054 ( \15771 , RI9921d48_600, RI9921dc0_599, RI9921e38_598, \9722 , RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14055 ( \15772 , RI89ec0a0_131, \15771 );
nor \U$14056 ( \15773 , \9719 , \9720 , \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14057 ( \15774 , RI89ec6b8_118, \15773 );
nor \U$14058 ( \15775 , RI9921d48_600, \9720 , \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14059 ( \15776 , RI9776ff8_105, \15775 );
nor \U$14060 ( \15777 , \9719 , RI9921dc0_599, \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14061 ( \15778 , RI98084f8_92, \15777 );
nor \U$14062 ( \15779 , RI9921d48_600, RI9921dc0_599, \9721 , RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14063 ( \15780 , RI9808b10_79, \15779 );
nor \U$14064 ( \15781 , \9719 , \9720 , RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14065 ( \15782 , RI98197a8_66, \15781 );
nor \U$14066 ( \15783 , RI9921d48_600, \9720 , RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14067 ( \15784 , RI98abcb0_53, \15783 );
nor \U$14068 ( \15785 , \9719 , RI9921dc0_599, RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14069 ( \15786 , RI98bc948_40, \15785 );
nor \U$14070 ( \15787 , RI9921d48_600, RI9921dc0_599, RI9921e38_598, RI9921eb0_597, RI9921f28_596, RI9921fa0_595, RI9922018_594, RI9922090_593, RI9922108_592, RI9922180_591, RI99221f8_590, RI9922270_589, RI99222e8_588);
and \U$14071 ( \15788 , RI994de48_27, \15787 );
or \U$14072 ( \15789 , \15756 , \15758 , \15760 , \15762 , \15764 , \15766 , \15768 , \15770 , \15772 , \15774 , \15776 , \15778 , \15780 , \15782 , \15784 , \15786 , \15788 );
buf \U$14073 ( \15790 , RI9921fa0_595);
buf \U$14074 ( \15791 , RI9922018_594);
buf \U$14075 ( \15792 , RI9922090_593);
buf \U$14076 ( \15793 , RI9922108_592);
buf \U$14077 ( \15794 , RI9922180_591);
buf \U$14078 ( \15795 , RI99221f8_590);
buf \U$14079 ( \15796 , RI9922270_589);
buf \U$14080 ( \15797 , RI99222e8_588);
buf \U$14081 ( \15798 , RI9921f28_596);
buf \U$14082 ( \15799 , RI9921d48_600);
buf \U$14083 ( \15800 , RI9921dc0_599);
buf \U$14084 ( \15801 , RI9921e38_598);
buf \U$14085 ( \15802 , RI9921eb0_597);
or \U$14086 ( \15803 , \15799 , \15800 , \15801 , \15802 );
and \U$14087 ( \15804 , \15798 , \15803 );
or \U$14088 ( \15805 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15804 );
buf \U$14089 ( \15806 , \15805 );
_DC g16b2 ( \15807_nG16b2 , \15789 , \15806 );
buf \U$14090 ( \15808 , \15807_nG16b2 );
not \U$14091 ( \15809 , \15808 );
nor \U$14092 ( \15810 , \12513 , \12517 , \12521 , \12525 , \12530 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14093 ( \15811 , RI995e4c8_235, \15810 );
nor \U$14094 ( \15812 , \12565 , \12566 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14095 ( \15813 , RI99670f0_222, \15812 );
nor \U$14096 ( \15814 , \12513 , \12566 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14097 ( \15815 , RI890f600_209, \15814 );
nor \U$14098 ( \15816 , \12565 , \12517 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14099 ( \15817 , RI89185e8_196, \15816 );
nor \U$14100 ( \15818 , \12513 , \12517 , \12567 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14101 ( \15819 , RI8924e10_183, \15818 );
nor \U$14102 ( \15820 , \12565 , \12566 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14103 ( \15821 , RI8930828_170, \15820 );
nor \U$14104 ( \15822 , \12513 , \12566 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14105 ( \15823 , RI8939810_157, \15822 );
nor \U$14106 ( \15824 , \12565 , \12517 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14107 ( \15825 , RI8946038_144, \15824 );
nor \U$14108 ( \15826 , \12513 , \12517 , \12521 , \12568 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14109 ( \15827 , RI89ec0a0_131, \15826 );
nor \U$14110 ( \15828 , \12565 , \12566 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14111 ( \15829 , RI89ec6b8_118, \15828 );
nor \U$14112 ( \15830 , \12513 , \12566 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14113 ( \15831 , RI9776ff8_105, \15830 );
nor \U$14114 ( \15832 , \12565 , \12517 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14115 ( \15833 , RI98084f8_92, \15832 );
nor \U$14116 ( \15834 , \12513 , \12517 , \12567 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14117 ( \15835 , RI9808b10_79, \15834 );
nor \U$14118 ( \15836 , \12565 , \12566 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14119 ( \15837 , RI98197a8_66, \15836 );
nor \U$14120 ( \15838 , \12513 , \12566 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14121 ( \15839 , RI98abcb0_53, \15838 );
nor \U$14122 ( \15840 , \12565 , \12517 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14123 ( \15841 , RI98bc948_40, \15840 );
nor \U$14124 ( \15842 , \12513 , \12517 , \12521 , \12525 , \12529 , \12534 , \12538 , \12542 , \12546 , \12550 , \12554 , \12558 , \12562 );
and \U$14125 ( \15843 , RI994de48_27, \15842 );
or \U$14126 ( \15844 , \15811 , \15813 , \15815 , \15817 , \15819 , \15821 , \15823 , \15825 , \15827 , \15829 , \15831 , \15833 , \15835 , \15837 , \15839 , \15841 , \15843 );
buf \U$14127 ( \15845 , \12534 );
buf \U$14128 ( \15846 , \12538 );
buf \U$14129 ( \15847 , \12542 );
buf \U$14130 ( \15848 , \12546 );
buf \U$14131 ( \15849 , \12550 );
buf \U$14132 ( \15850 , \12554 );
buf \U$14133 ( \15851 , \12558 );
buf \U$14134 ( \15852 , \12562 );
buf \U$14135 ( \15853 , \12529 );
buf \U$14136 ( \15854 , \12513 );
buf \U$14137 ( \15855 , \12517 );
buf \U$14138 ( \15856 , \12521 );
buf \U$14139 ( \15857 , \12525 );
or \U$14140 ( \15858 , \15854 , \15855 , \15856 , \15857 );
and \U$14141 ( \15859 , \15853 , \15858 );
or \U$14142 ( \15860 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15859 );
buf \U$14143 ( \15861 , \15860 );
_DC g16e9 ( \15862_nG16e9 , \15844 , \15861 );
buf \U$14144 ( \15863 , \15862_nG16e9 );
and \U$14145 ( \15864 , \15809 , \15863 );
and \U$14146 ( \15865 , RI995e450_236, \15755 );
and \U$14147 ( \15866 , RI9967078_223, \15757 );
and \U$14148 ( \15867 , RI9967690_210, \15759 );
and \U$14149 ( \15868 , RI890fba0_197, \15761 );
and \U$14150 ( \15869 , RI8918b88_184, \15763 );
and \U$14151 ( \15870 , RI89253b0_171, \15765 );
and \U$14152 ( \15871 , RI8930dc8_158, \15767 );
and \U$14153 ( \15872 , RI8939db0_145, \15769 );
and \U$14154 ( \15873 , RI89465d8_132, \15771 );
and \U$14155 ( \15874 , RI89ec640_119, \15773 );
and \U$14156 ( \15875 , RI9776f80_106, \15775 );
and \U$14157 ( \15876 , RI9808480_93, \15777 );
and \U$14158 ( \15877 , RI9808a98_80, \15779 );
and \U$14159 ( \15878 , RI9819730_67, \15781 );
and \U$14160 ( \15879 , RI98abc38_54, \15783 );
and \U$14161 ( \15880 , RI98bc8d0_41, \15785 );
and \U$14162 ( \15881 , RI994ddd0_28, \15787 );
or \U$14163 ( \15882 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 );
_DC g16fe ( \15883_nG16fe , \15882 , \15806 );
buf \U$14164 ( \15884 , \15883_nG16fe );
not \U$14165 ( \15885 , \15884 );
and \U$14166 ( \15886 , RI995e450_236, \15810 );
and \U$14167 ( \15887 , RI9967078_223, \15812 );
and \U$14168 ( \15888 , RI9967690_210, \15814 );
and \U$14169 ( \15889 , RI890fba0_197, \15816 );
and \U$14170 ( \15890 , RI8918b88_184, \15818 );
and \U$14171 ( \15891 , RI89253b0_171, \15820 );
and \U$14172 ( \15892 , RI8930dc8_158, \15822 );
and \U$14173 ( \15893 , RI8939db0_145, \15824 );
and \U$14174 ( \15894 , RI89465d8_132, \15826 );
and \U$14175 ( \15895 , RI89ec640_119, \15828 );
and \U$14176 ( \15896 , RI9776f80_106, \15830 );
and \U$14177 ( \15897 , RI9808480_93, \15832 );
and \U$14178 ( \15898 , RI9808a98_80, \15834 );
and \U$14179 ( \15899 , RI9819730_67, \15836 );
and \U$14180 ( \15900 , RI98abc38_54, \15838 );
and \U$14181 ( \15901 , RI98bc8d0_41, \15840 );
and \U$14182 ( \15902 , RI994ddd0_28, \15842 );
or \U$14183 ( \15903 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 );
_DC g1713 ( \15904_nG1713 , \15903 , \15861 );
buf \U$14184 ( \15905 , \15904_nG1713 );
and \U$14185 ( \15906 , \15885 , \15905 );
and \U$14186 ( \15907 , RI995e3d8_237, \15755 );
and \U$14187 ( \15908 , RI99669e8_224, \15757 );
and \U$14188 ( \15909 , RI9967618_211, \15759 );
and \U$14189 ( \15910 , RI890fb28_198, \15761 );
and \U$14190 ( \15911 , RI8918b10_185, \15763 );
and \U$14191 ( \15912 , RI8925338_172, \15765 );
and \U$14192 ( \15913 , RI8930d50_159, \15767 );
and \U$14193 ( \15914 , RI8939d38_146, \15769 );
and \U$14194 ( \15915 , RI8946560_133, \15771 );
and \U$14195 ( \15916 , RI89ec5c8_120, \15773 );
and \U$14196 ( \15917 , RI9776f08_107, \15775 );
and \U$14197 ( \15918 , RI9808408_94, \15777 );
and \U$14198 ( \15919 , RI9808a20_81, \15779 );
and \U$14199 ( \15920 , RI98196b8_68, \15781 );
and \U$14200 ( \15921 , RI98abbc0_55, \15783 );
and \U$14201 ( \15922 , RI98bc858_42, \15785 );
and \U$14202 ( \15923 , RI994dd58_29, \15787 );
or \U$14203 ( \15924 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 );
_DC g1728 ( \15925_nG1728 , \15924 , \15806 );
buf \U$14204 ( \15926 , \15925_nG1728 );
not \U$14205 ( \15927 , \15926 );
and \U$14206 ( \15928 , RI995e3d8_237, \15810 );
and \U$14207 ( \15929 , RI99669e8_224, \15812 );
and \U$14208 ( \15930 , RI9967618_211, \15814 );
and \U$14209 ( \15931 , RI890fb28_198, \15816 );
and \U$14210 ( \15932 , RI8918b10_185, \15818 );
and \U$14211 ( \15933 , RI8925338_172, \15820 );
and \U$14212 ( \15934 , RI8930d50_159, \15822 );
and \U$14213 ( \15935 , RI8939d38_146, \15824 );
and \U$14214 ( \15936 , RI8946560_133, \15826 );
and \U$14215 ( \15937 , RI89ec5c8_120, \15828 );
and \U$14216 ( \15938 , RI9776f08_107, \15830 );
and \U$14217 ( \15939 , RI9808408_94, \15832 );
and \U$14218 ( \15940 , RI9808a20_81, \15834 );
and \U$14219 ( \15941 , RI98196b8_68, \15836 );
and \U$14220 ( \15942 , RI98abbc0_55, \15838 );
and \U$14221 ( \15943 , RI98bc858_42, \15840 );
and \U$14222 ( \15944 , RI994dd58_29, \15842 );
or \U$14223 ( \15945 , \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 );
_DC g173d ( \15946_nG173d , \15945 , \15861 );
buf \U$14224 ( \15947 , \15946_nG173d );
and \U$14225 ( \15948 , \15927 , \15947 );
and \U$14226 ( \15949 , RI9959fe0_238, \15755 );
and \U$14227 ( \15950 , RI995e978_225, \15757 );
and \U$14228 ( \15951 , RI99675a0_212, \15759 );
and \U$14229 ( \15952 , RI890fab0_199, \15761 );
and \U$14230 ( \15953 , RI8918a98_186, \15763 );
and \U$14231 ( \15954 , RI89252c0_173, \15765 );
and \U$14232 ( \15955 , RI8930cd8_160, \15767 );
and \U$14233 ( \15956 , RI8939cc0_147, \15769 );
and \U$14234 ( \15957 , RI89464e8_134, \15771 );
and \U$14235 ( \15958 , RI89ec550_121, \15773 );
and \U$14236 ( \15959 , RI9776e90_108, \15775 );
and \U$14237 ( \15960 , RI9808390_95, \15777 );
and \U$14238 ( \15961 , RI98089a8_82, \15779 );
and \U$14239 ( \15962 , RI9819640_69, \15781 );
and \U$14240 ( \15963 , RI98abb48_56, \15783 );
and \U$14241 ( \15964 , RI98bc7e0_43, \15785 );
and \U$14242 ( \15965 , RI994dce0_30, \15787 );
or \U$14243 ( \15966 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 );
_DC g1752 ( \15967_nG1752 , \15966 , \15806 );
buf \U$14244 ( \15968 , \15967_nG1752 );
not \U$14245 ( \15969 , \15968 );
and \U$14246 ( \15970 , RI9959fe0_238, \15810 );
and \U$14247 ( \15971 , RI995e978_225, \15812 );
and \U$14248 ( \15972 , RI99675a0_212, \15814 );
and \U$14249 ( \15973 , RI890fab0_199, \15816 );
and \U$14250 ( \15974 , RI8918a98_186, \15818 );
and \U$14251 ( \15975 , RI89252c0_173, \15820 );
and \U$14252 ( \15976 , RI8930cd8_160, \15822 );
and \U$14253 ( \15977 , RI8939cc0_147, \15824 );
and \U$14254 ( \15978 , RI89464e8_134, \15826 );
and \U$14255 ( \15979 , RI89ec550_121, \15828 );
and \U$14256 ( \15980 , RI9776e90_108, \15830 );
and \U$14257 ( \15981 , RI9808390_95, \15832 );
and \U$14258 ( \15982 , RI98089a8_82, \15834 );
and \U$14259 ( \15983 , RI9819640_69, \15836 );
and \U$14260 ( \15984 , RI98abb48_56, \15838 );
and \U$14261 ( \15985 , RI98bc7e0_43, \15840 );
and \U$14262 ( \15986 , RI994dce0_30, \15842 );
or \U$14263 ( \15987 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 );
_DC g1767 ( \15988_nG1767 , \15987 , \15861 );
buf \U$14264 ( \15989 , \15988_nG1767 );
and \U$14265 ( \15990 , \15969 , \15989 );
and \U$14266 ( \15991 , RI9959f68_239, \15755 );
and \U$14267 ( \15992 , RI995e900_226, \15757 );
and \U$14268 ( \15993 , RI9967528_213, \15759 );
and \U$14269 ( \15994 , RI890fa38_200, \15761 );
and \U$14270 ( \15995 , RI8918a20_187, \15763 );
and \U$14271 ( \15996 , RI8925248_174, \15765 );
and \U$14272 ( \15997 , RI8930c60_161, \15767 );
and \U$14273 ( \15998 , RI8939c48_148, \15769 );
and \U$14274 ( \15999 , RI8946470_135, \15771 );
and \U$14275 ( \16000 , RI89ec4d8_122, \15773 );
and \U$14276 ( \16001 , RI9776e18_109, \15775 );
and \U$14277 ( \16002 , RI9808318_96, \15777 );
and \U$14278 ( \16003 , RI9808930_83, \15779 );
and \U$14279 ( \16004 , RI98195c8_70, \15781 );
and \U$14280 ( \16005 , RI98abad0_57, \15783 );
and \U$14281 ( \16006 , RI98bc768_44, \15785 );
and \U$14282 ( \16007 , RI994dc68_31, \15787 );
or \U$14283 ( \16008 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 );
_DC g177c ( \16009_nG177c , \16008 , \15806 );
buf \U$14284 ( \16010 , \16009_nG177c );
not \U$14285 ( \16011 , \16010 );
and \U$14286 ( \16012 , RI9959f68_239, \15810 );
and \U$14287 ( \16013 , RI995e900_226, \15812 );
and \U$14288 ( \16014 , RI9967528_213, \15814 );
and \U$14289 ( \16015 , RI890fa38_200, \15816 );
and \U$14290 ( \16016 , RI8918a20_187, \15818 );
and \U$14291 ( \16017 , RI8925248_174, \15820 );
and \U$14292 ( \16018 , RI8930c60_161, \15822 );
and \U$14293 ( \16019 , RI8939c48_148, \15824 );
and \U$14294 ( \16020 , RI8946470_135, \15826 );
and \U$14295 ( \16021 , RI89ec4d8_122, \15828 );
and \U$14296 ( \16022 , RI9776e18_109, \15830 );
and \U$14297 ( \16023 , RI9808318_96, \15832 );
and \U$14298 ( \16024 , RI9808930_83, \15834 );
and \U$14299 ( \16025 , RI98195c8_70, \15836 );
and \U$14300 ( \16026 , RI98abad0_57, \15838 );
and \U$14301 ( \16027 , RI98bc768_44, \15840 );
and \U$14302 ( \16028 , RI994dc68_31, \15842 );
or \U$14303 ( \16029 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 );
_DC g1791 ( \16030_nG1791 , \16029 , \15861 );
buf \U$14304 ( \16031 , \16030_nG1791 );
and \U$14305 ( \16032 , \16011 , \16031 );
and \U$14306 ( \16033 , RI9959860_240, \15755 );
and \U$14307 ( \16034 , RI995e888_227, \15757 );
and \U$14308 ( \16035 , RI99674b0_214, \15759 );
and \U$14309 ( \16036 , RI890f9c0_201, \15761 );
and \U$14310 ( \16037 , RI89189a8_188, \15763 );
and \U$14311 ( \16038 , RI89251d0_175, \15765 );
and \U$14312 ( \16039 , RI8930be8_162, \15767 );
and \U$14313 ( \16040 , RI8939bd0_149, \15769 );
and \U$14314 ( \16041 , RI89463f8_136, \15771 );
and \U$14315 ( \16042 , RI89ec460_123, \15773 );
and \U$14316 ( \16043 , RI9776da0_110, \15775 );
and \U$14317 ( \16044 , RI98082a0_97, \15777 );
and \U$14318 ( \16045 , RI98088b8_84, \15779 );
and \U$14319 ( \16046 , RI9819550_71, \15781 );
and \U$14320 ( \16047 , RI98aba58_58, \15783 );
and \U$14321 ( \16048 , RI98bc6f0_45, \15785 );
and \U$14322 ( \16049 , RI994dbf0_32, \15787 );
or \U$14323 ( \16050 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 );
_DC g17a6 ( \16051_nG17a6 , \16050 , \15806 );
buf \U$14324 ( \16052 , \16051_nG17a6 );
not \U$14325 ( \16053 , \16052 );
and \U$14326 ( \16054 , RI9959860_240, \15810 );
and \U$14327 ( \16055 , RI995e888_227, \15812 );
and \U$14328 ( \16056 , RI99674b0_214, \15814 );
and \U$14329 ( \16057 , RI890f9c0_201, \15816 );
and \U$14330 ( \16058 , RI89189a8_188, \15818 );
and \U$14331 ( \16059 , RI89251d0_175, \15820 );
and \U$14332 ( \16060 , RI8930be8_162, \15822 );
and \U$14333 ( \16061 , RI8939bd0_149, \15824 );
and \U$14334 ( \16062 , RI89463f8_136, \15826 );
and \U$14335 ( \16063 , RI89ec460_123, \15828 );
and \U$14336 ( \16064 , RI9776da0_110, \15830 );
and \U$14337 ( \16065 , RI98082a0_97, \15832 );
and \U$14338 ( \16066 , RI98088b8_84, \15834 );
and \U$14339 ( \16067 , RI9819550_71, \15836 );
and \U$14340 ( \16068 , RI98aba58_58, \15838 );
and \U$14341 ( \16069 , RI98bc6f0_45, \15840 );
and \U$14342 ( \16070 , RI994dbf0_32, \15842 );
or \U$14343 ( \16071 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 );
_DC g17bb ( \16072_nG17bb , \16071 , \15861 );
buf \U$14344 ( \16073 , \16072_nG17bb );
and \U$14345 ( \16074 , \16053 , \16073 );
and \U$14346 ( \16075 , RI994d998_241, \15755 );
and \U$14347 ( \16076 , RI995e810_228, \15757 );
and \U$14348 ( \16077 , RI9967438_215, \15759 );
and \U$14349 ( \16078 , RI890f948_202, \15761 );
and \U$14350 ( \16079 , RI8918930_189, \15763 );
and \U$14351 ( \16080 , RI8925158_176, \15765 );
and \U$14352 ( \16081 , RI8930b70_163, \15767 );
and \U$14353 ( \16082 , RI8939b58_150, \15769 );
and \U$14354 ( \16083 , RI8946380_137, \15771 );
and \U$14355 ( \16084 , RI89ec3e8_124, \15773 );
and \U$14356 ( \16085 , RI9776d28_111, \15775 );
and \U$14357 ( \16086 , RI9808228_98, \15777 );
and \U$14358 ( \16087 , RI9808840_85, \15779 );
and \U$14359 ( \16088 , RI98194d8_72, \15781 );
and \U$14360 ( \16089 , RI98ab9e0_59, \15783 );
and \U$14361 ( \16090 , RI98abff8_46, \15785 );
and \U$14362 ( \16091 , RI98bcc90_33, \15787 );
or \U$14363 ( \16092 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 );
_DC g17d0 ( \16093_nG17d0 , \16092 , \15806 );
buf \U$14364 ( \16094 , \16093_nG17d0 );
not \U$14365 ( \16095 , \16094 );
and \U$14366 ( \16096 , RI994d998_241, \15810 );
and \U$14367 ( \16097 , RI995e810_228, \15812 );
and \U$14368 ( \16098 , RI9967438_215, \15814 );
and \U$14369 ( \16099 , RI890f948_202, \15816 );
and \U$14370 ( \16100 , RI8918930_189, \15818 );
and \U$14371 ( \16101 , RI8925158_176, \15820 );
and \U$14372 ( \16102 , RI8930b70_163, \15822 );
and \U$14373 ( \16103 , RI8939b58_150, \15824 );
and \U$14374 ( \16104 , RI8946380_137, \15826 );
and \U$14375 ( \16105 , RI89ec3e8_124, \15828 );
and \U$14376 ( \16106 , RI9776d28_111, \15830 );
and \U$14377 ( \16107 , RI9808228_98, \15832 );
and \U$14378 ( \16108 , RI9808840_85, \15834 );
and \U$14379 ( \16109 , RI98194d8_72, \15836 );
and \U$14380 ( \16110 , RI98ab9e0_59, \15838 );
and \U$14381 ( \16111 , RI98abff8_46, \15840 );
and \U$14382 ( \16112 , RI98bcc90_33, \15842 );
or \U$14383 ( \16113 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 );
_DC g17e5 ( \16114_nG17e5 , \16113 , \15861 );
buf \U$14384 ( \16115 , \16114_nG17e5 );
and \U$14385 ( \16116 , \16095 , \16115 );
and \U$14386 ( \16117 , RI994d920_242, \15755 );
and \U$14387 ( \16118 , RI995e798_229, \15757 );
and \U$14388 ( \16119 , RI99673c0_216, \15759 );
and \U$14389 ( \16120 , RI890f8d0_203, \15761 );
and \U$14390 ( \16121 , RI89188b8_190, \15763 );
and \U$14391 ( \16122 , RI89250e0_177, \15765 );
and \U$14392 ( \16123 , RI8930af8_164, \15767 );
and \U$14393 ( \16124 , RI8939ae0_151, \15769 );
and \U$14394 ( \16125 , RI8946308_138, \15771 );
and \U$14395 ( \16126 , RI89ec370_125, \15773 );
and \U$14396 ( \16127 , RI89ec988_112, \15775 );
and \U$14397 ( \16128 , RI97772c8_99, \15777 );
and \U$14398 ( \16129 , RI98087c8_86, \15779 );
and \U$14399 ( \16130 , RI9819460_73, \15781 );
and \U$14400 ( \16131 , RI98ab968_60, \15783 );
and \U$14401 ( \16132 , RI98abf80_47, \15785 );
and \U$14402 ( \16133 , RI98bcc18_34, \15787 );
or \U$14403 ( \16134 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 );
_DC g17fa ( \16135_nG17fa , \16134 , \15806 );
buf \U$14404 ( \16136 , \16135_nG17fa );
not \U$14405 ( \16137 , \16136 );
and \U$14406 ( \16138 , RI994d920_242, \15810 );
and \U$14407 ( \16139 , RI995e798_229, \15812 );
and \U$14408 ( \16140 , RI99673c0_216, \15814 );
and \U$14409 ( \16141 , RI890f8d0_203, \15816 );
and \U$14410 ( \16142 , RI89188b8_190, \15818 );
and \U$14411 ( \16143 , RI89250e0_177, \15820 );
and \U$14412 ( \16144 , RI8930af8_164, \15822 );
and \U$14413 ( \16145 , RI8939ae0_151, \15824 );
and \U$14414 ( \16146 , RI8946308_138, \15826 );
and \U$14415 ( \16147 , RI89ec370_125, \15828 );
and \U$14416 ( \16148 , RI89ec988_112, \15830 );
and \U$14417 ( \16149 , RI97772c8_99, \15832 );
and \U$14418 ( \16150 , RI98087c8_86, \15834 );
and \U$14419 ( \16151 , RI9819460_73, \15836 );
and \U$14420 ( \16152 , RI98ab968_60, \15838 );
and \U$14421 ( \16153 , RI98abf80_47, \15840 );
and \U$14422 ( \16154 , RI98bcc18_34, \15842 );
or \U$14423 ( \16155 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 );
_DC g180f ( \16156_nG180f , \16155 , \15861 );
buf \U$14424 ( \16157 , \16156_nG180f );
and \U$14425 ( \16158 , \16137 , \16157 );
and \U$14426 ( \16159 , RI994d8a8_243, \15755 );
and \U$14427 ( \16160 , RI995e720_230, \15757 );
and \U$14428 ( \16161 , RI9967348_217, \15759 );
and \U$14429 ( \16162 , RI890f858_204, \15761 );
and \U$14430 ( \16163 , RI8918840_191, \15763 );
and \U$14431 ( \16164 , RI8925068_178, \15765 );
and \U$14432 ( \16165 , RI8930a80_165, \15767 );
and \U$14433 ( \16166 , RI8939a68_152, \15769 );
and \U$14434 ( \16167 , RI8946290_139, \15771 );
and \U$14435 ( \16168 , RI89ec2f8_126, \15773 );
and \U$14436 ( \16169 , RI89ec910_113, \15775 );
and \U$14437 ( \16170 , RI9777250_100, \15777 );
and \U$14438 ( \16171 , RI9808750_87, \15779 );
and \U$14439 ( \16172 , RI98193e8_74, \15781 );
and \U$14440 ( \16173 , RI98ab8f0_61, \15783 );
and \U$14441 ( \16174 , RI98abf08_48, \15785 );
and \U$14442 ( \16175 , RI98bcba0_35, \15787 );
or \U$14443 ( \16176 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 );
_DC g1824 ( \16177_nG1824 , \16176 , \15806 );
buf \U$14444 ( \16178 , \16177_nG1824 );
not \U$14445 ( \16179 , \16178 );
and \U$14446 ( \16180 , RI994d8a8_243, \15810 );
and \U$14447 ( \16181 , RI995e720_230, \15812 );
and \U$14448 ( \16182 , RI9967348_217, \15814 );
and \U$14449 ( \16183 , RI890f858_204, \15816 );
and \U$14450 ( \16184 , RI8918840_191, \15818 );
and \U$14451 ( \16185 , RI8925068_178, \15820 );
and \U$14452 ( \16186 , RI8930a80_165, \15822 );
and \U$14453 ( \16187 , RI8939a68_152, \15824 );
and \U$14454 ( \16188 , RI8946290_139, \15826 );
and \U$14455 ( \16189 , RI89ec2f8_126, \15828 );
and \U$14456 ( \16190 , RI89ec910_113, \15830 );
and \U$14457 ( \16191 , RI9777250_100, \15832 );
and \U$14458 ( \16192 , RI9808750_87, \15834 );
and \U$14459 ( \16193 , RI98193e8_74, \15836 );
and \U$14460 ( \16194 , RI98ab8f0_61, \15838 );
and \U$14461 ( \16195 , RI98abf08_48, \15840 );
and \U$14462 ( \16196 , RI98bcba0_35, \15842 );
or \U$14463 ( \16197 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 );
_DC g1839 ( \16198_nG1839 , \16197 , \15861 );
buf \U$14464 ( \16199 , \16198_nG1839 );
and \U$14465 ( \16200 , \16179 , \16199 );
and \U$14466 ( \16201 , RI994d830_244, \15755 );
and \U$14467 ( \16202 , RI995e6a8_231, \15757 );
and \U$14468 ( \16203 , RI99672d0_218, \15759 );
and \U$14469 ( \16204 , RI890f7e0_205, \15761 );
and \U$14470 ( \16205 , RI89187c8_192, \15763 );
and \U$14471 ( \16206 , RI8924ff0_179, \15765 );
and \U$14472 ( \16207 , RI8930a08_166, \15767 );
and \U$14473 ( \16208 , RI89399f0_153, \15769 );
and \U$14474 ( \16209 , RI8946218_140, \15771 );
and \U$14475 ( \16210 , RI89ec280_127, \15773 );
and \U$14476 ( \16211 , RI89ec898_114, \15775 );
and \U$14477 ( \16212 , RI97771d8_101, \15777 );
and \U$14478 ( \16213 , RI98086d8_88, \15779 );
and \U$14479 ( \16214 , RI9819370_75, \15781 );
and \U$14480 ( \16215 , RI98ab878_62, \15783 );
and \U$14481 ( \16216 , RI98abe90_49, \15785 );
and \U$14482 ( \16217 , RI98bcb28_36, \15787 );
or \U$14483 ( \16218 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 );
_DC g184e ( \16219_nG184e , \16218 , \15806 );
buf \U$14484 ( \16220 , \16219_nG184e );
not \U$14485 ( \16221 , \16220 );
and \U$14486 ( \16222 , RI994d830_244, \15810 );
and \U$14487 ( \16223 , RI995e6a8_231, \15812 );
and \U$14488 ( \16224 , RI99672d0_218, \15814 );
and \U$14489 ( \16225 , RI890f7e0_205, \15816 );
and \U$14490 ( \16226 , RI89187c8_192, \15818 );
and \U$14491 ( \16227 , RI8924ff0_179, \15820 );
and \U$14492 ( \16228 , RI8930a08_166, \15822 );
and \U$14493 ( \16229 , RI89399f0_153, \15824 );
and \U$14494 ( \16230 , RI8946218_140, \15826 );
and \U$14495 ( \16231 , RI89ec280_127, \15828 );
and \U$14496 ( \16232 , RI89ec898_114, \15830 );
and \U$14497 ( \16233 , RI97771d8_101, \15832 );
and \U$14498 ( \16234 , RI98086d8_88, \15834 );
and \U$14499 ( \16235 , RI9819370_75, \15836 );
and \U$14500 ( \16236 , RI98ab878_62, \15838 );
and \U$14501 ( \16237 , RI98abe90_49, \15840 );
and \U$14502 ( \16238 , RI98bcb28_36, \15842 );
or \U$14503 ( \16239 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 );
_DC g1863 ( \16240_nG1863 , \16239 , \15861 );
buf \U$14504 ( \16241 , \16240_nG1863 );
and \U$14505 ( \16242 , \16221 , \16241 );
and \U$14506 ( \16243 , RI994d7b8_245, \15755 );
and \U$14507 ( \16244 , RI995e630_232, \15757 );
and \U$14508 ( \16245 , RI9967258_219, \15759 );
and \U$14509 ( \16246 , RI890f768_206, \15761 );
and \U$14510 ( \16247 , RI8918750_193, \15763 );
and \U$14511 ( \16248 , RI8924f78_180, \15765 );
and \U$14512 ( \16249 , RI8930990_167, \15767 );
and \U$14513 ( \16250 , RI8939978_154, \15769 );
and \U$14514 ( \16251 , RI89461a0_141, \15771 );
and \U$14515 ( \16252 , RI89ec208_128, \15773 );
and \U$14516 ( \16253 , RI89ec820_115, \15775 );
and \U$14517 ( \16254 , RI9777160_102, \15777 );
and \U$14518 ( \16255 , RI9808660_89, \15779 );
and \U$14519 ( \16256 , RI98192f8_76, \15781 );
and \U$14520 ( \16257 , RI98ab800_63, \15783 );
and \U$14521 ( \16258 , RI98abe18_50, \15785 );
and \U$14522 ( \16259 , RI98bcab0_37, \15787 );
or \U$14523 ( \16260 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 );
_DC g1878 ( \16261_nG1878 , \16260 , \15806 );
buf \U$14524 ( \16262 , \16261_nG1878 );
not \U$14525 ( \16263 , \16262 );
and \U$14526 ( \16264 , RI994d7b8_245, \15810 );
and \U$14527 ( \16265 , RI995e630_232, \15812 );
and \U$14528 ( \16266 , RI9967258_219, \15814 );
and \U$14529 ( \16267 , RI890f768_206, \15816 );
and \U$14530 ( \16268 , RI8918750_193, \15818 );
and \U$14531 ( \16269 , RI8924f78_180, \15820 );
and \U$14532 ( \16270 , RI8930990_167, \15822 );
and \U$14533 ( \16271 , RI8939978_154, \15824 );
and \U$14534 ( \16272 , RI89461a0_141, \15826 );
and \U$14535 ( \16273 , RI89ec208_128, \15828 );
and \U$14536 ( \16274 , RI89ec820_115, \15830 );
and \U$14537 ( \16275 , RI9777160_102, \15832 );
and \U$14538 ( \16276 , RI9808660_89, \15834 );
and \U$14539 ( \16277 , RI98192f8_76, \15836 );
and \U$14540 ( \16278 , RI98ab800_63, \15838 );
and \U$14541 ( \16279 , RI98abe18_50, \15840 );
and \U$14542 ( \16280 , RI98bcab0_37, \15842 );
or \U$14543 ( \16281 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 );
_DC g188d ( \16282_nG188d , \16281 , \15861 );
buf \U$14544 ( \16283 , \16282_nG188d );
and \U$14545 ( \16284 , \16263 , \16283 );
and \U$14546 ( \16285 , RI994d740_246, \15755 );
and \U$14547 ( \16286 , RI995e5b8_233, \15757 );
and \U$14548 ( \16287 , RI99671e0_220, \15759 );
and \U$14549 ( \16288 , RI890f6f0_207, \15761 );
and \U$14550 ( \16289 , RI89186d8_194, \15763 );
and \U$14551 ( \16290 , RI8924f00_181, \15765 );
and \U$14552 ( \16291 , RI8930918_168, \15767 );
and \U$14553 ( \16292 , RI8939900_155, \15769 );
and \U$14554 ( \16293 , RI8946128_142, \15771 );
and \U$14555 ( \16294 , RI89ec190_129, \15773 );
and \U$14556 ( \16295 , RI89ec7a8_116, \15775 );
and \U$14557 ( \16296 , RI97770e8_103, \15777 );
and \U$14558 ( \16297 , RI98085e8_90, \15779 );
and \U$14559 ( \16298 , RI9819280_77, \15781 );
and \U$14560 ( \16299 , RI98ab788_64, \15783 );
and \U$14561 ( \16300 , RI98abda0_51, \15785 );
and \U$14562 ( \16301 , RI98bca38_38, \15787 );
or \U$14563 ( \16302 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 );
_DC g18a2 ( \16303_nG18a2 , \16302 , \15806 );
buf \U$14564 ( \16304 , \16303_nG18a2 );
not \U$14565 ( \16305 , \16304 );
and \U$14566 ( \16306 , RI994d740_246, \15810 );
and \U$14567 ( \16307 , RI995e5b8_233, \15812 );
and \U$14568 ( \16308 , RI99671e0_220, \15814 );
and \U$14569 ( \16309 , RI890f6f0_207, \15816 );
and \U$14570 ( \16310 , RI89186d8_194, \15818 );
and \U$14571 ( \16311 , RI8924f00_181, \15820 );
and \U$14572 ( \16312 , RI8930918_168, \15822 );
and \U$14573 ( \16313 , RI8939900_155, \15824 );
and \U$14574 ( \16314 , RI8946128_142, \15826 );
and \U$14575 ( \16315 , RI89ec190_129, \15828 );
and \U$14576 ( \16316 , RI89ec7a8_116, \15830 );
and \U$14577 ( \16317 , RI97770e8_103, \15832 );
and \U$14578 ( \16318 , RI98085e8_90, \15834 );
and \U$14579 ( \16319 , RI9819280_77, \15836 );
and \U$14580 ( \16320 , RI98ab788_64, \15838 );
and \U$14581 ( \16321 , RI98abda0_51, \15840 );
and \U$14582 ( \16322 , RI98bca38_38, \15842 );
or \U$14583 ( \16323 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 );
_DC g18b7 ( \16324_nG18b7 , \16323 , \15861 );
buf \U$14584 ( \16325 , \16324_nG18b7 );
and \U$14585 ( \16326 , \16305 , \16325 );
and \U$14586 ( \16327 , RI994d6c8_247, \15755 );
and \U$14587 ( \16328 , RI995e540_234, \15757 );
and \U$14588 ( \16329 , RI9967168_221, \15759 );
and \U$14589 ( \16330 , RI890f678_208, \15761 );
and \U$14590 ( \16331 , RI8918660_195, \15763 );
and \U$14591 ( \16332 , RI8924e88_182, \15765 );
and \U$14592 ( \16333 , RI89308a0_169, \15767 );
and \U$14593 ( \16334 , RI8939888_156, \15769 );
and \U$14594 ( \16335 , RI89460b0_143, \15771 );
and \U$14595 ( \16336 , RI89ec118_130, \15773 );
and \U$14596 ( \16337 , RI89ec730_117, \15775 );
and \U$14597 ( \16338 , RI9777070_104, \15777 );
and \U$14598 ( \16339 , RI9808570_91, \15779 );
and \U$14599 ( \16340 , RI9819208_78, \15781 );
and \U$14600 ( \16341 , RI98ab710_65, \15783 );
and \U$14601 ( \16342 , RI98abd28_52, \15785 );
and \U$14602 ( \16343 , RI98bc9c0_39, \15787 );
or \U$14603 ( \16344 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 );
_DC g18cc ( \16345_nG18cc , \16344 , \15806 );
buf \U$14604 ( \16346 , \16345_nG18cc );
not \U$14605 ( \16347 , \16346 );
and \U$14606 ( \16348 , RI994d6c8_247, \15810 );
and \U$14607 ( \16349 , RI995e540_234, \15812 );
and \U$14608 ( \16350 , RI9967168_221, \15814 );
and \U$14609 ( \16351 , RI890f678_208, \15816 );
and \U$14610 ( \16352 , RI8918660_195, \15818 );
and \U$14611 ( \16353 , RI8924e88_182, \15820 );
and \U$14612 ( \16354 , RI89308a0_169, \15822 );
and \U$14613 ( \16355 , RI8939888_156, \15824 );
and \U$14614 ( \16356 , RI89460b0_143, \15826 );
and \U$14615 ( \16357 , RI89ec118_130, \15828 );
and \U$14616 ( \16358 , RI89ec730_117, \15830 );
and \U$14617 ( \16359 , RI9777070_104, \15832 );
and \U$14618 ( \16360 , RI9808570_91, \15834 );
and \U$14619 ( \16361 , RI9819208_78, \15836 );
and \U$14620 ( \16362 , RI98ab710_65, \15838 );
and \U$14621 ( \16363 , RI98abd28_52, \15840 );
and \U$14622 ( \16364 , RI98bc9c0_39, \15842 );
or \U$14623 ( \16365 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 );
_DC g18e1 ( \16366_nG18e1 , \16365 , \15861 );
buf \U$14624 ( \16367 , \16366_nG18e1 );
and \U$14625 ( \16368 , \16347 , \16367 );
xnor \U$14626 ( \16369 , \16325 , \16304 );
and \U$14627 ( \16370 , \16368 , \16369 );
or \U$14628 ( \16371 , \16326 , \16370 );
xnor \U$14629 ( \16372 , \16283 , \16262 );
and \U$14630 ( \16373 , \16371 , \16372 );
or \U$14631 ( \16374 , \16284 , \16373 );
xnor \U$14632 ( \16375 , \16241 , \16220 );
and \U$14633 ( \16376 , \16374 , \16375 );
or \U$14634 ( \16377 , \16242 , \16376 );
xnor \U$14635 ( \16378 , \16199 , \16178 );
and \U$14636 ( \16379 , \16377 , \16378 );
or \U$14637 ( \16380 , \16200 , \16379 );
xnor \U$14638 ( \16381 , \16157 , \16136 );
and \U$14639 ( \16382 , \16380 , \16381 );
or \U$14640 ( \16383 , \16158 , \16382 );
xnor \U$14641 ( \16384 , \16115 , \16094 );
and \U$14642 ( \16385 , \16383 , \16384 );
or \U$14643 ( \16386 , \16116 , \16385 );
xnor \U$14644 ( \16387 , \16073 , \16052 );
and \U$14645 ( \16388 , \16386 , \16387 );
or \U$14646 ( \16389 , \16074 , \16388 );
xnor \U$14647 ( \16390 , \16031 , \16010 );
and \U$14648 ( \16391 , \16389 , \16390 );
or \U$14649 ( \16392 , \16032 , \16391 );
xnor \U$14650 ( \16393 , \15989 , \15968 );
and \U$14651 ( \16394 , \16392 , \16393 );
or \U$14652 ( \16395 , \15990 , \16394 );
xnor \U$14653 ( \16396 , \15947 , \15926 );
and \U$14654 ( \16397 , \16395 , \16396 );
or \U$14655 ( \16398 , \15948 , \16397 );
xnor \U$14656 ( \16399 , \15905 , \15884 );
and \U$14657 ( \16400 , \16398 , \16399 );
or \U$14658 ( \16401 , \15906 , \16400 );
xnor \U$14659 ( \16402 , \15863 , \15808 );
and \U$14660 ( \16403 , \16401 , \16402 );
or \U$14661 ( \16404 , \15864 , \16403 );
buf \U$14662 ( \16405 , \16404 );
and \U$14663 ( \16406 , \15754 , \16405 );
_HMUX g4ba1_GF_PartitionCandidate ( \16407_nG4ba1 , \12470_nG4b72 , \15316_nG4ba0 , \16406 );
buf \U$14664 ( \16408 , \16407_nG4ba1 );
not \U$14665 ( \16409 , \11933 );
nand \U$14666 ( \16410 , \12462 , \16409 );
nor \U$14667 ( \16411 , \12280 , \11116 );
nor \U$14668 ( \16412 , \11191 , \11268 );
nand \U$14669 ( \16413 , \16411 , \16412 );
nor \U$14670 ( \16414 , \11343 , \11420 );
nor \U$14671 ( \16415 , \11496 , \11569 );
nand \U$14672 ( \16416 , \16414 , \16415 );
nor \U$14673 ( \16417 , \16413 , \16416 );
nor \U$14674 ( \16418 , \11638 , \11702 );
nor \U$14675 ( \16419 , \11762 , \11819 );
nand \U$14676 ( \16420 , \16418 , \16419 );
nor \U$14677 ( \16421 , \11857 , \11889 );
nor \U$14678 ( \16422 , \11910 , \11926 );
nand \U$14679 ( \16423 , \16421 , \16422 );
nor \U$14680 ( \16424 , \16420 , \16423 );
nand \U$14681 ( \16425 , \16417 , \16424 );
nor \U$14682 ( \16426 , \12341 , \12045 );
nor \U$14683 ( \16427 , \12090 , \12142 );
nand \U$14684 ( \16428 , \16426 , \16427 );
nor \U$14685 ( \16429 , \12197 , \12236 );
nor \U$14686 ( \16430 , \12257 , \12273 );
nand \U$14687 ( \16431 , \16429 , \16430 );
nor \U$14688 ( \16432 , \16428 , \16431 );
nor \U$14689 ( \16433 , \12361 , \12316 );
nor \U$14690 ( \16434 , \12327 , \12338 );
nand \U$14691 ( \16435 , \16433 , \16434 );
nor \U$14692 ( \16436 , \12366 , \12358 );
not \U$14693 ( \16437 , \12374 );
and \U$14694 ( \16438 , \16436 , \16437 );
or \U$14695 ( \16439 , \12358 , \12376 );
nand \U$14696 ( \16440 , \16439 , \12379 );
nor \U$14697 ( \16441 , \16438 , \16440 );
or \U$14698 ( \16442 , \16435 , \16441 );
or \U$14699 ( \16443 , \12316 , \12381 );
nand \U$14700 ( \16444 , \16443 , \12385 );
and \U$14701 ( \16445 , \16434 , \16444 );
or \U$14702 ( \16446 , \12338 , \12387 );
nand \U$14703 ( \16447 , \16446 , \12390 );
nor \U$14704 ( \16448 , \16445 , \16447 );
nand \U$14705 ( \16449 , \16442 , \16448 );
and \U$14706 ( \16450 , \16432 , \16449 );
or \U$14707 ( \16451 , \12045 , \12392 );
nand \U$14708 ( \16452 , \16451 , \12397 );
and \U$14709 ( \16453 , \16427 , \16452 );
or \U$14710 ( \16454 , \12142 , \12399 );
nand \U$14711 ( \16455 , \16454 , \12402 );
nor \U$14712 ( \16456 , \16453 , \16455 );
or \U$14713 ( \16457 , \16431 , \16456 );
or \U$14714 ( \16458 , \12236 , \12404 );
nand \U$14715 ( \16459 , \16458 , \12408 );
and \U$14716 ( \16460 , \16430 , \16459 );
or \U$14717 ( \16461 , \12273 , \12410 );
nand \U$14718 ( \16462 , \16461 , \12413 );
nor \U$14719 ( \16463 , \16460 , \16462 );
nand \U$14720 ( \16464 , \16457 , \16463 );
nor \U$14721 ( \16465 , \16450 , \16464 );
or \U$14722 ( \16466 , \16425 , \16465 );
or \U$14723 ( \16467 , \11116 , \12415 );
nand \U$14724 ( \16468 , \16467 , \12421 );
and \U$14725 ( \16469 , \16412 , \16468 );
or \U$14726 ( \16470 , \11268 , \12423 );
nand \U$14727 ( \16471 , \16470 , \12426 );
nor \U$14728 ( \16472 , \16469 , \16471 );
or \U$14729 ( \16473 , \16416 , \16472 );
or \U$14730 ( \16474 , \11420 , \12428 );
nand \U$14731 ( \16475 , \16474 , \12432 );
and \U$14732 ( \16476 , \16415 , \16475 );
or \U$14733 ( \16477 , \11569 , \12434 );
nand \U$14734 ( \16478 , \16477 , \12437 );
nor \U$14735 ( \16479 , \16476 , \16478 );
nand \U$14736 ( \16480 , \16473 , \16479 );
and \U$14737 ( \16481 , \16424 , \16480 );
or \U$14738 ( \16482 , \11702 , \12439 );
nand \U$14739 ( \16483 , \16482 , \12444 );
and \U$14740 ( \16484 , \16419 , \16483 );
or \U$14741 ( \16485 , \11819 , \12446 );
nand \U$14742 ( \16486 , \16485 , \12449 );
nor \U$14743 ( \16487 , \16484 , \16486 );
or \U$14744 ( \16488 , \16423 , \16487 );
or \U$14745 ( \16489 , \11889 , \12451 );
nand \U$14746 ( \16490 , \16489 , \12455 );
and \U$14747 ( \16491 , \16422 , \16490 );
or \U$14748 ( \16492 , \11926 , \12457 );
nand \U$14749 ( \16493 , \16492 , \12460 );
nor \U$14750 ( \16494 , \16491 , \16493 );
nand \U$14751 ( \16495 , \16488 , \16494 );
nor \U$14752 ( \16496 , \16481 , \16495 );
nand \U$14753 ( \16497 , \16466 , \16496 );
not \U$14754 ( \16498 , \16497 );
xor \U$14755 ( \16499 , \16410 , \16498 );
buf g4b0f_GF_PartitionCandidate( \16500_nG4b0f , \16499 );
not \U$14756 ( \16501 , \14779 );
nand \U$14757 ( \16502 , \15308 , \16501 );
nor \U$14758 ( \16503 , \15126 , \13962 );
nor \U$14759 ( \16504 , \14037 , \14114 );
nand \U$14760 ( \16505 , \16503 , \16504 );
nor \U$14761 ( \16506 , \14189 , \14266 );
nor \U$14762 ( \16507 , \14342 , \14415 );
nand \U$14763 ( \16508 , \16506 , \16507 );
nor \U$14764 ( \16509 , \16505 , \16508 );
nor \U$14765 ( \16510 , \14484 , \14548 );
nor \U$14766 ( \16511 , \14608 , \14665 );
nand \U$14767 ( \16512 , \16510 , \16511 );
nor \U$14768 ( \16513 , \14703 , \14735 );
nor \U$14769 ( \16514 , \14756 , \14772 );
nand \U$14770 ( \16515 , \16513 , \16514 );
nor \U$14771 ( \16516 , \16512 , \16515 );
nand \U$14772 ( \16517 , \16509 , \16516 );
nor \U$14773 ( \16518 , \15187 , \14891 );
nor \U$14774 ( \16519 , \14936 , \14988 );
nand \U$14775 ( \16520 , \16518 , \16519 );
nor \U$14776 ( \16521 , \15043 , \15082 );
nor \U$14777 ( \16522 , \15103 , \15119 );
nand \U$14778 ( \16523 , \16521 , \16522 );
nor \U$14779 ( \16524 , \16520 , \16523 );
nor \U$14780 ( \16525 , \15207 , \15162 );
nor \U$14781 ( \16526 , \15173 , \15184 );
nand \U$14782 ( \16527 , \16525 , \16526 );
nor \U$14783 ( \16528 , \15212 , \15204 );
not \U$14784 ( \16529 , \15220 );
and \U$14785 ( \16530 , \16528 , \16529 );
or \U$14786 ( \16531 , \15204 , \15222 );
nand \U$14787 ( \16532 , \16531 , \15225 );
nor \U$14788 ( \16533 , \16530 , \16532 );
or \U$14789 ( \16534 , \16527 , \16533 );
or \U$14790 ( \16535 , \15162 , \15227 );
nand \U$14791 ( \16536 , \16535 , \15231 );
and \U$14792 ( \16537 , \16526 , \16536 );
or \U$14793 ( \16538 , \15184 , \15233 );
nand \U$14794 ( \16539 , \16538 , \15236 );
nor \U$14795 ( \16540 , \16537 , \16539 );
nand \U$14796 ( \16541 , \16534 , \16540 );
and \U$14797 ( \16542 , \16524 , \16541 );
or \U$14798 ( \16543 , \14891 , \15238 );
nand \U$14799 ( \16544 , \16543 , \15243 );
and \U$14800 ( \16545 , \16519 , \16544 );
or \U$14801 ( \16546 , \14988 , \15245 );
nand \U$14802 ( \16547 , \16546 , \15248 );
nor \U$14803 ( \16548 , \16545 , \16547 );
or \U$14804 ( \16549 , \16523 , \16548 );
or \U$14805 ( \16550 , \15082 , \15250 );
nand \U$14806 ( \16551 , \16550 , \15254 );
and \U$14807 ( \16552 , \16522 , \16551 );
or \U$14808 ( \16553 , \15119 , \15256 );
nand \U$14809 ( \16554 , \16553 , \15259 );
nor \U$14810 ( \16555 , \16552 , \16554 );
nand \U$14811 ( \16556 , \16549 , \16555 );
nor \U$14812 ( \16557 , \16542 , \16556 );
or \U$14813 ( \16558 , \16517 , \16557 );
or \U$14814 ( \16559 , \13962 , \15261 );
nand \U$14815 ( \16560 , \16559 , \15267 );
and \U$14816 ( \16561 , \16504 , \16560 );
or \U$14817 ( \16562 , \14114 , \15269 );
nand \U$14818 ( \16563 , \16562 , \15272 );
nor \U$14819 ( \16564 , \16561 , \16563 );
or \U$14820 ( \16565 , \16508 , \16564 );
or \U$14821 ( \16566 , \14266 , \15274 );
nand \U$14822 ( \16567 , \16566 , \15278 );
and \U$14823 ( \16568 , \16507 , \16567 );
or \U$14824 ( \16569 , \14415 , \15280 );
nand \U$14825 ( \16570 , \16569 , \15283 );
nor \U$14826 ( \16571 , \16568 , \16570 );
nand \U$14827 ( \16572 , \16565 , \16571 );
and \U$14828 ( \16573 , \16516 , \16572 );
or \U$14829 ( \16574 , \14548 , \15285 );
nand \U$14830 ( \16575 , \16574 , \15290 );
and \U$14831 ( \16576 , \16511 , \16575 );
or \U$14832 ( \16577 , \14665 , \15292 );
nand \U$14833 ( \16578 , \16577 , \15295 );
nor \U$14834 ( \16579 , \16576 , \16578 );
or \U$14835 ( \16580 , \16515 , \16579 );
or \U$14836 ( \16581 , \14735 , \15297 );
nand \U$14837 ( \16582 , \16581 , \15301 );
and \U$14838 ( \16583 , \16514 , \16582 );
or \U$14839 ( \16584 , \14772 , \15303 );
nand \U$14840 ( \16585 , \16584 , \15306 );
nor \U$14841 ( \16586 , \16583 , \16585 );
nand \U$14842 ( \16587 , \16580 , \16586 );
nor \U$14843 ( \16588 , \16573 , \16587 );
nand \U$14844 ( \16589 , \16558 , \16588 );
not \U$14845 ( \16590 , \16589 );
xor \U$14846 ( \16591 , \16502 , \16590 );
buf g4b43_GF_PartitionCandidate( \16592_nG4b43 , \16591 );
_HMUX g4b44_GF_PartitionCandidate ( \16593_nG4b44 , \16500_nG4b0f , \16592_nG4b43 , \16406 );
buf \U$14847 ( \16594 , \16593_nG4b44 );
not \U$14848 ( \16595 , \11926 );
nand \U$14849 ( \16596 , \12460 , \16595 );
nand \U$14850 ( \16597 , \12281 , \11192 );
nand \U$14851 ( \16598 , \11344 , \11497 );
nor \U$14852 ( \16599 , \16597 , \16598 );
nand \U$14853 ( \16600 , \11639 , \11763 );
nand \U$14854 ( \16601 , \11858 , \11911 );
nor \U$14855 ( \16602 , \16600 , \16601 );
nand \U$14856 ( \16603 , \16599 , \16602 );
nand \U$14857 ( \16604 , \12342 , \12091 );
nand \U$14858 ( \16605 , \12198 , \12258 );
nor \U$14859 ( \16606 , \16604 , \16605 );
nand \U$14860 ( \16607 , \12362 , \12328 );
not \U$14861 ( \16608 , \12377 );
or \U$14862 ( \16609 , \16607 , \16608 );
and \U$14863 ( \16610 , \12328 , \12382 );
nor \U$14864 ( \16611 , \16610 , \12388 );
nand \U$14865 ( \16612 , \16609 , \16611 );
and \U$14866 ( \16613 , \16606 , \16612 );
and \U$14867 ( \16614 , \12091 , \12393 );
nor \U$14868 ( \16615 , \16614 , \12400 );
or \U$14869 ( \16616 , \16605 , \16615 );
and \U$14870 ( \16617 , \12258 , \12405 );
nor \U$14871 ( \16618 , \16617 , \12411 );
nand \U$14872 ( \16619 , \16616 , \16618 );
nor \U$14873 ( \16620 , \16613 , \16619 );
or \U$14874 ( \16621 , \16603 , \16620 );
and \U$14875 ( \16622 , \11192 , \12416 );
nor \U$14876 ( \16623 , \16622 , \12424 );
or \U$14877 ( \16624 , \16598 , \16623 );
and \U$14878 ( \16625 , \11497 , \12429 );
nor \U$14879 ( \16626 , \16625 , \12435 );
nand \U$14880 ( \16627 , \16624 , \16626 );
and \U$14881 ( \16628 , \16602 , \16627 );
and \U$14882 ( \16629 , \11763 , \12440 );
nor \U$14883 ( \16630 , \16629 , \12447 );
or \U$14884 ( \16631 , \16601 , \16630 );
and \U$14885 ( \16632 , \11911 , \12452 );
nor \U$14886 ( \16633 , \16632 , \12458 );
nand \U$14887 ( \16634 , \16631 , \16633 );
nor \U$14888 ( \16635 , \16628 , \16634 );
nand \U$14889 ( \16636 , \16621 , \16635 );
not \U$14890 ( \16637 , \16636 );
xor \U$14891 ( \16638 , \16596 , \16637 );
buf g4aa0_GF_PartitionCandidate( \16639_nG4aa0 , \16638 );
not \U$14892 ( \16640 , \14772 );
nand \U$14893 ( \16641 , \15306 , \16640 );
nand \U$14894 ( \16642 , \15127 , \14038 );
nand \U$14895 ( \16643 , \14190 , \14343 );
nor \U$14896 ( \16644 , \16642 , \16643 );
nand \U$14897 ( \16645 , \14485 , \14609 );
nand \U$14898 ( \16646 , \14704 , \14757 );
nor \U$14899 ( \16647 , \16645 , \16646 );
nand \U$14900 ( \16648 , \16644 , \16647 );
nand \U$14901 ( \16649 , \15188 , \14937 );
nand \U$14902 ( \16650 , \15044 , \15104 );
nor \U$14903 ( \16651 , \16649 , \16650 );
nand \U$14904 ( \16652 , \15208 , \15174 );
not \U$14905 ( \16653 , \15223 );
or \U$14906 ( \16654 , \16652 , \16653 );
and \U$14907 ( \16655 , \15174 , \15228 );
nor \U$14908 ( \16656 , \16655 , \15234 );
nand \U$14909 ( \16657 , \16654 , \16656 );
and \U$14910 ( \16658 , \16651 , \16657 );
and \U$14911 ( \16659 , \14937 , \15239 );
nor \U$14912 ( \16660 , \16659 , \15246 );
or \U$14913 ( \16661 , \16650 , \16660 );
and \U$14914 ( \16662 , \15104 , \15251 );
nor \U$14915 ( \16663 , \16662 , \15257 );
nand \U$14916 ( \16664 , \16661 , \16663 );
nor \U$14917 ( \16665 , \16658 , \16664 );
or \U$14918 ( \16666 , \16648 , \16665 );
and \U$14919 ( \16667 , \14038 , \15262 );
nor \U$14920 ( \16668 , \16667 , \15270 );
or \U$14921 ( \16669 , \16643 , \16668 );
and \U$14922 ( \16670 , \14343 , \15275 );
nor \U$14923 ( \16671 , \16670 , \15281 );
nand \U$14924 ( \16672 , \16669 , \16671 );
and \U$14925 ( \16673 , \16647 , \16672 );
and \U$14926 ( \16674 , \14609 , \15286 );
nor \U$14927 ( \16675 , \16674 , \15293 );
or \U$14928 ( \16676 , \16646 , \16675 );
and \U$14929 ( \16677 , \14757 , \15298 );
nor \U$14930 ( \16678 , \16677 , \15304 );
nand \U$14931 ( \16679 , \16676 , \16678 );
nor \U$14932 ( \16680 , \16673 , \16679 );
nand \U$14933 ( \16681 , \16666 , \16680 );
not \U$14934 ( \16682 , \16681 );
xor \U$14935 ( \16683 , \16641 , \16682 );
buf g4ada_GF_PartitionCandidate( \16684_nG4ada , \16683 );
_HMUX g4adb_GF_PartitionCandidate ( \16685_nG4adb , \16639_nG4aa0 , \16684_nG4ada , \16406 );
buf \U$14936 ( \16686 , \16685_nG4adb );
not \U$14937 ( \16687 , \11910 );
nand \U$14938 ( \16688 , \12457 , \16687 );
nand \U$14939 ( \16689 , \16430 , \16411 );
nand \U$14940 ( \16690 , \16412 , \16414 );
nor \U$14941 ( \16691 , \16689 , \16690 );
nand \U$14942 ( \16692 , \16415 , \16418 );
nand \U$14943 ( \16693 , \16419 , \16421 );
nor \U$14944 ( \16694 , \16692 , \16693 );
nand \U$14945 ( \16695 , \16691 , \16694 );
nand \U$14946 ( \16696 , \16434 , \16426 );
nand \U$14947 ( \16697 , \16427 , \16429 );
nor \U$14948 ( \16698 , \16696 , \16697 );
nand \U$14949 ( \16699 , \16436 , \16433 );
or \U$14950 ( \16700 , \16699 , \12374 );
and \U$14951 ( \16701 , \16433 , \16440 );
nor \U$14952 ( \16702 , \16701 , \16444 );
nand \U$14953 ( \16703 , \16700 , \16702 );
and \U$14954 ( \16704 , \16698 , \16703 );
and \U$14955 ( \16705 , \16426 , \16447 );
nor \U$14956 ( \16706 , \16705 , \16452 );
or \U$14957 ( \16707 , \16697 , \16706 );
and \U$14958 ( \16708 , \16429 , \16455 );
nor \U$14959 ( \16709 , \16708 , \16459 );
nand \U$14960 ( \16710 , \16707 , \16709 );
nor \U$14961 ( \16711 , \16704 , \16710 );
or \U$14962 ( \16712 , \16695 , \16711 );
and \U$14963 ( \16713 , \16411 , \16462 );
nor \U$14964 ( \16714 , \16713 , \16468 );
or \U$14965 ( \16715 , \16690 , \16714 );
and \U$14966 ( \16716 , \16414 , \16471 );
nor \U$14967 ( \16717 , \16716 , \16475 );
nand \U$14968 ( \16718 , \16715 , \16717 );
and \U$14969 ( \16719 , \16694 , \16718 );
and \U$14970 ( \16720 , \16418 , \16478 );
nor \U$14971 ( \16721 , \16720 , \16483 );
or \U$14972 ( \16722 , \16693 , \16721 );
and \U$14973 ( \16723 , \16421 , \16486 );
nor \U$14974 ( \16724 , \16723 , \16490 );
nand \U$14975 ( \16725 , \16722 , \16724 );
nor \U$14976 ( \16726 , \16719 , \16725 );
nand \U$14977 ( \16727 , \16712 , \16726 );
not \U$14978 ( \16728 , \16727 );
xor \U$14979 ( \16729 , \16688 , \16728 );
buf g4a23_GF_PartitionCandidate( \16730_nG4a23 , \16729 );
not \U$14980 ( \16731 , \14756 );
nand \U$14981 ( \16732 , \15303 , \16731 );
nand \U$14982 ( \16733 , \16522 , \16503 );
nand \U$14983 ( \16734 , \16504 , \16506 );
nor \U$14984 ( \16735 , \16733 , \16734 );
nand \U$14985 ( \16736 , \16507 , \16510 );
nand \U$14986 ( \16737 , \16511 , \16513 );
nor \U$14987 ( \16738 , \16736 , \16737 );
nand \U$14988 ( \16739 , \16735 , \16738 );
nand \U$14989 ( \16740 , \16526 , \16518 );
nand \U$14990 ( \16741 , \16519 , \16521 );
nor \U$14991 ( \16742 , \16740 , \16741 );
nand \U$14992 ( \16743 , \16528 , \16525 );
or \U$14993 ( \16744 , \16743 , \15220 );
and \U$14994 ( \16745 , \16525 , \16532 );
nor \U$14995 ( \16746 , \16745 , \16536 );
nand \U$14996 ( \16747 , \16744 , \16746 );
and \U$14997 ( \16748 , \16742 , \16747 );
and \U$14998 ( \16749 , \16518 , \16539 );
nor \U$14999 ( \16750 , \16749 , \16544 );
or \U$15000 ( \16751 , \16741 , \16750 );
and \U$15001 ( \16752 , \16521 , \16547 );
nor \U$15002 ( \16753 , \16752 , \16551 );
nand \U$15003 ( \16754 , \16751 , \16753 );
nor \U$15004 ( \16755 , \16748 , \16754 );
or \U$15005 ( \16756 , \16739 , \16755 );
and \U$15006 ( \16757 , \16503 , \16554 );
nor \U$15007 ( \16758 , \16757 , \16560 );
or \U$15008 ( \16759 , \16734 , \16758 );
and \U$15009 ( \16760 , \16506 , \16563 );
nor \U$15010 ( \16761 , \16760 , \16567 );
nand \U$15011 ( \16762 , \16759 , \16761 );
and \U$15012 ( \16763 , \16738 , \16762 );
and \U$15013 ( \16764 , \16510 , \16570 );
nor \U$15014 ( \16765 , \16764 , \16575 );
or \U$15015 ( \16766 , \16737 , \16765 );
and \U$15016 ( \16767 , \16513 , \16578 );
nor \U$15017 ( \16768 , \16767 , \16582 );
nand \U$15018 ( \16769 , \16766 , \16768 );
nor \U$15019 ( \16770 , \16763 , \16769 );
nand \U$15020 ( \16771 , \16756 , \16770 );
not \U$15021 ( \16772 , \16771 );
xor \U$15022 ( \16773 , \16732 , \16772 );
buf g4a65_GF_PartitionCandidate( \16774_nG4a65 , \16773 );
_HMUX g4a66_GF_PartitionCandidate ( \16775_nG4a66 , \16730_nG4a23 , \16774_nG4a65 , \16406 );
buf \U$15023 ( \16776 , \16775_nG4a66 );
not \U$15024 ( \16777 , \11889 );
nand \U$15025 ( \16778 , \12455 , \16777 );
nor \U$15026 ( \16779 , \12282 , \11345 );
nor \U$15027 ( \16780 , \11640 , \11859 );
nand \U$15028 ( \16781 , \16779 , \16780 );
nor \U$15029 ( \16782 , \12343 , \12199 );
not \U$15030 ( \16783 , \12383 );
and \U$15031 ( \16784 , \16782 , \16783 );
or \U$15032 ( \16785 , \12199 , \12394 );
nand \U$15033 ( \16786 , \16785 , \12406 );
nor \U$15034 ( \16787 , \16784 , \16786 );
or \U$15035 ( \16788 , \16781 , \16787 );
or \U$15036 ( \16789 , \11345 , \12417 );
nand \U$15037 ( \16790 , \16789 , \12430 );
and \U$15038 ( \16791 , \16780 , \16790 );
or \U$15039 ( \16792 , \11859 , \12441 );
nand \U$15040 ( \16793 , \16792 , \12453 );
nor \U$15041 ( \16794 , \16791 , \16793 );
nand \U$15042 ( \16795 , \16788 , \16794 );
not \U$15043 ( \16796 , \16795 );
xor \U$15044 ( \16797 , \16778 , \16796 );
buf g499a_GF_PartitionCandidate( \16798_nG499a , \16797 );
not \U$15045 ( \16799 , \14735 );
nand \U$15046 ( \16800 , \15301 , \16799 );
nor \U$15047 ( \16801 , \15128 , \14191 );
nor \U$15048 ( \16802 , \14486 , \14705 );
nand \U$15049 ( \16803 , \16801 , \16802 );
nor \U$15050 ( \16804 , \15189 , \15045 );
not \U$15051 ( \16805 , \15229 );
and \U$15052 ( \16806 , \16804 , \16805 );
or \U$15053 ( \16807 , \15045 , \15240 );
nand \U$15054 ( \16808 , \16807 , \15252 );
nor \U$15055 ( \16809 , \16806 , \16808 );
or \U$15056 ( \16810 , \16803 , \16809 );
or \U$15057 ( \16811 , \14191 , \15263 );
nand \U$15058 ( \16812 , \16811 , \15276 );
and \U$15059 ( \16813 , \16802 , \16812 );
or \U$15060 ( \16814 , \14705 , \15287 );
nand \U$15061 ( \16815 , \16814 , \15299 );
nor \U$15062 ( \16816 , \16813 , \16815 );
nand \U$15063 ( \16817 , \16810 , \16816 );
not \U$15064 ( \16818 , \16817 );
xor \U$15065 ( \16819 , \16800 , \16818 );
buf g49e0_GF_PartitionCandidate( \16820_nG49e0 , \16819 );
_HMUX g49e1_GF_PartitionCandidate ( \16821_nG49e1 , \16798_nG499a , \16820_nG49e0 , \16406 );
buf \U$15066 ( \16822 , \16821_nG49e1 );
not \U$15067 ( \16823 , \11857 );
nand \U$15068 ( \16824 , \12451 , \16823 );
nor \U$15069 ( \16825 , \16431 , \16413 );
nor \U$15070 ( \16826 , \16416 , \16420 );
nand \U$15071 ( \16827 , \16825 , \16826 );
nor \U$15072 ( \16828 , \16435 , \16428 );
not \U$15073 ( \16829 , \16441 );
and \U$15074 ( \16830 , \16828 , \16829 );
or \U$15075 ( \16831 , \16428 , \16448 );
nand \U$15076 ( \16832 , \16831 , \16456 );
nor \U$15077 ( \16833 , \16830 , \16832 );
or \U$15078 ( \16834 , \16827 , \16833 );
or \U$15079 ( \16835 , \16413 , \16463 );
nand \U$15080 ( \16836 , \16835 , \16472 );
and \U$15081 ( \16837 , \16826 , \16836 );
or \U$15082 ( \16838 , \16420 , \16479 );
nand \U$15083 ( \16839 , \16838 , \16487 );
nor \U$15084 ( \16840 , \16837 , \16839 );
nand \U$15085 ( \16841 , \16834 , \16840 );
not \U$15086 ( \16842 , \16841 );
xor \U$15087 ( \16843 , \16824 , \16842 );
buf g490b_GF_PartitionCandidate( \16844_nG490b , \16843 );
not \U$15088 ( \16845 , \14703 );
nand \U$15089 ( \16846 , \15297 , \16845 );
nor \U$15090 ( \16847 , \16523 , \16505 );
nor \U$15091 ( \16848 , \16508 , \16512 );
nand \U$15092 ( \16849 , \16847 , \16848 );
nor \U$15093 ( \16850 , \16527 , \16520 );
not \U$15094 ( \16851 , \16533 );
and \U$15095 ( \16852 , \16850 , \16851 );
or \U$15096 ( \16853 , \16520 , \16540 );
nand \U$15097 ( \16854 , \16853 , \16548 );
nor \U$15098 ( \16855 , \16852 , \16854 );
or \U$15099 ( \16856 , \16849 , \16855 );
or \U$15100 ( \16857 , \16505 , \16555 );
nand \U$15101 ( \16858 , \16857 , \16564 );
and \U$15102 ( \16859 , \16848 , \16858 );
or \U$15103 ( \16860 , \16512 , \16571 );
nand \U$15104 ( \16861 , \16860 , \16579 );
nor \U$15105 ( \16862 , \16859 , \16861 );
nand \U$15106 ( \16863 , \16856 , \16862 );
not \U$15107 ( \16864 , \16863 );
xor \U$15108 ( \16865 , \16846 , \16864 );
buf g4953_GF_PartitionCandidate( \16866_nG4953 , \16865 );
_HMUX g4954_GF_PartitionCandidate ( \16867_nG4954 , \16844_nG490b , \16866_nG4953 , \16406 );
buf \U$15109 ( \16868 , \16867_nG4954 );
not \U$15110 ( \16869 , \11819 );
nand \U$15111 ( \16870 , \12449 , \16869 );
nor \U$15112 ( \16871 , \16605 , \16597 );
nor \U$15113 ( \16872 , \16598 , \16600 );
nand \U$15114 ( \16873 , \16871 , \16872 );
nor \U$15115 ( \16874 , \16607 , \16604 );
and \U$15116 ( \16875 , \16874 , \12377 );
or \U$15117 ( \16876 , \16604 , \16611 );
nand \U$15118 ( \16877 , \16876 , \16615 );
nor \U$15119 ( \16878 , \16875 , \16877 );
or \U$15120 ( \16879 , \16873 , \16878 );
or \U$15121 ( \16880 , \16597 , \16618 );
nand \U$15122 ( \16881 , \16880 , \16623 );
and \U$15123 ( \16882 , \16872 , \16881 );
or \U$15124 ( \16883 , \16600 , \16626 );
nand \U$15125 ( \16884 , \16883 , \16630 );
nor \U$15126 ( \16885 , \16882 , \16884 );
nand \U$15127 ( \16886 , \16879 , \16885 );
not \U$15128 ( \16887 , \16886 );
xor \U$15129 ( \16888 , \16870 , \16887 );
buf g4876_GF_PartitionCandidate( \16889_nG4876 , \16888 );
not \U$15130 ( \16890 , \14665 );
nand \U$15131 ( \16891 , \15295 , \16890 );
nor \U$15132 ( \16892 , \16650 , \16642 );
nor \U$15133 ( \16893 , \16643 , \16645 );
nand \U$15134 ( \16894 , \16892 , \16893 );
nor \U$15135 ( \16895 , \16652 , \16649 );
and \U$15136 ( \16896 , \16895 , \15223 );
or \U$15137 ( \16897 , \16649 , \16656 );
nand \U$15138 ( \16898 , \16897 , \16660 );
nor \U$15139 ( \16899 , \16896 , \16898 );
or \U$15140 ( \16900 , \16894 , \16899 );
or \U$15141 ( \16901 , \16642 , \16663 );
nand \U$15142 ( \16902 , \16901 , \16668 );
and \U$15143 ( \16903 , \16893 , \16902 );
or \U$15144 ( \16904 , \16645 , \16671 );
nand \U$15145 ( \16905 , \16904 , \16675 );
nor \U$15146 ( \16906 , \16903 , \16905 );
nand \U$15147 ( \16907 , \16900 , \16906 );
not \U$15148 ( \16908 , \16907 );
xor \U$15149 ( \16909 , \16891 , \16908 );
buf g48c2_GF_PartitionCandidate( \16910_nG48c2 , \16909 );
_HMUX g48c3_GF_PartitionCandidate ( \16911_nG48c3 , \16889_nG4876 , \16910_nG48c2 , \16406 );
buf \U$15150 ( \16912 , \16911_nG48c3 );
not \U$15151 ( \16913 , \11762 );
nand \U$15152 ( \16914 , \12446 , \16913 );
nor \U$15153 ( \16915 , \16697 , \16689 );
nor \U$15154 ( \16916 , \16690 , \16692 );
nand \U$15155 ( \16917 , \16915 , \16916 );
nor \U$15156 ( \16918 , \16699 , \16696 );
and \U$15157 ( \16919 , \16918 , \16437 );
or \U$15158 ( \16920 , \16696 , \16702 );
nand \U$15159 ( \16921 , \16920 , \16706 );
nor \U$15160 ( \16922 , \16919 , \16921 );
or \U$15161 ( \16923 , \16917 , \16922 );
or \U$15162 ( \16924 , \16689 , \16709 );
nand \U$15163 ( \16925 , \16924 , \16714 );
and \U$15164 ( \16926 , \16916 , \16925 );
or \U$15165 ( \16927 , \16692 , \16717 );
nand \U$15166 ( \16928 , \16927 , \16721 );
nor \U$15167 ( \16929 , \16926 , \16928 );
nand \U$15168 ( \16930 , \16923 , \16929 );
not \U$15169 ( \16931 , \16930 );
xor \U$15170 ( \16932 , \16914 , \16931 );
buf g47d9_GF_PartitionCandidate( \16933_nG47d9 , \16932 );
not \U$15171 ( \16934 , \14608 );
nand \U$15172 ( \16935 , \15292 , \16934 );
nor \U$15173 ( \16936 , \16741 , \16733 );
nor \U$15174 ( \16937 , \16734 , \16736 );
nand \U$15175 ( \16938 , \16936 , \16937 );
nor \U$15176 ( \16939 , \16743 , \16740 );
and \U$15177 ( \16940 , \16939 , \16529 );
or \U$15178 ( \16941 , \16740 , \16746 );
nand \U$15179 ( \16942 , \16941 , \16750 );
nor \U$15180 ( \16943 , \16940 , \16942 );
or \U$15181 ( \16944 , \16938 , \16943 );
or \U$15182 ( \16945 , \16733 , \16753 );
nand \U$15183 ( \16946 , \16945 , \16758 );
and \U$15184 ( \16947 , \16937 , \16946 );
or \U$15185 ( \16948 , \16736 , \16761 );
nand \U$15186 ( \16949 , \16948 , \16765 );
nor \U$15187 ( \16950 , \16947 , \16949 );
nand \U$15188 ( \16951 , \16944 , \16950 );
not \U$15189 ( \16952 , \16951 );
xor \U$15190 ( \16953 , \16935 , \16952 );
buf g4829_GF_PartitionCandidate( \16954_nG4829 , \16953 );
_HMUX g482a_GF_PartitionCandidate ( \16955_nG482a , \16933_nG47d9 , \16954_nG4829 , \16406 );
buf \U$15191 ( \16956 , \16955_nG482a );
not \U$15192 ( \16957 , \11702 );
nand \U$15193 ( \16958 , \12444 , \16957 );
nand \U$15194 ( \16959 , \12283 , \11641 );
not \U$15195 ( \16960 , \12395 );
or \U$15196 ( \16961 , \16959 , \16960 );
and \U$15197 ( \16962 , \11641 , \12418 );
nor \U$15198 ( \16963 , \16962 , \12442 );
nand \U$15199 ( \16964 , \16961 , \16963 );
not \U$15200 ( \16965 , \16964 );
xor \U$15201 ( \16966 , \16958 , \16965 );
buf g4737_GF_PartitionCandidate( \16967_nG4737 , \16966 );
not \U$15202 ( \16968 , \14548 );
nand \U$15203 ( \16969 , \15290 , \16968 );
nand \U$15204 ( \16970 , \15129 , \14487 );
not \U$15205 ( \16971 , \15241 );
or \U$15206 ( \16972 , \16970 , \16971 );
and \U$15207 ( \16973 , \14487 , \15264 );
nor \U$15208 ( \16974 , \16973 , \15288 );
nand \U$15209 ( \16975 , \16972 , \16974 );
not \U$15210 ( \16976 , \16975 );
xor \U$15211 ( \16977 , \16969 , \16976 );
buf g4788_GF_PartitionCandidate( \16978_nG4788 , \16977 );
_HMUX g4789_GF_PartitionCandidate ( \16979_nG4789 , \16967_nG4737 , \16978_nG4788 , \16406 );
buf \U$15212 ( \16980 , \16979_nG4789 );
not \U$15213 ( \16981 , \11638 );
nand \U$15214 ( \16982 , \12439 , \16981 );
nand \U$15215 ( \16983 , \16432 , \16417 );
not \U$15216 ( \16984 , \16449 );
or \U$15217 ( \16985 , \16983 , \16984 );
and \U$15218 ( \16986 , \16417 , \16464 );
nor \U$15219 ( \16987 , \16986 , \16480 );
nand \U$15220 ( \16988 , \16985 , \16987 );
not \U$15221 ( \16989 , \16988 );
xor \U$15222 ( \16990 , \16982 , \16989 );
buf g468c_GF_PartitionCandidate( \16991_nG468c , \16990 );
not \U$15223 ( \16992 , \14484 );
nand \U$15224 ( \16993 , \15285 , \16992 );
nand \U$15225 ( \16994 , \16524 , \16509 );
not \U$15226 ( \16995 , \16541 );
or \U$15227 ( \16996 , \16994 , \16995 );
and \U$15228 ( \16997 , \16509 , \16556 );
nor \U$15229 ( \16998 , \16997 , \16572 );
nand \U$15230 ( \16999 , \16996 , \16998 );
not \U$15231 ( \17000 , \16999 );
xor \U$15232 ( \17001 , \16993 , \17000 );
buf g46e5_GF_PartitionCandidate( \17002_nG46e5 , \17001 );
_HMUX g46e6_GF_PartitionCandidate ( \17003_nG46e6 , \16991_nG468c , \17002_nG46e5 , \16406 );
buf \U$15233 ( \17004 , \17003_nG46e6 );
not \U$15234 ( \17005 , \11569 );
nand \U$15235 ( \17006 , \12437 , \17005 );
nand \U$15236 ( \17007 , \16606 , \16599 );
not \U$15237 ( \17008 , \16612 );
or \U$15238 ( \17009 , \17007 , \17008 );
and \U$15239 ( \17010 , \16599 , \16619 );
nor \U$15240 ( \17011 , \17010 , \16627 );
nand \U$15241 ( \17012 , \17009 , \17011 );
not \U$15242 ( \17013 , \17012 );
xor \U$15243 ( \17014 , \17006 , \17013 );
buf g45d6_GF_PartitionCandidate( \17015_nG45d6 , \17014 );
not \U$15244 ( \17016 , \14415 );
nand \U$15245 ( \17017 , \15283 , \17016 );
nand \U$15246 ( \17018 , \16651 , \16644 );
not \U$15247 ( \17019 , \16657 );
or \U$15248 ( \17020 , \17018 , \17019 );
and \U$15249 ( \17021 , \16644 , \16664 );
nor \U$15250 ( \17022 , \17021 , \16672 );
nand \U$15251 ( \17023 , \17020 , \17022 );
not \U$15252 ( \17024 , \17023 );
xor \U$15253 ( \17025 , \17017 , \17024 );
buf g4632_GF_PartitionCandidate( \17026_nG4632 , \17025 );
_HMUX g4633_GF_PartitionCandidate ( \17027_nG4633 , \17015_nG45d6 , \17026_nG4632 , \16406 );
buf \U$15254 ( \17028 , \17027_nG4633 );
not \U$15255 ( \17029 , \11496 );
nand \U$15256 ( \17030 , \12434 , \17029 );
nand \U$15257 ( \17031 , \16698 , \16691 );
not \U$15258 ( \17032 , \16703 );
or \U$15259 ( \17033 , \17031 , \17032 );
and \U$15260 ( \17034 , \16691 , \16710 );
nor \U$15261 ( \17035 , \17034 , \16718 );
nand \U$15262 ( \17036 , \17033 , \17035 );
not \U$15263 ( \17037 , \17036 );
xor \U$15264 ( \17038 , \17030 , \17037 );
buf g4519_GF_PartitionCandidate( \17039_nG4519 , \17038 );
not \U$15265 ( \17040 , \14342 );
nand \U$15266 ( \17041 , \15280 , \17040 );
nand \U$15267 ( \17042 , \16742 , \16735 );
not \U$15268 ( \17043 , \16747 );
or \U$15269 ( \17044 , \17042 , \17043 );
and \U$15270 ( \17045 , \16735 , \16754 );
nor \U$15271 ( \17046 , \17045 , \16762 );
nand \U$15272 ( \17047 , \17044 , \17046 );
not \U$15273 ( \17048 , \17047 );
xor \U$15274 ( \17049 , \17041 , \17048 );
buf g4579_GF_PartitionCandidate( \17050_nG4579 , \17049 );
_HMUX g457a_GF_PartitionCandidate ( \17051_nG457a , \17039_nG4519 , \17050_nG4579 , \16406 );
buf \U$15275 ( \17052 , \17051_nG457a );
not \U$15276 ( \17053 , \11420 );
nand \U$15277 ( \17054 , \12432 , \17053 );
nand \U$15278 ( \17055 , \16782 , \16779 );
or \U$15279 ( \17056 , \17055 , \12383 );
and \U$15280 ( \17057 , \16779 , \16786 );
nor \U$15281 ( \17058 , \17057 , \16790 );
nand \U$15282 ( \17059 , \17056 , \17058 );
not \U$15283 ( \17060 , \17059 );
xor \U$15284 ( \17061 , \17054 , \17060 );
buf g4459_GF_PartitionCandidate( \17062_nG4459 , \17061 );
not \U$15285 ( \17063 , \14266 );
nand \U$15286 ( \17064 , \15278 , \17063 );
nand \U$15287 ( \17065 , \16804 , \16801 );
or \U$15288 ( \17066 , \17065 , \15229 );
and \U$15289 ( \17067 , \16801 , \16808 );
nor \U$15290 ( \17068 , \17067 , \16812 );
nand \U$15291 ( \17069 , \17066 , \17068 );
not \U$15292 ( \17070 , \17069 );
xor \U$15293 ( \17071 , \17064 , \17070 );
buf g44b8_GF_PartitionCandidate( \17072_nG44b8 , \17071 );
_HMUX g44b9_GF_PartitionCandidate ( \17073_nG44b9 , \17062_nG4459 , \17072_nG44b8 , \16406 );
buf \U$15294 ( \17074 , \17073_nG44b9 );
not \U$15295 ( \17075 , \11343 );
nand \U$15296 ( \17076 , \12428 , \17075 );
nand \U$15297 ( \17077 , \16828 , \16825 );
or \U$15298 ( \17078 , \17077 , \16441 );
and \U$15299 ( \17079 , \16825 , \16832 );
nor \U$15300 ( \17080 , \17079 , \16836 );
nand \U$15301 ( \17081 , \17078 , \17080 );
not \U$15302 ( \17082 , \17081 );
xor \U$15303 ( \17083 , \17076 , \17082 );
buf g439a_GF_PartitionCandidate( \17084_nG439a , \17083 );
not \U$15304 ( \17085 , \14189 );
nand \U$15305 ( \17086 , \15274 , \17085 );
nand \U$15306 ( \17087 , \16850 , \16847 );
or \U$15307 ( \17088 , \17087 , \16533 );
and \U$15308 ( \17089 , \16847 , \16854 );
nor \U$15309 ( \17090 , \17089 , \16858 );
nand \U$15310 ( \17091 , \17088 , \17090 );
not \U$15311 ( \17092 , \17091 );
xor \U$15312 ( \17093 , \17086 , \17092 );
buf g43f9_GF_PartitionCandidate( \17094_nG43f9 , \17093 );
_HMUX g43fa_GF_PartitionCandidate ( \17095_nG43fa , \17084_nG439a , \17094_nG43f9 , \16406 );
buf \U$15313 ( \17096 , \17095_nG43fa );
not \U$15314 ( \17097 , \11268 );
nand \U$15315 ( \17098 , \12426 , \17097 );
nand \U$15316 ( \17099 , \16874 , \16871 );
or \U$15317 ( \17100 , \17099 , \16608 );
and \U$15318 ( \17101 , \16871 , \16877 );
nor \U$15319 ( \17102 , \17101 , \16881 );
nand \U$15320 ( \17103 , \17100 , \17102 );
not \U$15321 ( \17104 , \17103 );
xor \U$15322 ( \17105 , \17098 , \17104 );
buf g42c6_GF_PartitionCandidate( \17106_nG42c6 , \17105 );
not \U$15323 ( \17107 , \14114 );
nand \U$15324 ( \17108 , \15272 , \17107 );
nand \U$15325 ( \17109 , \16895 , \16892 );
or \U$15326 ( \17110 , \17109 , \16653 );
and \U$15327 ( \17111 , \16892 , \16898 );
nor \U$15328 ( \17112 , \17111 , \16902 );
nand \U$15329 ( \17113 , \17110 , \17112 );
not \U$15330 ( \17114 , \17113 );
xor \U$15331 ( \17115 , \17108 , \17114 );
buf g433a_GF_PartitionCandidate( \17116_nG433a , \17115 );
_HMUX g433b_GF_PartitionCandidate ( \17117_nG433b , \17106_nG42c6 , \17116_nG433a , \16406 );
buf \U$15332 ( \17118 , \17117_nG433b );
not \U$15333 ( \17119 , \11191 );
nand \U$15334 ( \17120 , \12423 , \17119 );
nand \U$15335 ( \17121 , \16918 , \16915 );
or \U$15336 ( \17122 , \17121 , \12374 );
and \U$15337 ( \17123 , \16915 , \16921 );
nor \U$15338 ( \17124 , \17123 , \16925 );
nand \U$15339 ( \17125 , \17122 , \17124 );
not \U$15340 ( \17126 , \17125 );
xor \U$15341 ( \17127 , \17120 , \17126 );
buf g41de_GF_PartitionCandidate( \17128_nG41de , \17127 );
not \U$15342 ( \17129 , \14037 );
nand \U$15343 ( \17130 , \15269 , \17129 );
nand \U$15344 ( \17131 , \16939 , \16936 );
or \U$15345 ( \17132 , \17131 , \15220 );
and \U$15346 ( \17133 , \16936 , \16942 );
nor \U$15347 ( \17134 , \17133 , \16946 );
nand \U$15348 ( \17135 , \17132 , \17134 );
not \U$15349 ( \17136 , \17135 );
xor \U$15350 ( \17137 , \17130 , \17136 );
buf g4251_GF_PartitionCandidate( \17138_nG4251 , \17137 );
_HMUX g4252_GF_PartitionCandidate ( \17139_nG4252 , \17128_nG41de , \17138_nG4251 , \16406 );
buf \U$15351 ( \17140 , \17139_nG4252 );
not \U$15352 ( \17141 , \11116 );
nand \U$15353 ( \17142 , \12421 , \17141 );
xor \U$15354 ( \17143 , \17142 , \12419 );
buf g40fe_GF_PartitionCandidate( \17144_nG40fe , \17143 );
not \U$15355 ( \17145 , \13962 );
nand \U$15356 ( \17146 , \15267 , \17145 );
xor \U$15357 ( \17147 , \17146 , \15265 );
buf g416a_GF_PartitionCandidate( \17148_nG416a , \17147 );
_HMUX g416b_GF_PartitionCandidate ( \17149_nG416b , \17144_nG40fe , \17148_nG416a , \16406 );
buf \U$15358 ( \17150 , \17149_nG416b );
not \U$15359 ( \17151 , \12280 );
nand \U$15360 ( \17152 , \12415 , \17151 );
xor \U$15361 ( \17153 , \17152 , \16465 );
buf g4025_GF_PartitionCandidate( \17154_nG4025 , \17153 );
not \U$15362 ( \17155 , \15126 );
nand \U$15363 ( \17156 , \15261 , \17155 );
xor \U$15364 ( \17157 , \17156 , \16557 );
buf g4091_GF_PartitionCandidate( \17158_nG4091 , \17157 );
_HMUX g4092_GF_PartitionCandidate ( \17159_nG4092 , \17154_nG4025 , \17158_nG4091 , \16406 );
buf \U$15365 ( \17160 , \17159_nG4092 );
not \U$15366 ( \17161 , \12273 );
nand \U$15367 ( \17162 , \12413 , \17161 );
xor \U$15368 ( \17163 , \17162 , \16620 );
buf g3f50_GF_PartitionCandidate( \17164_nG3f50 , \17163 );
not \U$15369 ( \17165 , \15119 );
nand \U$15370 ( \17166 , \15259 , \17165 );
xor \U$15371 ( \17167 , \17166 , \16665 );
buf g3fb8_GF_PartitionCandidate( \17168_nG3fb8 , \17167 );
_HMUX g3fb9_GF_PartitionCandidate ( \17169_nG3fb9 , \17164_nG3f50 , \17168_nG3fb8 , \16406 );
buf \U$15372 ( \17170 , \17169_nG3fb9 );
not \U$15373 ( \17171 , \12257 );
nand \U$15374 ( \17172 , \12410 , \17171 );
xor \U$15375 ( \17173 , \17172 , \16711 );
buf g3e7d_GF_PartitionCandidate( \17174_nG3e7d , \17173 );
not \U$15376 ( \17175 , \15103 );
nand \U$15377 ( \17176 , \15256 , \17175 );
xor \U$15378 ( \17177 , \17176 , \16755 );
buf g3ee7_GF_PartitionCandidate( \17178_nG3ee7 , \17177 );
_HMUX g3ee8_GF_PartitionCandidate ( \17179_nG3ee8 , \17174_nG3e7d , \17178_nG3ee7 , \16406 );
buf \U$15379 ( \17180 , \17179_nG3ee8 );
not \U$15380 ( \17181 , \12236 );
nand \U$15381 ( \17182 , \12408 , \17181 );
xor \U$15382 ( \17183 , \17182 , \16787 );
buf g3dad_GF_PartitionCandidate( \17184_nG3dad , \17183 );
not \U$15383 ( \17185 , \15082 );
nand \U$15384 ( \17186 , \15254 , \17185 );
xor \U$15385 ( \17187 , \17186 , \16809 );
buf g3e12_GF_PartitionCandidate( \17188_nG3e12 , \17187 );
_HMUX g3e13_GF_PartitionCandidate ( \17189_nG3e13 , \17184_nG3dad , \17188_nG3e12 , \16406 );
buf \U$15386 ( \17190 , \17189_nG3e13 );
not \U$15387 ( \17191 , \12197 );
nand \U$15388 ( \17192 , \12404 , \17191 );
xor \U$15389 ( \17193 , \17192 , \16833 );
buf g3cbb_GF_PartitionCandidate( \17194_nG3cbb , \17193 );
not \U$15390 ( \17195 , \15043 );
nand \U$15391 ( \17196 , \15250 , \17195 );
xor \U$15392 ( \17197 , \17196 , \16855 );
buf g3d47_GF_PartitionCandidate( \17198_nG3d47 , \17197 );
_HMUX g3d48_GF_PartitionCandidate ( \17199_nG3d48 , \17194_nG3cbb , \17198_nG3d47 , \16406 );
buf \U$15393 ( \17200 , \17199_nG3d48 );
not \U$15394 ( \17201 , \12142 );
nand \U$15395 ( \17202 , \12402 , \17201 );
xor \U$15396 ( \17203 , \17202 , \16878 );
buf g3bd4_GF_PartitionCandidate( \17204_nG3bd4 , \17203 );
not \U$15397 ( \17205 , \14988 );
nand \U$15398 ( \17206 , \15248 , \17205 );
xor \U$15399 ( \17207 , \17206 , \16899 );
buf g3c2e_GF_PartitionCandidate( \17208_nG3c2e , \17207 );
_HMUX g3c2f_GF_PartitionCandidate ( \17209_nG3c2f , \17204_nG3bd4 , \17208_nG3c2e , \16406 );
buf \U$15400 ( \17210 , \17209_nG3c2f );
not \U$15401 ( \17211 , \12090 );
nand \U$15402 ( \17212 , \12399 , \17211 );
xor \U$15403 ( \17213 , \17212 , \16922 );
buf g3ae0_GF_PartitionCandidate( \17214_nG3ae0 , \17213 );
not \U$15404 ( \17215 , \14936 );
nand \U$15405 ( \17216 , \15245 , \17215 );
xor \U$15406 ( \17217 , \17216 , \16943 );
buf g3b79_GF_PartitionCandidate( \17218_nG3b79 , \17217 );
_HMUX g3b7a_GF_PartitionCandidate ( \17219_nG3b7a , \17214_nG3ae0 , \17218_nG3b79 , \16406 );
buf \U$15407 ( \17220 , \17219_nG3b7a );
not \U$15408 ( \17221 , \12045 );
nand \U$15409 ( \17222 , \12397 , \17221 );
xor \U$15410 ( \17223 , \17222 , \16960 );
buf g39f8_GF_PartitionCandidate( \17224_nG39f8 , \17223 );
not \U$15411 ( \17225 , \14891 );
nand \U$15412 ( \17226 , \15243 , \17225 );
xor \U$15413 ( \17227 , \17226 , \16971 );
buf g3a46_GF_PartitionCandidate( \17228_nG3a46 , \17227 );
_HMUX g3a47_GF_PartitionCandidate ( \17229_nG3a47 , \17224_nG39f8 , \17228_nG3a46 , \16406 );
buf \U$15414 ( \17230 , \17229_nG3a47 );
not \U$15415 ( \17231 , \12341 );
nand \U$15416 ( \17232 , \12392 , \17231 );
xor \U$15417 ( \17233 , \17232 , \16984 );
buf g391c_GF_PartitionCandidate( \17234_nG391c , \17233 );
not \U$15418 ( \17235 , \15187 );
nand \U$15419 ( \17236 , \15238 , \17235 );
xor \U$15420 ( \17237 , \17236 , \16995 );
buf g39a9_GF_PartitionCandidate( \17238_nG39a9 , \17237 );
_HMUX g39aa_GF_PartitionCandidate ( \17239_nG39aa , \17234_nG391c , \17238_nG39a9 , \16406 );
buf \U$15421 ( \17240 , \17239_nG39aa );
not \U$15422 ( \17241 , \12338 );
nand \U$15423 ( \17242 , \12390 , \17241 );
xor \U$15424 ( \17243 , \17242 , \17008 );
buf g384a_GF_PartitionCandidate( \17244_nG384a , \17243 );
not \U$15425 ( \17245 , \15184 );
nand \U$15426 ( \17246 , \15236 , \17245 );
xor \U$15427 ( \17247 , \17246 , \17019 );
buf g388e_GF_PartitionCandidate( \17248_nG388e , \17247 );
_HMUX g388f_GF_PartitionCandidate ( \17249_nG388f , \17244_nG384a , \17248_nG388e , \16406 );
buf \U$15428 ( \17250 , \17249_nG388f );
endmodule

