//
// Conformal-LEC Version 20.10-d130 (26-Jun-2020)
//
module top(RI2b5e785ebcf0_2,RI2b5e785ebc78_3,RI2b5e785ebc00_4,RI2b5e785ebb88_5,RI2b5e785ebb10_6,RI2b5e785eba98_7,RI2b5e785eba20_8,RI2b5e785eb9a8_9,RI2b5e785eb930_10,
        RI2b5e785eb8b8_11,RI2b5e785eb840_12,RI2b5e785daa40_28,RI2b5e785ae9b8_600,RI2b5e785aea30_599,RI2b5e785aeaa8_598,RI2b5e785aeb20_597,RI2b5e785aeb98_596,RI2b5e78549540_41,RI2b5e785388a8_54,
        RI2b5e784a6330_67,RI2b5e78495698_80,RI2b5e78495080_93,RI2b5e78403b80_106,RI2b5e775b1e60_119,RI2b5e7750bdf8_132,RI2b5e774ff5d0_145,RI2b5e774f65e8_158,RI2b5e774eabd0_171,RI2b5e774de3a8_184,
        RI2b5e774d53c0_197,RI2b5e785f4300_210,RI2b5e785f3ce8_223,RI2b5e785eb0c0_236,RI2b5e785da9c8_29,RI2b5e785494c8_42,RI2b5e78538830_55,RI2b5e784a62b8_68,RI2b5e78495620_81,RI2b5e78495008_94,
        RI2b5e78403b08_107,RI2b5e775b1de8_120,RI2b5e7750bd80_133,RI2b5e774ff558_146,RI2b5e774f6570_159,RI2b5e774eab58_172,RI2b5e774de330_185,RI2b5e774d5348_198,RI2b5e785f4288_211,RI2b5e785f3658_224,
        RI2b5e785eb048_237,RI2b5e785da950_30,RI2b5e78549450_43,RI2b5e785387b8_56,RI2b5e784a6240_69,RI2b5e784955a8_82,RI2b5e78494f90_95,RI2b5e78403a90_108,RI2b5e775b1d70_121,RI2b5e7750bd08_134,
        RI2b5e774ff4e0_147,RI2b5e774f64f8_160,RI2b5e774eaae0_173,RI2b5e774de2b8_186,RI2b5e774d52d0_199,RI2b5e785f4210_212,RI2b5e785eb5e8_225,RI2b5e785e6c50_238,RI2b5e785da8d8_31,RI2b5e785493d8_44,
        RI2b5e78538740_57,RI2b5e784a61c8_70,RI2b5e78495530_83,RI2b5e78494f18_96,RI2b5e78403a18_109,RI2b5e775b1cf8_122,RI2b5e7750bc90_135,RI2b5e774ff468_148,RI2b5e774f6480_161,RI2b5e774eaa68_174,
        RI2b5e774de240_187,RI2b5e774d5258_200,RI2b5e785f4198_213,RI2b5e785eb570_226,RI2b5e785e6bd8_239,RI2b5e785da860_32,RI2b5e78549360_45,RI2b5e785386c8_58,RI2b5e784a6150_71,RI2b5e784954b8_84,
        RI2b5e78494ea0_97,RI2b5e784039a0_110,RI2b5e775b1c80_123,RI2b5e7750bc18_136,RI2b5e774ff3f0_149,RI2b5e774f6408_162,RI2b5e774ea9f0_175,RI2b5e774de1c8_188,RI2b5e774d51e0_201,RI2b5e785f4120_214,
        RI2b5e785eb4f8_227,RI2b5e785e64d0_240,RI2b5e78549900_33,RI2b5e78538c68_46,RI2b5e78538650_59,RI2b5e784a60d8_72,RI2b5e78495440_85,RI2b5e78494e28_98,RI2b5e78403928_111,RI2b5e775b1c08_124,
        RI2b5e7750bba0_137,RI2b5e774ff378_150,RI2b5e774f6390_163,RI2b5e774ea978_176,RI2b5e774de150_189,RI2b5e774d5168_202,RI2b5e785f40a8_215,RI2b5e785eb480_228,RI2b5e785da608_241,RI2b5e78549888_34,
        RI2b5e78538bf0_47,RI2b5e785385d8_60,RI2b5e784a6060_73,RI2b5e784953c8_86,RI2b5e78403ec8_99,RI2b5e775b21a8_112,RI2b5e775b1b90_125,RI2b5e7750bb28_138,RI2b5e774ff300_151,RI2b5e774f6318_164,
        RI2b5e774ea900_177,RI2b5e774de0d8_190,RI2b5e774d50f0_203,RI2b5e785f4030_216,RI2b5e785eb408_229,RI2b5e785da590_242,RI2b5e78549810_35,RI2b5e78538b78_48,RI2b5e78538560_61,RI2b5e784a5fe8_74,
        RI2b5e78495350_87,RI2b5e78403e50_100,RI2b5e775b2130_113,RI2b5e775b1b18_126,RI2b5e7750bab0_139,RI2b5e774ff288_152,RI2b5e774f62a0_165,RI2b5e774ea888_178,RI2b5e774de060_191,RI2b5e774d5078_204,
        RI2b5e785f3fb8_217,RI2b5e785eb390_230,RI2b5e785da518_243,RI2b5e78549798_36,RI2b5e78538b00_49,RI2b5e785384e8_62,RI2b5e784a5f70_75,RI2b5e784952d8_88,RI2b5e78403dd8_101,RI2b5e775b20b8_114,
        RI2b5e775b1aa0_127,RI2b5e7750ba38_140,RI2b5e774ff210_153,RI2b5e774f6228_166,RI2b5e774ea810_179,RI2b5e774ddfe8_192,RI2b5e774d5000_205,RI2b5e785f3f40_218,RI2b5e785eb318_231,RI2b5e785da4a0_244,
        RI2b5e78549720_37,RI2b5e78538a88_50,RI2b5e78538470_63,RI2b5e784a5ef8_76,RI2b5e78495260_89,RI2b5e78403d60_102,RI2b5e775b2040_115,RI2b5e775b1a28_128,RI2b5e7750b9c0_141,RI2b5e774ff198_154,
        RI2b5e774f61b0_167,RI2b5e774ea798_180,RI2b5e774ddf70_193,RI2b5e774d4f88_206,RI2b5e785f3ec8_219,RI2b5e785eb2a0_232,RI2b5e785da428_245,RI2b5e785496a8_38,RI2b5e78538a10_51,RI2b5e785383f8_64,
        RI2b5e784a5e80_77,RI2b5e784951e8_90,RI2b5e78403ce8_103,RI2b5e775b1fc8_116,RI2b5e775b19b0_129,RI2b5e7750b948_142,RI2b5e774ff120_155,RI2b5e774f6138_168,RI2b5e774ea720_181,RI2b5e774ddef8_194,
        RI2b5e774d4f10_207,RI2b5e785f3e50_220,RI2b5e785eb228_233,RI2b5e785da3b0_246,RI2b5e785db148_13,RI2b5e78549630_39,RI2b5e78538998_52,RI2b5e78538380_65,RI2b5e784a5e08_78,RI2b5e78495170_91,
        RI2b5e78403c70_104,RI2b5e775b1f50_117,RI2b5e775b1938_130,RI2b5e7750b8d0_143,RI2b5e774ff0a8_156,RI2b5e774f60c0_169,RI2b5e774ea6a8_182,RI2b5e774dde80_195,RI2b5e774d4e98_208,RI2b5e785f3dd8_221,
        RI2b5e785eb1b0_234,RI2b5e785da338_247,RI2b5e785da248_249,RI2b5e785aec10_595,RI2b5e785aec88_594,RI2b5e785aed00_593,RI2b5e785aed78_592,RI2b5e785aedf0_591,RI2b5e785aee68_590,RI2b5e785aeee0_589,
        RI2b5e785aef58_588,RI2b5e785be750_269,RI2b5e785bc4a0_289,RI2b5e785bbb40_309,RI2b5e785b9c50_329,RI2b5e785b8120_349,RI2b5e785b77c0_369,RI2b5e785b6e60_389,RI2b5e785b56f0_409,RI2b5e785b4d90_429,
        RI2b5e785b39e0_449,RI2b5e785b3080_469,RI2b5e785b2720_489,RI2b5e785b1730_509,RI2b5e785b0dd0_529,RI2b5e785b0470_549,RI2b5e785af840_569,RI2b5e785ebd68_1,RI2b5e785daab8_27,RI2b5e785495b8_40,
        RI2b5e78538920_53,RI2b5e784a63a8_66,RI2b5e78495710_79,RI2b5e784950f8_92,RI2b5e78403bf8_105,RI2b5e775b1ed8_118,RI2b5e775b18c0_131,RI2b5e7750b858_144,RI2b5e774ff030_157,RI2b5e774f6048_170,
        RI2b5e774ea630_183,RI2b5e774dde08_196,RI2b5e774d4e20_209,RI2b5e785f3d60_222,RI2b5e785eb138_235,RI2b5e785da2c0_248,RI2b5e785be7c8_268,RI2b5e785bc518_288,RI2b5e785bbbb8_308,RI2b5e785b9cc8_328,
        RI2b5e785b9368_348,RI2b5e785b7838_368,RI2b5e785b6ed8_388,RI2b5e785b5768_408,RI2b5e785b4e08_428,RI2b5e785b3a58_448,RI2b5e785b30f8_468,RI2b5e785b2798_488,RI2b5e785b17a8_508,RI2b5e785b0e48_528,
        RI2b5e785b04e8_548,RI2b5e785afb88_568,RI2b5e785da1d0_250,RI2b5e785be6d8_270,RI2b5e785bc428_290,RI2b5e785bbac8_310,RI2b5e785b9bd8_330,RI2b5e785b80a8_350,RI2b5e785b7748_370,RI2b5e785b6de8_390,
        RI2b5e785b5678_410,RI2b5e785b4d18_430,RI2b5e785b3968_450,RI2b5e785b3008_470,RI2b5e785b26a8_490,RI2b5e785b16b8_510,RI2b5e785b0d58_530,RI2b5e785b03f8_550,RI2b5e785af7c8_570,RI2b5e785da0e0_252,
        RI2b5e785be5e8_272,RI2b5e785bc338_292,RI2b5e785bb9d8_312,RI2b5e785b9ae8_332,RI2b5e785b7fb8_352,RI2b5e785b7658_372,RI2b5e785b5ee8_392,RI2b5e785b5588_412,RI2b5e785b4c28_432,RI2b5e785b3878_452,
        RI2b5e785b2f18_472,RI2b5e785b25b8_492,RI2b5e785b15c8_512,RI2b5e785b0c68_532,RI2b5e785b0308_552,RI2b5e785af6d8_572,RI2b5e785da158_251,RI2b5e785be660_271,RI2b5e785bc3b0_291,RI2b5e785bba50_311,
        RI2b5e785b9b60_331,RI2b5e785b8030_351,RI2b5e785b76d0_371,RI2b5e785b6d70_391,RI2b5e785b5600_411,RI2b5e785b4ca0_431,RI2b5e785b38f0_451,RI2b5e785b2f90_471,RI2b5e785b2630_491,RI2b5e785b1640_511,
        RI2b5e785b0ce0_531,RI2b5e785b0380_551,RI2b5e785af750_571,RI2b5e785da068_253,RI2b5e785be570_273,RI2b5e785bc2c0_293,RI2b5e785bb960_313,RI2b5e785b9a70_333,RI2b5e785b7f40_353,RI2b5e785b75e0_373,
        RI2b5e785b5e70_393,RI2b5e785b5510_413,RI2b5e785b4bb0_433,RI2b5e785b3800_453,RI2b5e785b2ea0_473,RI2b5e785b2540_493,RI2b5e785b1550_513,RI2b5e785b0bf0_533,RI2b5e785b0290_553,RI2b5e785af660_573,
        RI2b5e785c2bc0_255,RI2b5e785be480_275,RI2b5e785bc1d0_295,RI2b5e785ba2e0_315,RI2b5e785b9980_335,RI2b5e785b7e50_355,RI2b5e785b74f0_375,RI2b5e785b5d80_395,RI2b5e785b5420_415,RI2b5e785b4ac0_435,
        RI2b5e785b3710_455,RI2b5e785b2db0_475,RI2b5e785b2450_495,RI2b5e785b1460_515,RI2b5e785b0b00_535,RI2b5e785b01a0_555,RI2b5e785af570_575,RI2b5e785c2c38_254,RI2b5e785be4f8_274,RI2b5e785bc248_294,
        RI2b5e785ba358_314,RI2b5e785b99f8_334,RI2b5e785b7ec8_354,RI2b5e785b7568_374,RI2b5e785b5df8_394,RI2b5e785b5498_414,RI2b5e785b4b38_434,RI2b5e785b3788_454,RI2b5e785b2e28_474,RI2b5e785b24c8_494,
        RI2b5e785b14d8_514,RI2b5e785b0b78_534,RI2b5e785b0218_554,RI2b5e785af5e8_574,RI2b5e785c0a00_257,RI2b5e785be390_277,RI2b5e785bc0e0_297,RI2b5e785ba1f0_317,RI2b5e785b9890_337,RI2b5e785b7d60_357,
        RI2b5e785b7400_377,RI2b5e785b5c90_397,RI2b5e785b5330_417,RI2b5e785b49d0_437,RI2b5e785b3620_457,RI2b5e785b2cc0_477,RI2b5e785b2360_497,RI2b5e785b1370_517,RI2b5e785b0a10_537,RI2b5e785b00b0_557,
        RI2b5e785af480_577,RI2b5e785c2b48_256,RI2b5e785be408_276,RI2b5e785bc158_296,RI2b5e785ba268_316,RI2b5e785b9908_336,RI2b5e785b7dd8_356,RI2b5e785b7478_376,RI2b5e785b5d08_396,RI2b5e785b53a8_416,
        RI2b5e785b4a48_436,RI2b5e785b3698_456,RI2b5e785b2d38_476,RI2b5e785b23d8_496,RI2b5e785b13e8_516,RI2b5e785b0a88_536,RI2b5e785b0128_556,RI2b5e785af4f8_576,RI2b5e785c0910_259,RI2b5e785be2a0_279,
        RI2b5e785bbff0_299,RI2b5e785ba100_319,RI2b5e785b97a0_339,RI2b5e785b7c70_359,RI2b5e785b7310_379,RI2b5e785b5ba0_399,RI2b5e785b5240_419,RI2b5e785b48e0_439,RI2b5e785b3530_459,RI2b5e785b2bd0_479,
        RI2b5e785b2270_499,RI2b5e785b1280_519,RI2b5e785b0920_539,RI2b5e785affc0_559,RI2b5e785af390_579,RI2b5e785c0988_258,RI2b5e785be318_278,RI2b5e785bc068_298,RI2b5e785ba178_318,RI2b5e785b9818_338,
        RI2b5e785b7ce8_358,RI2b5e785b7388_378,RI2b5e785b5c18_398,RI2b5e785b52b8_418,RI2b5e785b4958_438,RI2b5e785b35a8_458,RI2b5e785b2c48_478,RI2b5e785b22e8_498,RI2b5e785b12f8_518,RI2b5e785b0998_538,
        RI2b5e785b0038_558,RI2b5e785af408_578,RI2b5e785c0820_261,RI2b5e785be1b0_281,RI2b5e785bbf00_301,RI2b5e785ba010_321,RI2b5e785b96b0_341,RI2b5e785b7b80_361,RI2b5e785b7220_381,RI2b5e785b5ab0_401,
        RI2b5e785b5150_421,RI2b5e785b47f0_441,RI2b5e785b3440_461,RI2b5e785b2ae0_481,RI2b5e785b2180_501,RI2b5e785b1190_521,RI2b5e785b0830_541,RI2b5e785afed0_561,RI2b5e785af2a0_581,RI2b5e785c0898_260,
        RI2b5e785be228_280,RI2b5e785bbf78_300,RI2b5e785ba088_320,RI2b5e785b9728_340,RI2b5e785b7bf8_360,RI2b5e785b7298_380,RI2b5e785b5b28_400,RI2b5e785b51c8_420,RI2b5e785b4868_440,RI2b5e785b34b8_460,
        RI2b5e785b2b58_480,RI2b5e785b21f8_500,RI2b5e785b1208_520,RI2b5e785b08a8_540,RI2b5e785aff48_560,RI2b5e785af318_580,RI2b5e785c0730_263,RI2b5e785be0c0_283,RI2b5e785bbe10_303,RI2b5e785b9f20_323,
        RI2b5e785b95c0_343,RI2b5e785b7a90_363,RI2b5e785b7130_383,RI2b5e785b59c0_403,RI2b5e785b5060_423,RI2b5e785b3cb0_443,RI2b5e785b3350_463,RI2b5e785b29f0_483,RI2b5e785b1a00_503,RI2b5e785b10a0_523,
        RI2b5e785b0740_543,RI2b5e785afde0_563,RI2b5e785af1b0_583,RI2b5e785c07a8_262,RI2b5e785be138_282,RI2b5e785bbe88_302,RI2b5e785b9f98_322,RI2b5e785b9638_342,RI2b5e785b7b08_362,RI2b5e785b71a8_382,
        RI2b5e785b5a38_402,RI2b5e785b50d8_422,RI2b5e785b4778_442,RI2b5e785b33c8_462,RI2b5e785b2a68_482,RI2b5e785b1a78_502,RI2b5e785b1118_522,RI2b5e785b07b8_542,RI2b5e785afe58_562,RI2b5e785af228_582,
        RI2b5e785c0640_265,RI2b5e785bdfd0_285,RI2b5e785bbd20_305,RI2b5e785b9e30_325,RI2b5e785b94d0_345,RI2b5e785b79a0_365,RI2b5e785b7040_385,RI2b5e785b58d0_405,RI2b5e785b4f70_425,RI2b5e785b3bc0_445,
        RI2b5e785b3260_465,RI2b5e785b2900_485,RI2b5e785b1910_505,RI2b5e785b0fb0_525,RI2b5e785b0650_545,RI2b5e785afcf0_565,RI2b5e785af0c0_585,RI2b5e785c06b8_264,RI2b5e785be048_284,RI2b5e785bbd98_304,
        RI2b5e785b9ea8_324,RI2b5e785b9548_344,RI2b5e785b7a18_364,RI2b5e785b70b8_384,RI2b5e785b5948_404,RI2b5e785b4fe8_424,RI2b5e785b3c38_444,RI2b5e785b32d8_464,RI2b5e785b2978_484,RI2b5e785b1988_504,
        RI2b5e785b1028_524,RI2b5e785b06c8_544,RI2b5e785afd68_564,RI2b5e785af138_584,RI2b5e785c05c8_266,RI2b5e785bdf58_286,RI2b5e785bbca8_306,RI2b5e785b9db8_326,RI2b5e785b9458_346,RI2b5e785b7928_366,
        RI2b5e785b6fc8_386,RI2b5e785b5858_406,RI2b5e785b4ef8_426,RI2b5e785b3b48_446,RI2b5e785b31e8_466,RI2b5e785b2888_486,RI2b5e785b1898_506,RI2b5e785b0f38_526,RI2b5e785b05d8_546,RI2b5e785afc78_566,
        RI2b5e785af048_586,RI2b5e785c0550_267,RI2b5e785bc590_287,RI2b5e785bbc30_307,RI2b5e785b9d40_327,RI2b5e785b93e0_347,RI2b5e785b78b0_367,RI2b5e785b6f50_387,RI2b5e785b57e0_407,RI2b5e785b4e80_427,
        RI2b5e785b3ad0_447,RI2b5e785b3170_467,RI2b5e785b2810_487,RI2b5e785b1820_507,RI2b5e785b0ec0_527,RI2b5e785b0560_547,RI2b5e785afc00_567,RI2b5e785aefd0_587,RI2b5e785ae328_614,RI2b5e785db058_15,
        RI2b5e785dafe0_16,RI2b5e785daf68_17,RI2b5e785daef0_18,RI2b5e785dae78_19,RI2b5e785dae00_20,RI2b5e785dad88_21,RI2b5e785dad10_22,RI2b5e785dac98_23,RI2b5e785dac20_24,RI2b5e785daba8_25,
        RI2b5e785ae3a0_613,RI2b5e785ae418_612,RI2b5e785ae490_611,RI2b5e785ae508_610,RI2b5e785ae580_609,RI2b5e785dab30_26,RI2b5e785ae5f8_608,RI2b5e785ae670_607,RI2b5e785ae6e8_606,RI2b5e785ae760_605,
        RI2b5e785ae7d8_604,RI2b5e785ae850_603,RI2b5e785ae8c8_602,RI2b5e785ae940_601,RI2b5e785db0d0_14,R_267_b04ddc8,R_268_b04de70,R_269_b04df18,R_26a_b04dfc0,R_26b_b04e068,
        R_26c_b04e110,R_26d_b04e1b8,R_26e_b04e260,R_26f_b04e308,R_270_b04e3b0,R_271_b04e458,R_272_b04e500,R_273_b04e5a8,R_274_b04e650,R_275_b04e6f8,
        R_276_b04e7a0,R_277_b04e848,R_278_b04e8f0,R_279_b04e998,R_27a_b04ea40,R_27b_b04eae8,R_27c_b04eb90,R_27d_b04ec38,R_27e_b04ece0,R_27f_b04ed88,
        R_280_b04ee30,R_281_b04eed8,R_282_b04ef80,R_283_b04f028,R_284_b04f0d0,R_285_b04f178,R_286_b04f220,R_287_b04f2c8,R_288_b04f370,R_289_b04f418,
        R_28a_b04f4c0,R_28b_b04f568,R_28c_b04f610,R_28d_b04f6b8,R_28e_b04f760,R_28f_b04f808,R_290_b04f8b0,R_291_b04f958,R_292_b04fa00,R_293_b04faa8,
        R_294_b04fb50,R_295_b04fbf8,R_296_b04fca0,R_297_b04fd48,R_298_b04fdf0,R_299_b04fe98,R_29a_b04ff40,R_29b_b04ffe8,R_29c_b050090,R_29d_b050138,
        R_29e_b0501e0,R_29f_b050288,R_2a0_b050330,R_2a1_b0503d8,R_2a2_b050480,R_2a3_b050528,R_2a4_b0505d0,R_2a5_b050678,R_2a6_b050720,R_2a7_b0507c8,
        R_2a8_b050870,R_2a9_b050918,R_2aa_b0509c0);
input RI2b5e785ebcf0_2,RI2b5e785ebc78_3,RI2b5e785ebc00_4,RI2b5e785ebb88_5,RI2b5e785ebb10_6,RI2b5e785eba98_7,RI2b5e785eba20_8,RI2b5e785eb9a8_9,RI2b5e785eb930_10,
        RI2b5e785eb8b8_11,RI2b5e785eb840_12,RI2b5e785daa40_28,RI2b5e785ae9b8_600,RI2b5e785aea30_599,RI2b5e785aeaa8_598,RI2b5e785aeb20_597,RI2b5e785aeb98_596,RI2b5e78549540_41,RI2b5e785388a8_54,
        RI2b5e784a6330_67,RI2b5e78495698_80,RI2b5e78495080_93,RI2b5e78403b80_106,RI2b5e775b1e60_119,RI2b5e7750bdf8_132,RI2b5e774ff5d0_145,RI2b5e774f65e8_158,RI2b5e774eabd0_171,RI2b5e774de3a8_184,
        RI2b5e774d53c0_197,RI2b5e785f4300_210,RI2b5e785f3ce8_223,RI2b5e785eb0c0_236,RI2b5e785da9c8_29,RI2b5e785494c8_42,RI2b5e78538830_55,RI2b5e784a62b8_68,RI2b5e78495620_81,RI2b5e78495008_94,
        RI2b5e78403b08_107,RI2b5e775b1de8_120,RI2b5e7750bd80_133,RI2b5e774ff558_146,RI2b5e774f6570_159,RI2b5e774eab58_172,RI2b5e774de330_185,RI2b5e774d5348_198,RI2b5e785f4288_211,RI2b5e785f3658_224,
        RI2b5e785eb048_237,RI2b5e785da950_30,RI2b5e78549450_43,RI2b5e785387b8_56,RI2b5e784a6240_69,RI2b5e784955a8_82,RI2b5e78494f90_95,RI2b5e78403a90_108,RI2b5e775b1d70_121,RI2b5e7750bd08_134,
        RI2b5e774ff4e0_147,RI2b5e774f64f8_160,RI2b5e774eaae0_173,RI2b5e774de2b8_186,RI2b5e774d52d0_199,RI2b5e785f4210_212,RI2b5e785eb5e8_225,RI2b5e785e6c50_238,RI2b5e785da8d8_31,RI2b5e785493d8_44,
        RI2b5e78538740_57,RI2b5e784a61c8_70,RI2b5e78495530_83,RI2b5e78494f18_96,RI2b5e78403a18_109,RI2b5e775b1cf8_122,RI2b5e7750bc90_135,RI2b5e774ff468_148,RI2b5e774f6480_161,RI2b5e774eaa68_174,
        RI2b5e774de240_187,RI2b5e774d5258_200,RI2b5e785f4198_213,RI2b5e785eb570_226,RI2b5e785e6bd8_239,RI2b5e785da860_32,RI2b5e78549360_45,RI2b5e785386c8_58,RI2b5e784a6150_71,RI2b5e784954b8_84,
        RI2b5e78494ea0_97,RI2b5e784039a0_110,RI2b5e775b1c80_123,RI2b5e7750bc18_136,RI2b5e774ff3f0_149,RI2b5e774f6408_162,RI2b5e774ea9f0_175,RI2b5e774de1c8_188,RI2b5e774d51e0_201,RI2b5e785f4120_214,
        RI2b5e785eb4f8_227,RI2b5e785e64d0_240,RI2b5e78549900_33,RI2b5e78538c68_46,RI2b5e78538650_59,RI2b5e784a60d8_72,RI2b5e78495440_85,RI2b5e78494e28_98,RI2b5e78403928_111,RI2b5e775b1c08_124,
        RI2b5e7750bba0_137,RI2b5e774ff378_150,RI2b5e774f6390_163,RI2b5e774ea978_176,RI2b5e774de150_189,RI2b5e774d5168_202,RI2b5e785f40a8_215,RI2b5e785eb480_228,RI2b5e785da608_241,RI2b5e78549888_34,
        RI2b5e78538bf0_47,RI2b5e785385d8_60,RI2b5e784a6060_73,RI2b5e784953c8_86,RI2b5e78403ec8_99,RI2b5e775b21a8_112,RI2b5e775b1b90_125,RI2b5e7750bb28_138,RI2b5e774ff300_151,RI2b5e774f6318_164,
        RI2b5e774ea900_177,RI2b5e774de0d8_190,RI2b5e774d50f0_203,RI2b5e785f4030_216,RI2b5e785eb408_229,RI2b5e785da590_242,RI2b5e78549810_35,RI2b5e78538b78_48,RI2b5e78538560_61,RI2b5e784a5fe8_74,
        RI2b5e78495350_87,RI2b5e78403e50_100,RI2b5e775b2130_113,RI2b5e775b1b18_126,RI2b5e7750bab0_139,RI2b5e774ff288_152,RI2b5e774f62a0_165,RI2b5e774ea888_178,RI2b5e774de060_191,RI2b5e774d5078_204,
        RI2b5e785f3fb8_217,RI2b5e785eb390_230,RI2b5e785da518_243,RI2b5e78549798_36,RI2b5e78538b00_49,RI2b5e785384e8_62,RI2b5e784a5f70_75,RI2b5e784952d8_88,RI2b5e78403dd8_101,RI2b5e775b20b8_114,
        RI2b5e775b1aa0_127,RI2b5e7750ba38_140,RI2b5e774ff210_153,RI2b5e774f6228_166,RI2b5e774ea810_179,RI2b5e774ddfe8_192,RI2b5e774d5000_205,RI2b5e785f3f40_218,RI2b5e785eb318_231,RI2b5e785da4a0_244,
        RI2b5e78549720_37,RI2b5e78538a88_50,RI2b5e78538470_63,RI2b5e784a5ef8_76,RI2b5e78495260_89,RI2b5e78403d60_102,RI2b5e775b2040_115,RI2b5e775b1a28_128,RI2b5e7750b9c0_141,RI2b5e774ff198_154,
        RI2b5e774f61b0_167,RI2b5e774ea798_180,RI2b5e774ddf70_193,RI2b5e774d4f88_206,RI2b5e785f3ec8_219,RI2b5e785eb2a0_232,RI2b5e785da428_245,RI2b5e785496a8_38,RI2b5e78538a10_51,RI2b5e785383f8_64,
        RI2b5e784a5e80_77,RI2b5e784951e8_90,RI2b5e78403ce8_103,RI2b5e775b1fc8_116,RI2b5e775b19b0_129,RI2b5e7750b948_142,RI2b5e774ff120_155,RI2b5e774f6138_168,RI2b5e774ea720_181,RI2b5e774ddef8_194,
        RI2b5e774d4f10_207,RI2b5e785f3e50_220,RI2b5e785eb228_233,RI2b5e785da3b0_246,RI2b5e785db148_13,RI2b5e78549630_39,RI2b5e78538998_52,RI2b5e78538380_65,RI2b5e784a5e08_78,RI2b5e78495170_91,
        RI2b5e78403c70_104,RI2b5e775b1f50_117,RI2b5e775b1938_130,RI2b5e7750b8d0_143,RI2b5e774ff0a8_156,RI2b5e774f60c0_169,RI2b5e774ea6a8_182,RI2b5e774dde80_195,RI2b5e774d4e98_208,RI2b5e785f3dd8_221,
        RI2b5e785eb1b0_234,RI2b5e785da338_247,RI2b5e785da248_249,RI2b5e785aec10_595,RI2b5e785aec88_594,RI2b5e785aed00_593,RI2b5e785aed78_592,RI2b5e785aedf0_591,RI2b5e785aee68_590,RI2b5e785aeee0_589,
        RI2b5e785aef58_588,RI2b5e785be750_269,RI2b5e785bc4a0_289,RI2b5e785bbb40_309,RI2b5e785b9c50_329,RI2b5e785b8120_349,RI2b5e785b77c0_369,RI2b5e785b6e60_389,RI2b5e785b56f0_409,RI2b5e785b4d90_429,
        RI2b5e785b39e0_449,RI2b5e785b3080_469,RI2b5e785b2720_489,RI2b5e785b1730_509,RI2b5e785b0dd0_529,RI2b5e785b0470_549,RI2b5e785af840_569,RI2b5e785ebd68_1,RI2b5e785daab8_27,RI2b5e785495b8_40,
        RI2b5e78538920_53,RI2b5e784a63a8_66,RI2b5e78495710_79,RI2b5e784950f8_92,RI2b5e78403bf8_105,RI2b5e775b1ed8_118,RI2b5e775b18c0_131,RI2b5e7750b858_144,RI2b5e774ff030_157,RI2b5e774f6048_170,
        RI2b5e774ea630_183,RI2b5e774dde08_196,RI2b5e774d4e20_209,RI2b5e785f3d60_222,RI2b5e785eb138_235,RI2b5e785da2c0_248,RI2b5e785be7c8_268,RI2b5e785bc518_288,RI2b5e785bbbb8_308,RI2b5e785b9cc8_328,
        RI2b5e785b9368_348,RI2b5e785b7838_368,RI2b5e785b6ed8_388,RI2b5e785b5768_408,RI2b5e785b4e08_428,RI2b5e785b3a58_448,RI2b5e785b30f8_468,RI2b5e785b2798_488,RI2b5e785b17a8_508,RI2b5e785b0e48_528,
        RI2b5e785b04e8_548,RI2b5e785afb88_568,RI2b5e785da1d0_250,RI2b5e785be6d8_270,RI2b5e785bc428_290,RI2b5e785bbac8_310,RI2b5e785b9bd8_330,RI2b5e785b80a8_350,RI2b5e785b7748_370,RI2b5e785b6de8_390,
        RI2b5e785b5678_410,RI2b5e785b4d18_430,RI2b5e785b3968_450,RI2b5e785b3008_470,RI2b5e785b26a8_490,RI2b5e785b16b8_510,RI2b5e785b0d58_530,RI2b5e785b03f8_550,RI2b5e785af7c8_570,RI2b5e785da0e0_252,
        RI2b5e785be5e8_272,RI2b5e785bc338_292,RI2b5e785bb9d8_312,RI2b5e785b9ae8_332,RI2b5e785b7fb8_352,RI2b5e785b7658_372,RI2b5e785b5ee8_392,RI2b5e785b5588_412,RI2b5e785b4c28_432,RI2b5e785b3878_452,
        RI2b5e785b2f18_472,RI2b5e785b25b8_492,RI2b5e785b15c8_512,RI2b5e785b0c68_532,RI2b5e785b0308_552,RI2b5e785af6d8_572,RI2b5e785da158_251,RI2b5e785be660_271,RI2b5e785bc3b0_291,RI2b5e785bba50_311,
        RI2b5e785b9b60_331,RI2b5e785b8030_351,RI2b5e785b76d0_371,RI2b5e785b6d70_391,RI2b5e785b5600_411,RI2b5e785b4ca0_431,RI2b5e785b38f0_451,RI2b5e785b2f90_471,RI2b5e785b2630_491,RI2b5e785b1640_511,
        RI2b5e785b0ce0_531,RI2b5e785b0380_551,RI2b5e785af750_571,RI2b5e785da068_253,RI2b5e785be570_273,RI2b5e785bc2c0_293,RI2b5e785bb960_313,RI2b5e785b9a70_333,RI2b5e785b7f40_353,RI2b5e785b75e0_373,
        RI2b5e785b5e70_393,RI2b5e785b5510_413,RI2b5e785b4bb0_433,RI2b5e785b3800_453,RI2b5e785b2ea0_473,RI2b5e785b2540_493,RI2b5e785b1550_513,RI2b5e785b0bf0_533,RI2b5e785b0290_553,RI2b5e785af660_573,
        RI2b5e785c2bc0_255,RI2b5e785be480_275,RI2b5e785bc1d0_295,RI2b5e785ba2e0_315,RI2b5e785b9980_335,RI2b5e785b7e50_355,RI2b5e785b74f0_375,RI2b5e785b5d80_395,RI2b5e785b5420_415,RI2b5e785b4ac0_435,
        RI2b5e785b3710_455,RI2b5e785b2db0_475,RI2b5e785b2450_495,RI2b5e785b1460_515,RI2b5e785b0b00_535,RI2b5e785b01a0_555,RI2b5e785af570_575,RI2b5e785c2c38_254,RI2b5e785be4f8_274,RI2b5e785bc248_294,
        RI2b5e785ba358_314,RI2b5e785b99f8_334,RI2b5e785b7ec8_354,RI2b5e785b7568_374,RI2b5e785b5df8_394,RI2b5e785b5498_414,RI2b5e785b4b38_434,RI2b5e785b3788_454,RI2b5e785b2e28_474,RI2b5e785b24c8_494,
        RI2b5e785b14d8_514,RI2b5e785b0b78_534,RI2b5e785b0218_554,RI2b5e785af5e8_574,RI2b5e785c0a00_257,RI2b5e785be390_277,RI2b5e785bc0e0_297,RI2b5e785ba1f0_317,RI2b5e785b9890_337,RI2b5e785b7d60_357,
        RI2b5e785b7400_377,RI2b5e785b5c90_397,RI2b5e785b5330_417,RI2b5e785b49d0_437,RI2b5e785b3620_457,RI2b5e785b2cc0_477,RI2b5e785b2360_497,RI2b5e785b1370_517,RI2b5e785b0a10_537,RI2b5e785b00b0_557,
        RI2b5e785af480_577,RI2b5e785c2b48_256,RI2b5e785be408_276,RI2b5e785bc158_296,RI2b5e785ba268_316,RI2b5e785b9908_336,RI2b5e785b7dd8_356,RI2b5e785b7478_376,RI2b5e785b5d08_396,RI2b5e785b53a8_416,
        RI2b5e785b4a48_436,RI2b5e785b3698_456,RI2b5e785b2d38_476,RI2b5e785b23d8_496,RI2b5e785b13e8_516,RI2b5e785b0a88_536,RI2b5e785b0128_556,RI2b5e785af4f8_576,RI2b5e785c0910_259,RI2b5e785be2a0_279,
        RI2b5e785bbff0_299,RI2b5e785ba100_319,RI2b5e785b97a0_339,RI2b5e785b7c70_359,RI2b5e785b7310_379,RI2b5e785b5ba0_399,RI2b5e785b5240_419,RI2b5e785b48e0_439,RI2b5e785b3530_459,RI2b5e785b2bd0_479,
        RI2b5e785b2270_499,RI2b5e785b1280_519,RI2b5e785b0920_539,RI2b5e785affc0_559,RI2b5e785af390_579,RI2b5e785c0988_258,RI2b5e785be318_278,RI2b5e785bc068_298,RI2b5e785ba178_318,RI2b5e785b9818_338,
        RI2b5e785b7ce8_358,RI2b5e785b7388_378,RI2b5e785b5c18_398,RI2b5e785b52b8_418,RI2b5e785b4958_438,RI2b5e785b35a8_458,RI2b5e785b2c48_478,RI2b5e785b22e8_498,RI2b5e785b12f8_518,RI2b5e785b0998_538,
        RI2b5e785b0038_558,RI2b5e785af408_578,RI2b5e785c0820_261,RI2b5e785be1b0_281,RI2b5e785bbf00_301,RI2b5e785ba010_321,RI2b5e785b96b0_341,RI2b5e785b7b80_361,RI2b5e785b7220_381,RI2b5e785b5ab0_401,
        RI2b5e785b5150_421,RI2b5e785b47f0_441,RI2b5e785b3440_461,RI2b5e785b2ae0_481,RI2b5e785b2180_501,RI2b5e785b1190_521,RI2b5e785b0830_541,RI2b5e785afed0_561,RI2b5e785af2a0_581,RI2b5e785c0898_260,
        RI2b5e785be228_280,RI2b5e785bbf78_300,RI2b5e785ba088_320,RI2b5e785b9728_340,RI2b5e785b7bf8_360,RI2b5e785b7298_380,RI2b5e785b5b28_400,RI2b5e785b51c8_420,RI2b5e785b4868_440,RI2b5e785b34b8_460,
        RI2b5e785b2b58_480,RI2b5e785b21f8_500,RI2b5e785b1208_520,RI2b5e785b08a8_540,RI2b5e785aff48_560,RI2b5e785af318_580,RI2b5e785c0730_263,RI2b5e785be0c0_283,RI2b5e785bbe10_303,RI2b5e785b9f20_323,
        RI2b5e785b95c0_343,RI2b5e785b7a90_363,RI2b5e785b7130_383,RI2b5e785b59c0_403,RI2b5e785b5060_423,RI2b5e785b3cb0_443,RI2b5e785b3350_463,RI2b5e785b29f0_483,RI2b5e785b1a00_503,RI2b5e785b10a0_523,
        RI2b5e785b0740_543,RI2b5e785afde0_563,RI2b5e785af1b0_583,RI2b5e785c07a8_262,RI2b5e785be138_282,RI2b5e785bbe88_302,RI2b5e785b9f98_322,RI2b5e785b9638_342,RI2b5e785b7b08_362,RI2b5e785b71a8_382,
        RI2b5e785b5a38_402,RI2b5e785b50d8_422,RI2b5e785b4778_442,RI2b5e785b33c8_462,RI2b5e785b2a68_482,RI2b5e785b1a78_502,RI2b5e785b1118_522,RI2b5e785b07b8_542,RI2b5e785afe58_562,RI2b5e785af228_582,
        RI2b5e785c0640_265,RI2b5e785bdfd0_285,RI2b5e785bbd20_305,RI2b5e785b9e30_325,RI2b5e785b94d0_345,RI2b5e785b79a0_365,RI2b5e785b7040_385,RI2b5e785b58d0_405,RI2b5e785b4f70_425,RI2b5e785b3bc0_445,
        RI2b5e785b3260_465,RI2b5e785b2900_485,RI2b5e785b1910_505,RI2b5e785b0fb0_525,RI2b5e785b0650_545,RI2b5e785afcf0_565,RI2b5e785af0c0_585,RI2b5e785c06b8_264,RI2b5e785be048_284,RI2b5e785bbd98_304,
        RI2b5e785b9ea8_324,RI2b5e785b9548_344,RI2b5e785b7a18_364,RI2b5e785b70b8_384,RI2b5e785b5948_404,RI2b5e785b4fe8_424,RI2b5e785b3c38_444,RI2b5e785b32d8_464,RI2b5e785b2978_484,RI2b5e785b1988_504,
        RI2b5e785b1028_524,RI2b5e785b06c8_544,RI2b5e785afd68_564,RI2b5e785af138_584,RI2b5e785c05c8_266,RI2b5e785bdf58_286,RI2b5e785bbca8_306,RI2b5e785b9db8_326,RI2b5e785b9458_346,RI2b5e785b7928_366,
        RI2b5e785b6fc8_386,RI2b5e785b5858_406,RI2b5e785b4ef8_426,RI2b5e785b3b48_446,RI2b5e785b31e8_466,RI2b5e785b2888_486,RI2b5e785b1898_506,RI2b5e785b0f38_526,RI2b5e785b05d8_546,RI2b5e785afc78_566,
        RI2b5e785af048_586,RI2b5e785c0550_267,RI2b5e785bc590_287,RI2b5e785bbc30_307,RI2b5e785b9d40_327,RI2b5e785b93e0_347,RI2b5e785b78b0_367,RI2b5e785b6f50_387,RI2b5e785b57e0_407,RI2b5e785b4e80_427,
        RI2b5e785b3ad0_447,RI2b5e785b3170_467,RI2b5e785b2810_487,RI2b5e785b1820_507,RI2b5e785b0ec0_527,RI2b5e785b0560_547,RI2b5e785afc00_567,RI2b5e785aefd0_587,RI2b5e785ae328_614,RI2b5e785db058_15,
        RI2b5e785dafe0_16,RI2b5e785daf68_17,RI2b5e785daef0_18,RI2b5e785dae78_19,RI2b5e785dae00_20,RI2b5e785dad88_21,RI2b5e785dad10_22,RI2b5e785dac98_23,RI2b5e785dac20_24,RI2b5e785daba8_25,
        RI2b5e785ae3a0_613,RI2b5e785ae418_612,RI2b5e785ae490_611,RI2b5e785ae508_610,RI2b5e785ae580_609,RI2b5e785dab30_26,RI2b5e785ae5f8_608,RI2b5e785ae670_607,RI2b5e785ae6e8_606,RI2b5e785ae760_605,
        RI2b5e785ae7d8_604,RI2b5e785ae850_603,RI2b5e785ae8c8_602,RI2b5e785ae940_601,RI2b5e785db0d0_14;
output R_267_b04ddc8,R_268_b04de70,R_269_b04df18,R_26a_b04dfc0,R_26b_b04e068,R_26c_b04e110,R_26d_b04e1b8,R_26e_b04e260,R_26f_b04e308,
        R_270_b04e3b0,R_271_b04e458,R_272_b04e500,R_273_b04e5a8,R_274_b04e650,R_275_b04e6f8,R_276_b04e7a0,R_277_b04e848,R_278_b04e8f0,R_279_b04e998,
        R_27a_b04ea40,R_27b_b04eae8,R_27c_b04eb90,R_27d_b04ec38,R_27e_b04ece0,R_27f_b04ed88,R_280_b04ee30,R_281_b04eed8,R_282_b04ef80,R_283_b04f028,
        R_284_b04f0d0,R_285_b04f178,R_286_b04f220,R_287_b04f2c8,R_288_b04f370,R_289_b04f418,R_28a_b04f4c0,R_28b_b04f568,R_28c_b04f610,R_28d_b04f6b8,
        R_28e_b04f760,R_28f_b04f808,R_290_b04f8b0,R_291_b04f958,R_292_b04fa00,R_293_b04faa8,R_294_b04fb50,R_295_b04fbf8,R_296_b04fca0,R_297_b04fd48,
        R_298_b04fdf0,R_299_b04fe98,R_29a_b04ff40,R_29b_b04ffe8,R_29c_b050090,R_29d_b050138,R_29e_b0501e0,R_29f_b050288,R_2a0_b050330,R_2a1_b0503d8,
        R_2a2_b050480,R_2a3_b050528,R_2a4_b0505d0,R_2a5_b050678,R_2a6_b050720,R_2a7_b0507c8,R_2a8_b050870,R_2a9_b050918,R_2aa_b0509c0;

wire \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 ,
         \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 ,
         \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 ,
         \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 ,
         \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 ,
         \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 ,
         \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 ,
         \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 ,
         \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 ,
         \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 ,
         \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 ,
         \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 ,
         \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 ,
         \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 ,
         \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 ,
         \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 ,
         \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 ,
         \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 ,
         \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 ,
         \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 ,
         \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 ,
         \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 ,
         \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 ,
         \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 ,
         \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 ,
         \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 ,
         \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 ,
         \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 ,
         \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 ,
         \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 ,
         \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 ,
         \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 ,
         \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 ,
         \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 ,
         \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 ,
         \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 ,
         \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 ,
         \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 ,
         \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 ,
         \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 ,
         \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 ,
         \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 ,
         \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 ,
         \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 ,
         \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 ,
         \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 ,
         \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 ,
         \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 ,
         \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 ,
         \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 ,
         \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 ,
         \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 ,
         \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 ,
         \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 ,
         \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 ,
         \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 ,
         \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 ,
         \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 ,
         \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 ,
         \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 ,
         \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 ,
         \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 ,
         \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 ,
         \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 ,
         \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 ,
         \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
         \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 ,
         \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 ,
         \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 ,
         \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 ,
         \1382 , \1383 , \1384 , \1385 , \1386 , \1387_N$1 , \1388_N$2 , \1389_N$3 , \1390_N$4 , \1391_N$5 ,
         \1392_N$6 , \1393_N$7 , \1394_N$8 , \1395_N$9 , \1396_N$10 , \1397_N$11 , \1398_N$12 , \1399_N$13 , \1400_N$14 , \1401_N$15 ,
         \1402_N$16 , \1403_N$17 , \1404_N$18 , \1405_N$20 , \1406_N$21 , \1407_N$22 , \1408_N$23 , \1409_N$24 , \1410_N$25 , \1411_N$26 ,
         \1412_N$27 , \1413_N$28 , \1414_N$29 , \1415_N$30 , \1416_N$31 , \1417_N$32 , \1418_N$33 , \1419_N$34 , \1420_N$35 , \1421_N$36 ,
         \1422_N$37 , \1423_N$38 , \1424_N$39 , \1425_N$40 , \1426_N$41 , \1427_N$42 , \1428_N$43 , \1429_N$45 , \1430_N$46 , \1431_N$47 ,
         \1432_N$48 , \1433_N$49 , \1434_N$50 , \1435_N$51 , \1436_N$52 , \1437_N$53 , \1438_N$54 , \1439_N$55 , \1440_N$56 , \1441_N$57 ,
         \1442_N$58 , \1443_N$59 , \1444_N$60 , \1445_N$61 , \1446_N$62 , \1447_N$63 , \1448_N$64 , \1449_N$65 , \1450_N$66 , \1451_N$67 ,
         \1452_N$68 , \1453_N$69 , \1454_N$70 , \1455_N$71 , \1456_N$72 , \1457_N$73 , \1458_N$74 , \1459_N$75 , \1460_N$76 , \1461_N$77 ,
         \1462_N$78 , \1463_N$79 , \1464_N$80 , \1465_N$81 , \1466_N$82 , \1467_N$83 , \1468_N$85 , \1469_N$86 , \1470_N$87 , \1471_N$88 ,
         \1472_N$90 , \1473_N$91 , \1474_N$92 , \1475_N$93 , \1476_N$94 , \1477_N$95 , \1478_N$96 , \1479_N$98 , \1480_N$99 , \1481_N$100 ,
         \1482_N$101 , \1483_N$102 , \1484_N$103 , \1485_N$104 , \1486_N$105 , \1487_N$106 , \1488_N$107 , \1489_N$108 , \1490_N$109 , \1491_N$110 ,
         \1492_N$111 , \1493_N$112 , \1494_N$113 , \1495_N$114 , \1496_N$115 , \1497_N$116 , \1498_N$117 , \1499_N$118 , \1500_N$119 , \1501_N$120 ,
         \1502_N$121 , \1503_N$122 , \1504_N$123 , \1505_N$124 , \1506_N$125 , \1507_N$126 , \1508_N$127 , \1509_N$128 , \1510_N$129 , \1511_N$130 ,
         \1512_N$131 , \1513_N$132 , \1514_N$133 , \1515_N$134 , \1516_N$135 , \1517_N$137 , \1518_N$138 , \1519_N$139 , \1520_N$140 , \1521_N$141 ,
         \1522_N$142 , \1523_N$143 , \1524_N$144 , \1525_N$145 , \1526_N$146 , \1527_N$147 , \1528_N$148 , \1529_N$149 , \1530_N$150 , \1531_N$151 ,
         \1532_N$152 , \1533_N$153 , \1534_N$154 , \1535_N$155 , \1536_N$156 , \1537_N$157 , \1538_N$158 , \1539_N$159 , \1540_N$160 , \1541_N$161 ,
         \1542_N$162 , \1543_N$163 , \1544_N$164 , \1545_N$165 , \1546_N$166 , \1547_N$167 , \1548_N$168 , \1549_N$169 , \1550_N$171 , \1551_N$172 ,
         \1552_N$173 , \1553_N$174 , \1554_N$175 , \1555_N$176 , \1556_N$177 , \1557_N$178 , \1558_N$179 , \1559_N$180 , \1560_N$181 , \1561_N$182 ,
         \1562_N$183 , \1563_N$184 , \1564_N$185 , \1565_N$186 , \1566_N$187 , \1567_N$188 , \1568_N$189 , \1569_N$190 , \1570_N$191 , \1571_N$192 ,
         \1572_N$193 , \1573_N$194 , \1574_N$195 , \1575_N$196 , \1576_N$197 , \1577_N$198 , \1578_N$199 , \1579_N$200 , \1580_N$201 , \1581_N$203 ,
         \1582_N$204 , \1583_N$205 , \1584_N$206 , \1585_N$207 , \1586_N$208 , \1587_N$209 , \1588_N$210 , \1589_N$211 , \1590_N$212 , \1591_N$213 ,
         \1592_N$214 , \1593_N$215 , \1594_N$216 , \1595_N$217 , \1596_N$218 , \1597_N$219 , \1598_N$220 , \1599_N$221 , \1600_N$222 , \1601_N$223 ,
         \1602_N$224 , \1603_N$225 , \1604_N$226 , \1605_N$228 , \1606_N$229 , \1607_N$230 , \1608_N$231 , \1609_N$232 , \1610_N$233 , \1611_N$234 ,
         \1612_N$235 , \1613_N$236 , \1614_N$237 , \1615_N$238 , \1616_N$239 , \1617_N$240 , \1618_N$241 , \1619_N$242 , \1620_N$243 , \1621_N$244 ,
         \1622_N$245 , \1623_N$246 , \1624_N$247 , \1625_N$248 , \1626_N$249 , \1627_N$250 , \1628_N$251 , \1629_N$252 , \1630_N$253 , \1631_N$254 ,
         \1632_N$255 , \1633_N$256 , \1634_N$257 , \1635_N$258 , \1636_N$259 , \1637_N$260 , \1638_N$261 , \1639_N$262 , \1640_N$263 , \1641_N$264 ,
         \1642_N$265 , \1643_N$266 , \1644_N$268 , \1645_N$269 , \1646_N$270 , \1647_N$271 , \1648_N$273 , \1649_N$274 , \1650_N$275 , \1651_N$276 ,
         \1652_N$277 , \1653_N$278 , \1654_N$279 , \1655_N$281 , \1656_N$282 , \1657_N$283 , \1658_N$284 , \1659_N$285 , \1660_N$286 , \1661_N$287 ,
         \1662_N$288 , \1663_N$289 , \1664_N$290 , \1665_N$291 , \1666_N$292 , \1667_N$293 , \1668_N$294 , \1669_N$295 , \1670_N$296 , \1671_N$297 ,
         \1672_N$298 , \1673_N$299 , \1674_N$300 , \1675_N$301 , \1676_N$302 , \1677_N$303 , \1678_N$304 , \1679_N$305 , \1680_N$306 , \1681_N$307 ,
         \1682_N$308 , \1683_N$309 , \1684_N$310 , \1685_N$311 , \1686_N$312 , \1687_N$313 , \1688_N$314 , \1689_N$315 , \1690_N$316 , \1691_N$317 ,
         \1692_N$318 , \1693_N$320 , \1694_N$321 , \1695_N$322 , \1696_N$323 , \1697_N$324 , \1698_N$325 , \1699_N$326 , \1700_N$327 , \1701_N$328 ,
         \1702_N$329 , \1703_N$330 , \1704_N$331 , \1705_N$332 , \1706_N$333 , \1707_N$334 , \1708_N$335 , \1709_N$336 , \1710_N$337 , \1711_N$338 ,
         \1712_N$339 , \1713_N$340 , \1714_N$341 , \1715_N$342 , \1716_N$343 , \1717_N$344 , \1718_N$345 , \1719_N$346 , \1720_N$347 , \1721_N$348 ,
         \1722_N$349 , \1723_N$350 , \1724_N$351 , \1725_N$352 , \1726_N$354 , \1727_N$355 , \1728_N$356 , \1729_N$357 , \1730_N$358 , \1731_N$359 ,
         \1732_N$360 , \1733_N$361 , \1734_N$362 , \1735_N$363 , \1736_N$364 , \1737_N$365 , \1738_N$366 , \1739_N$367 , \1740_N$368 , \1741_N$369 ,
         \1742_N$370 , \1743_N$371 , \1744_N$372 , \1745_N$373 , \1746_N$374 , \1747_N$375 , \1748_N$376 , \1749_N$377 , \1750_N$378 , \1751_N$379 ,
         \1752_N$380 , \1753_N$381 , \1754_N$382 , \1755_N$383 , \1756_N$384 , \1757_N$386 , \1758_N$387 , \1759_N$388 , \1760_N$389 , \1761_N$390 ,
         \1762_N$391 , \1763_N$392 , \1764_N$393 , \1765_N$394 , \1766_N$395 , \1767_N$396 , \1768_N$397 , \1769_N$398 , \1770_N$399 , \1771_N$400 ,
         \1772_N$401 , \1773_N$402 , \1774_N$403 , \1775_N$404 , \1776_N$405 , \1777_N$406 , \1778_N$407 , \1779_N$408 , \1780_N$409 , \1781_N$411 ,
         \1782_N$412 , \1783_N$413 , \1784_N$414 , \1785_N$415 , \1786_N$416 , \1787_N$417 , \1788_N$418 , \1789_N$419 , \1790_N$420 , \1791_N$421 ,
         \1792_N$422 , \1793_N$423 , \1794_N$424 , \1795_N$425 , \1796_N$426 , \1797_N$427 , \1798_N$428 , \1799_N$429 , \1800_N$430 , \1801_N$431 ,
         \1802_N$432 , \1803_N$433 , \1804_N$434 , \1805_N$435 , \1806_N$436 , \1807_N$437 , \1808_N$438 , \1809_N$439 , \1810_N$440 , \1811_N$441 ,
         \1812_N$442 , \1813_N$443 , \1814_N$444 , \1815_N$445 , \1816_N$446 , \1817_N$447 , \1818_N$448 , \1819_N$449 , \1820_N$451 , \1821_N$452 ,
         \1822_N$453 , \1823_N$454 , \1824_N$456 , \1825_N$457 , \1826_N$458 , \1827_N$459 , \1828_N$460 , \1829_N$461 , \1830_N$462 , \1831_N$464 ,
         \1832_N$465 , \1833_N$466 , \1834_N$467 , \1835_N$468 , \1836_N$469 , \1837_N$470 , \1838_N$471 , \1839_N$472 , \1840_N$473 , \1841_N$474 ,
         \1842_N$475 , \1843_N$476 , \1844_N$477 , \1845_N$478 , \1846_N$479 , \1847_N$480 , \1848_N$481 , \1849_N$482 , \1850_N$483 , \1851_N$484 ,
         \1852_N$485 , \1853_N$486 , \1854_N$487 , \1855_N$488 , \1856_N$489 , \1857_N$490 , \1858_N$491 , \1859_N$492 , \1860_N$493 , \1861_N$494 ,
         \1862_N$495 , \1863_N$496 , \1864_N$497 , \1865_N$498 , \1866_N$499 , \1867_N$500 , \1868_N$501 , \1869_N$503 , \1870_N$504 , \1871_N$505 ,
         \1872_N$506 , \1873_N$507 , \1874_N$508 , \1875_N$509 , \1876_N$510 , \1877_N$511 , \1878_N$512 , \1879_N$513 , \1880_N$514 , \1881_N$515 ,
         \1882_N$516 , \1883_N$517 , \1884_N$518 , \1885_N$519 , \1886_N$520 , \1887_N$521 , \1888_N$522 , \1889_N$523 , \1890_N$524 , \1891_N$525 ,
         \1892_N$526 , \1893_N$527 , \1894_N$528 , \1895_N$529 , \1896_N$530 , \1897_N$531 , \1898_N$532 , \1899_N$533 , \1900_N$534 , \1901_N$535 ,
         \1902_N$537 , \1903_N$538 , \1904_N$539 , \1905_N$540 , \1906_N$541 , \1907_N$542 , \1908_N$543 , \1909_N$544 , \1910_N$545 , \1911_N$546 ,
         \1912_N$547 , \1913_N$548 , \1914_N$549 , \1915_N$550 , \1916_N$551 , \1917_N$552 , \1918_N$553 , \1919_N$554 , \1920_N$555 , \1921_N$556 ,
         \1922_N$557 , \1923_N$558 , \1924_N$559 , \1925_N$560 , \1926_N$561 , \1927_N$562 , \1928_N$563 , \1929_N$564 , \1930_N$565 , \1931_N$566 ,
         \1932_N$567 , \1933_N$569 , \1934_N$570 , \1935_N$571 , \1936_N$572 , \1937_N$573 , \1938_N$574 , \1939_N$575 , \1940_N$576 , \1941_N$577 ,
         \1942_N$578 , \1943_N$579 , \1944_N$580 , \1945_N$581 , \1946_N$582 , \1947_N$583 , \1948_N$584 , \1949_N$585 , \1950_N$586 , \1951_N$587 ,
         \1952_N$588 , \1953_N$589 , \1954_N$590 , \1955_N$591 , \1956_N$592 , \1957_N$594 , \1958_N$595 , \1959_N$596 , \1960_N$597 , \1961_N$598 ,
         \1962_N$599 , \1963_N$600 , \1964_N$601 , \1965_N$602 , \1966_N$603 , \1967_N$604 , \1968_N$605 , \1969_N$606 , \1970_N$607 , \1971_N$608 ,
         \1972_N$609 , \1973_N$610 , \1974_N$611 , \1975_N$612 , \1976_N$613 , \1977_N$614 , \1978_N$615 , \1979_N$616 , \1980_N$617 , \1981_N$618 ,
         \1982_N$619 , \1983_N$620 , \1984_N$621 , \1985_N$622 , \1986_N$623 , \1987_N$624 , \1988_N$625 , \1989_N$626 , \1990_N$627 , \1991_N$628 ,
         \1992_N$629 , \1993_N$630 , \1994_N$631 , \1995_N$632 , \1996_N$634 , \1997_N$635 , \1998_N$636 , \1999_N$637 , \2000_N$639 , \2001_N$640 ,
         \2002_N$641 , \2003_N$642 , \2004_N$643 , \2005_N$644 , \2006_N$645 , \2007_N$647 , \2008_N$648 , \2009_N$649 , \2010_N$650 , \2011_N$651 ,
         \2012_N$652 , \2013_N$653 , \2014_N$654 , \2015_N$655 , \2016_N$656 , \2017_N$657 , \2018_N$658 , \2019_N$659 , \2020_N$660 , \2021_N$661 ,
         \2022_N$662 , \2023_N$663 , \2024_N$664 , \2025_N$665 , \2026_N$666 , \2027_N$667 , \2028_N$668 , \2029_N$669 , \2030_N$670 , \2031_N$671 ,
         \2032_N$672 , \2033_N$673 , \2034_N$674 , \2035_N$675 , \2036_N$676 , \2037_N$677 , \2038_N$678 , \2039_N$679 , \2040_N$680 , \2041_N$681 ,
         \2042_N$682 , \2043_N$683 , \2044_N$684 , \2045_N$686 , \2046_N$687 , \2047_N$688 , \2048_N$689 , \2049_N$690 , \2050_N$691 , \2051_N$692 ,
         \2052_N$693 , \2053_N$694 , \2054_N$695 , \2055_N$696 , \2056_N$697 , \2057_N$698 , \2058_N$699 , \2059_N$700 , \2060_N$701 , \2061_N$702 ,
         \2062_N$703 , \2063_N$704 , \2064_N$705 , \2065_N$706 , \2066_N$707 , \2067_N$708 , \2068_N$709 , \2069_N$710 , \2070_N$711 , \2071_N$712 ,
         \2072_N$713 , \2073_N$714 , \2074_N$715 , \2075_N$716 , \2076_N$717 , \2077_N$718 , \2078_N$720 , \2079_N$721 , \2080_N$722 , \2081_N$723 ,
         \2082_N$724 , \2083_N$725 , \2084_N$726 , \2085_N$727 , \2086_N$728 , \2087_N$729 , \2088_N$730 , \2089_N$731 , \2090_N$732 , \2091_ZERO ,
         \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 ,
         \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 ,
         \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120_N$19 , \2121_N$44 ,
         \2122_N$84 , \2123_N$89 , \2124_N$97 , \2125_N$136 , \2126_N$170 , \2127_N$202 , \2128_N$227 , \2129_N$267 , \2130_N$272 , \2131_N$280 ,
         \2132_N$319 , \2133_N$353 , \2134_N$385 , \2135_N$410 , \2136_N$450 , \2137_N$455 , \2138_N$463 , \2139_N$502 , \2140_N$536 , \2141_N$568 ,
         \2142_N$593 , \2143_N$633 , \2144_N$638 , \2145_N$646 , \2146_N$685 , \2147_N$719 , \2148_ONE , \2149 , \2150 , \2151 ,
         \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 ,
         \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 ,
         \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 ,
         \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 ,
         \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 ,
         \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 ,
         \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219_nR2049 , \2220 , \2221 ,
         \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 ,
         \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 ,
         \2242 , \2243 , \2244_nR2025 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 ,
         \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 ,
         \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269_nR1e9e , \2270 , \2271 ,
         \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 ,
         \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 ,
         \2292 , \2293 , \2294_nR1e7a , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 ,
         \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 ,
         \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319_nR1d05 , \2320 , \2321 ,
         \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 ,
         \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 ,
         \2342 , \2343 , \2344_nR1ce1 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 ,
         \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 ,
         \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369_nR1ba3 , \2370 , \2371 ,
         \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 ,
         \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 ,
         \2392 , \2393 , \2394_nR1b7f , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 ,
         \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 ,
         \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419_nR1a72 , \2420 , \2421 ,
         \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 ,
         \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 ,
         \2442 , \2443 , \2444_nR1a8b , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 ,
         \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 ,
         \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469_nR1968 , \2470 , \2471 ,
         \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 ,
         \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 ,
         \2492 , \2493_nR194c , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 ,
         \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 ,
         \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 ,
         \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 ,
         \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 ,
         \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 ,
         \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 ,
         \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 ,
         \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 ,
         \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 ,
         \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 ,
         \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 ,
         \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620_nR2749 , \2621 ,
         \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 ,
         \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 ,
         \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648_nR2211 , \2649 , \2650 , \2651 ,
         \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 ,
         \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 ,
         \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 ,
         \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689_nR283d , \2690 , \2691 ,
         \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 ,
         \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 ,
         \2712 , \2713 , \2714 , \2715 , \2716_nR2687 , \2717 , \2718 , \2719 , \2720 , \2721 ,
         \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 ,
         \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 ,
         \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 ,
         \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 ,
         \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 ,
         \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 ,
         \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 ,
         \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 ,
         \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 ,
         \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 ,
         \2822 , \2823 , \2824 , \2825 , \2826 , \2827_nR24ec , \2828 , \2829 , \2830 , \2831 ,
         \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 ,
         \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848_nR25c6 , \2849 , \2850 , \2851 ,
         \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 ,
         \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871_nR2401 ,
         \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 ,
         \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 ,
         \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 ,
         \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 ,
         \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 ,
         \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 ,
         \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 ,
         \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 ,
         \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 ,
         \2962 , \2963 , \2964_nR224e , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 ,
         \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 ,
         \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 ,
         \2992 , \2993 , \2994 , \2995 , \2996 , \2997_nR2322 , \2998 , \2999 , \3000 , \3001 ,
         \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 ,
         \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 ,
         \3022 , \3023 , \3024_nR2081 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 ,
         \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 ,
         \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 ,
         \3052 , \3053 , \3054 , \3055 , \3056 , \3057_nR2158 , \3058 , \3059 , \3060 , \3061 ,
         \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 ,
         \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 ,
         \3082 , \3083 , \3084 , \3085 , \3086_nR1ec2 , \3087 , \3088 , \3089 , \3090 , \3091 ,
         \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 ,
         \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 ,
         \3112 , \3113 , \3114 , \3115_nR1f8b , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 ,
         \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 ,
         \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141_nR1d29 ,
         \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 ,
         \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 ,
         \3162_nR1ddc , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 ,
         \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 ,
         \3182 , \3183 , \3184 , \3185 , \3186_nR1bc5 , \3187 , \3188 , \3189 , \3190 , \3191 ,
         \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 ,
         \3202 , \3203 , \3204 , \3205 , \3206 , \3207_nR1c6c , \3208 , \3209 , \3210 , \3211 ,
         \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 ,
         \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 ,
         \3232 , \3233 , \3234_nR1a55 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 ,
         \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 ,
         \3252 , \3253 , \3254 , \3255_nR1b26 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 ,
         \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 ,
         \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278_nR1a13 , \3279 , \3280 , \3281 ,
         \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 ,
         \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 ,
         \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 ,
         \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 ,
         \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 ,
         \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 ,
         \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 ,
         \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 ,
         \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 ,
         \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 ,
         \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 ,
         \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 ,
         \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411_nR191b ,
         \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 ,
         \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 ,
         \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 ,
         \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 ,
         \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 ,
         \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 ,
         \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 ,
         \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 ,
         \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 ,
         \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 ,
         \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 ,
         \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 ,
         \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 ,
         \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 ,
         \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 ,
         \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 ,
         \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 ,
         \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 ,
         \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 ,
         \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 ,
         \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 ,
         \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 ,
         \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 ,
         \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 ,
         \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 ,
         \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 ,
         \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 ,
         \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 ,
         \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 ,
         \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 ,
         \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 ,
         \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 ,
         \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 ,
         \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 ,
         \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 ,
         \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 ,
         \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 ,
         \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 ,
         \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 ,
         \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 ,
         \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 ,
         \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 ,
         \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 ,
         \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 ,
         \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 ,
         \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 ,
         \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 ,
         \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 ,
         \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 ,
         \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 ,
         \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 ,
         \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 ,
         \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 ,
         \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 ,
         \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 ,
         \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 ,
         \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 ,
         \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 ,
         \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 ,
         \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 ,
         \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 ,
         \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 ,
         \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 ,
         \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 ,
         \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 ,
         \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 ,
         \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 ,
         \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 ,
         \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 ,
         \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 ,
         \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 ,
         \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 ,
         \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 ,
         \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 ,
         \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 ,
         \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 ,
         \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 ,
         \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 ,
         \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 ,
         \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 ,
         \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 ,
         \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 ,
         \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 ,
         \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 ,
         \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 ,
         \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 ,
         \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 ,
         \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 ,
         \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 ,
         \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 ,
         \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 ,
         \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 ,
         \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 ,
         \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 ,
         \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 ,
         \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 ,
         \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 ,
         \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 ,
         \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 ,
         \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 ,
         \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 ,
         \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 ,
         \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 ,
         \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 ,
         \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 ,
         \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 ,
         \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 ,
         \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 ,
         \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 ,
         \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 ,
         \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 ,
         \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 ,
         \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 ,
         \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 ,
         \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 ,
         \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 ,
         \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 ,
         \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 ,
         \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 ,
         \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 ,
         \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 ,
         \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 ,
         \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 ,
         \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 ,
         \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 ,
         \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 ,
         \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 ,
         \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 ,
         \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 ,
         \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 ,
         \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 ,
         \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 ,
         \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 ,
         \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 ,
         \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 ,
         \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 ,
         \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 ,
         \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 ,
         \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 ,
         \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 ,
         \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 ,
         \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 ,
         \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 ,
         \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 ,
         \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 ,
         \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 ,
         \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 ,
         \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 ,
         \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 ,
         \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 ,
         \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 ,
         \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 ,
         \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 ,
         \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 ,
         \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 ,
         \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 ,
         \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981_nR20e2 ,
         \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 ,
         \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 ,
         \5002 , \5003 , \5004 , \5005 , \5006_nR20be , \5007 , \5008 , \5009 , \5010 , \5011 ,
         \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 ,
         \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031_nR1f2b ,
         \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 ,
         \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 ,
         \5052 , \5053 , \5054 , \5055 , \5056_nR1f07 , \5057 , \5058 , \5059 , \5060 , \5061 ,
         \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 ,
         \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081_nR1d88 ,
         \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 ,
         \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 ,
         \5102 , \5103 , \5104 , \5105 , \5106_nR1d64 , \5107 , \5108 , \5109 , \5110 , \5111 ,
         \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 ,
         \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131_nR1c19 ,
         \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 ,
         \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 ,
         \5152 , \5153 , \5154 , \5155 , \5156_nR1bf5 , \5157 , \5158 , \5159 , \5160 , \5161 ,
         \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 ,
         \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181_nR1ada ,
         \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 ,
         \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 ,
         \5202 , \5203 , \5204 , \5205 , \5206_nR1af3 , \5207 , \5208 , \5209 , \5210 , \5211 ,
         \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 ,
         \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231_nR19f0 ,
         \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 ,
         \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 ,
         \5252 , \5253 , \5254 , \5255_nR19d4 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 ,
         \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 ,
         \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 ,
         \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 ,
         \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 ,
         \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 ,
         \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 ,
         \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 ,
         \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 ,
         \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 ,
         \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 ,
         \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 ,
         \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 ,
         \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 ,
         \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 ,
         \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 ,
         \5412 , \5413 , \5414_nR27bc , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 ,
         \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 ,
         \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 ,
         \5442_nR229d , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 ,
         \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 ,
         \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 ,
         \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 ,
         \5482 , \5483_nR28b1 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 ,
         \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 ,
         \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510_nR26f3 , \5511 ,
         \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 ,
         \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 ,
         \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 ,
         \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 ,
         \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 ,
         \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 ,
         \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 ,
         \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 ,
         \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 ,
         \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 ,
         \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621_nR2554 ,
         \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 ,
         \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 ,
         \5642_nR2632 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 ,
         \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 ,
         \5662 , \5663 , \5664 , \5665_nR246b , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 ,
         \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 ,
         \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 ,
         \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 ,
         \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 ,
         \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 ,
         \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 ,
         \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 ,
         \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 ,
         \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758_nR22da , \5759 , \5760 , \5761 ,
         \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 ,
         \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 ,
         \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791_nR2387 ,
         \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 ,
         \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 ,
         \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818_nR211a , \5819 , \5820 , \5821 ,
         \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 ,
         \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 ,
         \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851_nR21b2 ,
         \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 ,
         \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 ,
         \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880_nR1f4f , \5881 ,
         \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 ,
         \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 ,
         \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909_nR1fd9 , \5910 , \5911 ,
         \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 ,
         \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 ,
         \5932 , \5933 , \5934 , \5935_nR1dac , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 ,
         \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 ,
         \5952 , \5953 , \5954 , \5955 , \5956_nR1e20 , \5957 , \5958 , \5959 , \5960 , \5961 ,
         \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 ,
         \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980_nR1c3b , \5981 ,
         \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 ,
         \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001_nR1ca2 ,
         \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 ,
         \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 ,
         \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028_nR1abd , \6029 , \6030 , \6031 ,
         \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 ,
         \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049_nR1b50 , \6050 , \6051 ,
         \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 ,
         \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 ,
         \6072_nR1a35 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 ,
         \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 ,
         \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 ,
         \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 ,
         \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 ,
         \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 ,
         \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 ,
         \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 ,
         \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 ,
         \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 ,
         \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 ,
         \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 ,
         \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 ,
         \6202 , \6203 , \6204 , \6205_nR19a3 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 ,
         \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 ,
         \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 ,
         \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 ,
         \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 ,
         \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 ,
         \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 ,
         \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 ,
         \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 ,
         \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 ,
         \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 ,
         \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 ,
         \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 ,
         \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 ,
         \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 ,
         \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 ,
         \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 ,
         \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 ,
         \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 ,
         \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 ,
         \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 ,
         \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 ,
         \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 ,
         \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 ,
         \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 ,
         \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 ,
         \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 ,
         \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 ,
         \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 ,
         \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 ,
         \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 ,
         \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 ,
         \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 ,
         \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 ,
         \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 ,
         \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 ,
         \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 ,
         \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 ,
         \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 ,
         \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 ,
         \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 ,
         \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 ,
         \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 ,
         \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 ,
         \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 ,
         \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 ,
         \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 ,
         \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 ,
         \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 ,
         \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 ,
         \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 ,
         \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 ,
         \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 ,
         \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 ,
         \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 ,
         \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 ,
         \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 ,
         \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 ,
         \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 ,
         \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 ,
         \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 ,
         \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 ,
         \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 ,
         \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 ,
         \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 ,
         \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 ,
         \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 ,
         \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 ,
         \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 ,
         \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 ,
         \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 ,
         \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 ,
         \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 ,
         \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 ,
         \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 ,
         \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 ,
         \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 ,
         \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 ,
         \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 ,
         \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 ,
         \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 ,
         \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 ,
         \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 ,
         \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 ,
         \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 ,
         \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 ,
         \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 ,
         \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 ,
         \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 ,
         \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 ,
         \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 ,
         \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 ,
         \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 ,
         \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 ,
         \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 ,
         \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 ,
         \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 ,
         \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 ,
         \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 ,
         \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 ,
         \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 ,
         \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 ,
         \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 ,
         \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 ,
         \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 ,
         \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 ,
         \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 ,
         \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 ,
         \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 ,
         \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 ,
         \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 ,
         \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 ,
         \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 ,
         \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 ,
         \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 ,
         \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 ,
         \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 ,
         \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 ,
         \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 ,
         \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 ,
         \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 ,
         \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 ,
         \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 ,
         \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 ,
         \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 ,
         \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 ,
         \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 ,
         \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 ,
         \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 ,
         \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 ,
         \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 ,
         \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
         \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 ,
         \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 ,
         \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 ,
         \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 ,
         \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 ,
         \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 ,
         \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 ,
         \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 ,
         \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 ,
         \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 ,
         \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 ,
         \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 ,
         \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 ,
         \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 ,
         \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 ,
         \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 ,
         \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 ,
         \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 ,
         \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 ,
         \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 ,
         \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 ,
         \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741_nRfe6 ,
         \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 ,
         \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 ,
         \7762 , \7763 , \7764 , \7765 , \7766_nRfff , \7767 , \7768 , \7769 , \7770 , \7771 ,
         \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 ,
         \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791_nR1018 ,
         \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 ,
         \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 ,
         \7812 , \7813 , \7814 , \7815 , \7816_nR1031 , \7817 , \7818 , \7819 , \7820 , \7821 ,
         \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 ,
         \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841_nR104a ,
         \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 ,
         \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 ,
         \7862 , \7863 , \7864 , \7865 , \7866_nR1063 , \7867 , \7868 , \7869 , \7870 , \7871 ,
         \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 ,
         \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891_nR107c ,
         \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 ,
         \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 ,
         \7912 , \7913 , \7914 , \7915 , \7916_nR1095 , \7917 , \7918 , \7919 , \7920 , \7921 ,
         \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 ,
         \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941_nR10ae ,
         \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 ,
         \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 ,
         \7962 , \7963 , \7964 , \7965 , \7966_nR10c7 , \7967 , \7968 , \7969 , \7970 , \7971 ,
         \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 ,
         \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991_nR10e0 ,
         \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 ,
         \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 ,
         \8012 , \8013 , \8014 , \8015 , \8016_nR10f9 , \8017 , \8018 , \8019 , \8020 , \8021 ,
         \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 ,
         \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040_nR1113 , \8041 ,
         \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 ,
         \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 ,
         \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 ,
         \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 ,
         \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 ,
         \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 ,
         \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 ,
         \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 ,
         \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 ,
         \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141_nR117c ,
         \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 ,
         \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 ,
         \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 ,
         \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 ,
         \8182 , \8183 , \8184 , \8185 , \8186 , \8187_nR11aa , \8188 , \8189 , \8190 , \8191 ,
         \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 ,
         \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208_nR11bf , \8209 , \8210 , \8211 ,
         \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 ,
         \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229_nR11d4 , \8230 , \8231 ,
         \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 ,
         \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250_nR11e9 , \8251 ,
         \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 ,
         \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271_nR11fe ,
         \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 ,
         \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 ,
         \8292_nR1213 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 ,
         \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 ,
         \8312 , \8313_nR1228 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 ,
         \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 ,
         \8332 , \8333 , \8334_nR123d , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 ,
         \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 ,
         \8352 , \8353 , \8354 , \8355_nR1252 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 ,
         \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 ,
         \8372 , \8373 , \8374 , \8375 , \8376_nR1267 , \8377 , \8378 , \8379 , \8380 , \8381 ,
         \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 ,
         \8392 , \8393 , \8394 , \8395 , \8396 , \8397_nR127c , \8398 , \8399 , \8400 , \8401 ,
         \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 ,
         \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418_nR1291 , \8419 , \8420 , \8421 ,
         \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 ,
         \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439_nR12a6 , \8440 , \8441 ,
         \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 ,
         \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460_nR12bb , \8461 ,
         \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 ,
         \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481_nR12d0 ,
         \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 ,
         \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 ,
         \8502_nR12e5 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 ,
         \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 ,
         \8522 , \8523_nR12fa , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 ,
         \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 ,
         \8542 , \8543 , \8544_nR130f , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 ,
         \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 ,
         \8562 , \8563 , \8564 , \8565_nR1324 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 ,
         \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 ,
         \8582 , \8583 , \8584 , \8585 , \8586_nR1339 , \8587 , \8588 , \8589 , \8590 , \8591 ,
         \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 ,
         \8602 , \8603 , \8604 , \8605 , \8606 , \8607_nR134e , \8608 , \8609 , \8610 , \8611 ,
         \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 ,
         \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628_nR1363 , \8629 , \8630 , \8631 ,
         \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 ,
         \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649_nR1378 , \8650 , \8651 ,
         \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 ,
         \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670_nR138d , \8671 ,
         \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 ,
         \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691_nR13a2 ,
         \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 ,
         \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 ,
         \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 ,
         \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 ,
         \8732_nR3163 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 ,
         \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 ,
         \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 ,
         \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 ,
         \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 ,
         \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 ,
         \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 ,
         \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 ,
         \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 ,
         \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 ,
         \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 ,
         \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 ,
         \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 ,
         \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 ,
         \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 ,
         \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 ,
         \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 ,
         \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 ,
         \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918_nR3106 , \8919 , \8920 , \8921 ,
         \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 ,
         \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 ,
         \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 ,
         \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 ,
         \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 ,
         \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 ,
         \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 ,
         \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 ,
         \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010_nR309d , \9011 ,
         \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 ,
         \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 ,
         \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 ,
         \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 ,
         \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 ,
         \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 ,
         \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 ,
         \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 ,
         \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100_nR3028 , \9101 ,
         \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 ,
         \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 ,
         \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 ,
         \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 ,
         \9142 , \9143 , \9144 , \9145 , \9146_nR2fa3 , \9147 , \9148 , \9149 , \9150 , \9151 ,
         \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 ,
         \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 ,
         \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 ,
         \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 ,
         \9192_nR2f16 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 ,
         \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 ,
         \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 ,
         \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 ,
         \9232 , \9233 , \9234 , \9235 , \9236_nR2e85 , \9237 , \9238 , \9239 , \9240 , \9241 ,
         \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 ,
         \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 ,
         \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 ,
         \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280_nR2dec , \9281 ,
         \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 ,
         \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 ,
         \9302 , \9303 , \9304_nR2d4b , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 ,
         \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 ,
         \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328_nR2ca8 , \9329 , \9330 , \9331 ,
         \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 ,
         \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 ,
         \9352_nR2bf5 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 ,
         \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 ,
         \9372 , \9373 , \9374 , \9375 , \9376_nR2b3c , \9377 , \9378 , \9379 , \9380 , \9381 ,
         \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 ,
         \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398_nR2a7b , \9399 , \9400 , \9401 ,
         \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 ,
         \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420_nR29bc , \9421 ,
         \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 ,
         \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 ,
         \9442_nR28fd , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 ,
         \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 ,
         \9462 , \9463 , \9464_nR2814 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 ,
         \9472 , \9473 , \9474_nR272d , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 ,
         \9482 , \9483 , \9484_nR2654 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 ,
         \9492 , \9493 , \9494_nR257b , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 ,
         \9502 , \9503 , \9504_nR24aa , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 ,
         \9512 , \9513 , \9514_nR23d5 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 ,
         \9522 , \9523 , \9524_nR230a , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 ,
         \9532 , \9533 , \9534_nR21f1 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 ,
         \9542 , \9543 , \9544_nR213c , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 ,
         \9552 , \9553 , \9554_nR2009 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 ,
         \9562 , \9563 , \9564_nR1f6c , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 ,
         \9572 , \9573 , \9574_nR1e51 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 ,
         \9582 , \9583 , \9584_nR1dc8 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 ,
         \9592 , \9593 , \9594_nR1cc1 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 ,
         \9602 , \9603 , \9604_nR1c54 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 ,
         \9612 , \9613 , \9614_nR1b67 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 ,
         \9622 , \9623 , \9624_nR1b12 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 ,
         \9632 , \9633 , \9634 , \9635 , \9636_nR1a41 , \9637 , \9638 , \9639 , \9640 , \9641 ,
         \9642_nR19fc , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 ,
         \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 ,
         \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 ,
         \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 ,
         \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 ,
         \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 ,
         \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 ,
         \9712 , \9713 , \9714_nR3911 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 ,
         \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 ,
         \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739_nR38ed , \9740 , \9741 ,
         \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 ,
         \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 ,
         \9762 , \9763 , \9764_nR3766 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 ,
         \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 ,
         \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789_nR3742 , \9790 , \9791 ,
         \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 ,
         \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 ,
         \9812 , \9813 , \9814_nR35cd , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 ,
         \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 ,
         \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839_nR35a9 , \9840 , \9841 ,
         \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 ,
         \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 ,
         \9862 , \9863 , \9864_nR346b , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 ,
         \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 ,
         \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889_nR3447 , \9890 , \9891 ,
         \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 ,
         \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 ,
         \9912 , \9913 , \9914_nR333a , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 ,
         \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 ,
         \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939_nR3353 , \9940 , \9941 ,
         \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 ,
         \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 ,
         \9962 , \9963 , \9964_nR3230 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 ,
         \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 ,
         \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988_nR3214 , \9989 , \9990 , \9991 ,
         \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 ,
         \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 ,
         \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 ,
         \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 ,
         \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 ,
         \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 ,
         \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 ,
         \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 ,
         \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 ,
         \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 ,
         \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 ,
         \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 ,
         \10112 , \10113 , \10114 , \10115_nR4011 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 ,
         \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 ,
         \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 ,
         \10142 , \10143_nR3ad9 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 ,
         \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 ,
         \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 ,
         \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 ,
         \10182 , \10183 , \10184_nR4105 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 ,
         \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 ,
         \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211_nR3f4f ,
         \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 ,
         \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 ,
         \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 ,
         \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 ,
         \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 ,
         \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 ,
         \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 ,
         \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 ,
         \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 ,
         \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 ,
         \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 ,
         \10322_nR3db4 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 ,
         \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 ,
         \10342 , \10343_nR3e8e , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 ,
         \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 ,
         \10362 , \10363 , \10364 , \10365 , \10366_nR3cc9 , \10367 , \10368 , \10369 , \10370 , \10371 ,
         \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 ,
         \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 ,
         \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 ,
         \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 ,
         \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 ,
         \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 ,
         \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 ,
         \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 ,
         \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459_nR3b16 , \10460 , \10461 ,
         \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 ,
         \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 ,
         \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 ,
         \10492_nR3bea , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 ,
         \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 ,
         \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519_nR3949 , \10520 , \10521 ,
         \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 ,
         \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 ,
         \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 ,
         \10552_nR3a20 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 ,
         \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 ,
         \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581_nR378a ,
         \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 ,
         \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 ,
         \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610_nR3853 , \10611 ,
         \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 ,
         \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 ,
         \10632 , \10633 , \10634 , \10635 , \10636_nR35f1 , \10637 , \10638 , \10639 , \10640 , \10641 ,
         \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 ,
         \10652 , \10653 , \10654 , \10655 , \10656 , \10657_nR36a4 , \10658 , \10659 , \10660 , \10661 ,
         \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 ,
         \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681_nR348d ,
         \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 ,
         \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 ,
         \10702_nR3534 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 ,
         \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 ,
         \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729_nR331d , \10730 , \10731 ,
         \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 ,
         \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750_nR33ee , \10751 ,
         \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 ,
         \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 ,
         \10772 , \10773_nR32db , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 ,
         \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 ,
         \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 ,
         \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 ,
         \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 ,
         \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 ,
         \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 ,
         \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 ,
         \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 ,
         \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 ,
         \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 ,
         \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 ,
         \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 ,
         \10902 , \10903 , \10904 , \10905 , \10906_nR31e3 , \10907 , \10908 , \10909 , \10910 , \10911 ,
         \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 ,
         \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 ,
         \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 ,
         \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 ,
         \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 ,
         \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 ,
         \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 ,
         \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 ,
         \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 ,
         \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 ,
         \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 ,
         \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 ,
         \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 ,
         \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 ,
         \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 ,
         \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 ,
         \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 ,
         \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 ,
         \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 ,
         \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 ,
         \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 ,
         \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 ,
         \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 ,
         \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 ,
         \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 ,
         \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 ,
         \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 ,
         \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 ,
         \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 ,
         \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 ,
         \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 ,
         \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 ,
         \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 ,
         \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 ,
         \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 ,
         \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 ,
         \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 ,
         \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 ,
         \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 ,
         \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 ,
         \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 ,
         \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 ,
         \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 ,
         \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 ,
         \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 ,
         \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 ,
         \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 ,
         \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 ,
         \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 ,
         \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 ,
         \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 ,
         \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 ,
         \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 ,
         \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 ,
         \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 ,
         \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 ,
         \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 ,
         \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 ,
         \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 ,
         \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 ,
         \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 ,
         \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 ,
         \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 ,
         \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 ,
         \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 ,
         \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 ,
         \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 ,
         \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 ,
         \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 ,
         \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 ,
         \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 ,
         \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 ,
         \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 ,
         \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 ,
         \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 ,
         \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 ,
         \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 ,
         \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 ,
         \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 ,
         \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 ,
         \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 ,
         \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 ,
         \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 ,
         \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 ,
         \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 ,
         \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 ,
         \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 ,
         \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 ,
         \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 ,
         \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 ,
         \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 ,
         \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 ,
         \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 ,
         \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 ,
         \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 ,
         \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 ,
         \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 ,
         \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 ,
         \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 ,
         \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 ,
         \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 ,
         \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 ,
         \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 ,
         \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 ,
         \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 ,
         \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 ,
         \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 ,
         \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 ,
         \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 ,
         \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 ,
         \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 ,
         \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 ,
         \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 ,
         \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 ,
         \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 ,
         \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 ,
         \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 ,
         \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 ,
         \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 ,
         \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 ,
         \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 ,
         \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 ,
         \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 ,
         \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 ,
         \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 ,
         \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 ,
         \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 ,
         \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 ,
         \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 ,
         \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 ,
         \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 ,
         \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 ,
         \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 ,
         \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 ,
         \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 ,
         \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 ,
         \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 ,
         \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 ,
         \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 ,
         \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 ,
         \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 ,
         \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 ,
         \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 ,
         \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 ,
         \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 ,
         \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 ,
         \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 ,
         \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 ,
         \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 ,
         \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 ,
         \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 ,
         \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 ,
         \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 ,
         \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 ,
         \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 ,
         \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 ,
         \12472 , \12473 , \12474 , \12475 , \12476_nR39aa , \12477 , \12478 , \12479 , \12480 , \12481 ,
         \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 ,
         \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501_nR3986 ,
         \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 ,
         \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 ,
         \12522 , \12523 , \12524 , \12525 , \12526_nR37f3 , \12527 , \12528 , \12529 , \12530 , \12531 ,
         \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 ,
         \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551_nR37cf ,
         \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 ,
         \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 ,
         \12572 , \12573 , \12574 , \12575 , \12576_nR3650 , \12577 , \12578 , \12579 , \12580 , \12581 ,
         \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 ,
         \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601_nR362c ,
         \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 ,
         \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 ,
         \12622 , \12623 , \12624 , \12625 , \12626_nR34e1 , \12627 , \12628 , \12629 , \12630 , \12631 ,
         \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 ,
         \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651_nR34bd ,
         \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 ,
         \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 ,
         \12672 , \12673 , \12674 , \12675 , \12676_nR33a2 , \12677 , \12678 , \12679 , \12680 , \12681 ,
         \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 ,
         \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701_nR33bb ,
         \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 ,
         \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 ,
         \12722 , \12723 , \12724 , \12725 , \12726_nR32b8 , \12727 , \12728 , \12729 , \12730 , \12731 ,
         \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 ,
         \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750_nR329c , \12751 ,
         \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 ,
         \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 ,
         \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 ,
         \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 ,
         \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 ,
         \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 ,
         \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 ,
         \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 ,
         \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 ,
         \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 ,
         \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 ,
         \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 ,
         \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 ,
         \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 ,
         \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 ,
         \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909_nR4084 , \12910 , \12911 ,
         \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 ,
         \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 ,
         \12932 , \12933 , \12934 , \12935 , \12936 , \12937_nR3b65 , \12938 , \12939 , \12940 , \12941 ,
         \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 ,
         \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 ,
         \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 ,
         \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978_nR4179 , \12979 , \12980 , \12981 ,
         \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 ,
         \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 ,
         \13002 , \13003 , \13004 , \13005_nR3fbb , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 ,
         \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 ,
         \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 ,
         \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 ,
         \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 ,
         \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 ,
         \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 ,
         \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 ,
         \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 ,
         \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 ,
         \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 ,
         \13112 , \13113 , \13114 , \13115 , \13116_nR3e1c , \13117 , \13118 , \13119 , \13120 , \13121 ,
         \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 ,
         \13132 , \13133 , \13134 , \13135 , \13136 , \13137_nR3efa , \13138 , \13139 , \13140 , \13141 ,
         \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 ,
         \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160_nR3d33 , \13161 ,
         \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 ,
         \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 ,
         \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 ,
         \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 ,
         \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 ,
         \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 ,
         \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 ,
         \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 ,
         \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 ,
         \13252 , \13253_nR3ba2 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 ,
         \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 ,
         \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 ,
         \13282 , \13283 , \13284 , \13285 , \13286_nR3c4f , \13287 , \13288 , \13289 , \13290 , \13291 ,
         \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 ,
         \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 ,
         \13312 , \13313_nR39e2 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 ,
         \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 ,
         \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 ,
         \13342 , \13343 , \13344 , \13345 , \13346_nR3a7a , \13347 , \13348 , \13349 , \13350 , \13351 ,
         \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 ,
         \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 ,
         \13372 , \13373 , \13374 , \13375_nR3817 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 ,
         \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 ,
         \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 ,
         \13402 , \13403 , \13404_nR38a1 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 ,
         \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 ,
         \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430_nR3674 , \13431 ,
         \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 ,
         \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451_nR36e8 ,
         \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 ,
         \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 ,
         \13472 , \13473 , \13474 , \13475_nR3503 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 ,
         \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 ,
         \13492 , \13493 , \13494 , \13495 , \13496_nR356a , \13497 , \13498 , \13499 , \13500 , \13501 ,
         \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 ,
         \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 ,
         \13522 , \13523_nR3385 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 ,
         \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 ,
         \13542 , \13543 , \13544_nR3418 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 ,
         \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 ,
         \13562 , \13563 , \13564 , \13565 , \13566 , \13567_nR32fd , \13568 , \13569 , \13570 , \13571 ,
         \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 ,
         \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 ,
         \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 ,
         \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 ,
         \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 ,
         \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 ,
         \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 ,
         \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 ,
         \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 ,
         \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 ,
         \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 ,
         \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 ,
         \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700_nR326b , \13701 ,
         \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 ,
         \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 ,
         \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 ,
         \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 ,
         \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 ,
         \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 ,
         \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 ,
         \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 ,
         \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 ,
         \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 ,
         \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 ,
         \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 ,
         \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 ,
         \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 ,
         \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 ,
         \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 ,
         \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 ,
         \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 ,
         \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 ,
         \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 ,
         \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 ,
         \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 ,
         \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 ,
         \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 ,
         \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 ,
         \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 ,
         \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 ,
         \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 ,
         \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 ,
         \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 ,
         \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 ,
         \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 ,
         \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 ,
         \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 ,
         \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 ,
         \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 ,
         \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 ,
         \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 ,
         \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 ,
         \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 ,
         \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 ,
         \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 ,
         \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 ,
         \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 ,
         \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 ,
         \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 ,
         \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 ,
         \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 ,
         \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 ,
         \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 ,
         \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 ,
         \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 ,
         \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 ,
         \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 ,
         \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 ,
         \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 ,
         \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 ,
         \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 ,
         \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 ,
         \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 ,
         \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 ,
         \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 ,
         \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 ,
         \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 ,
         \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 ,
         \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 ,
         \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 ,
         \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 ,
         \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 ,
         \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 ,
         \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 ,
         \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 ,
         \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 ,
         \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 ,
         \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 ,
         \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 ,
         \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 ,
         \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 ,
         \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 ,
         \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 ,
         \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 ,
         \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 ,
         \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 ,
         \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 ,
         \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 ,
         \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 ,
         \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 ,
         \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 ,
         \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 ,
         \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 ,
         \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 ,
         \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 ,
         \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 ,
         \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 ,
         \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 ,
         \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 ,
         \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 ,
         \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 ,
         \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 ,
         \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 ,
         \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 ,
         \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 ,
         \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 ,
         \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 ,
         \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 ,
         \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 ,
         \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 ,
         \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 ,
         \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 ,
         \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 ,
         \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 ,
         \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 ,
         \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 ,
         \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 ,
         \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 ,
         \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 ,
         \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 ,
         \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 ,
         \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 ,
         \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 ,
         \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 ,
         \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 ,
         \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 ,
         \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 ,
         \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 ,
         \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 ,
         \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 ,
         \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 ,
         \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 ,
         \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 ,
         \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 ,
         \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 ,
         \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 ,
         \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 ,
         \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 ,
         \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 ,
         \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 ,
         \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 ,
         \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 ,
         \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 ,
         \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 ,
         \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 ,
         \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 ,
         \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 ,
         \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 ,
         \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 ,
         \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 ,
         \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 ,
         \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 ,
         \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 ,
         \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 ,
         \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 ,
         \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 ,
         \15232 , \15233 , \15234 , \15235 , \15236_nR143b , \15237 , \15238 , \15239 , \15240 , \15241 ,
         \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 ,
         \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261_nR1454 ,
         \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 ,
         \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 ,
         \15282 , \15283 , \15284 , \15285 , \15286_nR146d , \15287 , \15288 , \15289 , \15290 , \15291 ,
         \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 ,
         \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311_nR1486 ,
         \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 ,
         \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 ,
         \15332 , \15333 , \15334 , \15335 , \15336_nR149f , \15337 , \15338 , \15339 , \15340 , \15341 ,
         \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 ,
         \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361_nR14b8 ,
         \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 ,
         \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 ,
         \15382 , \15383 , \15384 , \15385 , \15386_nR14d1 , \15387 , \15388 , \15389 , \15390 , \15391 ,
         \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 ,
         \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411_nR14ea ,
         \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 ,
         \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 ,
         \15432 , \15433 , \15434 , \15435 , \15436_nR1503 , \15437 , \15438 , \15439 , \15440 , \15441 ,
         \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 ,
         \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461_nR151c ,
         \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 ,
         \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 ,
         \15482 , \15483 , \15484 , \15485 , \15486_nR1535 , \15487 , \15488 , \15489 , \15490 , \15491 ,
         \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 ,
         \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511_nR154e ,
         \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 ,
         \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 ,
         \15532 , \15533 , \15534 , \15535_nR1568 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 ,
         \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 ,
         \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 ,
         \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 ,
         \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 ,
         \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 ,
         \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 ,
         \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 ,
         \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 ,
         \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 ,
         \15632 , \15633 , \15634 , \15635 , \15636_nR15d1 , \15637 , \15638 , \15639 , \15640 , \15641 ,
         \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 ,
         \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 ,
         \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 ,
         \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 ,
         \15682_nR15ff , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 ,
         \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 ,
         \15702 , \15703_nR1614 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 ,
         \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 ,
         \15722 , \15723 , \15724_nR1629 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 ,
         \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 ,
         \15742 , \15743 , \15744 , \15745_nR163e , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 ,
         \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 ,
         \15762 , \15763 , \15764 , \15765 , \15766_nR1653 , \15767 , \15768 , \15769 , \15770 , \15771 ,
         \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 ,
         \15782 , \15783 , \15784 , \15785 , \15786 , \15787_nR1668 , \15788 , \15789 , \15790 , \15791 ,
         \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 ,
         \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808_nR167d , \15809 , \15810 , \15811 ,
         \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 ,
         \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829_nR1692 , \15830 , \15831 ,
         \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 ,
         \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850_nR16a7 , \15851 ,
         \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 ,
         \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871_nR16bc ,
         \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 ,
         \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 ,
         \15892_nR16d1 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 ,
         \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 ,
         \15912 , \15913_nR16e6 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 ,
         \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 ,
         \15932 , \15933 , \15934_nR16fb , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 ,
         \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 ,
         \15952 , \15953 , \15954 , \15955_nR1710 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 ,
         \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 ,
         \15972 , \15973 , \15974 , \15975 , \15976_nR1725 , \15977 , \15978 , \15979 , \15980 , \15981 ,
         \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 ,
         \15992 , \15993 , \15994 , \15995 , \15996 , \15997_nR173a , \15998 , \15999 , \16000 , \16001 ,
         \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 ,
         \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018_nR174f , \16019 , \16020 , \16021 ,
         \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 ,
         \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039_nR1764 , \16040 , \16041 ,
         \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 ,
         \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060_nR1779 , \16061 ,
         \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 ,
         \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081_nR178e ,
         \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 ,
         \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 ,
         \16102_nR17a3 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 ,
         \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 ,
         \16122 , \16123_nR17b8 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 ,
         \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 ,
         \16142 , \16143 , \16144_nR17cd , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 ,
         \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 ,
         \16162 , \16163 , \16164 , \16165_nR17e2 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 ,
         \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 ,
         \16182 , \16183 , \16184 , \16185 , \16186_nR17f7 , \16187 , \16188 , \16189 , \16190 , \16191 ,
         \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 ,
         \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 ,
         \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 ,
         \16222 , \16223 , \16224 , \16225 , \16226 , \16227_nR4a2b , \16228 , \16229 , \16230 , \16231 ,
         \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 ,
         \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 ,
         \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 ,
         \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 ,
         \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 ,
         \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 ,
         \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 ,
         \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 ,
         \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 ,
         \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 ,
         \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 ,
         \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 ,
         \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 ,
         \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 ,
         \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 ,
         \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 ,
         \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 ,
         \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 ,
         \16412 , \16413_nR49ce , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 ,
         \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 ,
         \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 ,
         \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 ,
         \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 ,
         \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 ,
         \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 ,
         \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 ,
         \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 ,
         \16502 , \16503 , \16504 , \16505_nR4965 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 ,
         \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 ,
         \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 ,
         \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 ,
         \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 ,
         \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 ,
         \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 ,
         \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 ,
         \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 ,
         \16592 , \16593 , \16594 , \16595_nR48f0 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 ,
         \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 ,
         \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 ,
         \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 ,
         \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641_nR486b ,
         \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 ,
         \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 ,
         \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 ,
         \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 ,
         \16682 , \16683 , \16684 , \16685 , \16686 , \16687_nR47de , \16688 , \16689 , \16690 , \16691 ,
         \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 ,
         \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 ,
         \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 ,
         \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731_nR474d ,
         \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 ,
         \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 ,
         \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 ,
         \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 ,
         \16772 , \16773 , \16774 , \16775_nR46b4 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 ,
         \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 ,
         \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799_nR4613 , \16800 , \16801 ,
         \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 ,
         \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 ,
         \16822 , \16823_nR4570 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 ,
         \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 ,
         \16842 , \16843 , \16844 , \16845 , \16846 , \16847_nR44bd , \16848 , \16849 , \16850 , \16851 ,
         \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 ,
         \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871_nR4404 ,
         \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 ,
         \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 ,
         \16892 , \16893_nR4343 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 ,
         \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 ,
         \16912 , \16913 , \16914 , \16915_nR4284 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 ,
         \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 ,
         \16932 , \16933 , \16934 , \16935 , \16936 , \16937_nR41c5 , \16938 , \16939 , \16940 , \16941 ,
         \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 ,
         \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959_nR40dc , \16960 , \16961 ,
         \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969_nR3ff5 , \16970 , \16971 ,
         \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979_nR3f1c , \16980 , \16981 ,
         \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989_nR3e43 , \16990 , \16991 ,
         \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999_nR3d72 , \17000 , \17001 ,
         \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009_nR3c9d , \17010 , \17011 ,
         \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019_nR3bd2 , \17020 , \17021 ,
         \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029_nR3ab9 , \17030 , \17031 ,
         \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039_nR3a04 , \17040 , \17041 ,
         \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049_nR38d1 , \17050 , \17051 ,
         \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059_nR3834 , \17060 , \17061 ,
         \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069_nR3719 , \17070 , \17071 ,
         \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079_nR3690 , \17080 , \17081 ,
         \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089_nR3589 , \17090 , \17091 ,
         \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099_nR351c , \17100 , \17101 ,
         \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109_nR342f , \17110 , \17111 ,
         \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119_nR33da , \17120 , \17121 ,
         \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131_nR3309 ,
         \17132 , \17133 , \17134 , \17135 , \17136 , \17137_nR32c4 , \17138 ;
buf \U$labaj1789 ( R_267_b04ddc8, \8733 );
buf \U$labaj1790 ( R_268_b04de70, \8919 );
buf \U$labaj1791 ( R_269_b04df18, \9011 );
buf \U$labaj1792 ( R_26a_b04dfc0, \9101 );
buf \U$labaj1793 ( R_26b_b04e068, \9147 );
buf \U$labaj1794 ( R_26c_b04e110, \9193 );
buf \U$labaj1795 ( R_26d_b04e1b8, \9237 );
buf \U$labaj1796 ( R_26e_b04e260, \9281 );
buf \U$labaj1797 ( R_26f_b04e308, \9305 );
buf \U$labaj1798 ( R_270_b04e3b0, \9329 );
buf \U$labaj1799 ( R_271_b04e458, \9353 );
buf \U$labaj1800 ( R_272_b04e500, \9377 );
buf \U$labaj1801 ( R_273_b04e5a8, \9399 );
buf \U$labaj1802 ( R_274_b04e650, \9421 );
buf \U$labaj1803 ( R_275_b04e6f8, \9443 );
buf \U$labaj1804 ( R_276_b04e7a0, \9465 );
buf \U$labaj1805 ( R_277_b04e848, \9475 );
buf \U$labaj1806 ( R_278_b04e8f0, \9485 );
buf \U$labaj1807 ( R_279_b04e998, \9495 );
buf \U$labaj1808 ( R_27a_b04ea40, \9505 );
buf \U$labaj1809 ( R_27b_b04eae8, \9515 );
buf \U$labaj1810 ( R_27c_b04eb90, \9525 );
buf \U$labaj1811 ( R_27d_b04ec38, \9535 );
buf \U$labaj1812 ( R_27e_b04ece0, \9545 );
buf \U$labaj1813 ( R_27f_b04ed88, \9555 );
buf \U$labaj1814 ( R_280_b04ee30, \9565 );
buf \U$labaj1815 ( R_281_b04eed8, \9575 );
buf \U$labaj1816 ( R_282_b04ef80, \9585 );
buf \U$labaj1817 ( R_283_b04f028, \9595 );
buf \U$labaj1818 ( R_284_b04f0d0, \9605 );
buf \U$labaj1819 ( R_285_b04f178, \9615 );
buf \U$labaj1820 ( R_286_b04f220, \9625 );
buf \U$labaj1821 ( R_287_b04f2c8, \9637 );
buf \U$labaj1822 ( R_288_b04f370, \9643 );
buf \U$labaj1823 ( R_289_b04f418, \16228 );
buf \U$labaj1824 ( R_28a_b04f4c0, \16414 );
buf \U$labaj1825 ( R_28b_b04f568, \16506 );
buf \U$labaj1826 ( R_28c_b04f610, \16596 );
buf \U$labaj1827 ( R_28d_b04f6b8, \16642 );
buf \U$labaj1828 ( R_28e_b04f760, \16688 );
buf \U$labaj1829 ( R_28f_b04f808, \16732 );
buf \U$labaj1830 ( R_290_b04f8b0, \16776 );
buf \U$labaj1831 ( R_291_b04f958, \16800 );
buf \U$labaj1832 ( R_292_b04fa00, \16824 );
buf \U$labaj1833 ( R_293_b04faa8, \16848 );
buf \U$labaj1834 ( R_294_b04fb50, \16872 );
buf \U$labaj1835 ( R_295_b04fbf8, \16894 );
buf \U$labaj1836 ( R_296_b04fca0, \16916 );
buf \U$labaj1837 ( R_297_b04fd48, \16938 );
buf \U$labaj1838 ( R_298_b04fdf0, \16960 );
buf \U$labaj1839 ( R_299_b04fe98, \16970 );
buf \U$labaj1840 ( R_29a_b04ff40, \16980 );
buf \U$labaj1841 ( R_29b_b04ffe8, \16990 );
buf \U$labaj1842 ( R_29c_b050090, \17000 );
buf \U$labaj1843 ( R_29d_b050138, \17010 );
buf \U$labaj1844 ( R_29e_b0501e0, \17020 );
buf \U$labaj1845 ( R_29f_b050288, \17030 );
buf \U$labaj1846 ( R_2a0_b050330, \17040 );
buf \U$labaj1847 ( R_2a1_b0503d8, \17050 );
buf \U$labaj1848 ( R_2a2_b050480, \17060 );
buf \U$labaj1849 ( R_2a3_b050528, \17070 );
buf \U$labaj1850 ( R_2a4_b0505d0, \17080 );
buf \U$labaj1851 ( R_2a5_b050678, \17090 );
buf \U$labaj1852 ( R_2a6_b050720, \17100 );
buf \U$labaj1853 ( R_2a7_b0507c8, \17110 );
buf \U$labaj1854 ( R_2a8_b050870, \17120 );
buf \U$labaj1855 ( R_2a9_b050918, \17132 );
buf \U$labaj1856 ( R_2aa_b0509c0, \17138 );
buf \U$5 ( \2149 , RI2b5e785ebcf0_2);
buf \U$6 ( \2150 , RI2b5e785ebc78_3);
buf \U$7 ( \2151 , RI2b5e785ebc00_4);
buf \U$8 ( \2152 , RI2b5e785ebb88_5);
buf \U$9 ( \2153 , RI2b5e785ebb10_6);
buf \U$10 ( \2154 , RI2b5e785eba98_7);
buf \U$11 ( \2155 , RI2b5e785eba20_8);
buf \U$12 ( \2156 , RI2b5e785eb9a8_9);
buf \U$13 ( \2157 , RI2b5e785eb930_10);
buf \U$14 ( \2158 , RI2b5e785eb8b8_11);
buf \U$15 ( \2159 , RI2b5e785eb840_12);
and \U$16 ( \2160 , \2158 , \2159 );
and \U$17 ( \2161 , \2157 , \2160 );
and \U$18 ( \2162 , \2156 , \2161 );
and \U$19 ( \2163 , \2155 , \2162 );
and \U$20 ( \2164 , \2154 , \2163 );
and \U$21 ( \2165 , \2153 , \2164 );
and \U$22 ( \2166 , \2152 , \2165 );
and \U$23 ( \2167 , \2151 , \2166 );
and \U$24 ( \2168 , \2150 , \2167 );
xor \U$25 ( \2169 , \2149 , \2168 );
buf \U$26 ( \2170 , \2169 );
buf \U$27 ( \2171 , \2170 );
not \U$28 ( \2172 , RI2b5e785aeb98_596);
nor \U$29 ( \2173 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$30 ( \2174 , RI2b5e785daa40_28, \2173 );
and \U$31 ( \2175 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$32 ( \2176 , RI2b5e78549540_41, \2175 );
not \U$33 ( \2177 , RI2b5e785ae9b8_600);
and \U$34 ( \2178 , \2177 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$35 ( \2179 , RI2b5e785388a8_54, \2178 );
not \U$36 ( \2180 , RI2b5e785aea30_599);
and \U$37 ( \2181 , RI2b5e785ae9b8_600, \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$38 ( \2182 , RI2b5e784a6330_67, \2181 );
and \U$39 ( \2183 , \2177 , \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$40 ( \2184 , RI2b5e78495698_80, \2183 );
not \U$41 ( \2185 , RI2b5e785aeaa8_598);
and \U$42 ( \2186 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, \2172 );
and \U$43 ( \2187 , RI2b5e78495080_93, \2186 );
and \U$44 ( \2188 , \2177 , RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, \2172 );
and \U$45 ( \2189 , RI2b5e78403b80_106, \2188 );
and \U$46 ( \2190 , RI2b5e785ae9b8_600, \2180 , \2185 , RI2b5e785aeb20_597, \2172 );
and \U$47 ( \2191 , RI2b5e775b1e60_119, \2190 );
and \U$48 ( \2192 , \2177 , \2180 , \2185 , RI2b5e785aeb20_597, \2172 );
and \U$49 ( \2193 , RI2b5e7750bdf8_132, \2192 );
nor \U$50 ( \2194 , \2177 , \2180 , \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$51 ( \2195 , RI2b5e774ff5d0_145, \2194 );
nor \U$52 ( \2196 , RI2b5e785ae9b8_600, \2180 , \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$53 ( \2197 , RI2b5e774f65e8_158, \2196 );
nor \U$54 ( \2198 , \2177 , RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$55 ( \2199 , RI2b5e774eabd0_171, \2198 );
nor \U$56 ( \2200 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$57 ( \2201 , RI2b5e774de3a8_184, \2200 );
nor \U$58 ( \2202 , \2177 , \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$59 ( \2203 , RI2b5e774d53c0_197, \2202 );
nor \U$60 ( \2204 , RI2b5e785ae9b8_600, \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$61 ( \2205 , RI2b5e785f4300_210, \2204 );
nor \U$62 ( \2206 , \2177 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$63 ( \2207 , RI2b5e785f3ce8_223, \2206 );
nor \U$64 ( \2208 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$65 ( \2209 , RI2b5e785eb0c0_236, \2208 );
or \U$66 ( \2210 , \2174 , \2176 , \2179 , \2182 , \2184 , \2187 , \2189 , \2191 , \2193 , \2195 , \2197 , \2199 , \2201 , \2203 , \2205 , \2207 , \2209 );
buf \U$67 ( \2211 , RI2b5e785aeb98_596);
buf \U$68 ( \2212 , RI2b5e785ae9b8_600);
buf \U$69 ( \2213 , RI2b5e785aea30_599);
buf \U$70 ( \2214 , RI2b5e785aeaa8_598);
buf \U$71 ( \2215 , RI2b5e785aeb20_597);
or \U$72 ( \2216 , \2212 , \2213 , \2214 , \2215 );
and \U$73 ( \2217 , \2211 , \2216 );
buf \U$74 ( \2218 , \2217 );
_DC r2049 ( \2219_nR2049 , \2210 , \2218 );
buf \U$75 ( \2220 , \2219_nR2049 );
not \U$76 ( \2221 , \2220 );
xor \U$77 ( \2222 , \2171 , \2221 );
xor \U$78 ( \2223 , \2150 , \2167 );
buf \U$79 ( \2224 , \2223 );
buf \U$80 ( \2225 , \2224 );
and \U$81 ( \2226 , RI2b5e785da9c8_29, \2173 );
and \U$82 ( \2227 , RI2b5e785494c8_42, \2175 );
and \U$83 ( \2228 , RI2b5e78538830_55, \2178 );
and \U$84 ( \2229 , RI2b5e784a62b8_68, \2181 );
and \U$85 ( \2230 , RI2b5e78495620_81, \2183 );
and \U$86 ( \2231 , RI2b5e78495008_94, \2186 );
and \U$87 ( \2232 , RI2b5e78403b08_107, \2188 );
and \U$88 ( \2233 , RI2b5e775b1de8_120, \2190 );
and \U$89 ( \2234 , RI2b5e7750bd80_133, \2192 );
and \U$90 ( \2235 , RI2b5e774ff558_146, \2194 );
and \U$91 ( \2236 , RI2b5e774f6570_159, \2196 );
and \U$92 ( \2237 , RI2b5e774eab58_172, \2198 );
and \U$93 ( \2238 , RI2b5e774de330_185, \2200 );
and \U$94 ( \2239 , RI2b5e774d5348_198, \2202 );
and \U$95 ( \2240 , RI2b5e785f4288_211, \2204 );
and \U$96 ( \2241 , RI2b5e785f3658_224, \2206 );
and \U$97 ( \2242 , RI2b5e785eb048_237, \2208 );
or \U$98 ( \2243 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 );
_DC r2025 ( \2244_nR2025 , \2243 , \2218 );
buf \U$99 ( \2245 , \2244_nR2025 );
not \U$100 ( \2246 , \2245 );
and \U$101 ( \2247 , \2225 , \2246 );
xor \U$102 ( \2248 , \2151 , \2166 );
buf \U$103 ( \2249 , \2248 );
buf \U$104 ( \2250 , \2249 );
and \U$105 ( \2251 , RI2b5e785da950_30, \2173 );
and \U$106 ( \2252 , RI2b5e78549450_43, \2175 );
and \U$107 ( \2253 , RI2b5e785387b8_56, \2178 );
and \U$108 ( \2254 , RI2b5e784a6240_69, \2181 );
and \U$109 ( \2255 , RI2b5e784955a8_82, \2183 );
and \U$110 ( \2256 , RI2b5e78494f90_95, \2186 );
and \U$111 ( \2257 , RI2b5e78403a90_108, \2188 );
and \U$112 ( \2258 , RI2b5e775b1d70_121, \2190 );
and \U$113 ( \2259 , RI2b5e7750bd08_134, \2192 );
and \U$114 ( \2260 , RI2b5e774ff4e0_147, \2194 );
and \U$115 ( \2261 , RI2b5e774f64f8_160, \2196 );
and \U$116 ( \2262 , RI2b5e774eaae0_173, \2198 );
and \U$117 ( \2263 , RI2b5e774de2b8_186, \2200 );
and \U$118 ( \2264 , RI2b5e774d52d0_199, \2202 );
and \U$119 ( \2265 , RI2b5e785f4210_212, \2204 );
and \U$120 ( \2266 , RI2b5e785eb5e8_225, \2206 );
and \U$121 ( \2267 , RI2b5e785e6c50_238, \2208 );
or \U$122 ( \2268 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 );
_DC r1e9e ( \2269_nR1e9e , \2268 , \2218 );
buf \U$123 ( \2270 , \2269_nR1e9e );
not \U$124 ( \2271 , \2270 );
and \U$125 ( \2272 , \2250 , \2271 );
xor \U$126 ( \2273 , \2152 , \2165 );
buf \U$127 ( \2274 , \2273 );
buf \U$128 ( \2275 , \2274 );
and \U$129 ( \2276 , RI2b5e785da8d8_31, \2173 );
and \U$130 ( \2277 , RI2b5e785493d8_44, \2175 );
and \U$131 ( \2278 , RI2b5e78538740_57, \2178 );
and \U$132 ( \2279 , RI2b5e784a61c8_70, \2181 );
and \U$133 ( \2280 , RI2b5e78495530_83, \2183 );
and \U$134 ( \2281 , RI2b5e78494f18_96, \2186 );
and \U$135 ( \2282 , RI2b5e78403a18_109, \2188 );
and \U$136 ( \2283 , RI2b5e775b1cf8_122, \2190 );
and \U$137 ( \2284 , RI2b5e7750bc90_135, \2192 );
and \U$138 ( \2285 , RI2b5e774ff468_148, \2194 );
and \U$139 ( \2286 , RI2b5e774f6480_161, \2196 );
and \U$140 ( \2287 , RI2b5e774eaa68_174, \2198 );
and \U$141 ( \2288 , RI2b5e774de240_187, \2200 );
and \U$142 ( \2289 , RI2b5e774d5258_200, \2202 );
and \U$143 ( \2290 , RI2b5e785f4198_213, \2204 );
and \U$144 ( \2291 , RI2b5e785eb570_226, \2206 );
and \U$145 ( \2292 , RI2b5e785e6bd8_239, \2208 );
or \U$146 ( \2293 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 );
_DC r1e7a ( \2294_nR1e7a , \2293 , \2218 );
buf \U$147 ( \2295 , \2294_nR1e7a );
not \U$148 ( \2296 , \2295 );
and \U$149 ( \2297 , \2275 , \2296 );
xor \U$150 ( \2298 , \2153 , \2164 );
buf \U$151 ( \2299 , \2298 );
buf \U$152 ( \2300 , \2299 );
and \U$153 ( \2301 , RI2b5e785da860_32, \2173 );
and \U$154 ( \2302 , RI2b5e78549360_45, \2175 );
and \U$155 ( \2303 , RI2b5e785386c8_58, \2178 );
and \U$156 ( \2304 , RI2b5e784a6150_71, \2181 );
and \U$157 ( \2305 , RI2b5e784954b8_84, \2183 );
and \U$158 ( \2306 , RI2b5e78494ea0_97, \2186 );
and \U$159 ( \2307 , RI2b5e784039a0_110, \2188 );
and \U$160 ( \2308 , RI2b5e775b1c80_123, \2190 );
and \U$161 ( \2309 , RI2b5e7750bc18_136, \2192 );
and \U$162 ( \2310 , RI2b5e774ff3f0_149, \2194 );
and \U$163 ( \2311 , RI2b5e774f6408_162, \2196 );
and \U$164 ( \2312 , RI2b5e774ea9f0_175, \2198 );
and \U$165 ( \2313 , RI2b5e774de1c8_188, \2200 );
and \U$166 ( \2314 , RI2b5e774d51e0_201, \2202 );
and \U$167 ( \2315 , RI2b5e785f4120_214, \2204 );
and \U$168 ( \2316 , RI2b5e785eb4f8_227, \2206 );
and \U$169 ( \2317 , RI2b5e785e64d0_240, \2208 );
or \U$170 ( \2318 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 );
_DC r1d05 ( \2319_nR1d05 , \2318 , \2218 );
buf \U$171 ( \2320 , \2319_nR1d05 );
not \U$172 ( \2321 , \2320 );
and \U$173 ( \2322 , \2300 , \2321 );
xor \U$174 ( \2323 , \2154 , \2163 );
buf \U$175 ( \2324 , \2323 );
buf \U$176 ( \2325 , \2324 );
and \U$177 ( \2326 , RI2b5e78549900_33, \2173 );
and \U$178 ( \2327 , RI2b5e78538c68_46, \2175 );
and \U$179 ( \2328 , RI2b5e78538650_59, \2178 );
and \U$180 ( \2329 , RI2b5e784a60d8_72, \2181 );
and \U$181 ( \2330 , RI2b5e78495440_85, \2183 );
and \U$182 ( \2331 , RI2b5e78494e28_98, \2186 );
and \U$183 ( \2332 , RI2b5e78403928_111, \2188 );
and \U$184 ( \2333 , RI2b5e775b1c08_124, \2190 );
and \U$185 ( \2334 , RI2b5e7750bba0_137, \2192 );
and \U$186 ( \2335 , RI2b5e774ff378_150, \2194 );
and \U$187 ( \2336 , RI2b5e774f6390_163, \2196 );
and \U$188 ( \2337 , RI2b5e774ea978_176, \2198 );
and \U$189 ( \2338 , RI2b5e774de150_189, \2200 );
and \U$190 ( \2339 , RI2b5e774d5168_202, \2202 );
and \U$191 ( \2340 , RI2b5e785f40a8_215, \2204 );
and \U$192 ( \2341 , RI2b5e785eb480_228, \2206 );
and \U$193 ( \2342 , RI2b5e785da608_241, \2208 );
or \U$194 ( \2343 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 );
_DC r1ce1 ( \2344_nR1ce1 , \2343 , \2218 );
buf \U$195 ( \2345 , \2344_nR1ce1 );
not \U$196 ( \2346 , \2345 );
and \U$197 ( \2347 , \2325 , \2346 );
xor \U$198 ( \2348 , \2155 , \2162 );
buf \U$199 ( \2349 , \2348 );
buf \U$200 ( \2350 , \2349 );
and \U$201 ( \2351 , RI2b5e78549888_34, \2173 );
and \U$202 ( \2352 , RI2b5e78538bf0_47, \2175 );
and \U$203 ( \2353 , RI2b5e785385d8_60, \2178 );
and \U$204 ( \2354 , RI2b5e784a6060_73, \2181 );
and \U$205 ( \2355 , RI2b5e784953c8_86, \2183 );
and \U$206 ( \2356 , RI2b5e78403ec8_99, \2186 );
and \U$207 ( \2357 , RI2b5e775b21a8_112, \2188 );
and \U$208 ( \2358 , RI2b5e775b1b90_125, \2190 );
and \U$209 ( \2359 , RI2b5e7750bb28_138, \2192 );
and \U$210 ( \2360 , RI2b5e774ff300_151, \2194 );
and \U$211 ( \2361 , RI2b5e774f6318_164, \2196 );
and \U$212 ( \2362 , RI2b5e774ea900_177, \2198 );
and \U$213 ( \2363 , RI2b5e774de0d8_190, \2200 );
and \U$214 ( \2364 , RI2b5e774d50f0_203, \2202 );
and \U$215 ( \2365 , RI2b5e785f4030_216, \2204 );
and \U$216 ( \2366 , RI2b5e785eb408_229, \2206 );
and \U$217 ( \2367 , RI2b5e785da590_242, \2208 );
or \U$218 ( \2368 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 );
_DC r1ba3 ( \2369_nR1ba3 , \2368 , \2218 );
buf \U$219 ( \2370 , \2369_nR1ba3 );
not \U$220 ( \2371 , \2370 );
and \U$221 ( \2372 , \2350 , \2371 );
xor \U$222 ( \2373 , \2156 , \2161 );
buf \U$223 ( \2374 , \2373 );
buf \U$224 ( \2375 , \2374 );
and \U$225 ( \2376 , RI2b5e78549810_35, \2173 );
and \U$226 ( \2377 , RI2b5e78538b78_48, \2175 );
and \U$227 ( \2378 , RI2b5e78538560_61, \2178 );
and \U$228 ( \2379 , RI2b5e784a5fe8_74, \2181 );
and \U$229 ( \2380 , RI2b5e78495350_87, \2183 );
and \U$230 ( \2381 , RI2b5e78403e50_100, \2186 );
and \U$231 ( \2382 , RI2b5e775b2130_113, \2188 );
and \U$232 ( \2383 , RI2b5e775b1b18_126, \2190 );
and \U$233 ( \2384 , RI2b5e7750bab0_139, \2192 );
and \U$234 ( \2385 , RI2b5e774ff288_152, \2194 );
and \U$235 ( \2386 , RI2b5e774f62a0_165, \2196 );
and \U$236 ( \2387 , RI2b5e774ea888_178, \2198 );
and \U$237 ( \2388 , RI2b5e774de060_191, \2200 );
and \U$238 ( \2389 , RI2b5e774d5078_204, \2202 );
and \U$239 ( \2390 , RI2b5e785f3fb8_217, \2204 );
and \U$240 ( \2391 , RI2b5e785eb390_230, \2206 );
and \U$241 ( \2392 , RI2b5e785da518_243, \2208 );
or \U$242 ( \2393 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 );
_DC r1b7f ( \2394_nR1b7f , \2393 , \2218 );
buf \U$243 ( \2395 , \2394_nR1b7f );
not \U$244 ( \2396 , \2395 );
and \U$245 ( \2397 , \2375 , \2396 );
xor \U$246 ( \2398 , \2157 , \2160 );
buf \U$247 ( \2399 , \2398 );
buf \U$248 ( \2400 , \2399 );
and \U$249 ( \2401 , RI2b5e78549798_36, \2173 );
and \U$250 ( \2402 , RI2b5e78538b00_49, \2175 );
and \U$251 ( \2403 , RI2b5e785384e8_62, \2178 );
and \U$252 ( \2404 , RI2b5e784a5f70_75, \2181 );
and \U$253 ( \2405 , RI2b5e784952d8_88, \2183 );
and \U$254 ( \2406 , RI2b5e78403dd8_101, \2186 );
and \U$255 ( \2407 , RI2b5e775b20b8_114, \2188 );
and \U$256 ( \2408 , RI2b5e775b1aa0_127, \2190 );
and \U$257 ( \2409 , RI2b5e7750ba38_140, \2192 );
and \U$258 ( \2410 , RI2b5e774ff210_153, \2194 );
and \U$259 ( \2411 , RI2b5e774f6228_166, \2196 );
and \U$260 ( \2412 , RI2b5e774ea810_179, \2198 );
and \U$261 ( \2413 , RI2b5e774ddfe8_192, \2200 );
and \U$262 ( \2414 , RI2b5e774d5000_205, \2202 );
and \U$263 ( \2415 , RI2b5e785f3f40_218, \2204 );
and \U$264 ( \2416 , RI2b5e785eb318_231, \2206 );
and \U$265 ( \2417 , RI2b5e785da4a0_244, \2208 );
or \U$266 ( \2418 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 );
_DC r1a72 ( \2419_nR1a72 , \2418 , \2218 );
buf \U$267 ( \2420 , \2419_nR1a72 );
not \U$268 ( \2421 , \2420 );
and \U$269 ( \2422 , \2400 , \2421 );
xor \U$270 ( \2423 , \2158 , \2159 );
buf \U$271 ( \2424 , \2423 );
buf \U$272 ( \2425 , \2424 );
and \U$273 ( \2426 , RI2b5e78549720_37, \2173 );
and \U$274 ( \2427 , RI2b5e78538a88_50, \2175 );
and \U$275 ( \2428 , RI2b5e78538470_63, \2178 );
and \U$276 ( \2429 , RI2b5e784a5ef8_76, \2181 );
and \U$277 ( \2430 , RI2b5e78495260_89, \2183 );
and \U$278 ( \2431 , RI2b5e78403d60_102, \2186 );
and \U$279 ( \2432 , RI2b5e775b2040_115, \2188 );
and \U$280 ( \2433 , RI2b5e775b1a28_128, \2190 );
and \U$281 ( \2434 , RI2b5e7750b9c0_141, \2192 );
and \U$282 ( \2435 , RI2b5e774ff198_154, \2194 );
and \U$283 ( \2436 , RI2b5e774f61b0_167, \2196 );
and \U$284 ( \2437 , RI2b5e774ea798_180, \2198 );
and \U$285 ( \2438 , RI2b5e774ddf70_193, \2200 );
and \U$286 ( \2439 , RI2b5e774d4f88_206, \2202 );
and \U$287 ( \2440 , RI2b5e785f3ec8_219, \2204 );
and \U$288 ( \2441 , RI2b5e785eb2a0_232, \2206 );
and \U$289 ( \2442 , RI2b5e785da428_245, \2208 );
or \U$290 ( \2443 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 );
_DC r1a8b ( \2444_nR1a8b , \2443 , \2218 );
buf \U$291 ( \2445 , \2444_nR1a8b );
not \U$292 ( \2446 , \2445 );
and \U$293 ( \2447 , \2425 , \2446 );
not \U$294 ( \2448 , \2159 );
buf \U$295 ( \2449 , \2448 );
buf \U$296 ( \2450 , \2449 );
and \U$297 ( \2451 , RI2b5e785496a8_38, \2173 );
and \U$298 ( \2452 , RI2b5e78538a10_51, \2175 );
and \U$299 ( \2453 , RI2b5e785383f8_64, \2178 );
and \U$300 ( \2454 , RI2b5e784a5e80_77, \2181 );
and \U$301 ( \2455 , RI2b5e784951e8_90, \2183 );
and \U$302 ( \2456 , RI2b5e78403ce8_103, \2186 );
and \U$303 ( \2457 , RI2b5e775b1fc8_116, \2188 );
and \U$304 ( \2458 , RI2b5e775b19b0_129, \2190 );
and \U$305 ( \2459 , RI2b5e7750b948_142, \2192 );
and \U$306 ( \2460 , RI2b5e774ff120_155, \2194 );
and \U$307 ( \2461 , RI2b5e774f6138_168, \2196 );
and \U$308 ( \2462 , RI2b5e774ea720_181, \2198 );
and \U$309 ( \2463 , RI2b5e774ddef8_194, \2200 );
and \U$310 ( \2464 , RI2b5e774d4f10_207, \2202 );
and \U$311 ( \2465 , RI2b5e785f3e50_220, \2204 );
and \U$312 ( \2466 , RI2b5e785eb228_233, \2206 );
and \U$313 ( \2467 , RI2b5e785da3b0_246, \2208 );
or \U$314 ( \2468 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 );
_DC r1968 ( \2469_nR1968 , \2468 , \2218 );
buf \U$315 ( \2470 , \2469_nR1968 );
not \U$316 ( \2471 , \2470 );
and \U$317 ( \2472 , \2450 , \2471 );
buf \U$318 ( \2473 , RI2b5e785db148_13);
buf \U$321 ( \2474 , \2473 );
and \U$322 ( \2475 , RI2b5e78549630_39, \2173 );
and \U$323 ( \2476 , RI2b5e78538998_52, \2175 );
and \U$324 ( \2477 , RI2b5e78538380_65, \2178 );
and \U$325 ( \2478 , RI2b5e784a5e08_78, \2181 );
and \U$326 ( \2479 , RI2b5e78495170_91, \2183 );
and \U$327 ( \2480 , RI2b5e78403c70_104, \2186 );
and \U$328 ( \2481 , RI2b5e775b1f50_117, \2188 );
and \U$329 ( \2482 , RI2b5e775b1938_130, \2190 );
and \U$330 ( \2483 , RI2b5e7750b8d0_143, \2192 );
and \U$331 ( \2484 , RI2b5e774ff0a8_156, \2194 );
and \U$332 ( \2485 , RI2b5e774f60c0_169, \2196 );
and \U$333 ( \2486 , RI2b5e774ea6a8_182, \2198 );
and \U$334 ( \2487 , RI2b5e774dde80_195, \2200 );
and \U$335 ( \2488 , RI2b5e774d4e98_208, \2202 );
and \U$336 ( \2489 , RI2b5e785f3dd8_221, \2204 );
and \U$337 ( \2490 , RI2b5e785eb1b0_234, \2206 );
and \U$338 ( \2491 , RI2b5e785da338_247, \2208 );
or \U$339 ( \2492 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 );
_DC r194c ( \2493_nR194c , \2492 , \2218 );
buf \U$340 ( \2494 , \2493_nR194c );
not \U$341 ( \2495 , \2494 );
or \U$342 ( \2496 , \2474 , \2495 );
and \U$343 ( \2497 , \2471 , \2496 );
and \U$344 ( \2498 , \2450 , \2496 );
or \U$345 ( \2499 , \2472 , \2497 , \2498 );
and \U$346 ( \2500 , \2446 , \2499 );
and \U$347 ( \2501 , \2425 , \2499 );
or \U$348 ( \2502 , \2447 , \2500 , \2501 );
and \U$349 ( \2503 , \2421 , \2502 );
and \U$350 ( \2504 , \2400 , \2502 );
or \U$351 ( \2505 , \2422 , \2503 , \2504 );
and \U$352 ( \2506 , \2396 , \2505 );
and \U$353 ( \2507 , \2375 , \2505 );
or \U$354 ( \2508 , \2397 , \2506 , \2507 );
and \U$355 ( \2509 , \2371 , \2508 );
and \U$356 ( \2510 , \2350 , \2508 );
or \U$357 ( \2511 , \2372 , \2509 , \2510 );
and \U$358 ( \2512 , \2346 , \2511 );
and \U$359 ( \2513 , \2325 , \2511 );
or \U$360 ( \2514 , \2347 , \2512 , \2513 );
and \U$361 ( \2515 , \2321 , \2514 );
and \U$362 ( \2516 , \2300 , \2514 );
or \U$363 ( \2517 , \2322 , \2515 , \2516 );
and \U$364 ( \2518 , \2296 , \2517 );
and \U$365 ( \2519 , \2275 , \2517 );
or \U$366 ( \2520 , \2297 , \2518 , \2519 );
and \U$367 ( \2521 , \2271 , \2520 );
and \U$368 ( \2522 , \2250 , \2520 );
or \U$369 ( \2523 , \2272 , \2521 , \2522 );
and \U$370 ( \2524 , \2246 , \2523 );
and \U$371 ( \2525 , \2225 , \2523 );
or \U$372 ( \2526 , \2247 , \2524 , \2525 );
xor \U$373 ( \2527 , \2222 , \2526 );
buf \U$374 ( \2528 , \2527 );
buf \U$375 ( \2529 , \2528 );
xor \U$376 ( \2530 , \2225 , \2246 );
xor \U$377 ( \2531 , \2530 , \2523 );
buf \U$378 ( \2532 , \2531 );
buf \U$379 ( \2533 , \2532 );
xor \U$380 ( \2534 , \2250 , \2271 );
xor \U$381 ( \2535 , \2534 , \2520 );
buf \U$382 ( \2536 , \2535 );
buf \U$383 ( \2537 , \2536 );
and \U$384 ( \2538 , \2533 , \2537 );
not \U$385 ( \2539 , \2538 );
and \U$386 ( \2540 , \2529 , \2539 );
not \U$387 ( \2541 , \2540 );
buf \U$388 ( \2542 , RI2b5e785ae9b8_600);
buf \U$389 ( \2543 , RI2b5e785aec10_595);
buf \U$390 ( \2544 , RI2b5e785aec88_594);
buf \U$391 ( \2545 , RI2b5e785aed00_593);
buf \U$392 ( \2546 , RI2b5e785aed78_592);
buf \U$393 ( \2547 , RI2b5e785aedf0_591);
buf \U$394 ( \2548 , RI2b5e785aee68_590);
buf \U$395 ( \2549 , RI2b5e785aeee0_589);
buf \U$396 ( \2550 , RI2b5e785aef58_588);
buf \U$397 ( \2551 , RI2b5e785aeb98_596);
nor \U$398 ( \2552 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 );
buf \U$399 ( \2553 , \2552 );
buf \U$400 ( \2554 , \2553 );
xor \U$401 ( \2555 , \2542 , \2554 );
buf \U$402 ( \2556 , \2555 );
buf \U$403 ( \2557 , RI2b5e785aea30_599);
and \U$404 ( \2558 , \2542 , \2554 );
xor \U$405 ( \2559 , \2557 , \2558 );
buf \U$406 ( \2560 , \2559 );
buf \U$407 ( \2561 , RI2b5e785aeaa8_598);
and \U$408 ( \2562 , \2557 , \2558 );
xor \U$409 ( \2563 , \2561 , \2562 );
buf \U$410 ( \2564 , \2563 );
buf \U$411 ( \2565 , RI2b5e785aeb20_597);
and \U$412 ( \2566 , \2561 , \2562 );
xor \U$413 ( \2567 , \2565 , \2566 );
buf \U$414 ( \2568 , \2567 );
buf \U$415 ( \2569 , RI2b5e785aeb98_596);
and \U$416 ( \2570 , \2565 , \2566 );
xor \U$417 ( \2571 , \2569 , \2570 );
buf \U$418 ( \2572 , \2571 );
not \U$419 ( \2573 , \2572 );
nor \U$420 ( \2574 , \2556 , \2560 , \2564 , \2568 , \2573 );
and \U$421 ( \2575 , RI2b5e785da248_249, \2574 );
and \U$422 ( \2576 , \2556 , \2560 , \2564 , \2568 , \2573 );
and \U$423 ( \2577 , RI2b5e785be750_269, \2576 );
not \U$424 ( \2578 , \2556 );
and \U$425 ( \2579 , \2578 , \2560 , \2564 , \2568 , \2573 );
and \U$426 ( \2580 , RI2b5e785bc4a0_289, \2579 );
not \U$427 ( \2581 , \2560 );
and \U$428 ( \2582 , \2556 , \2581 , \2564 , \2568 , \2573 );
and \U$429 ( \2583 , RI2b5e785bbb40_309, \2582 );
and \U$430 ( \2584 , \2578 , \2581 , \2564 , \2568 , \2573 );
and \U$431 ( \2585 , RI2b5e785b9c50_329, \2584 );
not \U$432 ( \2586 , \2564 );
and \U$433 ( \2587 , \2556 , \2560 , \2586 , \2568 , \2573 );
and \U$434 ( \2588 , RI2b5e785b8120_349, \2587 );
and \U$435 ( \2589 , \2578 , \2560 , \2586 , \2568 , \2573 );
and \U$436 ( \2590 , RI2b5e785b77c0_369, \2589 );
and \U$437 ( \2591 , \2556 , \2581 , \2586 , \2568 , \2573 );
and \U$438 ( \2592 , RI2b5e785b6e60_389, \2591 );
and \U$439 ( \2593 , \2578 , \2581 , \2586 , \2568 , \2573 );
and \U$440 ( \2594 , RI2b5e785b56f0_409, \2593 );
nor \U$441 ( \2595 , \2578 , \2581 , \2586 , \2568 , \2572 );
and \U$442 ( \2596 , RI2b5e785b4d90_429, \2595 );
nor \U$443 ( \2597 , \2556 , \2581 , \2586 , \2568 , \2572 );
and \U$444 ( \2598 , RI2b5e785b39e0_449, \2597 );
nor \U$445 ( \2599 , \2578 , \2560 , \2586 , \2568 , \2572 );
and \U$446 ( \2600 , RI2b5e785b3080_469, \2599 );
nor \U$447 ( \2601 , \2556 , \2560 , \2586 , \2568 , \2572 );
and \U$448 ( \2602 , RI2b5e785b2720_489, \2601 );
nor \U$449 ( \2603 , \2578 , \2581 , \2564 , \2568 , \2572 );
and \U$450 ( \2604 , RI2b5e785b1730_509, \2603 );
nor \U$451 ( \2605 , \2556 , \2581 , \2564 , \2568 , \2572 );
and \U$452 ( \2606 , RI2b5e785b0dd0_529, \2605 );
nor \U$453 ( \2607 , \2578 , \2560 , \2564 , \2568 , \2572 );
and \U$454 ( \2608 , RI2b5e785b0470_549, \2607 );
nor \U$455 ( \2609 , \2556 , \2560 , \2564 , \2568 , \2572 );
and \U$456 ( \2610 , RI2b5e785af840_569, \2609 );
or \U$457 ( \2611 , \2575 , \2577 , \2580 , \2583 , \2585 , \2588 , \2590 , \2592 , \2594 , \2596 , \2598 , \2600 , \2602 , \2604 , \2606 , \2608 , \2610 );
buf \U$458 ( \2612 , \2572 );
buf \U$459 ( \2613 , \2556 );
buf \U$460 ( \2614 , \2560 );
buf \U$461 ( \2615 , \2564 );
buf \U$462 ( \2616 , \2568 );
or \U$463 ( \2617 , \2613 , \2614 , \2615 , \2616 );
and \U$464 ( \2618 , \2612 , \2617 );
buf \U$465 ( \2619 , \2618 );
_DC r2749 ( \2620_nR2749 , \2611 , \2619 );
buf \U$466 ( \2621 , \2620_nR2749 );
buf \U$467 ( \2622 , RI2b5e785ebd68_1);
and \U$468 ( \2623 , \2149 , \2168 );
and \U$469 ( \2624 , \2622 , \2623 );
buf \U$470 ( \2625 , \2624 );
buf \U$471 ( \2626 , \2625 );
xor \U$472 ( \2627 , \2622 , \2623 );
buf \U$473 ( \2628 , \2627 );
buf \U$474 ( \2629 , \2628 );
and \U$475 ( \2630 , RI2b5e785daab8_27, \2173 );
and \U$476 ( \2631 , RI2b5e785495b8_40, \2175 );
and \U$477 ( \2632 , RI2b5e78538920_53, \2178 );
and \U$478 ( \2633 , RI2b5e784a63a8_66, \2181 );
and \U$479 ( \2634 , RI2b5e78495710_79, \2183 );
and \U$480 ( \2635 , RI2b5e784950f8_92, \2186 );
and \U$481 ( \2636 , RI2b5e78403bf8_105, \2188 );
and \U$482 ( \2637 , RI2b5e775b1ed8_118, \2190 );
and \U$483 ( \2638 , RI2b5e775b18c0_131, \2192 );
and \U$484 ( \2639 , RI2b5e7750b858_144, \2194 );
and \U$485 ( \2640 , RI2b5e774ff030_157, \2196 );
and \U$486 ( \2641 , RI2b5e774f6048_170, \2198 );
and \U$487 ( \2642 , RI2b5e774ea630_183, \2200 );
and \U$488 ( \2643 , RI2b5e774dde08_196, \2202 );
and \U$489 ( \2644 , RI2b5e774d4e20_209, \2204 );
and \U$490 ( \2645 , RI2b5e785f3d60_222, \2206 );
and \U$491 ( \2646 , RI2b5e785eb138_235, \2208 );
or \U$492 ( \2647 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 );
_DC r2211 ( \2648_nR2211 , \2647 , \2218 );
buf \U$493 ( \2649 , \2648_nR2211 );
not \U$494 ( \2650 , \2649 );
and \U$495 ( \2651 , \2629 , \2650 );
and \U$496 ( \2652 , \2171 , \2221 );
and \U$497 ( \2653 , \2221 , \2526 );
and \U$498 ( \2654 , \2171 , \2526 );
or \U$499 ( \2655 , \2652 , \2653 , \2654 );
and \U$500 ( \2656 , \2650 , \2655 );
and \U$501 ( \2657 , \2629 , \2655 );
or \U$502 ( \2658 , \2651 , \2656 , \2657 );
xnor \U$503 ( \2659 , \2626 , \2658 );
buf \U$504 ( \2660 , \2659 );
buf \U$505 ( \2661 , \2660 );
xor \U$506 ( \2662 , \2629 , \2650 );
xor \U$507 ( \2663 , \2662 , \2655 );
buf \U$508 ( \2664 , \2663 );
buf \U$509 ( \2665 , \2664 );
xor \U$510 ( \2666 , \2661 , \2665 );
xor \U$511 ( \2667 , \2665 , \2529 );
not \U$512 ( \2668 , \2667 );
and \U$513 ( \2669 , \2666 , \2668 );
and \U$514 ( \2670 , \2621 , \2669 );
and \U$515 ( \2671 , RI2b5e785da2c0_248, \2574 );
and \U$516 ( \2672 , RI2b5e785be7c8_268, \2576 );
and \U$517 ( \2673 , RI2b5e785bc518_288, \2579 );
and \U$518 ( \2674 , RI2b5e785bbbb8_308, \2582 );
and \U$519 ( \2675 , RI2b5e785b9cc8_328, \2584 );
and \U$520 ( \2676 , RI2b5e785b9368_348, \2587 );
and \U$521 ( \2677 , RI2b5e785b7838_368, \2589 );
and \U$522 ( \2678 , RI2b5e785b6ed8_388, \2591 );
and \U$523 ( \2679 , RI2b5e785b5768_408, \2593 );
and \U$524 ( \2680 , RI2b5e785b4e08_428, \2595 );
and \U$525 ( \2681 , RI2b5e785b3a58_448, \2597 );
and \U$526 ( \2682 , RI2b5e785b30f8_468, \2599 );
and \U$527 ( \2683 , RI2b5e785b2798_488, \2601 );
and \U$528 ( \2684 , RI2b5e785b17a8_508, \2603 );
and \U$529 ( \2685 , RI2b5e785b0e48_528, \2605 );
and \U$530 ( \2686 , RI2b5e785b04e8_548, \2607 );
and \U$531 ( \2687 , RI2b5e785afb88_568, \2609 );
or \U$532 ( \2688 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 );
_DC r283d ( \2689_nR283d , \2688 , \2619 );
buf \U$533 ( \2690 , \2689_nR283d );
and \U$534 ( \2691 , \2690 , \2667 );
nor \U$535 ( \2692 , \2670 , \2691 );
and \U$536 ( \2693 , \2665 , \2529 );
not \U$537 ( \2694 , \2693 );
and \U$538 ( \2695 , \2661 , \2694 );
xnor \U$539 ( \2696 , \2692 , \2695 );
xor \U$540 ( \2697 , \2541 , \2696 );
and \U$542 ( \2698 , RI2b5e785da1d0_250, \2574 );
and \U$543 ( \2699 , RI2b5e785be6d8_270, \2576 );
and \U$544 ( \2700 , RI2b5e785bc428_290, \2579 );
and \U$545 ( \2701 , RI2b5e785bbac8_310, \2582 );
and \U$546 ( \2702 , RI2b5e785b9bd8_330, \2584 );
and \U$547 ( \2703 , RI2b5e785b80a8_350, \2587 );
and \U$548 ( \2704 , RI2b5e785b7748_370, \2589 );
and \U$549 ( \2705 , RI2b5e785b6de8_390, \2591 );
and \U$550 ( \2706 , RI2b5e785b5678_410, \2593 );
and \U$551 ( \2707 , RI2b5e785b4d18_430, \2595 );
and \U$552 ( \2708 , RI2b5e785b3968_450, \2597 );
and \U$553 ( \2709 , RI2b5e785b3008_470, \2599 );
and \U$554 ( \2710 , RI2b5e785b26a8_490, \2601 );
and \U$555 ( \2711 , RI2b5e785b16b8_510, \2603 );
and \U$556 ( \2712 , RI2b5e785b0d58_530, \2605 );
and \U$557 ( \2713 , RI2b5e785b03f8_550, \2607 );
and \U$558 ( \2714 , RI2b5e785af7c8_570, \2609 );
or \U$559 ( \2715 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 );
_DC r2687 ( \2716_nR2687 , \2715 , \2619 );
buf \U$560 ( \2717 , \2716_nR2687 );
or \U$561 ( \2718 , \2626 , \2658 );
not \U$562 ( \2719 , \2718 );
buf \U$563 ( \2720 , \2719 );
buf \U$564 ( \2721 , \2720 );
xor \U$565 ( \2722 , \2721 , \2661 );
and \U$566 ( \2723 , \2717 , \2722 );
nor \U$567 ( \2724 , 1'b0 , \2723 );
xnor \U$569 ( \2725 , \2724 , 1'b0 );
xor \U$570 ( \2726 , \2697 , \2725 );
xor \U$571 ( \2727 , 1'b0 , \2726 );
xor \U$573 ( \2728 , \2529 , \2533 );
xor \U$574 ( \2729 , \2533 , \2537 );
not \U$575 ( \2730 , \2729 );
and \U$576 ( \2731 , \2728 , \2730 );
and \U$577 ( \2732 , \2690 , \2731 );
not \U$578 ( \2733 , \2732 );
xnor \U$579 ( \2734 , \2733 , \2540 );
and \U$580 ( \2735 , \2717 , \2669 );
and \U$581 ( \2736 , \2621 , \2667 );
nor \U$582 ( \2737 , \2735 , \2736 );
xnor \U$583 ( \2738 , \2737 , \2695 );
and \U$584 ( \2739 , \2734 , \2738 );
or \U$586 ( \2740 , 1'b0 , \2739 , 1'b0 );
xor \U$588 ( \2741 , \2740 , 1'b0 );
xor \U$590 ( \2742 , \2741 , 1'b0 );
and \U$591 ( \2743 , \2727 , \2742 );
or \U$592 ( \2744 , 1'b0 , 1'b0 , \2743 );
and \U$595 ( \2745 , \2690 , \2669 );
not \U$596 ( \2746 , \2745 );
xnor \U$597 ( \2747 , \2746 , \2695 );
xor \U$598 ( \2748 , 1'b0 , \2747 );
and \U$600 ( \2749 , \2621 , \2722 );
nor \U$601 ( \2750 , 1'b0 , \2749 );
xnor \U$602 ( \2751 , \2750 , 1'b0 );
xor \U$603 ( \2752 , \2748 , \2751 );
xor \U$604 ( \2753 , 1'b0 , \2752 );
xor \U$606 ( \2754 , \2753 , 1'b1 );
and \U$607 ( \2755 , \2541 , \2696 );
and \U$608 ( \2756 , \2696 , \2725 );
and \U$609 ( \2757 , \2541 , \2725 );
or \U$610 ( \2758 , \2755 , \2756 , \2757 );
xor \U$612 ( \2759 , \2758 , 1'b0 );
xor \U$614 ( \2760 , \2759 , 1'b0 );
xor \U$615 ( \2761 , \2754 , \2760 );
and \U$616 ( \2762 , \2744 , \2761 );
or \U$618 ( \2763 , 1'b0 , \2762 , 1'b0 );
xor \U$620 ( \2764 , \2763 , 1'b0 );
and \U$622 ( \2765 , \2753 , 1'b1 );
and \U$623 ( \2766 , 1'b1 , \2760 );
and \U$624 ( \2767 , \2753 , \2760 );
or \U$625 ( \2768 , \2765 , \2766 , \2767 );
xor \U$626 ( \2769 , 1'b0 , \2768 );
not \U$628 ( \2770 , \2695 );
and \U$630 ( \2771 , \2690 , \2722 );
nor \U$631 ( \2772 , 1'b0 , \2771 );
xnor \U$632 ( \2773 , \2772 , 1'b0 );
xor \U$633 ( \2774 , \2770 , \2773 );
xor \U$635 ( \2775 , \2774 , 1'b0 );
xor \U$636 ( \2776 , 1'b0 , \2775 );
xor \U$638 ( \2777 , \2776 , 1'b0 );
and \U$640 ( \2778 , \2747 , \2751 );
or \U$642 ( \2779 , 1'b0 , \2778 , 1'b0 );
xor \U$644 ( \2780 , \2779 , 1'b0 );
xor \U$646 ( \2781 , \2780 , 1'b0 );
xor \U$647 ( \2782 , \2777 , \2781 );
xor \U$648 ( \2783 , \2769 , \2782 );
xor \U$649 ( \2784 , \2764 , \2783 );
xor \U$655 ( \2785 , \2275 , \2296 );
xor \U$656 ( \2786 , \2785 , \2517 );
buf \U$657 ( \2787 , \2786 );
buf \U$658 ( \2788 , \2787 );
xor \U$659 ( \2789 , \2537 , \2788 );
xor \U$660 ( \2790 , \2300 , \2321 );
xor \U$661 ( \2791 , \2790 , \2514 );
buf \U$662 ( \2792 , \2791 );
buf \U$663 ( \2793 , \2792 );
xor \U$664 ( \2794 , \2788 , \2793 );
not \U$665 ( \2795 , \2794 );
and \U$666 ( \2796 , \2789 , \2795 );
and \U$667 ( \2797 , \2690 , \2796 );
not \U$668 ( \2798 , \2797 );
and \U$669 ( \2799 , \2788 , \2793 );
not \U$670 ( \2800 , \2799 );
and \U$671 ( \2801 , \2537 , \2800 );
xnor \U$672 ( \2802 , \2798 , \2801 );
and \U$673 ( \2803 , \2717 , \2731 );
and \U$674 ( \2804 , \2621 , \2729 );
nor \U$675 ( \2805 , \2803 , \2804 );
xnor \U$676 ( \2806 , \2805 , \2540 );
and \U$677 ( \2807 , \2802 , \2806 );
or \U$679 ( \2808 , 1'b0 , \2807 , 1'b0 );
and \U$680 ( \2809 , RI2b5e785da0e0_252, \2574 );
and \U$681 ( \2810 , RI2b5e785be5e8_272, \2576 );
and \U$682 ( \2811 , RI2b5e785bc338_292, \2579 );
and \U$683 ( \2812 , RI2b5e785bb9d8_312, \2582 );
and \U$684 ( \2813 , RI2b5e785b9ae8_332, \2584 );
and \U$685 ( \2814 , RI2b5e785b7fb8_352, \2587 );
and \U$686 ( \2815 , RI2b5e785b7658_372, \2589 );
and \U$687 ( \2816 , RI2b5e785b5ee8_392, \2591 );
and \U$688 ( \2817 , RI2b5e785b5588_412, \2593 );
and \U$689 ( \2818 , RI2b5e785b4c28_432, \2595 );
and \U$690 ( \2819 , RI2b5e785b3878_452, \2597 );
and \U$691 ( \2820 , RI2b5e785b2f18_472, \2599 );
and \U$692 ( \2821 , RI2b5e785b25b8_492, \2601 );
and \U$693 ( \2822 , RI2b5e785b15c8_512, \2603 );
and \U$694 ( \2823 , RI2b5e785b0c68_532, \2605 );
and \U$695 ( \2824 , RI2b5e785b0308_552, \2607 );
and \U$696 ( \2825 , RI2b5e785af6d8_572, \2609 );
or \U$697 ( \2826 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 );
_DC r24ec ( \2827_nR24ec , \2826 , \2619 );
buf \U$698 ( \2828 , \2827_nR24ec );
and \U$699 ( \2829 , \2828 , \2669 );
and \U$700 ( \2830 , RI2b5e785da158_251, \2574 );
and \U$701 ( \2831 , RI2b5e785be660_271, \2576 );
and \U$702 ( \2832 , RI2b5e785bc3b0_291, \2579 );
and \U$703 ( \2833 , RI2b5e785bba50_311, \2582 );
and \U$704 ( \2834 , RI2b5e785b9b60_331, \2584 );
and \U$705 ( \2835 , RI2b5e785b8030_351, \2587 );
and \U$706 ( \2836 , RI2b5e785b76d0_371, \2589 );
and \U$707 ( \2837 , RI2b5e785b6d70_391, \2591 );
and \U$708 ( \2838 , RI2b5e785b5600_411, \2593 );
and \U$709 ( \2839 , RI2b5e785b4ca0_431, \2595 );
and \U$710 ( \2840 , RI2b5e785b38f0_451, \2597 );
and \U$711 ( \2841 , RI2b5e785b2f90_471, \2599 );
and \U$712 ( \2842 , RI2b5e785b2630_491, \2601 );
and \U$713 ( \2843 , RI2b5e785b1640_511, \2603 );
and \U$714 ( \2844 , RI2b5e785b0ce0_531, \2605 );
and \U$715 ( \2845 , RI2b5e785b0380_551, \2607 );
and \U$716 ( \2846 , RI2b5e785af750_571, \2609 );
or \U$717 ( \2847 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 );
_DC r25c6 ( \2848_nR25c6 , \2847 , \2619 );
buf \U$718 ( \2849 , \2848_nR25c6 );
and \U$719 ( \2850 , \2849 , \2667 );
nor \U$720 ( \2851 , \2829 , \2850 );
xnor \U$721 ( \2852 , \2851 , \2695 );
and \U$723 ( \2853 , RI2b5e785da068_253, \2574 );
and \U$724 ( \2854 , RI2b5e785be570_273, \2576 );
and \U$725 ( \2855 , RI2b5e785bc2c0_293, \2579 );
and \U$726 ( \2856 , RI2b5e785bb960_313, \2582 );
and \U$727 ( \2857 , RI2b5e785b9a70_333, \2584 );
and \U$728 ( \2858 , RI2b5e785b7f40_353, \2587 );
and \U$729 ( \2859 , RI2b5e785b75e0_373, \2589 );
and \U$730 ( \2860 , RI2b5e785b5e70_393, \2591 );
and \U$731 ( \2861 , RI2b5e785b5510_413, \2593 );
and \U$732 ( \2862 , RI2b5e785b4bb0_433, \2595 );
and \U$733 ( \2863 , RI2b5e785b3800_453, \2597 );
and \U$734 ( \2864 , RI2b5e785b2ea0_473, \2599 );
and \U$735 ( \2865 , RI2b5e785b2540_493, \2601 );
and \U$736 ( \2866 , RI2b5e785b1550_513, \2603 );
and \U$737 ( \2867 , RI2b5e785b0bf0_533, \2605 );
and \U$738 ( \2868 , RI2b5e785b0290_553, \2607 );
and \U$739 ( \2869 , RI2b5e785af660_573, \2609 );
or \U$740 ( \2870 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 );
_DC r2401 ( \2871_nR2401 , \2870 , \2619 );
buf \U$741 ( \2872 , \2871_nR2401 );
and \U$742 ( \2873 , \2872 , \2722 );
nor \U$743 ( \2874 , 1'b0 , \2873 );
xnor \U$744 ( \2875 , \2874 , 1'b0 );
and \U$745 ( \2876 , \2852 , \2875 );
or \U$748 ( \2877 , \2876 , 1'b0 , 1'b0 );
and \U$749 ( \2878 , \2808 , \2877 );
or \U$752 ( \2879 , \2878 , 1'b0 , 1'b0 );
and \U$755 ( \2880 , \2828 , \2722 );
nor \U$756 ( \2881 , 1'b0 , \2880 );
xnor \U$757 ( \2882 , \2881 , 1'b0 );
xor \U$759 ( \2883 , \2882 , 1'b0 );
xor \U$761 ( \2884 , \2883 , 1'b0 );
not \U$762 ( \2885 , \2801 );
and \U$763 ( \2886 , \2621 , \2731 );
and \U$764 ( \2887 , \2690 , \2729 );
nor \U$765 ( \2888 , \2886 , \2887 );
xnor \U$766 ( \2889 , \2888 , \2540 );
xor \U$767 ( \2890 , \2885 , \2889 );
and \U$768 ( \2891 , \2849 , \2669 );
and \U$769 ( \2892 , \2717 , \2667 );
nor \U$770 ( \2893 , \2891 , \2892 );
xnor \U$771 ( \2894 , \2893 , \2695 );
xor \U$772 ( \2895 , \2890 , \2894 );
and \U$773 ( \2896 , \2884 , \2895 );
or \U$775 ( \2897 , 1'b0 , \2896 , 1'b0 );
and \U$776 ( \2898 , \2879 , \2897 );
or \U$777 ( \2899 , 1'b0 , 1'b0 , \2898 );
and \U$779 ( \2900 , \2849 , \2722 );
nor \U$780 ( \2901 , 1'b0 , \2900 );
xnor \U$781 ( \2902 , \2901 , 1'b0 );
xor \U$783 ( \2903 , \2902 , 1'b0 );
xor \U$785 ( \2904 , \2903 , 1'b0 );
xor \U$787 ( \2905 , 1'b0 , \2734 );
xor \U$788 ( \2906 , \2905 , \2738 );
xor \U$789 ( \2907 , \2904 , \2906 );
and \U$791 ( \2908 , \2907 , 1'b1 );
and \U$792 ( \2909 , \2885 , \2889 );
and \U$793 ( \2910 , \2889 , \2894 );
and \U$794 ( \2911 , \2885 , \2894 );
or \U$795 ( \2912 , \2909 , \2910 , \2911 );
xor \U$797 ( \2913 , \2912 , 1'b0 );
xor \U$799 ( \2914 , \2913 , 1'b0 );
and \U$800 ( \2915 , 1'b1 , \2914 );
and \U$801 ( \2916 , \2907 , \2914 );
or \U$802 ( \2917 , \2908 , \2915 , \2916 );
and \U$803 ( \2918 , \2899 , \2917 );
xor \U$805 ( \2919 , \2727 , 1'b0 );
xor \U$806 ( \2920 , \2919 , \2742 );
and \U$807 ( \2921 , \2917 , \2920 );
and \U$808 ( \2922 , \2899 , \2920 );
or \U$809 ( \2923 , \2918 , \2921 , \2922 );
xor \U$811 ( \2924 , 1'b0 , \2744 );
xor \U$812 ( \2925 , \2924 , \2761 );
and \U$813 ( \2926 , \2923 , \2925 );
or \U$814 ( \2927 , 1'b0 , 1'b0 , \2926 );
nand \U$815 ( \2928 , \2784 , \2927 );
nor \U$816 ( \2929 , \2784 , \2927 );
not \U$817 ( \2930 , \2929 );
nand \U$818 ( \2931 , \2928 , \2930 );
xor \U$819 ( \2932 , \2450 , \2471 );
xor \U$820 ( \2933 , \2932 , \2496 );
buf \U$821 ( \2934 , \2933 );
buf \U$822 ( \2935 , \2934 );
xor \U$823 ( \2936 , \2474 , \2494 );
buf \U$824 ( \2937 , \2936 );
buf \U$825 ( \2938 , \2937 );
xor \U$826 ( \2939 , \2935 , \2938 );
not \U$827 ( \2940 , \2938 );
and \U$828 ( \2941 , \2939 , \2940 );
and \U$829 ( \2942 , \2872 , \2941 );
and \U$830 ( \2943 , \2828 , \2938 );
nor \U$831 ( \2944 , \2942 , \2943 );
xnor \U$832 ( \2945 , \2944 , \2935 );
and \U$833 ( \2946 , RI2b5e785c2bc0_255, \2574 );
and \U$834 ( \2947 , RI2b5e785be480_275, \2576 );
and \U$835 ( \2948 , RI2b5e785bc1d0_295, \2579 );
and \U$836 ( \2949 , RI2b5e785ba2e0_315, \2582 );
and \U$837 ( \2950 , RI2b5e785b9980_335, \2584 );
and \U$838 ( \2951 , RI2b5e785b7e50_355, \2587 );
and \U$839 ( \2952 , RI2b5e785b74f0_375, \2589 );
and \U$840 ( \2953 , RI2b5e785b5d80_395, \2591 );
and \U$841 ( \2954 , RI2b5e785b5420_415, \2593 );
and \U$842 ( \2955 , RI2b5e785b4ac0_435, \2595 );
and \U$843 ( \2956 , RI2b5e785b3710_455, \2597 );
and \U$844 ( \2957 , RI2b5e785b2db0_475, \2599 );
and \U$845 ( \2958 , RI2b5e785b2450_495, \2601 );
and \U$846 ( \2959 , RI2b5e785b1460_515, \2603 );
and \U$847 ( \2960 , RI2b5e785b0b00_535, \2605 );
and \U$848 ( \2961 , RI2b5e785b01a0_555, \2607 );
and \U$849 ( \2962 , RI2b5e785af570_575, \2609 );
or \U$850 ( \2963 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 );
_DC r224e ( \2964_nR224e , \2963 , \2619 );
buf \U$851 ( \2965 , \2964_nR224e );
xor \U$852 ( \2966 , \2400 , \2421 );
xor \U$853 ( \2967 , \2966 , \2502 );
buf \U$854 ( \2968 , \2967 );
buf \U$855 ( \2969 , \2968 );
xor \U$856 ( \2970 , \2425 , \2446 );
xor \U$857 ( \2971 , \2970 , \2499 );
buf \U$858 ( \2972 , \2971 );
buf \U$859 ( \2973 , \2972 );
xor \U$860 ( \2974 , \2969 , \2973 );
xor \U$861 ( \2975 , \2973 , \2935 );
not \U$862 ( \2976 , \2975 );
and \U$863 ( \2977 , \2974 , \2976 );
and \U$864 ( \2978 , \2965 , \2977 );
and \U$865 ( \2979 , RI2b5e785c2c38_254, \2574 );
and \U$866 ( \2980 , RI2b5e785be4f8_274, \2576 );
and \U$867 ( \2981 , RI2b5e785bc248_294, \2579 );
and \U$868 ( \2982 , RI2b5e785ba358_314, \2582 );
and \U$869 ( \2983 , RI2b5e785b99f8_334, \2584 );
and \U$870 ( \2984 , RI2b5e785b7ec8_354, \2587 );
and \U$871 ( \2985 , RI2b5e785b7568_374, \2589 );
and \U$872 ( \2986 , RI2b5e785b5df8_394, \2591 );
and \U$873 ( \2987 , RI2b5e785b5498_414, \2593 );
and \U$874 ( \2988 , RI2b5e785b4b38_434, \2595 );
and \U$875 ( \2989 , RI2b5e785b3788_454, \2597 );
and \U$876 ( \2990 , RI2b5e785b2e28_474, \2599 );
and \U$877 ( \2991 , RI2b5e785b24c8_494, \2601 );
and \U$878 ( \2992 , RI2b5e785b14d8_514, \2603 );
and \U$879 ( \2993 , RI2b5e785b0b78_534, \2605 );
and \U$880 ( \2994 , RI2b5e785b0218_554, \2607 );
and \U$881 ( \2995 , RI2b5e785af5e8_574, \2609 );
or \U$882 ( \2996 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 );
_DC r2322 ( \2997_nR2322 , \2996 , \2619 );
buf \U$883 ( \2998 , \2997_nR2322 );
and \U$884 ( \2999 , \2998 , \2975 );
nor \U$885 ( \3000 , \2978 , \2999 );
and \U$886 ( \3001 , \2973 , \2935 );
not \U$887 ( \3002 , \3001 );
and \U$888 ( \3003 , \2969 , \3002 );
xnor \U$889 ( \3004 , \3000 , \3003 );
and \U$890 ( \3005 , \2945 , \3004 );
and \U$891 ( \3006 , RI2b5e785c0a00_257, \2574 );
and \U$892 ( \3007 , RI2b5e785be390_277, \2576 );
and \U$893 ( \3008 , RI2b5e785bc0e0_297, \2579 );
and \U$894 ( \3009 , RI2b5e785ba1f0_317, \2582 );
and \U$895 ( \3010 , RI2b5e785b9890_337, \2584 );
and \U$896 ( \3011 , RI2b5e785b7d60_357, \2587 );
and \U$897 ( \3012 , RI2b5e785b7400_377, \2589 );
and \U$898 ( \3013 , RI2b5e785b5c90_397, \2591 );
and \U$899 ( \3014 , RI2b5e785b5330_417, \2593 );
and \U$900 ( \3015 , RI2b5e785b49d0_437, \2595 );
and \U$901 ( \3016 , RI2b5e785b3620_457, \2597 );
and \U$902 ( \3017 , RI2b5e785b2cc0_477, \2599 );
and \U$903 ( \3018 , RI2b5e785b2360_497, \2601 );
and \U$904 ( \3019 , RI2b5e785b1370_517, \2603 );
and \U$905 ( \3020 , RI2b5e785b0a10_537, \2605 );
and \U$906 ( \3021 , RI2b5e785b00b0_557, \2607 );
and \U$907 ( \3022 , RI2b5e785af480_577, \2609 );
or \U$908 ( \3023 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 );
_DC r2081 ( \3024_nR2081 , \3023 , \2619 );
buf \U$909 ( \3025 , \3024_nR2081 );
xor \U$910 ( \3026 , \2350 , \2371 );
xor \U$911 ( \3027 , \3026 , \2508 );
buf \U$912 ( \3028 , \3027 );
buf \U$913 ( \3029 , \3028 );
xor \U$914 ( \3030 , \2375 , \2396 );
xor \U$915 ( \3031 , \3030 , \2505 );
buf \U$916 ( \3032 , \3031 );
buf \U$917 ( \3033 , \3032 );
xor \U$918 ( \3034 , \3029 , \3033 );
xor \U$919 ( \3035 , \3033 , \2969 );
not \U$920 ( \3036 , \3035 );
and \U$921 ( \3037 , \3034 , \3036 );
and \U$922 ( \3038 , \3025 , \3037 );
and \U$923 ( \3039 , RI2b5e785c2b48_256, \2574 );
and \U$924 ( \3040 , RI2b5e785be408_276, \2576 );
and \U$925 ( \3041 , RI2b5e785bc158_296, \2579 );
and \U$926 ( \3042 , RI2b5e785ba268_316, \2582 );
and \U$927 ( \3043 , RI2b5e785b9908_336, \2584 );
and \U$928 ( \3044 , RI2b5e785b7dd8_356, \2587 );
and \U$929 ( \3045 , RI2b5e785b7478_376, \2589 );
and \U$930 ( \3046 , RI2b5e785b5d08_396, \2591 );
and \U$931 ( \3047 , RI2b5e785b53a8_416, \2593 );
and \U$932 ( \3048 , RI2b5e785b4a48_436, \2595 );
and \U$933 ( \3049 , RI2b5e785b3698_456, \2597 );
and \U$934 ( \3050 , RI2b5e785b2d38_476, \2599 );
and \U$935 ( \3051 , RI2b5e785b23d8_496, \2601 );
and \U$936 ( \3052 , RI2b5e785b13e8_516, \2603 );
and \U$937 ( \3053 , RI2b5e785b0a88_536, \2605 );
and \U$938 ( \3054 , RI2b5e785b0128_556, \2607 );
and \U$939 ( \3055 , RI2b5e785af4f8_576, \2609 );
or \U$940 ( \3056 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 );
_DC r2158 ( \3057_nR2158 , \3056 , \2619 );
buf \U$941 ( \3058 , \3057_nR2158 );
and \U$942 ( \3059 , \3058 , \3035 );
nor \U$943 ( \3060 , \3038 , \3059 );
and \U$944 ( \3061 , \3033 , \2969 );
not \U$945 ( \3062 , \3061 );
and \U$946 ( \3063 , \3029 , \3062 );
xnor \U$947 ( \3064 , \3060 , \3063 );
and \U$948 ( \3065 , \3004 , \3064 );
and \U$949 ( \3066 , \2945 , \3064 );
or \U$950 ( \3067 , \3005 , \3065 , \3066 );
and \U$951 ( \3068 , RI2b5e785c0910_259, \2574 );
and \U$952 ( \3069 , RI2b5e785be2a0_279, \2576 );
and \U$953 ( \3070 , RI2b5e785bbff0_299, \2579 );
and \U$954 ( \3071 , RI2b5e785ba100_319, \2582 );
and \U$955 ( \3072 , RI2b5e785b97a0_339, \2584 );
and \U$956 ( \3073 , RI2b5e785b7c70_359, \2587 );
and \U$957 ( \3074 , RI2b5e785b7310_379, \2589 );
and \U$958 ( \3075 , RI2b5e785b5ba0_399, \2591 );
and \U$959 ( \3076 , RI2b5e785b5240_419, \2593 );
and \U$960 ( \3077 , RI2b5e785b48e0_439, \2595 );
and \U$961 ( \3078 , RI2b5e785b3530_459, \2597 );
and \U$962 ( \3079 , RI2b5e785b2bd0_479, \2599 );
and \U$963 ( \3080 , RI2b5e785b2270_499, \2601 );
and \U$964 ( \3081 , RI2b5e785b1280_519, \2603 );
and \U$965 ( \3082 , RI2b5e785b0920_539, \2605 );
and \U$966 ( \3083 , RI2b5e785affc0_559, \2607 );
and \U$967 ( \3084 , RI2b5e785af390_579, \2609 );
or \U$968 ( \3085 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 );
_DC r1ec2 ( \3086_nR1ec2 , \3085 , \2619 );
buf \U$969 ( \3087 , \3086_nR1ec2 );
xor \U$970 ( \3088 , \2325 , \2346 );
xor \U$971 ( \3089 , \3088 , \2511 );
buf \U$972 ( \3090 , \3089 );
buf \U$973 ( \3091 , \3090 );
xor \U$974 ( \3092 , \2793 , \3091 );
xor \U$975 ( \3093 , \3091 , \3029 );
not \U$976 ( \3094 , \3093 );
and \U$977 ( \3095 , \3092 , \3094 );
and \U$978 ( \3096 , \3087 , \3095 );
and \U$979 ( \3097 , RI2b5e785c0988_258, \2574 );
and \U$980 ( \3098 , RI2b5e785be318_278, \2576 );
and \U$981 ( \3099 , RI2b5e785bc068_298, \2579 );
and \U$982 ( \3100 , RI2b5e785ba178_318, \2582 );
and \U$983 ( \3101 , RI2b5e785b9818_338, \2584 );
and \U$984 ( \3102 , RI2b5e785b7ce8_358, \2587 );
and \U$985 ( \3103 , RI2b5e785b7388_378, \2589 );
and \U$986 ( \3104 , RI2b5e785b5c18_398, \2591 );
and \U$987 ( \3105 , RI2b5e785b52b8_418, \2593 );
and \U$988 ( \3106 , RI2b5e785b4958_438, \2595 );
and \U$989 ( \3107 , RI2b5e785b35a8_458, \2597 );
and \U$990 ( \3108 , RI2b5e785b2c48_478, \2599 );
and \U$991 ( \3109 , RI2b5e785b22e8_498, \2601 );
and \U$992 ( \3110 , RI2b5e785b12f8_518, \2603 );
and \U$993 ( \3111 , RI2b5e785b0998_538, \2605 );
and \U$994 ( \3112 , RI2b5e785b0038_558, \2607 );
and \U$995 ( \3113 , RI2b5e785af408_578, \2609 );
or \U$996 ( \3114 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 );
_DC r1f8b ( \3115_nR1f8b , \3114 , \2619 );
buf \U$997 ( \3116 , \3115_nR1f8b );
and \U$998 ( \3117 , \3116 , \3093 );
nor \U$999 ( \3118 , \3096 , \3117 );
and \U$1000 ( \3119 , \3091 , \3029 );
not \U$1001 ( \3120 , \3119 );
and \U$1002 ( \3121 , \2793 , \3120 );
xnor \U$1003 ( \3122 , \3118 , \3121 );
and \U$1004 ( \3123 , RI2b5e785c0820_261, \2574 );
and \U$1005 ( \3124 , RI2b5e785be1b0_281, \2576 );
and \U$1006 ( \3125 , RI2b5e785bbf00_301, \2579 );
and \U$1007 ( \3126 , RI2b5e785ba010_321, \2582 );
and \U$1008 ( \3127 , RI2b5e785b96b0_341, \2584 );
and \U$1009 ( \3128 , RI2b5e785b7b80_361, \2587 );
and \U$1010 ( \3129 , RI2b5e785b7220_381, \2589 );
and \U$1011 ( \3130 , RI2b5e785b5ab0_401, \2591 );
and \U$1012 ( \3131 , RI2b5e785b5150_421, \2593 );
and \U$1013 ( \3132 , RI2b5e785b47f0_441, \2595 );
and \U$1014 ( \3133 , RI2b5e785b3440_461, \2597 );
and \U$1015 ( \3134 , RI2b5e785b2ae0_481, \2599 );
and \U$1016 ( \3135 , RI2b5e785b2180_501, \2601 );
and \U$1017 ( \3136 , RI2b5e785b1190_521, \2603 );
and \U$1018 ( \3137 , RI2b5e785b0830_541, \2605 );
and \U$1019 ( \3138 , RI2b5e785afed0_561, \2607 );
and \U$1020 ( \3139 , RI2b5e785af2a0_581, \2609 );
or \U$1021 ( \3140 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 );
_DC r1d29 ( \3141_nR1d29 , \3140 , \2619 );
buf \U$1022 ( \3142 , \3141_nR1d29 );
and \U$1023 ( \3143 , \3142 , \2796 );
and \U$1024 ( \3144 , RI2b5e785c0898_260, \2574 );
and \U$1025 ( \3145 , RI2b5e785be228_280, \2576 );
and \U$1026 ( \3146 , RI2b5e785bbf78_300, \2579 );
and \U$1027 ( \3147 , RI2b5e785ba088_320, \2582 );
and \U$1028 ( \3148 , RI2b5e785b9728_340, \2584 );
and \U$1029 ( \3149 , RI2b5e785b7bf8_360, \2587 );
and \U$1030 ( \3150 , RI2b5e785b7298_380, \2589 );
and \U$1031 ( \3151 , RI2b5e785b5b28_400, \2591 );
and \U$1032 ( \3152 , RI2b5e785b51c8_420, \2593 );
and \U$1033 ( \3153 , RI2b5e785b4868_440, \2595 );
and \U$1034 ( \3154 , RI2b5e785b34b8_460, \2597 );
and \U$1035 ( \3155 , RI2b5e785b2b58_480, \2599 );
and \U$1036 ( \3156 , RI2b5e785b21f8_500, \2601 );
and \U$1037 ( \3157 , RI2b5e785b1208_520, \2603 );
and \U$1038 ( \3158 , RI2b5e785b08a8_540, \2605 );
and \U$1039 ( \3159 , RI2b5e785aff48_560, \2607 );
and \U$1040 ( \3160 , RI2b5e785af318_580, \2609 );
or \U$1041 ( \3161 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 );
_DC r1ddc ( \3162_nR1ddc , \3161 , \2619 );
buf \U$1042 ( \3163 , \3162_nR1ddc );
and \U$1043 ( \3164 , \3163 , \2794 );
nor \U$1044 ( \3165 , \3143 , \3164 );
xnor \U$1045 ( \3166 , \3165 , \2801 );
and \U$1046 ( \3167 , \3122 , \3166 );
and \U$1047 ( \3168 , RI2b5e785c0730_263, \2574 );
and \U$1048 ( \3169 , RI2b5e785be0c0_283, \2576 );
and \U$1049 ( \3170 , RI2b5e785bbe10_303, \2579 );
and \U$1050 ( \3171 , RI2b5e785b9f20_323, \2582 );
and \U$1051 ( \3172 , RI2b5e785b95c0_343, \2584 );
and \U$1052 ( \3173 , RI2b5e785b7a90_363, \2587 );
and \U$1053 ( \3174 , RI2b5e785b7130_383, \2589 );
and \U$1054 ( \3175 , RI2b5e785b59c0_403, \2591 );
and \U$1055 ( \3176 , RI2b5e785b5060_423, \2593 );
and \U$1056 ( \3177 , RI2b5e785b3cb0_443, \2595 );
and \U$1057 ( \3178 , RI2b5e785b3350_463, \2597 );
and \U$1058 ( \3179 , RI2b5e785b29f0_483, \2599 );
and \U$1059 ( \3180 , RI2b5e785b1a00_503, \2601 );
and \U$1060 ( \3181 , RI2b5e785b10a0_523, \2603 );
and \U$1061 ( \3182 , RI2b5e785b0740_543, \2605 );
and \U$1062 ( \3183 , RI2b5e785afde0_563, \2607 );
and \U$1063 ( \3184 , RI2b5e785af1b0_583, \2609 );
or \U$1064 ( \3185 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 );
_DC r1bc5 ( \3186_nR1bc5 , \3185 , \2619 );
buf \U$1065 ( \3187 , \3186_nR1bc5 );
and \U$1066 ( \3188 , \3187 , \2731 );
and \U$1067 ( \3189 , RI2b5e785c07a8_262, \2574 );
and \U$1068 ( \3190 , RI2b5e785be138_282, \2576 );
and \U$1069 ( \3191 , RI2b5e785bbe88_302, \2579 );
and \U$1070 ( \3192 , RI2b5e785b9f98_322, \2582 );
and \U$1071 ( \3193 , RI2b5e785b9638_342, \2584 );
and \U$1072 ( \3194 , RI2b5e785b7b08_362, \2587 );
and \U$1073 ( \3195 , RI2b5e785b71a8_382, \2589 );
and \U$1074 ( \3196 , RI2b5e785b5a38_402, \2591 );
and \U$1075 ( \3197 , RI2b5e785b50d8_422, \2593 );
and \U$1076 ( \3198 , RI2b5e785b4778_442, \2595 );
and \U$1077 ( \3199 , RI2b5e785b33c8_462, \2597 );
and \U$1078 ( \3200 , RI2b5e785b2a68_482, \2599 );
and \U$1079 ( \3201 , RI2b5e785b1a78_502, \2601 );
and \U$1080 ( \3202 , RI2b5e785b1118_522, \2603 );
and \U$1081 ( \3203 , RI2b5e785b07b8_542, \2605 );
and \U$1082 ( \3204 , RI2b5e785afe58_562, \2607 );
and \U$1083 ( \3205 , RI2b5e785af228_582, \2609 );
or \U$1084 ( \3206 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 );
_DC r1c6c ( \3207_nR1c6c , \3206 , \2619 );
buf \U$1085 ( \3208 , \3207_nR1c6c );
and \U$1086 ( \3209 , \3208 , \2729 );
nor \U$1087 ( \3210 , \3188 , \3209 );
xnor \U$1088 ( \3211 , \3210 , \2540 );
and \U$1089 ( \3212 , \3166 , \3211 );
and \U$1090 ( \3213 , \3122 , \3211 );
or \U$1091 ( \3214 , \3167 , \3212 , \3213 );
and \U$1092 ( \3215 , \3067 , \3214 );
and \U$1093 ( \3216 , RI2b5e785c0640_265, \2574 );
and \U$1094 ( \3217 , RI2b5e785bdfd0_285, \2576 );
and \U$1095 ( \3218 , RI2b5e785bbd20_305, \2579 );
and \U$1096 ( \3219 , RI2b5e785b9e30_325, \2582 );
and \U$1097 ( \3220 , RI2b5e785b94d0_345, \2584 );
and \U$1098 ( \3221 , RI2b5e785b79a0_365, \2587 );
and \U$1099 ( \3222 , RI2b5e785b7040_385, \2589 );
and \U$1100 ( \3223 , RI2b5e785b58d0_405, \2591 );
and \U$1101 ( \3224 , RI2b5e785b4f70_425, \2593 );
and \U$1102 ( \3225 , RI2b5e785b3bc0_445, \2595 );
and \U$1103 ( \3226 , RI2b5e785b3260_465, \2597 );
and \U$1104 ( \3227 , RI2b5e785b2900_485, \2599 );
and \U$1105 ( \3228 , RI2b5e785b1910_505, \2601 );
and \U$1106 ( \3229 , RI2b5e785b0fb0_525, \2603 );
and \U$1107 ( \3230 , RI2b5e785b0650_545, \2605 );
and \U$1108 ( \3231 , RI2b5e785afcf0_565, \2607 );
and \U$1109 ( \3232 , RI2b5e785af0c0_585, \2609 );
or \U$1110 ( \3233 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 );
_DC r1a55 ( \3234_nR1a55 , \3233 , \2619 );
buf \U$1111 ( \3235 , \3234_nR1a55 );
and \U$1112 ( \3236 , \3235 , \2669 );
and \U$1113 ( \3237 , RI2b5e785c06b8_264, \2574 );
and \U$1114 ( \3238 , RI2b5e785be048_284, \2576 );
and \U$1115 ( \3239 , RI2b5e785bbd98_304, \2579 );
and \U$1116 ( \3240 , RI2b5e785b9ea8_324, \2582 );
and \U$1117 ( \3241 , RI2b5e785b9548_344, \2584 );
and \U$1118 ( \3242 , RI2b5e785b7a18_364, \2587 );
and \U$1119 ( \3243 , RI2b5e785b70b8_384, \2589 );
and \U$1120 ( \3244 , RI2b5e785b5948_404, \2591 );
and \U$1121 ( \3245 , RI2b5e785b4fe8_424, \2593 );
and \U$1122 ( \3246 , RI2b5e785b3c38_444, \2595 );
and \U$1123 ( \3247 , RI2b5e785b32d8_464, \2597 );
and \U$1124 ( \3248 , RI2b5e785b2978_484, \2599 );
and \U$1125 ( \3249 , RI2b5e785b1988_504, \2601 );
and \U$1126 ( \3250 , RI2b5e785b1028_524, \2603 );
and \U$1127 ( \3251 , RI2b5e785b06c8_544, \2605 );
and \U$1128 ( \3252 , RI2b5e785afd68_564, \2607 );
and \U$1129 ( \3253 , RI2b5e785af138_584, \2609 );
or \U$1130 ( \3254 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 );
_DC r1b26 ( \3255_nR1b26 , \3254 , \2619 );
buf \U$1131 ( \3256 , \3255_nR1b26 );
and \U$1132 ( \3257 , \3256 , \2667 );
nor \U$1133 ( \3258 , \3236 , \3257 );
xnor \U$1134 ( \3259 , \3258 , \2695 );
and \U$1136 ( \3260 , RI2b5e785c05c8_266, \2574 );
and \U$1137 ( \3261 , RI2b5e785bdf58_286, \2576 );
and \U$1138 ( \3262 , RI2b5e785bbca8_306, \2579 );
and \U$1139 ( \3263 , RI2b5e785b9db8_326, \2582 );
and \U$1140 ( \3264 , RI2b5e785b9458_346, \2584 );
and \U$1141 ( \3265 , RI2b5e785b7928_366, \2587 );
and \U$1142 ( \3266 , RI2b5e785b6fc8_386, \2589 );
and \U$1143 ( \3267 , RI2b5e785b5858_406, \2591 );
and \U$1144 ( \3268 , RI2b5e785b4ef8_426, \2593 );
and \U$1145 ( \3269 , RI2b5e785b3b48_446, \2595 );
and \U$1146 ( \3270 , RI2b5e785b31e8_466, \2597 );
and \U$1147 ( \3271 , RI2b5e785b2888_486, \2599 );
and \U$1148 ( \3272 , RI2b5e785b1898_506, \2601 );
and \U$1149 ( \3273 , RI2b5e785b0f38_526, \2603 );
and \U$1150 ( \3274 , RI2b5e785b05d8_546, \2605 );
and \U$1151 ( \3275 , RI2b5e785afc78_566, \2607 );
and \U$1152 ( \3276 , RI2b5e785af048_586, \2609 );
or \U$1153 ( \3277 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 );
_DC r1a13 ( \3278_nR1a13 , \3277 , \2619 );
buf \U$1154 ( \3279 , \3278_nR1a13 );
and \U$1155 ( \3280 , \3279 , \2722 );
nor \U$1156 ( \3281 , 1'b0 , \3280 );
xnor \U$1157 ( \3282 , \3281 , 1'b0 );
and \U$1158 ( \3283 , \3259 , \3282 );
and \U$1159 ( \3284 , \3214 , \3283 );
and \U$1160 ( \3285 , \3067 , \3283 );
or \U$1161 ( \3286 , \3215 , \3284 , \3285 );
and \U$1163 ( \3287 , \3208 , \2731 );
and \U$1164 ( \3288 , \3142 , \2729 );
nor \U$1165 ( \3289 , \3287 , \3288 );
xnor \U$1166 ( \3290 , \3289 , \2540 );
and \U$1167 ( \3291 , \3256 , \2669 );
and \U$1168 ( \3292 , \3187 , \2667 );
nor \U$1169 ( \3293 , \3291 , \3292 );
xnor \U$1170 ( \3294 , \3293 , \2695 );
xor \U$1171 ( \3295 , \3290 , \3294 );
and \U$1173 ( \3296 , \3235 , \2722 );
nor \U$1174 ( \3297 , 1'b0 , \3296 );
xnor \U$1175 ( \3298 , \3297 , 1'b0 );
xor \U$1176 ( \3299 , \3295 , \3298 );
and \U$1177 ( \3300 , \3058 , \3037 );
and \U$1178 ( \3301 , \2965 , \3035 );
nor \U$1179 ( \3302 , \3300 , \3301 );
xnor \U$1180 ( \3303 , \3302 , \3063 );
and \U$1181 ( \3304 , \3116 , \3095 );
and \U$1182 ( \3305 , \3025 , \3093 );
nor \U$1183 ( \3306 , \3304 , \3305 );
xnor \U$1184 ( \3307 , \3306 , \3121 );
xor \U$1185 ( \3308 , \3303 , \3307 );
and \U$1186 ( \3309 , \3163 , \2796 );
and \U$1187 ( \3310 , \3087 , \2794 );
nor \U$1188 ( \3311 , \3309 , \3310 );
xnor \U$1189 ( \3312 , \3311 , \2801 );
xor \U$1190 ( \3313 , \3308 , \3312 );
and \U$1191 ( \3314 , \3299 , \3313 );
or \U$1193 ( \3315 , 1'b0 , \3314 , 1'b0 );
xor \U$1194 ( \3316 , \3286 , \3315 );
and \U$1195 ( \3317 , \3187 , \2669 );
and \U$1196 ( \3318 , \3208 , \2667 );
nor \U$1197 ( \3319 , \3317 , \3318 );
xnor \U$1198 ( \3320 , \3319 , \2695 );
and \U$1200 ( \3321 , \3256 , \2722 );
nor \U$1201 ( \3322 , 1'b0 , \3321 );
xnor \U$1202 ( \3323 , \3322 , 1'b0 );
xor \U$1203 ( \3324 , \3320 , \3323 );
xor \U$1205 ( \3325 , \3324 , 1'b0 );
and \U$1206 ( \3326 , \3025 , \3095 );
and \U$1207 ( \3327 , \3058 , \3093 );
nor \U$1208 ( \3328 , \3326 , \3327 );
xnor \U$1209 ( \3329 , \3328 , \3121 );
and \U$1210 ( \3330 , \3087 , \2796 );
and \U$1211 ( \3331 , \3116 , \2794 );
nor \U$1212 ( \3332 , \3330 , \3331 );
xnor \U$1213 ( \3333 , \3332 , \2801 );
xor \U$1214 ( \3334 , \3329 , \3333 );
and \U$1215 ( \3335 , \3142 , \2731 );
and \U$1216 ( \3336 , \3163 , \2729 );
nor \U$1217 ( \3337 , \3335 , \3336 );
xnor \U$1218 ( \3338 , \3337 , \2540 );
xor \U$1219 ( \3339 , \3334 , \3338 );
xor \U$1220 ( \3340 , \3325 , \3339 );
and \U$1221 ( \3341 , \2849 , \2941 );
and \U$1222 ( \3342 , \2717 , \2938 );
nor \U$1223 ( \3343 , \3341 , \3342 );
xnor \U$1224 ( \3344 , \3343 , \2935 );
and \U$1225 ( \3345 , \2872 , \2977 );
and \U$1226 ( \3346 , \2828 , \2975 );
nor \U$1227 ( \3347 , \3345 , \3346 );
xnor \U$1228 ( \3348 , \3347 , \3003 );
xor \U$1229 ( \3349 , \3344 , \3348 );
and \U$1230 ( \3350 , \2965 , \3037 );
and \U$1231 ( \3351 , \2998 , \3035 );
nor \U$1232 ( \3352 , \3350 , \3351 );
xnor \U$1233 ( \3353 , \3352 , \3063 );
xor \U$1234 ( \3354 , \3349 , \3353 );
xor \U$1235 ( \3355 , \3340 , \3354 );
xor \U$1236 ( \3356 , \3316 , \3355 );
and \U$1238 ( \3357 , \2998 , \2941 );
and \U$1239 ( \3358 , \2872 , \2938 );
nor \U$1240 ( \3359 , \3357 , \3358 );
xnor \U$1241 ( \3360 , \3359 , \2935 );
and \U$1242 ( \3361 , \3058 , \2977 );
and \U$1243 ( \3362 , \2965 , \2975 );
nor \U$1244 ( \3363 , \3361 , \3362 );
xnor \U$1245 ( \3364 , \3363 , \3003 );
and \U$1246 ( \3365 , \3360 , \3364 );
or \U$1248 ( \3366 , 1'b0 , \3365 , 1'b0 );
and \U$1249 ( \3367 , \3116 , \3037 );
and \U$1250 ( \3368 , \3025 , \3035 );
nor \U$1251 ( \3369 , \3367 , \3368 );
xnor \U$1252 ( \3370 , \3369 , \3063 );
and \U$1253 ( \3371 , \3163 , \3095 );
and \U$1254 ( \3372 , \3087 , \3093 );
nor \U$1255 ( \3373 , \3371 , \3372 );
xnor \U$1256 ( \3374 , \3373 , \3121 );
and \U$1257 ( \3375 , \3370 , \3374 );
and \U$1258 ( \3376 , \3208 , \2796 );
and \U$1259 ( \3377 , \3142 , \2794 );
nor \U$1260 ( \3378 , \3376 , \3377 );
xnor \U$1261 ( \3379 , \3378 , \2801 );
and \U$1262 ( \3380 , \3374 , \3379 );
and \U$1263 ( \3381 , \3370 , \3379 );
or \U$1264 ( \3382 , \3375 , \3380 , \3381 );
and \U$1265 ( \3383 , \3366 , \3382 );
and \U$1266 ( \3384 , \3256 , \2731 );
and \U$1267 ( \3385 , \3187 , \2729 );
nor \U$1268 ( \3386 , \3384 , \3385 );
xnor \U$1269 ( \3387 , \3386 , \2540 );
and \U$1270 ( \3388 , \3279 , \2669 );
and \U$1271 ( \3389 , \3235 , \2667 );
nor \U$1272 ( \3390 , \3388 , \3389 );
xnor \U$1273 ( \3391 , \3390 , \2695 );
and \U$1274 ( \3392 , \3387 , \3391 );
and \U$1275 ( \3393 , RI2b5e785c0550_267, \2574 );
and \U$1276 ( \3394 , RI2b5e785bc590_287, \2576 );
and \U$1277 ( \3395 , RI2b5e785bbc30_307, \2579 );
and \U$1278 ( \3396 , RI2b5e785b9d40_327, \2582 );
and \U$1279 ( \3397 , RI2b5e785b93e0_347, \2584 );
and \U$1280 ( \3398 , RI2b5e785b78b0_367, \2587 );
and \U$1281 ( \3399 , RI2b5e785b6f50_387, \2589 );
and \U$1282 ( \3400 , RI2b5e785b57e0_407, \2591 );
and \U$1283 ( \3401 , RI2b5e785b4e80_427, \2593 );
and \U$1284 ( \3402 , RI2b5e785b3ad0_447, \2595 );
and \U$1285 ( \3403 , RI2b5e785b3170_467, \2597 );
and \U$1286 ( \3404 , RI2b5e785b2810_487, \2599 );
and \U$1287 ( \3405 , RI2b5e785b1820_507, \2601 );
and \U$1288 ( \3406 , RI2b5e785b0ec0_527, \2603 );
and \U$1289 ( \3407 , RI2b5e785b0560_547, \2605 );
and \U$1290 ( \3408 , RI2b5e785afc00_567, \2607 );
and \U$1291 ( \3409 , RI2b5e785aefd0_587, \2609 );
or \U$1292 ( \3410 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 );
_DC r191b ( \3411_nR191b , \3410 , \2619 );
buf \U$1293 ( \3412 , \3411_nR191b );
nand \U$1294 ( \3413 , \3412 , \2722 );
xnor \U$1295 ( \3414 , \3413 , 1'b0 );
and \U$1296 ( \3415 , \3391 , \3414 );
and \U$1297 ( \3416 , \3387 , \3414 );
or \U$1298 ( \3417 , \3392 , \3415 , \3416 );
and \U$1299 ( \3418 , \3382 , \3417 );
and \U$1300 ( \3419 , \3366 , \3417 );
or \U$1301 ( \3420 , \3383 , \3418 , \3419 );
xor \U$1302 ( \3421 , \3259 , \3282 );
xor \U$1303 ( \3422 , \3122 , \3166 );
xor \U$1304 ( \3423 , \3422 , \3211 );
and \U$1305 ( \3424 , \3421 , \3423 );
xor \U$1306 ( \3425 , \2945 , \3004 );
xor \U$1307 ( \3426 , \3425 , \3064 );
and \U$1308 ( \3427 , \3423 , \3426 );
and \U$1309 ( \3428 , \3421 , \3426 );
or \U$1310 ( \3429 , \3424 , \3427 , \3428 );
and \U$1311 ( \3430 , \3420 , \3429 );
and \U$1313 ( \3431 , \2828 , \2941 );
and \U$1314 ( \3432 , \2849 , \2938 );
nor \U$1315 ( \3433 , \3431 , \3432 );
xnor \U$1316 ( \3434 , \3433 , \2935 );
xor \U$1317 ( \3435 , 1'b0 , \3434 );
and \U$1318 ( \3436 , \2998 , \2977 );
and \U$1319 ( \3437 , \2872 , \2975 );
nor \U$1320 ( \3438 , \3436 , \3437 );
xnor \U$1321 ( \3439 , \3438 , \3003 );
xor \U$1322 ( \3440 , \3435 , \3439 );
and \U$1323 ( \3441 , \3429 , \3440 );
and \U$1324 ( \3442 , \3420 , \3440 );
or \U$1325 ( \3443 , \3430 , \3441 , \3442 );
xor \U$1327 ( \3444 , 1'b0 , \3299 );
xor \U$1328 ( \3445 , \3444 , \3313 );
xor \U$1329 ( \3446 , \3067 , \3214 );
xor \U$1330 ( \3447 , \3446 , \3283 );
and \U$1331 ( \3448 , \3445 , \3447 );
xor \U$1332 ( \3449 , \3443 , \3448 );
and \U$1334 ( \3450 , \3434 , \3439 );
or \U$1336 ( \3451 , 1'b0 , \3450 , 1'b0 );
and \U$1337 ( \3452 , \3303 , \3307 );
and \U$1338 ( \3453 , \3307 , \3312 );
and \U$1339 ( \3454 , \3303 , \3312 );
or \U$1340 ( \3455 , \3452 , \3453 , \3454 );
xor \U$1341 ( \3456 , \3451 , \3455 );
and \U$1342 ( \3457 , \3290 , \3294 );
and \U$1343 ( \3458 , \3294 , \3298 );
and \U$1344 ( \3459 , \3290 , \3298 );
or \U$1345 ( \3460 , \3457 , \3458 , \3459 );
xor \U$1346 ( \3461 , \3456 , \3460 );
xor \U$1347 ( \3462 , \3449 , \3461 );
xor \U$1348 ( \3463 , \3356 , \3462 );
and \U$1349 ( \3464 , \2965 , \2941 );
and \U$1350 ( \3465 , \2998 , \2938 );
nor \U$1351 ( \3466 , \3464 , \3465 );
xnor \U$1352 ( \3467 , \3466 , \2935 );
and \U$1353 ( \3468 , \3025 , \2977 );
and \U$1354 ( \3469 , \3058 , \2975 );
nor \U$1355 ( \3470 , \3468 , \3469 );
xnor \U$1356 ( \3471 , \3470 , \3003 );
and \U$1357 ( \3472 , \3467 , \3471 );
and \U$1358 ( \3473 , \3087 , \3037 );
and \U$1359 ( \3474 , \3116 , \3035 );
nor \U$1360 ( \3475 , \3473 , \3474 );
xnor \U$1361 ( \3476 , \3475 , \3063 );
and \U$1362 ( \3477 , \3471 , \3476 );
and \U$1363 ( \3478 , \3467 , \3476 );
or \U$1364 ( \3479 , \3472 , \3477 , \3478 );
and \U$1365 ( \3480 , \3142 , \3095 );
and \U$1366 ( \3481 , \3163 , \3093 );
nor \U$1367 ( \3482 , \3480 , \3481 );
xnor \U$1368 ( \3483 , \3482 , \3121 );
and \U$1369 ( \3484 , \3187 , \2796 );
and \U$1370 ( \3485 , \3208 , \2794 );
nor \U$1371 ( \3486 , \3484 , \3485 );
xnor \U$1372 ( \3487 , \3486 , \2801 );
and \U$1373 ( \3488 , \3483 , \3487 );
and \U$1374 ( \3489 , \3235 , \2731 );
and \U$1375 ( \3490 , \3256 , \2729 );
nor \U$1376 ( \3491 , \3489 , \3490 );
xnor \U$1377 ( \3492 , \3491 , \2540 );
and \U$1378 ( \3493 , \3487 , \3492 );
and \U$1379 ( \3494 , \3483 , \3492 );
or \U$1380 ( \3495 , \3488 , \3493 , \3494 );
and \U$1381 ( \3496 , \3479 , \3495 );
xor \U$1382 ( \3497 , \3387 , \3391 );
xor \U$1383 ( \3498 , \3497 , \3414 );
and \U$1384 ( \3499 , \3495 , \3498 );
and \U$1385 ( \3500 , \3479 , \3498 );
or \U$1386 ( \3501 , \3496 , \3499 , \3500 );
xor \U$1387 ( \3502 , \3370 , \3374 );
xor \U$1388 ( \3503 , \3502 , \3379 );
xor \U$1389 ( \3504 , 1'b0 , \3360 );
xor \U$1390 ( \3505 , \3504 , \3364 );
and \U$1391 ( \3506 , \3503 , \3505 );
and \U$1392 ( \3507 , \3501 , \3506 );
xor \U$1393 ( \3508 , \3421 , \3423 );
xor \U$1394 ( \3509 , \3508 , \3426 );
and \U$1395 ( \3510 , \3506 , \3509 );
and \U$1396 ( \3511 , \3501 , \3509 );
or \U$1397 ( \3512 , \3507 , \3510 , \3511 );
xor \U$1398 ( \3513 , \3445 , \3447 );
and \U$1399 ( \3514 , \3512 , \3513 );
xor \U$1400 ( \3515 , \3420 , \3429 );
xor \U$1401 ( \3516 , \3515 , \3440 );
and \U$1402 ( \3517 , \3513 , \3516 );
and \U$1403 ( \3518 , \3512 , \3516 );
or \U$1404 ( \3519 , \3514 , \3517 , \3518 );
nor \U$1405 ( \3520 , \3463 , \3519 );
and \U$1406 ( \3521 , \3443 , \3448 );
and \U$1407 ( \3522 , \3448 , \3461 );
and \U$1408 ( \3523 , \3443 , \3461 );
or \U$1409 ( \3524 , \3521 , \3522 , \3523 );
and \U$1410 ( \3525 , \3286 , \3315 );
and \U$1411 ( \3526 , \3315 , \3355 );
and \U$1412 ( \3527 , \3286 , \3355 );
or \U$1413 ( \3528 , \3525 , \3526 , \3527 );
and \U$1415 ( \3529 , \2717 , \2941 );
and \U$1416 ( \3530 , \2621 , \2938 );
nor \U$1417 ( \3531 , \3529 , \3530 );
xnor \U$1418 ( \3532 , \3531 , \2935 );
xor \U$1419 ( \3533 , 1'b0 , \3532 );
and \U$1420 ( \3534 , \2828 , \2977 );
and \U$1421 ( \3535 , \2849 , \2975 );
nor \U$1422 ( \3536 , \3534 , \3535 );
xnor \U$1423 ( \3537 , \3536 , \3003 );
xor \U$1424 ( \3538 , \3533 , \3537 );
and \U$1426 ( \3539 , \3163 , \2731 );
and \U$1427 ( \3540 , \3087 , \2729 );
nor \U$1428 ( \3541 , \3539 , \3540 );
xnor \U$1429 ( \3542 , \3541 , \2540 );
and \U$1430 ( \3543 , \3208 , \2669 );
and \U$1431 ( \3544 , \3142 , \2667 );
nor \U$1432 ( \3545 , \3543 , \3544 );
xnor \U$1433 ( \3546 , \3545 , \2695 );
xor \U$1434 ( \3547 , \3542 , \3546 );
and \U$1436 ( \3548 , \3187 , \2722 );
nor \U$1437 ( \3549 , 1'b0 , \3548 );
xnor \U$1438 ( \3550 , \3549 , 1'b0 );
xor \U$1439 ( \3551 , \3547 , \3550 );
xor \U$1440 ( \3552 , 1'b0 , \3551 );
xor \U$1441 ( \3553 , \3538 , \3552 );
and \U$1442 ( \3554 , \3344 , \3348 );
and \U$1443 ( \3555 , \3348 , \3353 );
and \U$1444 ( \3556 , \3344 , \3353 );
or \U$1445 ( \3557 , \3554 , \3555 , \3556 );
and \U$1446 ( \3558 , \3329 , \3333 );
and \U$1447 ( \3559 , \3333 , \3338 );
and \U$1448 ( \3560 , \3329 , \3338 );
or \U$1449 ( \3561 , \3558 , \3559 , \3560 );
xor \U$1450 ( \3562 , \3557 , \3561 );
and \U$1451 ( \3563 , \3320 , \3323 );
or \U$1454 ( \3564 , \3563 , 1'b0 , 1'b0 );
xor \U$1455 ( \3565 , \3562 , \3564 );
xor \U$1456 ( \3566 , \3553 , \3565 );
xor \U$1457 ( \3567 , \3528 , \3566 );
and \U$1458 ( \3568 , \3451 , \3455 );
and \U$1459 ( \3569 , \3455 , \3460 );
and \U$1460 ( \3570 , \3451 , \3460 );
or \U$1461 ( \3571 , \3568 , \3569 , \3570 );
and \U$1462 ( \3572 , \3325 , \3339 );
and \U$1463 ( \3573 , \3339 , \3354 );
and \U$1464 ( \3574 , \3325 , \3354 );
or \U$1465 ( \3575 , \3572 , \3573 , \3574 );
xor \U$1466 ( \3576 , \3571 , \3575 );
and \U$1467 ( \3577 , \2998 , \3037 );
and \U$1468 ( \3578 , \2872 , \3035 );
nor \U$1469 ( \3579 , \3577 , \3578 );
xnor \U$1470 ( \3580 , \3579 , \3063 );
and \U$1471 ( \3581 , \3058 , \3095 );
and \U$1472 ( \3582 , \2965 , \3093 );
nor \U$1473 ( \3583 , \3581 , \3582 );
xnor \U$1474 ( \3584 , \3583 , \3121 );
xor \U$1475 ( \3585 , \3580 , \3584 );
and \U$1476 ( \3586 , \3116 , \2796 );
and \U$1477 ( \3587 , \3025 , \2794 );
nor \U$1478 ( \3588 , \3586 , \3587 );
xnor \U$1479 ( \3589 , \3588 , \2801 );
xor \U$1480 ( \3590 , \3585 , \3589 );
xor \U$1481 ( \3591 , \3576 , \3590 );
xor \U$1482 ( \3592 , \3567 , \3591 );
xor \U$1483 ( \3593 , \3524 , \3592 );
and \U$1484 ( \3594 , \3356 , \3462 );
nor \U$1485 ( \3595 , \3593 , \3594 );
nor \U$1486 ( \3596 , \3520 , \3595 );
and \U$1487 ( \3597 , \3528 , \3566 );
and \U$1488 ( \3598 , \3566 , \3591 );
and \U$1489 ( \3599 , \3528 , \3591 );
or \U$1490 ( \3600 , \3597 , \3598 , \3599 );
and \U$1492 ( \3601 , \3532 , \3537 );
or \U$1494 ( \3602 , 1'b0 , \3601 , 1'b0 );
and \U$1495 ( \3603 , \3580 , \3584 );
and \U$1496 ( \3604 , \3584 , \3589 );
and \U$1497 ( \3605 , \3580 , \3589 );
or \U$1498 ( \3606 , \3603 , \3604 , \3605 );
xor \U$1499 ( \3607 , \3602 , \3606 );
and \U$1500 ( \3608 , \3542 , \3546 );
and \U$1501 ( \3609 , \3546 , \3550 );
and \U$1502 ( \3610 , \3542 , \3550 );
or \U$1503 ( \3611 , \3608 , \3609 , \3610 );
xor \U$1504 ( \3612 , \3607 , \3611 );
and \U$1505 ( \3613 , \3557 , \3561 );
and \U$1506 ( \3614 , \3561 , \3564 );
and \U$1507 ( \3615 , \3557 , \3564 );
or \U$1508 ( \3616 , \3613 , \3614 , \3615 );
xor \U$1510 ( \3617 , \3616 , 1'b0 );
and \U$1511 ( \3618 , \2621 , \2941 );
and \U$1512 ( \3619 , \2690 , \2938 );
nor \U$1513 ( \3620 , \3618 , \3619 );
xnor \U$1514 ( \3621 , \3620 , \2935 );
and \U$1515 ( \3622 , \2849 , \2977 );
and \U$1516 ( \3623 , \2717 , \2975 );
nor \U$1517 ( \3624 , \3622 , \3623 );
xnor \U$1518 ( \3625 , \3624 , \3003 );
xor \U$1519 ( \3626 , \3621 , \3625 );
and \U$1520 ( \3627 , \2872 , \3037 );
and \U$1521 ( \3628 , \2828 , \3035 );
nor \U$1522 ( \3629 , \3627 , \3628 );
xnor \U$1523 ( \3630 , \3629 , \3063 );
xor \U$1524 ( \3631 , \3626 , \3630 );
xor \U$1525 ( \3632 , \3617 , \3631 );
xor \U$1526 ( \3633 , \3612 , \3632 );
xor \U$1527 ( \3634 , \3600 , \3633 );
and \U$1528 ( \3635 , \3571 , \3575 );
and \U$1529 ( \3636 , \3575 , \3590 );
and \U$1530 ( \3637 , \3571 , \3590 );
or \U$1531 ( \3638 , \3635 , \3636 , \3637 );
and \U$1532 ( \3639 , \3538 , \3552 );
and \U$1533 ( \3640 , \3552 , \3565 );
and \U$1534 ( \3641 , \3538 , \3565 );
or \U$1535 ( \3642 , \3639 , \3640 , \3641 );
xor \U$1536 ( \3643 , \3638 , \3642 );
and \U$1538 ( \3644 , \3142 , \2669 );
and \U$1539 ( \3645 , \3163 , \2667 );
nor \U$1540 ( \3646 , \3644 , \3645 );
xnor \U$1541 ( \3647 , \3646 , \2695 );
and \U$1543 ( \3648 , \3208 , \2722 );
nor \U$1544 ( \3649 , 1'b0 , \3648 );
xnor \U$1545 ( \3650 , \3649 , 1'b0 );
xor \U$1546 ( \3651 , \3647 , \3650 );
xor \U$1548 ( \3652 , \3651 , 1'b0 );
xor \U$1549 ( \3653 , 1'b0 , \3652 );
and \U$1550 ( \3654 , \2965 , \3095 );
and \U$1551 ( \3655 , \2998 , \3093 );
nor \U$1552 ( \3656 , \3654 , \3655 );
xnor \U$1553 ( \3657 , \3656 , \3121 );
and \U$1554 ( \3658 , \3025 , \2796 );
and \U$1555 ( \3659 , \3058 , \2794 );
nor \U$1556 ( \3660 , \3658 , \3659 );
xnor \U$1557 ( \3661 , \3660 , \2801 );
xor \U$1558 ( \3662 , \3657 , \3661 );
and \U$1559 ( \3663 , \3087 , \2731 );
and \U$1560 ( \3664 , \3116 , \2729 );
nor \U$1561 ( \3665 , \3663 , \3664 );
xnor \U$1562 ( \3666 , \3665 , \2540 );
xor \U$1563 ( \3667 , \3662 , \3666 );
xor \U$1564 ( \3668 , \3653 , \3667 );
xor \U$1565 ( \3669 , \3643 , \3668 );
xor \U$1566 ( \3670 , \3634 , \3669 );
and \U$1567 ( \3671 , \3524 , \3592 );
nor \U$1568 ( \3672 , \3670 , \3671 );
and \U$1569 ( \3673 , \3638 , \3642 );
and \U$1570 ( \3674 , \3642 , \3668 );
and \U$1571 ( \3675 , \3638 , \3668 );
or \U$1572 ( \3676 , \3673 , \3674 , \3675 );
and \U$1573 ( \3677 , \3612 , \3632 );
xor \U$1574 ( \3678 , \3676 , \3677 );
and \U$1577 ( \3679 , \3616 , \3631 );
or \U$1578 ( \3680 , 1'b0 , 1'b0 , \3679 );
and \U$1580 ( \3681 , \3116 , \2731 );
and \U$1581 ( \3682 , \3025 , \2729 );
nor \U$1582 ( \3683 , \3681 , \3682 );
xnor \U$1583 ( \3684 , \3683 , \2540 );
and \U$1584 ( \3685 , \3163 , \2669 );
and \U$1585 ( \3686 , \3087 , \2667 );
nor \U$1586 ( \3687 , \3685 , \3686 );
xnor \U$1587 ( \3688 , \3687 , \2695 );
xor \U$1588 ( \3689 , \3684 , \3688 );
and \U$1590 ( \3690 , \3142 , \2722 );
nor \U$1591 ( \3691 , 1'b0 , \3690 );
xnor \U$1592 ( \3692 , \3691 , 1'b0 );
xor \U$1593 ( \3693 , \3689 , \3692 );
xor \U$1594 ( \3694 , 1'b0 , \3693 );
and \U$1595 ( \3695 , \2828 , \3037 );
and \U$1596 ( \3696 , \2849 , \3035 );
nor \U$1597 ( \3697 , \3695 , \3696 );
xnor \U$1598 ( \3698 , \3697 , \3063 );
and \U$1599 ( \3699 , \2998 , \3095 );
and \U$1600 ( \3700 , \2872 , \3093 );
nor \U$1601 ( \3701 , \3699 , \3700 );
xnor \U$1602 ( \3702 , \3701 , \3121 );
xor \U$1603 ( \3703 , \3698 , \3702 );
and \U$1604 ( \3704 , \3058 , \2796 );
and \U$1605 ( \3705 , \2965 , \2794 );
nor \U$1606 ( \3706 , \3704 , \3705 );
xnor \U$1607 ( \3707 , \3706 , \2801 );
xor \U$1608 ( \3708 , \3703 , \3707 );
xor \U$1609 ( \3709 , \3694 , \3708 );
and \U$1610 ( \3710 , \3621 , \3625 );
and \U$1611 ( \3711 , \3625 , \3630 );
and \U$1612 ( \3712 , \3621 , \3630 );
or \U$1613 ( \3713 , \3710 , \3711 , \3712 );
and \U$1614 ( \3714 , \3657 , \3661 );
and \U$1615 ( \3715 , \3661 , \3666 );
and \U$1616 ( \3716 , \3657 , \3666 );
or \U$1617 ( \3717 , \3714 , \3715 , \3716 );
xor \U$1618 ( \3718 , \3713 , \3717 );
and \U$1619 ( \3719 , \3647 , \3650 );
or \U$1622 ( \3720 , \3719 , 1'b0 , 1'b0 );
xor \U$1623 ( \3721 , \3718 , \3720 );
xor \U$1624 ( \3722 , \3709 , \3721 );
xor \U$1625 ( \3723 , \3680 , \3722 );
and \U$1626 ( \3724 , \3602 , \3606 );
and \U$1627 ( \3725 , \3606 , \3611 );
and \U$1628 ( \3726 , \3602 , \3611 );
or \U$1629 ( \3727 , \3724 , \3725 , \3726 );
and \U$1631 ( \3728 , \3652 , \3667 );
or \U$1633 ( \3729 , 1'b0 , \3728 , 1'b0 );
xor \U$1634 ( \3730 , \3727 , \3729 );
and \U$1636 ( \3731 , \2690 , \2941 );
not \U$1637 ( \3732 , \3731 );
xnor \U$1638 ( \3733 , \3732 , \2935 );
xor \U$1639 ( \3734 , 1'b0 , \3733 );
and \U$1640 ( \3735 , \2717 , \2977 );
and \U$1641 ( \3736 , \2621 , \2975 );
nor \U$1642 ( \3737 , \3735 , \3736 );
xnor \U$1643 ( \3738 , \3737 , \3003 );
xor \U$1644 ( \3739 , \3734 , \3738 );
xor \U$1645 ( \3740 , \3730 , \3739 );
xor \U$1646 ( \3741 , \3723 , \3740 );
xor \U$1647 ( \3742 , \3678 , \3741 );
and \U$1648 ( \3743 , \3600 , \3633 );
and \U$1649 ( \3744 , \3633 , \3669 );
and \U$1650 ( \3745 , \3600 , \3669 );
or \U$1651 ( \3746 , \3743 , \3744 , \3745 );
nor \U$1652 ( \3747 , \3742 , \3746 );
nor \U$1653 ( \3748 , \3672 , \3747 );
nand \U$1654 ( \3749 , \3596 , \3748 );
and \U$1655 ( \3750 , \3680 , \3722 );
and \U$1656 ( \3751 , \3722 , \3740 );
and \U$1657 ( \3752 , \3680 , \3740 );
or \U$1658 ( \3753 , \3750 , \3751 , \3752 );
and \U$1659 ( \3754 , \3713 , \3717 );
and \U$1660 ( \3755 , \3717 , \3720 );
and \U$1661 ( \3756 , \3713 , \3720 );
or \U$1662 ( \3757 , \3754 , \3755 , \3756 );
and \U$1664 ( \3758 , \3693 , \3708 );
or \U$1666 ( \3759 , 1'b0 , \3758 , 1'b0 );
xor \U$1667 ( \3760 , \3757 , \3759 );
and \U$1668 ( \3761 , \2872 , \3095 );
and \U$1669 ( \3762 , \2828 , \3093 );
nor \U$1670 ( \3763 , \3761 , \3762 );
xnor \U$1671 ( \3764 , \3763 , \3121 );
and \U$1672 ( \3765 , \2965 , \2796 );
and \U$1673 ( \3766 , \2998 , \2794 );
nor \U$1674 ( \3767 , \3765 , \3766 );
xnor \U$1675 ( \3768 , \3767 , \2801 );
xor \U$1676 ( \3769 , \3764 , \3768 );
and \U$1677 ( \3770 , \3025 , \2731 );
and \U$1678 ( \3771 , \3058 , \2729 );
nor \U$1679 ( \3772 , \3770 , \3771 );
xnor \U$1680 ( \3773 , \3772 , \2540 );
xor \U$1681 ( \3774 , \3769 , \3773 );
xor \U$1682 ( \3775 , \3760 , \3774 );
xor \U$1683 ( \3776 , \3753 , \3775 );
and \U$1684 ( \3777 , \3727 , \3729 );
and \U$1685 ( \3778 , \3729 , \3739 );
and \U$1686 ( \3779 , \3727 , \3739 );
or \U$1687 ( \3780 , \3777 , \3778 , \3779 );
and \U$1688 ( \3781 , \3709 , \3721 );
xor \U$1689 ( \3782 , \3780 , \3781 );
not \U$1690 ( \3783 , \2935 );
and \U$1691 ( \3784 , \2621 , \2977 );
and \U$1692 ( \3785 , \2690 , \2975 );
nor \U$1693 ( \3786 , \3784 , \3785 );
xnor \U$1694 ( \3787 , \3786 , \3003 );
xor \U$1695 ( \3788 , \3783 , \3787 );
and \U$1696 ( \3789 , \2849 , \3037 );
and \U$1697 ( \3790 , \2717 , \3035 );
nor \U$1698 ( \3791 , \3789 , \3790 );
xnor \U$1699 ( \3792 , \3791 , \3063 );
xor \U$1700 ( \3793 , \3788 , \3792 );
and \U$1702 ( \3794 , \3087 , \2669 );
and \U$1703 ( \3795 , \3116 , \2667 );
nor \U$1704 ( \3796 , \3794 , \3795 );
xnor \U$1705 ( \3797 , \3796 , \2695 );
and \U$1707 ( \3798 , \3163 , \2722 );
nor \U$1708 ( \3799 , 1'b0 , \3798 );
xnor \U$1709 ( \3800 , \3799 , 1'b0 );
xor \U$1710 ( \3801 , \3797 , \3800 );
xor \U$1712 ( \3802 , \3801 , 1'b0 );
xor \U$1713 ( \3803 , 1'b1 , \3802 );
xor \U$1714 ( \3804 , \3793 , \3803 );
and \U$1716 ( \3805 , \3733 , \3738 );
or \U$1718 ( \3806 , 1'b0 , \3805 , 1'b0 );
and \U$1719 ( \3807 , \3698 , \3702 );
and \U$1720 ( \3808 , \3702 , \3707 );
and \U$1721 ( \3809 , \3698 , \3707 );
or \U$1722 ( \3810 , \3807 , \3808 , \3809 );
xor \U$1723 ( \3811 , \3806 , \3810 );
and \U$1724 ( \3812 , \3684 , \3688 );
and \U$1725 ( \3813 , \3688 , \3692 );
and \U$1726 ( \3814 , \3684 , \3692 );
or \U$1727 ( \3815 , \3812 , \3813 , \3814 );
xor \U$1728 ( \3816 , \3811 , \3815 );
xor \U$1729 ( \3817 , \3804 , \3816 );
xor \U$1730 ( \3818 , \3782 , \3817 );
xor \U$1731 ( \3819 , \3776 , \3818 );
and \U$1732 ( \3820 , \3676 , \3677 );
and \U$1733 ( \3821 , \3677 , \3741 );
and \U$1734 ( \3822 , \3676 , \3741 );
or \U$1735 ( \3823 , \3820 , \3821 , \3822 );
nor \U$1736 ( \3824 , \3819 , \3823 );
and \U$1737 ( \3825 , \3780 , \3781 );
and \U$1738 ( \3826 , \3781 , \3817 );
and \U$1739 ( \3827 , \3780 , \3817 );
or \U$1740 ( \3828 , \3825 , \3826 , \3827 );
and \U$1741 ( \3829 , \3783 , \3787 );
and \U$1742 ( \3830 , \3787 , \3792 );
and \U$1743 ( \3831 , \3783 , \3792 );
or \U$1744 ( \3832 , \3829 , \3830 , \3831 );
and \U$1745 ( \3833 , \3764 , \3768 );
and \U$1746 ( \3834 , \3768 , \3773 );
and \U$1747 ( \3835 , \3764 , \3773 );
or \U$1748 ( \3836 , \3833 , \3834 , \3835 );
xor \U$1749 ( \3837 , \3832 , \3836 );
and \U$1750 ( \3838 , \3797 , \3800 );
or \U$1753 ( \3839 , \3838 , 1'b0 , 1'b0 );
xor \U$1754 ( \3840 , \3837 , \3839 );
and \U$1755 ( \3841 , \3806 , \3810 );
and \U$1756 ( \3842 , \3810 , \3815 );
and \U$1757 ( \3843 , \3806 , \3815 );
or \U$1758 ( \3844 , \3841 , \3842 , \3843 );
and \U$1761 ( \3845 , 1'b1 , \3802 );
or \U$1763 ( \3846 , 1'b0 , \3845 , 1'b0 );
xor \U$1764 ( \3847 , \3844 , \3846 );
and \U$1765 ( \3848 , \3116 , \2669 );
and \U$1766 ( \3849 , \3025 , \2667 );
nor \U$1767 ( \3850 , \3848 , \3849 );
xnor \U$1768 ( \3851 , \3850 , \2695 );
and \U$1770 ( \3852 , \3087 , \2722 );
nor \U$1771 ( \3853 , 1'b0 , \3852 );
xnor \U$1772 ( \3854 , \3853 , 1'b0 );
xor \U$1773 ( \3855 , \3851 , \3854 );
xor \U$1775 ( \3856 , \3855 , 1'b0 );
and \U$1776 ( \3857 , \2828 , \3095 );
and \U$1777 ( \3858 , \2849 , \3093 );
nor \U$1778 ( \3859 , \3857 , \3858 );
xnor \U$1779 ( \3860 , \3859 , \3121 );
and \U$1780 ( \3861 , \2998 , \2796 );
and \U$1781 ( \3862 , \2872 , \2794 );
nor \U$1782 ( \3863 , \3861 , \3862 );
xnor \U$1783 ( \3864 , \3863 , \2801 );
xor \U$1784 ( \3865 , \3860 , \3864 );
and \U$1785 ( \3866 , \3058 , \2731 );
and \U$1786 ( \3867 , \2965 , \2729 );
nor \U$1787 ( \3868 , \3866 , \3867 );
xnor \U$1788 ( \3869 , \3868 , \2540 );
xor \U$1789 ( \3870 , \3865 , \3869 );
xor \U$1790 ( \3871 , \3856 , \3870 );
and \U$1792 ( \3872 , \2690 , \2977 );
not \U$1793 ( \3873 , \3872 );
xnor \U$1794 ( \3874 , \3873 , \3003 );
xor \U$1795 ( \3875 , 1'b0 , \3874 );
and \U$1796 ( \3876 , \2717 , \3037 );
and \U$1797 ( \3877 , \2621 , \3035 );
nor \U$1798 ( \3878 , \3876 , \3877 );
xnor \U$1799 ( \3879 , \3878 , \3063 );
xor \U$1800 ( \3880 , \3875 , \3879 );
xor \U$1801 ( \3881 , \3871 , \3880 );
xor \U$1802 ( \3882 , \3847 , \3881 );
xor \U$1803 ( \3883 , \3840 , \3882 );
xor \U$1804 ( \3884 , \3828 , \3883 );
and \U$1805 ( \3885 , \3757 , \3759 );
and \U$1806 ( \3886 , \3759 , \3774 );
and \U$1807 ( \3887 , \3757 , \3774 );
or \U$1808 ( \3888 , \3885 , \3886 , \3887 );
and \U$1809 ( \3889 , \3793 , \3803 );
and \U$1810 ( \3890 , \3803 , \3816 );
and \U$1811 ( \3891 , \3793 , \3816 );
or \U$1812 ( \3892 , \3889 , \3890 , \3891 );
xor \U$1813 ( \3893 , \3888 , \3892 );
xor \U$1815 ( \3894 , \3893 , 1'b1 );
xor \U$1816 ( \3895 , \3884 , \3894 );
and \U$1817 ( \3896 , \3753 , \3775 );
and \U$1818 ( \3897 , \3775 , \3818 );
and \U$1819 ( \3898 , \3753 , \3818 );
or \U$1820 ( \3899 , \3896 , \3897 , \3898 );
nor \U$1821 ( \3900 , \3895 , \3899 );
nor \U$1822 ( \3901 , \3824 , \3900 );
and \U$1823 ( \3902 , \3888 , \3892 );
and \U$1824 ( \3903 , \3892 , 1'b1 );
and \U$1825 ( \3904 , \3888 , 1'b1 );
or \U$1826 ( \3905 , \3902 , \3903 , \3904 );
and \U$1827 ( \3906 , \3840 , \3882 );
xor \U$1828 ( \3907 , \3905 , \3906 );
and \U$1829 ( \3908 , \3844 , \3846 );
and \U$1830 ( \3909 , \3846 , \3881 );
and \U$1831 ( \3910 , \3844 , \3881 );
or \U$1832 ( \3911 , \3908 , \3909 , \3910 );
and \U$1834 ( \3912 , \3116 , \2722 );
nor \U$1835 ( \3913 , 1'b0 , \3912 );
xnor \U$1836 ( \3914 , \3913 , 1'b0 );
xor \U$1838 ( \3915 , \3914 , 1'b0 );
xor \U$1840 ( \3916 , \3915 , 1'b0 );
and \U$1841 ( \3917 , \2872 , \2796 );
and \U$1842 ( \3918 , \2828 , \2794 );
nor \U$1843 ( \3919 , \3917 , \3918 );
xnor \U$1844 ( \3920 , \3919 , \2801 );
and \U$1845 ( \3921 , \2965 , \2731 );
and \U$1846 ( \3922 , \2998 , \2729 );
nor \U$1847 ( \3923 , \3921 , \3922 );
xnor \U$1848 ( \3924 , \3923 , \2540 );
xor \U$1849 ( \3925 , \3920 , \3924 );
and \U$1850 ( \3926 , \3025 , \2669 );
and \U$1851 ( \3927 , \3058 , \2667 );
nor \U$1852 ( \3928 , \3926 , \3927 );
xnor \U$1853 ( \3929 , \3928 , \2695 );
xor \U$1854 ( \3930 , \3925 , \3929 );
xor \U$1855 ( \3931 , \3916 , \3930 );
not \U$1856 ( \3932 , \3003 );
and \U$1857 ( \3933 , \2621 , \3037 );
and \U$1858 ( \3934 , \2690 , \3035 );
nor \U$1859 ( \3935 , \3933 , \3934 );
xnor \U$1860 ( \3936 , \3935 , \3063 );
xor \U$1861 ( \3937 , \3932 , \3936 );
and \U$1862 ( \3938 , \2849 , \3095 );
and \U$1863 ( \3939 , \2717 , \3093 );
nor \U$1864 ( \3940 , \3938 , \3939 );
xnor \U$1865 ( \3941 , \3940 , \3121 );
xor \U$1866 ( \3942 , \3937 , \3941 );
xor \U$1867 ( \3943 , \3931 , \3942 );
xor \U$1869 ( \3944 , \3943 , 1'b0 );
and \U$1871 ( \3945 , \3874 , \3879 );
or \U$1873 ( \3946 , 1'b0 , \3945 , 1'b0 );
and \U$1874 ( \3947 , \3860 , \3864 );
and \U$1875 ( \3948 , \3864 , \3869 );
and \U$1876 ( \3949 , \3860 , \3869 );
or \U$1877 ( \3950 , \3947 , \3948 , \3949 );
xor \U$1878 ( \3951 , \3946 , \3950 );
and \U$1879 ( \3952 , \3851 , \3854 );
or \U$1882 ( \3953 , \3952 , 1'b0 , 1'b0 );
xor \U$1883 ( \3954 , \3951 , \3953 );
xor \U$1884 ( \3955 , \3944 , \3954 );
xor \U$1885 ( \3956 , \3911 , \3955 );
and \U$1886 ( \3957 , \3832 , \3836 );
and \U$1887 ( \3958 , \3836 , \3839 );
and \U$1888 ( \3959 , \3832 , \3839 );
or \U$1889 ( \3960 , \3957 , \3958 , \3959 );
xor \U$1891 ( \3961 , \3960 , 1'b0 );
and \U$1892 ( \3962 , \3856 , \3870 );
and \U$1893 ( \3963 , \3870 , \3880 );
and \U$1894 ( \3964 , \3856 , \3880 );
or \U$1895 ( \3965 , \3962 , \3963 , \3964 );
xor \U$1896 ( \3966 , \3961 , \3965 );
xor \U$1897 ( \3967 , \3956 , \3966 );
xor \U$1898 ( \3968 , \3907 , \3967 );
and \U$1899 ( \3969 , \3828 , \3883 );
and \U$1900 ( \3970 , \3883 , \3894 );
and \U$1901 ( \3971 , \3828 , \3894 );
or \U$1902 ( \3972 , \3969 , \3970 , \3971 );
nor \U$1903 ( \3973 , \3968 , \3972 );
and \U$1904 ( \3974 , \3911 , \3955 );
and \U$1905 ( \3975 , \3955 , \3966 );
and \U$1906 ( \3976 , \3911 , \3966 );
or \U$1907 ( \3977 , \3974 , \3975 , \3976 );
and \U$1908 ( \3978 , \3946 , \3950 );
and \U$1909 ( \3979 , \3950 , \3953 );
and \U$1910 ( \3980 , \3946 , \3953 );
or \U$1911 ( \3981 , \3978 , \3979 , \3980 );
xor \U$1913 ( \3982 , \3981 , 1'b0 );
and \U$1914 ( \3983 , \3916 , \3930 );
and \U$1915 ( \3984 , \3930 , \3942 );
and \U$1916 ( \3985 , \3916 , \3942 );
or \U$1917 ( \3986 , \3983 , \3984 , \3985 );
xor \U$1918 ( \3987 , \3982 , \3986 );
xor \U$1919 ( \3988 , \3977 , \3987 );
and \U$1922 ( \3989 , \3960 , \3965 );
or \U$1923 ( \3990 , 1'b0 , 1'b0 , \3989 );
and \U$1926 ( \3991 , \3943 , \3954 );
or \U$1927 ( \3992 , 1'b0 , 1'b0 , \3991 );
xor \U$1928 ( \3993 , \3990 , \3992 );
and \U$1929 ( \3994 , \2828 , \2796 );
and \U$1930 ( \3995 , \2849 , \2794 );
nor \U$1931 ( \3996 , \3994 , \3995 );
xnor \U$1932 ( \3997 , \3996 , \2801 );
and \U$1933 ( \3998 , \2998 , \2731 );
and \U$1934 ( \3999 , \2872 , \2729 );
nor \U$1935 ( \4000 , \3998 , \3999 );
xnor \U$1936 ( \4001 , \4000 , \2540 );
xor \U$1937 ( \4002 , \3997 , \4001 );
and \U$1938 ( \4003 , \3058 , \2669 );
and \U$1939 ( \4004 , \2965 , \2667 );
nor \U$1940 ( \4005 , \4003 , \4004 );
xnor \U$1941 ( \4006 , \4005 , \2695 );
xor \U$1942 ( \4007 , \4002 , \4006 );
and \U$1944 ( \4008 , \2690 , \3037 );
not \U$1945 ( \4009 , \4008 );
xnor \U$1946 ( \4010 , \4009 , \3063 );
xor \U$1947 ( \4011 , 1'b0 , \4010 );
and \U$1948 ( \4012 , \2717 , \3095 );
and \U$1949 ( \4013 , \2621 , \3093 );
nor \U$1950 ( \4014 , \4012 , \4013 );
xnor \U$1951 ( \4015 , \4014 , \3121 );
xor \U$1952 ( \4016 , \4011 , \4015 );
xor \U$1953 ( \4017 , \4007 , \4016 );
and \U$1956 ( \4018 , \3025 , \2722 );
nor \U$1957 ( \4019 , 1'b0 , \4018 );
xnor \U$1958 ( \4020 , \4019 , 1'b0 );
xor \U$1960 ( \4021 , \4020 , 1'b0 );
xor \U$1962 ( \4022 , \4021 , 1'b0 );
xnor \U$1963 ( \4023 , 1'b0 , \4022 );
xor \U$1964 ( \4024 , \4017 , \4023 );
and \U$1965 ( \4025 , \3932 , \3936 );
and \U$1966 ( \4026 , \3936 , \3941 );
and \U$1967 ( \4027 , \3932 , \3941 );
or \U$1968 ( \4028 , \4025 , \4026 , \4027 );
and \U$1969 ( \4029 , \3920 , \3924 );
and \U$1970 ( \4030 , \3924 , \3929 );
and \U$1971 ( \4031 , \3920 , \3929 );
or \U$1972 ( \4032 , \4029 , \4030 , \4031 );
xor \U$1973 ( \4033 , \4028 , \4032 );
xor \U$1975 ( \4034 , \4033 , 1'b0 );
xor \U$1976 ( \4035 , \4024 , \4034 );
xor \U$1977 ( \4036 , \3993 , \4035 );
xor \U$1978 ( \4037 , \3988 , \4036 );
and \U$1979 ( \4038 , \3905 , \3906 );
and \U$1980 ( \4039 , \3906 , \3967 );
and \U$1981 ( \4040 , \3905 , \3967 );
or \U$1982 ( \4041 , \4038 , \4039 , \4040 );
nor \U$1983 ( \4042 , \4037 , \4041 );
nor \U$1984 ( \4043 , \3973 , \4042 );
nand \U$1985 ( \4044 , \3901 , \4043 );
nor \U$1986 ( \4045 , \3749 , \4044 );
and \U$1987 ( \4046 , \3990 , \3992 );
and \U$1988 ( \4047 , \3992 , \4035 );
and \U$1989 ( \4048 , \3990 , \4035 );
or \U$1990 ( \4049 , \4046 , \4047 , \4048 );
and \U$1991 ( \4050 , \4028 , \4032 );
or \U$1994 ( \4051 , \4050 , 1'b0 , 1'b0 );
or \U$1995 ( \4052 , 1'b0 , \4022 );
xor \U$1996 ( \4053 , \4051 , \4052 );
and \U$1997 ( \4054 , \4007 , \4016 );
xor \U$1998 ( \4055 , \4053 , \4054 );
xor \U$1999 ( \4056 , \4049 , \4055 );
and \U$2002 ( \4057 , \3981 , \3986 );
or \U$2003 ( \4058 , 1'b0 , 1'b0 , \4057 );
and \U$2004 ( \4059 , \4017 , \4023 );
and \U$2005 ( \4060 , \4023 , \4034 );
and \U$2006 ( \4061 , \4017 , \4034 );
or \U$2007 ( \4062 , \4059 , \4060 , \4061 );
xor \U$2008 ( \4063 , \4058 , \4062 );
and \U$2010 ( \4064 , \2872 , \2731 );
and \U$2011 ( \4065 , \2828 , \2729 );
nor \U$2012 ( \4066 , \4064 , \4065 );
xnor \U$2013 ( \4067 , \4066 , \2540 );
and \U$2014 ( \4068 , \2965 , \2669 );
and \U$2015 ( \4069 , \2998 , \2667 );
nor \U$2016 ( \4070 , \4068 , \4069 );
xnor \U$2017 ( \4071 , \4070 , \2695 );
xor \U$2018 ( \4072 , \4067 , \4071 );
and \U$2020 ( \4073 , \3058 , \2722 );
nor \U$2021 ( \4074 , 1'b0 , \4073 );
xnor \U$2022 ( \4075 , \4074 , 1'b0 );
xor \U$2023 ( \4076 , \4072 , \4075 );
xor \U$2024 ( \4077 , 1'b0 , \4076 );
not \U$2025 ( \4078 , \3063 );
and \U$2026 ( \4079 , \2621 , \3095 );
and \U$2027 ( \4080 , \2690 , \3093 );
nor \U$2028 ( \4081 , \4079 , \4080 );
xnor \U$2029 ( \4082 , \4081 , \3121 );
xor \U$2030 ( \4083 , \4078 , \4082 );
and \U$2031 ( \4084 , \2849 , \2796 );
and \U$2032 ( \4085 , \2717 , \2794 );
nor \U$2033 ( \4086 , \4084 , \4085 );
xnor \U$2034 ( \4087 , \4086 , \2801 );
xor \U$2035 ( \4088 , \4083 , \4087 );
xor \U$2036 ( \4089 , \4077 , \4088 );
xor \U$2038 ( \4090 , \4089 , 1'b0 );
and \U$2040 ( \4091 , \4010 , \4015 );
or \U$2042 ( \4092 , 1'b0 , \4091 , 1'b0 );
and \U$2043 ( \4093 , \3997 , \4001 );
and \U$2044 ( \4094 , \4001 , \4006 );
and \U$2045 ( \4095 , \3997 , \4006 );
or \U$2046 ( \4096 , \4093 , \4094 , \4095 );
xor \U$2047 ( \4097 , \4092 , \4096 );
xor \U$2049 ( \4098 , \4097 , 1'b0 );
xor \U$2050 ( \4099 , \4090 , \4098 );
xor \U$2051 ( \4100 , \4063 , \4099 );
xor \U$2052 ( \4101 , \4056 , \4100 );
and \U$2053 ( \4102 , \3977 , \3987 );
and \U$2054 ( \4103 , \3987 , \4036 );
and \U$2055 ( \4104 , \3977 , \4036 );
or \U$2056 ( \4105 , \4102 , \4103 , \4104 );
nor \U$2057 ( \4106 , \4101 , \4105 );
and \U$2058 ( \4107 , \4058 , \4062 );
and \U$2059 ( \4108 , \4062 , \4099 );
and \U$2060 ( \4109 , \4058 , \4099 );
or \U$2061 ( \4110 , \4107 , \4108 , \4109 );
and \U$2062 ( \4111 , \4092 , \4096 );
or \U$2065 ( \4112 , \4111 , 1'b0 , 1'b0 );
xor \U$2067 ( \4113 , \4112 , 1'b0 );
and \U$2069 ( \4114 , \4076 , \4088 );
or \U$2071 ( \4115 , 1'b0 , \4114 , 1'b0 );
xor \U$2072 ( \4116 , \4113 , \4115 );
xor \U$2073 ( \4117 , \4110 , \4116 );
and \U$2074 ( \4118 , \4051 , \4052 );
and \U$2075 ( \4119 , \4052 , \4054 );
and \U$2076 ( \4120 , \4051 , \4054 );
or \U$2077 ( \4121 , \4118 , \4119 , \4120 );
and \U$2080 ( \4122 , \4089 , \4098 );
or \U$2081 ( \4123 , 1'b0 , 1'b0 , \4122 );
xor \U$2082 ( \4124 , \4121 , \4123 );
and \U$2083 ( \4125 , \2828 , \2731 );
and \U$2084 ( \4126 , \2849 , \2729 );
nor \U$2085 ( \4127 , \4125 , \4126 );
xnor \U$2086 ( \4128 , \4127 , \2540 );
and \U$2087 ( \4129 , \2998 , \2669 );
and \U$2088 ( \4130 , \2872 , \2667 );
nor \U$2089 ( \4131 , \4129 , \4130 );
xnor \U$2090 ( \4132 , \4131 , \2695 );
xor \U$2091 ( \4133 , \4128 , \4132 );
and \U$2093 ( \4134 , \2965 , \2722 );
nor \U$2094 ( \4135 , 1'b0 , \4134 );
xnor \U$2095 ( \4136 , \4135 , 1'b0 );
xor \U$2096 ( \4137 , \4133 , \4136 );
and \U$2098 ( \4138 , \2690 , \3095 );
not \U$2099 ( \4139 , \4138 );
xnor \U$2100 ( \4140 , \4139 , \3121 );
xor \U$2101 ( \4141 , 1'b0 , \4140 );
and \U$2102 ( \4142 , \2717 , \2796 );
and \U$2103 ( \4143 , \2621 , \2794 );
nor \U$2104 ( \4144 , \4142 , \4143 );
xnor \U$2105 ( \4145 , \4144 , \2801 );
xor \U$2106 ( \4146 , \4141 , \4145 );
xor \U$2107 ( \4147 , \4137 , \4146 );
xor \U$2109 ( \4148 , \4147 , 1'b1 );
and \U$2110 ( \4149 , \4078 , \4082 );
and \U$2111 ( \4150 , \4082 , \4087 );
and \U$2112 ( \4151 , \4078 , \4087 );
or \U$2113 ( \4152 , \4149 , \4150 , \4151 );
and \U$2114 ( \4153 , \4067 , \4071 );
and \U$2115 ( \4154 , \4071 , \4075 );
and \U$2116 ( \4155 , \4067 , \4075 );
or \U$2117 ( \4156 , \4153 , \4154 , \4155 );
xor \U$2118 ( \4157 , \4152 , \4156 );
xor \U$2120 ( \4158 , \4157 , 1'b0 );
xor \U$2121 ( \4159 , \4148 , \4158 );
xor \U$2122 ( \4160 , \4124 , \4159 );
xor \U$2123 ( \4161 , \4117 , \4160 );
and \U$2124 ( \4162 , \4049 , \4055 );
and \U$2125 ( \4163 , \4055 , \4100 );
and \U$2126 ( \4164 , \4049 , \4100 );
or \U$2127 ( \4165 , \4162 , \4163 , \4164 );
nor \U$2128 ( \4166 , \4161 , \4165 );
nor \U$2129 ( \4167 , \4106 , \4166 );
and \U$2130 ( \4168 , \4121 , \4123 );
and \U$2131 ( \4169 , \4123 , \4159 );
and \U$2132 ( \4170 , \4121 , \4159 );
or \U$2133 ( \4171 , \4168 , \4169 , \4170 );
and \U$2134 ( \4172 , \4152 , \4156 );
or \U$2137 ( \4173 , \4172 , 1'b0 , 1'b0 );
xor \U$2139 ( \4174 , \4173 , 1'b0 );
and \U$2140 ( \4175 , \4137 , \4146 );
xor \U$2141 ( \4176 , \4174 , \4175 );
xor \U$2142 ( \4177 , \4171 , \4176 );
and \U$2145 ( \4178 , \4112 , \4115 );
or \U$2146 ( \4179 , 1'b0 , 1'b0 , \4178 );
and \U$2147 ( \4180 , \4147 , 1'b1 );
and \U$2148 ( \4181 , 1'b1 , \4158 );
and \U$2149 ( \4182 , \4147 , \4158 );
or \U$2150 ( \4183 , \4180 , \4181 , \4182 );
xor \U$2151 ( \4184 , \4179 , \4183 );
and \U$2153 ( \4185 , \2872 , \2669 );
and \U$2154 ( \4186 , \2828 , \2667 );
nor \U$2155 ( \4187 , \4185 , \4186 );
xnor \U$2156 ( \4188 , \4187 , \2695 );
and \U$2158 ( \4189 , \2998 , \2722 );
nor \U$2159 ( \4190 , 1'b0 , \4189 );
xnor \U$2160 ( \4191 , \4190 , 1'b0 );
xor \U$2161 ( \4192 , \4188 , \4191 );
xor \U$2163 ( \4193 , \4192 , 1'b0 );
xor \U$2164 ( \4194 , 1'b0 , \4193 );
not \U$2165 ( \4195 , \3121 );
and \U$2166 ( \4196 , \2621 , \2796 );
and \U$2167 ( \4197 , \2690 , \2794 );
nor \U$2168 ( \4198 , \4196 , \4197 );
xnor \U$2169 ( \4199 , \4198 , \2801 );
xor \U$2170 ( \4200 , \4195 , \4199 );
and \U$2171 ( \4201 , \2849 , \2731 );
and \U$2172 ( \4202 , \2717 , \2729 );
nor \U$2173 ( \4203 , \4201 , \4202 );
xnor \U$2174 ( \4204 , \4203 , \2540 );
xor \U$2175 ( \4205 , \4200 , \4204 );
xor \U$2176 ( \4206 , \4194 , \4205 );
xor \U$2178 ( \4207 , \4206 , 1'b0 );
and \U$2180 ( \4208 , \4140 , \4145 );
or \U$2182 ( \4209 , 1'b0 , \4208 , 1'b0 );
and \U$2183 ( \4210 , \4128 , \4132 );
and \U$2184 ( \4211 , \4132 , \4136 );
and \U$2185 ( \4212 , \4128 , \4136 );
or \U$2186 ( \4213 , \4210 , \4211 , \4212 );
xor \U$2187 ( \4214 , \4209 , \4213 );
xor \U$2189 ( \4215 , \4214 , 1'b0 );
xor \U$2190 ( \4216 , \4207 , \4215 );
xor \U$2191 ( \4217 , \4184 , \4216 );
xor \U$2192 ( \4218 , \4177 , \4217 );
and \U$2193 ( \4219 , \4110 , \4116 );
and \U$2194 ( \4220 , \4116 , \4160 );
and \U$2195 ( \4221 , \4110 , \4160 );
or \U$2196 ( \4222 , \4219 , \4220 , \4221 );
nor \U$2197 ( \4223 , \4218 , \4222 );
and \U$2198 ( \4224 , \4179 , \4183 );
and \U$2199 ( \4225 , \4183 , \4216 );
and \U$2200 ( \4226 , \4179 , \4216 );
or \U$2201 ( \4227 , \4224 , \4225 , \4226 );
and \U$2202 ( \4228 , \4209 , \4213 );
or \U$2205 ( \4229 , \4228 , 1'b0 , 1'b0 );
xor \U$2207 ( \4230 , \4229 , 1'b0 );
and \U$2209 ( \4231 , \4193 , \4205 );
or \U$2211 ( \4232 , 1'b0 , \4231 , 1'b0 );
xor \U$2212 ( \4233 , \4230 , \4232 );
xor \U$2213 ( \4234 , \4227 , \4233 );
and \U$2216 ( \4235 , \4173 , \4175 );
or \U$2217 ( \4236 , 1'b0 , 1'b0 , \4235 );
and \U$2220 ( \4237 , \4206 , \4215 );
or \U$2221 ( \4238 , 1'b0 , 1'b0 , \4237 );
xor \U$2222 ( \4239 , \4236 , \4238 );
xor \U$2223 ( \4240 , \2852 , \2875 );
xor \U$2225 ( \4241 , \4240 , 1'b0 );
xor \U$2227 ( \4242 , 1'b0 , \2802 );
xor \U$2228 ( \4243 , \4242 , \2806 );
xor \U$2229 ( \4244 , \4241 , \4243 );
xor \U$2231 ( \4245 , \4244 , 1'b1 );
and \U$2232 ( \4246 , \4195 , \4199 );
and \U$2233 ( \4247 , \4199 , \4204 );
and \U$2234 ( \4248 , \4195 , \4204 );
or \U$2235 ( \4249 , \4246 , \4247 , \4248 );
and \U$2236 ( \4250 , \4188 , \4191 );
or \U$2239 ( \4251 , \4250 , 1'b0 , 1'b0 );
xor \U$2240 ( \4252 , \4249 , \4251 );
xor \U$2242 ( \4253 , \4252 , 1'b0 );
xor \U$2243 ( \4254 , \4245 , \4253 );
xor \U$2244 ( \4255 , \4239 , \4254 );
xor \U$2245 ( \4256 , \4234 , \4255 );
and \U$2246 ( \4257 , \4171 , \4176 );
and \U$2247 ( \4258 , \4176 , \4217 );
and \U$2248 ( \4259 , \4171 , \4217 );
or \U$2249 ( \4260 , \4257 , \4258 , \4259 );
nor \U$2250 ( \4261 , \4256 , \4260 );
nor \U$2251 ( \4262 , \4223 , \4261 );
nand \U$2252 ( \4263 , \4167 , \4262 );
and \U$2253 ( \4264 , \4236 , \4238 );
and \U$2254 ( \4265 , \4238 , \4254 );
and \U$2255 ( \4266 , \4236 , \4254 );
or \U$2256 ( \4267 , \4264 , \4265 , \4266 );
and \U$2257 ( \4268 , \4249 , \4251 );
or \U$2260 ( \4269 , \4268 , 1'b0 , 1'b0 );
xor \U$2262 ( \4270 , \4269 , 1'b0 );
and \U$2263 ( \4271 , \4241 , \4243 );
xor \U$2264 ( \4272 , \4270 , \4271 );
xor \U$2265 ( \4273 , \4267 , \4272 );
and \U$2268 ( \4274 , \4229 , \4232 );
or \U$2269 ( \4275 , 1'b0 , 1'b0 , \4274 );
and \U$2270 ( \4276 , \4244 , 1'b1 );
and \U$2271 ( \4277 , 1'b1 , \4253 );
and \U$2272 ( \4278 , \4244 , \4253 );
or \U$2273 ( \4279 , \4276 , \4277 , \4278 );
xor \U$2274 ( \4280 , \4275 , \4279 );
xor \U$2276 ( \4281 , 1'b0 , \2884 );
xor \U$2277 ( \4282 , \4281 , \2895 );
xor \U$2279 ( \4283 , \4282 , 1'b0 );
xor \U$2280 ( \4284 , \2808 , \2877 );
xor \U$2282 ( \4285 , \4284 , 1'b0 );
xor \U$2283 ( \4286 , \4283 , \4285 );
xor \U$2284 ( \4287 , \4280 , \4286 );
xor \U$2285 ( \4288 , \4273 , \4287 );
and \U$2286 ( \4289 , \4227 , \4233 );
and \U$2287 ( \4290 , \4233 , \4255 );
and \U$2288 ( \4291 , \4227 , \4255 );
or \U$2289 ( \4292 , \4289 , \4290 , \4291 );
nor \U$2290 ( \4293 , \4288 , \4292 );
and \U$2291 ( \4294 , \4275 , \4279 );
and \U$2292 ( \4295 , \4279 , \4286 );
and \U$2293 ( \4296 , \4275 , \4286 );
or \U$2294 ( \4297 , \4294 , \4295 , \4296 );
xor \U$2296 ( \4298 , \2879 , 1'b0 );
xor \U$2297 ( \4299 , \4298 , \2897 );
xor \U$2298 ( \4300 , \4297 , \4299 );
and \U$2301 ( \4301 , \4269 , \4271 );
or \U$2302 ( \4302 , 1'b0 , 1'b0 , \4301 );
and \U$2305 ( \4303 , \4282 , \4285 );
or \U$2306 ( \4304 , 1'b0 , 1'b0 , \4303 );
xor \U$2307 ( \4305 , \4302 , \4304 );
xor \U$2308 ( \4306 , \2907 , 1'b1 );
xor \U$2309 ( \4307 , \4306 , \2914 );
xor \U$2310 ( \4308 , \4305 , \4307 );
xor \U$2311 ( \4309 , \4300 , \4308 );
and \U$2312 ( \4310 , \4267 , \4272 );
and \U$2313 ( \4311 , \4272 , \4287 );
and \U$2314 ( \4312 , \4267 , \4287 );
or \U$2315 ( \4313 , \4310 , \4311 , \4312 );
nor \U$2316 ( \4314 , \4309 , \4313 );
nor \U$2317 ( \4315 , \4293 , \4314 );
and \U$2318 ( \4316 , \4302 , \4304 );
and \U$2319 ( \4317 , \4304 , \4307 );
and \U$2320 ( \4318 , \4302 , \4307 );
or \U$2321 ( \4319 , \4316 , \4317 , \4318 );
and \U$2323 ( \4320 , \2904 , \2906 );
xor \U$2324 ( \4321 , 1'b0 , \4320 );
xor \U$2325 ( \4322 , \4319 , \4321 );
xor \U$2326 ( \4323 , \2899 , \2917 );
xor \U$2327 ( \4324 , \4323 , \2920 );
xor \U$2328 ( \4325 , \4322 , \4324 );
and \U$2329 ( \4326 , \4297 , \4299 );
and \U$2330 ( \4327 , \4299 , \4308 );
and \U$2331 ( \4328 , \4297 , \4308 );
or \U$2332 ( \4329 , \4326 , \4327 , \4328 );
nor \U$2333 ( \4330 , \4325 , \4329 );
xor \U$2335 ( \4331 , \2923 , 1'b0 );
xor \U$2336 ( \4332 , \4331 , \2925 );
and \U$2337 ( \4333 , \4319 , \4321 );
and \U$2338 ( \4334 , \4321 , \4324 );
and \U$2339 ( \4335 , \4319 , \4324 );
or \U$2340 ( \4336 , \4333 , \4334 , \4335 );
nor \U$2341 ( \4337 , \4332 , \4336 );
nor \U$2342 ( \4338 , \4330 , \4337 );
nand \U$2343 ( \4339 , \4315 , \4338 );
nor \U$2344 ( \4340 , \4263 , \4339 );
nand \U$2345 ( \4341 , \4045 , \4340 );
and \U$2346 ( \4342 , \3142 , \2941 );
and \U$2347 ( \4343 , \3163 , \2938 );
nor \U$2348 ( \4344 , \4342 , \4343 );
xnor \U$2349 ( \4345 , \4344 , \2935 );
and \U$2350 ( \4346 , \3187 , \2977 );
and \U$2351 ( \4347 , \3208 , \2975 );
nor \U$2352 ( \4348 , \4346 , \4347 );
xnor \U$2353 ( \4349 , \4348 , \3003 );
and \U$2354 ( \4350 , \4345 , \4349 );
and \U$2355 ( \4351 , \3235 , \3037 );
and \U$2356 ( \4352 , \3256 , \3035 );
nor \U$2357 ( \4353 , \4351 , \4352 );
xnor \U$2358 ( \4354 , \4353 , \3063 );
and \U$2359 ( \4355 , \4349 , \4354 );
and \U$2360 ( \4356 , \4345 , \4354 );
or \U$2361 ( \4357 , \4350 , \4355 , \4356 );
and \U$2362 ( \4358 , \3256 , \3037 );
and \U$2363 ( \4359 , \3187 , \3035 );
nor \U$2364 ( \4360 , \4358 , \4359 );
xnor \U$2365 ( \4361 , \4360 , \3063 );
and \U$2366 ( \4362 , \3279 , \3095 );
and \U$2367 ( \4363 , \3235 , \3093 );
nor \U$2368 ( \4364 , \4362 , \4363 );
xnor \U$2369 ( \4365 , \4364 , \3121 );
xor \U$2370 ( \4366 , \4361 , \4365 );
nand \U$2371 ( \4367 , \3412 , \2794 );
xnor \U$2372 ( \4368 , \4367 , \2801 );
xor \U$2373 ( \4369 , \4366 , \4368 );
and \U$2374 ( \4370 , \4357 , \4369 );
and \U$2375 ( \4371 , \3163 , \2941 );
and \U$2376 ( \4372 , \3087 , \2938 );
nor \U$2377 ( \4373 , \4371 , \4372 );
xnor \U$2378 ( \4374 , \4373 , \2935 );
xor \U$2379 ( \4375 , \2801 , \4374 );
and \U$2380 ( \4376 , \3208 , \2977 );
and \U$2381 ( \4377 , \3142 , \2975 );
nor \U$2382 ( \4378 , \4376 , \4377 );
xnor \U$2383 ( \4379 , \4378 , \3003 );
xor \U$2384 ( \4380 , \4375 , \4379 );
and \U$2385 ( \4381 , \4369 , \4380 );
and \U$2386 ( \4382 , \4357 , \4380 );
or \U$2387 ( \4383 , \4370 , \4381 , \4382 );
and \U$2388 ( \4384 , \3412 , \2796 );
and \U$2389 ( \4385 , \3279 , \2794 );
nor \U$2390 ( \4386 , \4384 , \4385 );
xnor \U$2391 ( \4387 , \4386 , \2801 );
and \U$2392 ( \4388 , \3087 , \2941 );
and \U$2393 ( \4389 , \3116 , \2938 );
nor \U$2394 ( \4390 , \4388 , \4389 );
xnor \U$2395 ( \4391 , \4390 , \2935 );
and \U$2396 ( \4392 , \3142 , \2977 );
and \U$2397 ( \4393 , \3163 , \2975 );
nor \U$2398 ( \4394 , \4392 , \4393 );
xnor \U$2399 ( \4395 , \4394 , \3003 );
xor \U$2400 ( \4396 , \4391 , \4395 );
and \U$2401 ( \4397 , \3187 , \3037 );
and \U$2402 ( \4398 , \3208 , \3035 );
nor \U$2403 ( \4399 , \4397 , \4398 );
xnor \U$2404 ( \4400 , \4399 , \3063 );
xor \U$2405 ( \4401 , \4396 , \4400 );
xor \U$2406 ( \4402 , \4387 , \4401 );
xor \U$2407 ( \4403 , \4383 , \4402 );
and \U$2408 ( \4404 , \2801 , \4374 );
and \U$2409 ( \4405 , \4374 , \4379 );
and \U$2410 ( \4406 , \2801 , \4379 );
or \U$2411 ( \4407 , \4404 , \4405 , \4406 );
and \U$2412 ( \4408 , \4361 , \4365 );
and \U$2413 ( \4409 , \4365 , \4368 );
and \U$2414 ( \4410 , \4361 , \4368 );
or \U$2415 ( \4411 , \4408 , \4409 , \4410 );
xor \U$2416 ( \4412 , \4407 , \4411 );
and \U$2417 ( \4413 , \3235 , \3095 );
and \U$2418 ( \4414 , \3256 , \3093 );
nor \U$2419 ( \4415 , \4413 , \4414 );
xnor \U$2420 ( \4416 , \4415 , \3121 );
xor \U$2421 ( \4417 , \4412 , \4416 );
xor \U$2422 ( \4418 , \4403 , \4417 );
and \U$2423 ( \4419 , \3208 , \2941 );
and \U$2424 ( \4420 , \3142 , \2938 );
nor \U$2425 ( \4421 , \4419 , \4420 );
xnor \U$2426 ( \4422 , \4421 , \2935 );
and \U$2427 ( \4423 , \3121 , \4422 );
and \U$2428 ( \4424 , \3256 , \2977 );
and \U$2429 ( \4425 , \3187 , \2975 );
nor \U$2430 ( \4426 , \4424 , \4425 );
xnor \U$2431 ( \4427 , \4426 , \3003 );
and \U$2432 ( \4428 , \4422 , \4427 );
and \U$2433 ( \4429 , \3121 , \4427 );
or \U$2434 ( \4430 , \4423 , \4428 , \4429 );
and \U$2435 ( \4431 , \3279 , \3037 );
and \U$2436 ( \4432 , \3235 , \3035 );
nor \U$2437 ( \4433 , \4431 , \4432 );
xnor \U$2438 ( \4434 , \4433 , \3063 );
nand \U$2439 ( \4435 , \3412 , \3093 );
xnor \U$2440 ( \4436 , \4435 , \3121 );
and \U$2441 ( \4437 , \4434 , \4436 );
and \U$2442 ( \4438 , \4430 , \4437 );
and \U$2443 ( \4439 , \3412 , \3095 );
and \U$2444 ( \4440 , \3279 , \3093 );
nor \U$2445 ( \4441 , \4439 , \4440 );
xnor \U$2446 ( \4442 , \4441 , \3121 );
and \U$2447 ( \4443 , \4437 , \4442 );
and \U$2448 ( \4444 , \4430 , \4442 );
or \U$2449 ( \4445 , \4438 , \4443 , \4444 );
xor \U$2450 ( \4446 , \4357 , \4369 );
xor \U$2451 ( \4447 , \4446 , \4380 );
and \U$2452 ( \4448 , \4445 , \4447 );
nor \U$2453 ( \4449 , \4418 , \4448 );
and \U$2454 ( \4450 , \4391 , \4395 );
and \U$2455 ( \4451 , \4395 , \4400 );
and \U$2456 ( \4452 , \4391 , \4400 );
or \U$2457 ( \4453 , \4450 , \4451 , \4452 );
nand \U$2458 ( \4454 , \3412 , \2729 );
xnor \U$2459 ( \4455 , \4454 , \2540 );
xor \U$2460 ( \4456 , \4453 , \4455 );
and \U$2461 ( \4457 , \3208 , \3037 );
and \U$2462 ( \4458 , \3142 , \3035 );
nor \U$2463 ( \4459 , \4457 , \4458 );
xnor \U$2464 ( \4460 , \4459 , \3063 );
and \U$2465 ( \4461 , \3256 , \3095 );
and \U$2466 ( \4462 , \3187 , \3093 );
nor \U$2467 ( \4463 , \4461 , \4462 );
xnor \U$2468 ( \4464 , \4463 , \3121 );
xor \U$2469 ( \4465 , \4460 , \4464 );
and \U$2470 ( \4466 , \3279 , \2796 );
and \U$2471 ( \4467 , \3235 , \2794 );
nor \U$2472 ( \4468 , \4466 , \4467 );
xnor \U$2473 ( \4469 , \4468 , \2801 );
xor \U$2474 ( \4470 , \4465 , \4469 );
xor \U$2475 ( \4471 , \4456 , \4470 );
and \U$2476 ( \4472 , \4407 , \4411 );
and \U$2477 ( \4473 , \4411 , \4416 );
and \U$2478 ( \4474 , \4407 , \4416 );
or \U$2479 ( \4475 , \4472 , \4473 , \4474 );
and \U$2480 ( \4476 , \4387 , \4401 );
xor \U$2481 ( \4477 , \4475 , \4476 );
and \U$2482 ( \4478 , \3116 , \2941 );
and \U$2483 ( \4479 , \3025 , \2938 );
nor \U$2484 ( \4480 , \4478 , \4479 );
xnor \U$2485 ( \4481 , \4480 , \2935 );
xor \U$2486 ( \4482 , \2540 , \4481 );
and \U$2487 ( \4483 , \3163 , \2977 );
and \U$2488 ( \4484 , \3087 , \2975 );
nor \U$2489 ( \4485 , \4483 , \4484 );
xnor \U$2490 ( \4486 , \4485 , \3003 );
xor \U$2491 ( \4487 , \4482 , \4486 );
xor \U$2492 ( \4488 , \4477 , \4487 );
xor \U$2493 ( \4489 , \4471 , \4488 );
and \U$2494 ( \4490 , \4383 , \4402 );
and \U$2495 ( \4491 , \4402 , \4417 );
and \U$2496 ( \4492 , \4383 , \4417 );
or \U$2497 ( \4493 , \4490 , \4491 , \4492 );
nor \U$2498 ( \4494 , \4489 , \4493 );
nor \U$2499 ( \4495 , \4449 , \4494 );
and \U$2500 ( \4496 , \4475 , \4476 );
and \U$2501 ( \4497 , \4476 , \4487 );
and \U$2502 ( \4498 , \4475 , \4487 );
or \U$2503 ( \4499 , \4496 , \4497 , \4498 );
and \U$2504 ( \4500 , \4453 , \4455 );
and \U$2505 ( \4501 , \4455 , \4470 );
and \U$2506 ( \4502 , \4453 , \4470 );
or \U$2507 ( \4503 , \4500 , \4501 , \4502 );
and \U$2508 ( \4504 , \3025 , \2941 );
and \U$2509 ( \4505 , \3058 , \2938 );
nor \U$2510 ( \4506 , \4504 , \4505 );
xnor \U$2511 ( \4507 , \4506 , \2935 );
and \U$2512 ( \4508 , \3087 , \2977 );
and \U$2513 ( \4509 , \3116 , \2975 );
nor \U$2514 ( \4510 , \4508 , \4509 );
xnor \U$2515 ( \4511 , \4510 , \3003 );
xor \U$2516 ( \4512 , \4507 , \4511 );
and \U$2517 ( \4513 , \3142 , \3037 );
and \U$2518 ( \4514 , \3163 , \3035 );
nor \U$2519 ( \4515 , \4513 , \4514 );
xnor \U$2520 ( \4516 , \4515 , \3063 );
xor \U$2521 ( \4517 , \4512 , \4516 );
xor \U$2522 ( \4518 , \4503 , \4517 );
and \U$2523 ( \4519 , \2540 , \4481 );
and \U$2524 ( \4520 , \4481 , \4486 );
and \U$2525 ( \4521 , \2540 , \4486 );
or \U$2526 ( \4522 , \4519 , \4520 , \4521 );
and \U$2527 ( \4523 , \4460 , \4464 );
and \U$2528 ( \4524 , \4464 , \4469 );
and \U$2529 ( \4525 , \4460 , \4469 );
or \U$2530 ( \4526 , \4523 , \4524 , \4525 );
xor \U$2531 ( \4527 , \4522 , \4526 );
and \U$2532 ( \4528 , \3187 , \3095 );
and \U$2533 ( \4529 , \3208 , \3093 );
nor \U$2534 ( \4530 , \4528 , \4529 );
xnor \U$2535 ( \4531 , \4530 , \3121 );
and \U$2536 ( \4532 , \3235 , \2796 );
and \U$2537 ( \4533 , \3256 , \2794 );
nor \U$2538 ( \4534 , \4532 , \4533 );
xnor \U$2539 ( \4535 , \4534 , \2801 );
xor \U$2540 ( \4536 , \4531 , \4535 );
and \U$2541 ( \4537 , \3412 , \2731 );
and \U$2542 ( \4538 , \3279 , \2729 );
nor \U$2543 ( \4539 , \4537 , \4538 );
xnor \U$2544 ( \4540 , \4539 , \2540 );
xor \U$2545 ( \4541 , \4536 , \4540 );
xor \U$2546 ( \4542 , \4527 , \4541 );
xor \U$2547 ( \4543 , \4518 , \4542 );
xor \U$2548 ( \4544 , \4499 , \4543 );
and \U$2549 ( \4545 , \4471 , \4488 );
nor \U$2550 ( \4546 , \4544 , \4545 );
and \U$2551 ( \4547 , \4503 , \4517 );
and \U$2552 ( \4548 , \4517 , \4542 );
and \U$2553 ( \4549 , \4503 , \4542 );
or \U$2554 ( \4550 , \4547 , \4548 , \4549 );
and \U$2555 ( \4551 , \4522 , \4526 );
and \U$2556 ( \4552 , \4526 , \4541 );
and \U$2557 ( \4553 , \4522 , \4541 );
or \U$2558 ( \4554 , \4551 , \4552 , \4553 );
nand \U$2559 ( \4555 , \3412 , \2667 );
xnor \U$2560 ( \4556 , \4555 , \2695 );
and \U$2561 ( \4557 , \3163 , \3037 );
and \U$2562 ( \4558 , \3087 , \3035 );
nor \U$2563 ( \4559 , \4557 , \4558 );
xnor \U$2564 ( \4560 , \4559 , \3063 );
and \U$2565 ( \4561 , \3208 , \3095 );
and \U$2566 ( \4562 , \3142 , \3093 );
nor \U$2567 ( \4563 , \4561 , \4562 );
xnor \U$2568 ( \4564 , \4563 , \3121 );
xor \U$2569 ( \4565 , \4560 , \4564 );
and \U$2570 ( \4566 , \3256 , \2796 );
and \U$2571 ( \4567 , \3187 , \2794 );
nor \U$2572 ( \4568 , \4566 , \4567 );
xnor \U$2573 ( \4569 , \4568 , \2801 );
xor \U$2574 ( \4570 , \4565 , \4569 );
xor \U$2575 ( \4571 , \4556 , \4570 );
and \U$2576 ( \4572 , \3058 , \2941 );
and \U$2577 ( \4573 , \2965 , \2938 );
nor \U$2578 ( \4574 , \4572 , \4573 );
xnor \U$2579 ( \4575 , \4574 , \2935 );
xor \U$2580 ( \4576 , \2695 , \4575 );
and \U$2581 ( \4577 , \3116 , \2977 );
and \U$2582 ( \4578 , \3025 , \2975 );
nor \U$2583 ( \4579 , \4577 , \4578 );
xnor \U$2584 ( \4580 , \4579 , \3003 );
xor \U$2585 ( \4581 , \4576 , \4580 );
xor \U$2586 ( \4582 , \4571 , \4581 );
xor \U$2587 ( \4583 , \4554 , \4582 );
and \U$2588 ( \4584 , \4507 , \4511 );
and \U$2589 ( \4585 , \4511 , \4516 );
and \U$2590 ( \4586 , \4507 , \4516 );
or \U$2591 ( \4587 , \4584 , \4585 , \4586 );
and \U$2592 ( \4588 , \4531 , \4535 );
and \U$2593 ( \4589 , \4535 , \4540 );
and \U$2594 ( \4590 , \4531 , \4540 );
or \U$2595 ( \4591 , \4588 , \4589 , \4590 );
xor \U$2596 ( \4592 , \4587 , \4591 );
and \U$2597 ( \4593 , \3279 , \2731 );
and \U$2598 ( \4594 , \3235 , \2729 );
nor \U$2599 ( \4595 , \4593 , \4594 );
xnor \U$2600 ( \4596 , \4595 , \2540 );
xor \U$2601 ( \4597 , \4592 , \4596 );
xor \U$2602 ( \4598 , \4583 , \4597 );
xor \U$2603 ( \4599 , \4550 , \4598 );
and \U$2604 ( \4600 , \4499 , \4543 );
nor \U$2605 ( \4601 , \4599 , \4600 );
nor \U$2606 ( \4602 , \4546 , \4601 );
nand \U$2607 ( \4603 , \4495 , \4602 );
and \U$2608 ( \4604 , \4554 , \4582 );
and \U$2609 ( \4605 , \4582 , \4597 );
and \U$2610 ( \4606 , \4554 , \4597 );
or \U$2611 ( \4607 , \4604 , \4605 , \4606 );
xor \U$2612 ( \4608 , \3467 , \3471 );
xor \U$2613 ( \4609 , \4608 , \3476 );
and \U$2614 ( \4610 , \2695 , \4575 );
and \U$2615 ( \4611 , \4575 , \4580 );
and \U$2616 ( \4612 , \2695 , \4580 );
or \U$2617 ( \4613 , \4610 , \4611 , \4612 );
and \U$2618 ( \4614 , \4560 , \4564 );
and \U$2619 ( \4615 , \4564 , \4569 );
and \U$2620 ( \4616 , \4560 , \4569 );
or \U$2621 ( \4617 , \4614 , \4615 , \4616 );
xor \U$2622 ( \4618 , \4613 , \4617 );
and \U$2623 ( \4619 , \3412 , \2669 );
and \U$2624 ( \4620 , \3279 , \2667 );
nor \U$2625 ( \4621 , \4619 , \4620 );
xnor \U$2626 ( \4622 , \4621 , \2695 );
xor \U$2627 ( \4623 , \4618 , \4622 );
xor \U$2628 ( \4624 , \4609 , \4623 );
xor \U$2629 ( \4625 , \4607 , \4624 );
and \U$2630 ( \4626 , \4587 , \4591 );
and \U$2631 ( \4627 , \4591 , \4596 );
and \U$2632 ( \4628 , \4587 , \4596 );
or \U$2633 ( \4629 , \4626 , \4627 , \4628 );
and \U$2634 ( \4630 , \4556 , \4570 );
and \U$2635 ( \4631 , \4570 , \4581 );
and \U$2636 ( \4632 , \4556 , \4581 );
or \U$2637 ( \4633 , \4630 , \4631 , \4632 );
xor \U$2638 ( \4634 , \4629 , \4633 );
xor \U$2639 ( \4635 , \3483 , \3487 );
xor \U$2640 ( \4636 , \4635 , \3492 );
xor \U$2641 ( \4637 , \4634 , \4636 );
xor \U$2642 ( \4638 , \4625 , \4637 );
and \U$2643 ( \4639 , \4550 , \4598 );
nor \U$2644 ( \4640 , \4638 , \4639 );
and \U$2645 ( \4641 , \4629 , \4633 );
and \U$2646 ( \4642 , \4633 , \4636 );
and \U$2647 ( \4643 , \4629 , \4636 );
or \U$2648 ( \4644 , \4641 , \4642 , \4643 );
and \U$2649 ( \4645 , \4609 , \4623 );
xor \U$2650 ( \4646 , \4644 , \4645 );
and \U$2651 ( \4647 , \4613 , \4617 );
and \U$2652 ( \4648 , \4617 , \4622 );
and \U$2653 ( \4649 , \4613 , \4622 );
or \U$2654 ( \4650 , \4647 , \4648 , \4649 );
xor \U$2655 ( \4651 , \3503 , \3505 );
xor \U$2656 ( \4652 , \4650 , \4651 );
xor \U$2657 ( \4653 , \3479 , \3495 );
xor \U$2658 ( \4654 , \4653 , \3498 );
xor \U$2659 ( \4655 , \4652 , \4654 );
xor \U$2660 ( \4656 , \4646 , \4655 );
and \U$2661 ( \4657 , \4607 , \4624 );
and \U$2662 ( \4658 , \4624 , \4637 );
and \U$2663 ( \4659 , \4607 , \4637 );
or \U$2664 ( \4660 , \4657 , \4658 , \4659 );
nor \U$2665 ( \4661 , \4656 , \4660 );
nor \U$2666 ( \4662 , \4640 , \4661 );
and \U$2667 ( \4663 , \4650 , \4651 );
and \U$2668 ( \4664 , \4651 , \4654 );
and \U$2669 ( \4665 , \4650 , \4654 );
or \U$2670 ( \4666 , \4663 , \4664 , \4665 );
xor \U$2671 ( \4667 , \3366 , \3382 );
xor \U$2672 ( \4668 , \4667 , \3417 );
xor \U$2673 ( \4669 , \4666 , \4668 );
xor \U$2674 ( \4670 , \3501 , \3506 );
xor \U$2675 ( \4671 , \4670 , \3509 );
xor \U$2676 ( \4672 , \4669 , \4671 );
and \U$2677 ( \4673 , \4644 , \4645 );
and \U$2678 ( \4674 , \4645 , \4655 );
and \U$2679 ( \4675 , \4644 , \4655 );
or \U$2680 ( \4676 , \4673 , \4674 , \4675 );
nor \U$2681 ( \4677 , \4672 , \4676 );
xor \U$2682 ( \4678 , \3512 , \3513 );
xor \U$2683 ( \4679 , \4678 , \3516 );
and \U$2684 ( \4680 , \4666 , \4668 );
and \U$2685 ( \4681 , \4668 , \4671 );
and \U$2686 ( \4682 , \4666 , \4671 );
or \U$2687 ( \4683 , \4680 , \4681 , \4682 );
nor \U$2688 ( \4684 , \4679 , \4683 );
nor \U$2689 ( \4685 , \4677 , \4684 );
nand \U$2690 ( \4686 , \4662 , \4685 );
nor \U$2691 ( \4687 , \4603 , \4686 );
and \U$2692 ( \4688 , \3256 , \2941 );
and \U$2693 ( \4689 , \3187 , \2938 );
nor \U$2694 ( \4690 , \4688 , \4689 );
xnor \U$2695 ( \4691 , \4690 , \2935 );
and \U$2696 ( \4692 , \3063 , \4691 );
and \U$2697 ( \4693 , \3279 , \2977 );
and \U$2698 ( \4694 , \3235 , \2975 );
nor \U$2699 ( \4695 , \4693 , \4694 );
xnor \U$2700 ( \4696 , \4695 , \3003 );
and \U$2701 ( \4697 , \4691 , \4696 );
and \U$2702 ( \4698 , \3063 , \4696 );
or \U$2703 ( \4699 , \4692 , \4697 , \4698 );
and \U$2704 ( \4700 , \3187 , \2941 );
and \U$2705 ( \4701 , \3208 , \2938 );
nor \U$2706 ( \4702 , \4700 , \4701 );
xnor \U$2707 ( \4703 , \4702 , \2935 );
and \U$2708 ( \4704 , \3235 , \2977 );
and \U$2709 ( \4705 , \3256 , \2975 );
nor \U$2710 ( \4706 , \4704 , \4705 );
xnor \U$2711 ( \4707 , \4706 , \3003 );
xor \U$2712 ( \4708 , \4703 , \4707 );
and \U$2713 ( \4709 , \3412 , \3037 );
and \U$2714 ( \4710 , \3279 , \3035 );
nor \U$2715 ( \4711 , \4709 , \4710 );
xnor \U$2716 ( \4712 , \4711 , \3063 );
xor \U$2717 ( \4713 , \4708 , \4712 );
xor \U$2718 ( \4714 , \4699 , \4713 );
nand \U$2719 ( \4715 , \3412 , \3035 );
xnor \U$2720 ( \4716 , \4715 , \3063 );
xor \U$2721 ( \4717 , \3063 , \4691 );
xor \U$2722 ( \4718 , \4717 , \4696 );
and \U$2723 ( \4719 , \4716 , \4718 );
nor \U$2724 ( \4720 , \4714 , \4719 );
and \U$2725 ( \4721 , \4703 , \4707 );
and \U$2726 ( \4722 , \4707 , \4712 );
and \U$2727 ( \4723 , \4703 , \4712 );
or \U$2728 ( \4724 , \4721 , \4722 , \4723 );
xor \U$2729 ( \4725 , \4434 , \4436 );
xor \U$2730 ( \4726 , \4724 , \4725 );
xor \U$2731 ( \4727 , \3121 , \4422 );
xor \U$2732 ( \4728 , \4727 , \4427 );
xor \U$2733 ( \4729 , \4726 , \4728 );
and \U$2734 ( \4730 , \4699 , \4713 );
nor \U$2735 ( \4731 , \4729 , \4730 );
nor \U$2736 ( \4732 , \4720 , \4731 );
xor \U$2737 ( \4733 , \4345 , \4349 );
xor \U$2738 ( \4734 , \4733 , \4354 );
xor \U$2739 ( \4735 , \4430 , \4437 );
xor \U$2740 ( \4736 , \4735 , \4442 );
xor \U$2741 ( \4737 , \4734 , \4736 );
and \U$2742 ( \4738 , \4724 , \4725 );
and \U$2743 ( \4739 , \4725 , \4728 );
and \U$2744 ( \4740 , \4724 , \4728 );
or \U$2745 ( \4741 , \4738 , \4739 , \4740 );
nor \U$2746 ( \4742 , \4737 , \4741 );
xor \U$2747 ( \4743 , \4445 , \4447 );
and \U$2748 ( \4744 , \4734 , \4736 );
nor \U$2749 ( \4745 , \4743 , \4744 );
nor \U$2750 ( \4746 , \4742 , \4745 );
nand \U$2751 ( \4747 , \4732 , \4746 );
and \U$2752 ( \4748 , \3235 , \2941 );
and \U$2753 ( \4749 , \3256 , \2938 );
nor \U$2754 ( \4750 , \4748 , \4749 );
xnor \U$2755 ( \4751 , \4750 , \2935 );
and \U$2756 ( \4752 , \3412 , \2977 );
and \U$2757 ( \4753 , \3279 , \2975 );
nor \U$2758 ( \4754 , \4752 , \4753 );
xnor \U$2759 ( \4755 , \4754 , \3003 );
xor \U$2760 ( \4756 , \4751 , \4755 );
and \U$2761 ( \4757 , \3279 , \2941 );
and \U$2762 ( \4758 , \3235 , \2938 );
nor \U$2763 ( \4759 , \4757 , \4758 );
xnor \U$2764 ( \4760 , \4759 , \2935 );
and \U$2765 ( \4761 , \4760 , \3003 );
nor \U$2766 ( \4762 , \4756 , \4761 );
xor \U$2767 ( \4763 , \4716 , \4718 );
and \U$2768 ( \4764 , \4751 , \4755 );
nor \U$2769 ( \4765 , \4763 , \4764 );
nor \U$2770 ( \4766 , \4762 , \4765 );
xor \U$2771 ( \4767 , \4760 , \3003 );
nand \U$2772 ( \4768 , \3412 , \2975 );
xnor \U$2773 ( \4769 , \4768 , \3003 );
nor \U$2774 ( \4770 , \4767 , \4769 );
and \U$2775 ( \4771 , \3412 , \2941 );
and \U$2776 ( \4772 , \3279 , \2938 );
nor \U$2777 ( \4773 , \4771 , \4772 );
xnor \U$2778 ( \4774 , \4773 , \2935 );
nand \U$2779 ( \4775 , \3412 , \2938 );
xnor \U$2780 ( \4776 , \4775 , \2935 );
and \U$2781 ( \4777 , \4776 , \2935 );
nand \U$2782 ( \4778 , \4774 , \4777 );
or \U$2783 ( \4779 , \4770 , \4778 );
nand \U$2784 ( \4780 , \4767 , \4769 );
nand \U$2785 ( \4781 , \4779 , \4780 );
and \U$2786 ( \4782 , \4766 , \4781 );
nand \U$2787 ( \4783 , \4756 , \4761 );
or \U$2788 ( \4784 , \4765 , \4783 );
nand \U$2789 ( \4785 , \4763 , \4764 );
nand \U$2790 ( \4786 , \4784 , \4785 );
nor \U$2791 ( \4787 , \4782 , \4786 );
or \U$2792 ( \4788 , \4747 , \4787 );
nand \U$2793 ( \4789 , \4714 , \4719 );
or \U$2794 ( \4790 , \4731 , \4789 );
nand \U$2795 ( \4791 , \4729 , \4730 );
nand \U$2796 ( \4792 , \4790 , \4791 );
and \U$2797 ( \4793 , \4746 , \4792 );
nand \U$2798 ( \4794 , \4737 , \4741 );
or \U$2799 ( \4795 , \4745 , \4794 );
nand \U$2800 ( \4796 , \4743 , \4744 );
nand \U$2801 ( \4797 , \4795 , \4796 );
nor \U$2802 ( \4798 , \4793 , \4797 );
nand \U$2803 ( \4799 , \4788 , \4798 );
and \U$2804 ( \4800 , \4687 , \4799 );
nand \U$2805 ( \4801 , \4418 , \4448 );
or \U$2806 ( \4802 , \4494 , \4801 );
nand \U$2807 ( \4803 , \4489 , \4493 );
nand \U$2808 ( \4804 , \4802 , \4803 );
and \U$2809 ( \4805 , \4602 , \4804 );
nand \U$2810 ( \4806 , \4544 , \4545 );
or \U$2811 ( \4807 , \4601 , \4806 );
nand \U$2812 ( \4808 , \4599 , \4600 );
nand \U$2813 ( \4809 , \4807 , \4808 );
nor \U$2814 ( \4810 , \4805 , \4809 );
or \U$2815 ( \4811 , \4686 , \4810 );
nand \U$2816 ( \4812 , \4638 , \4639 );
or \U$2817 ( \4813 , \4661 , \4812 );
nand \U$2818 ( \4814 , \4656 , \4660 );
nand \U$2819 ( \4815 , \4813 , \4814 );
and \U$2820 ( \4816 , \4685 , \4815 );
nand \U$2821 ( \4817 , \4672 , \4676 );
or \U$2822 ( \4818 , \4684 , \4817 );
nand \U$2823 ( \4819 , \4679 , \4683 );
nand \U$2824 ( \4820 , \4818 , \4819 );
nor \U$2825 ( \4821 , \4816 , \4820 );
nand \U$2826 ( \4822 , \4811 , \4821 );
nor \U$2827 ( \4823 , \4800 , \4822 );
or \U$2828 ( \4824 , \4341 , \4823 );
nand \U$2829 ( \4825 , \3463 , \3519 );
or \U$2830 ( \4826 , \3595 , \4825 );
nand \U$2831 ( \4827 , \3593 , \3594 );
nand \U$2832 ( \4828 , \4826 , \4827 );
and \U$2833 ( \4829 , \3748 , \4828 );
nand \U$2834 ( \4830 , \3670 , \3671 );
or \U$2835 ( \4831 , \3747 , \4830 );
nand \U$2836 ( \4832 , \3742 , \3746 );
nand \U$2837 ( \4833 , \4831 , \4832 );
nor \U$2838 ( \4834 , \4829 , \4833 );
or \U$2839 ( \4835 , \4044 , \4834 );
nand \U$2840 ( \4836 , \3819 , \3823 );
or \U$2841 ( \4837 , \3900 , \4836 );
nand \U$2842 ( \4838 , \3895 , \3899 );
nand \U$2843 ( \4839 , \4837 , \4838 );
and \U$2844 ( \4840 , \4043 , \4839 );
nand \U$2845 ( \4841 , \3968 , \3972 );
or \U$2846 ( \4842 , \4042 , \4841 );
nand \U$2847 ( \4843 , \4037 , \4041 );
nand \U$2848 ( \4844 , \4842 , \4843 );
nor \U$2849 ( \4845 , \4840 , \4844 );
nand \U$2850 ( \4846 , \4835 , \4845 );
and \U$2851 ( \4847 , \4340 , \4846 );
nand \U$2852 ( \4848 , \4101 , \4105 );
or \U$2853 ( \4849 , \4166 , \4848 );
nand \U$2854 ( \4850 , \4161 , \4165 );
nand \U$2855 ( \4851 , \4849 , \4850 );
and \U$2856 ( \4852 , \4262 , \4851 );
nand \U$2857 ( \4853 , \4218 , \4222 );
or \U$2858 ( \4854 , \4261 , \4853 );
nand \U$2859 ( \4855 , \4256 , \4260 );
nand \U$2860 ( \4856 , \4854 , \4855 );
nor \U$2861 ( \4857 , \4852 , \4856 );
or \U$2862 ( \4858 , \4339 , \4857 );
nand \U$2863 ( \4859 , \4288 , \4292 );
or \U$2864 ( \4860 , \4314 , \4859 );
nand \U$2865 ( \4861 , \4309 , \4313 );
nand \U$2866 ( \4862 , \4860 , \4861 );
and \U$2867 ( \4863 , \4338 , \4862 );
nand \U$2868 ( \4864 , \4325 , \4329 );
or \U$2869 ( \4865 , \4337 , \4864 );
nand \U$2870 ( \4866 , \4332 , \4336 );
nand \U$2871 ( \4867 , \4865 , \4866 );
nor \U$2872 ( \4868 , \4863 , \4867 );
nand \U$2873 ( \4869 , \4858 , \4868 );
nor \U$2874 ( \4870 , \4847 , \4869 );
nand \U$2875 ( \4871 , \4824 , \4870 );
not \U$2876 ( \4872 , \4871 );
xor \U$2877 ( \4873 , \2931 , \4872 );
buf \U$2878 ( \4874 , \4873 );
buf \U$2883 ( \4875 , RI2b5e785ebcf0_2);
buf \U$2884 ( \4876 , RI2b5e785ebc78_3);
buf \U$2885 ( \4877 , RI2b5e785ebc00_4);
buf \U$2886 ( \4878 , RI2b5e785ebb88_5);
buf \U$2887 ( \4879 , RI2b5e785ebb10_6);
buf \U$2888 ( \4880 , RI2b5e785eba98_7);
buf \U$2889 ( \4881 , RI2b5e785eba20_8);
buf \U$2890 ( \4882 , RI2b5e785eb9a8_9);
buf \U$2891 ( \4883 , RI2b5e785eb930_10);
buf \U$2892 ( \4884 , RI2b5e785eb8b8_11);
buf \U$2893 ( \4885 , RI2b5e785eb840_12);
and \U$2894 ( \4886 , \4884 , \4885 );
and \U$2895 ( \4887 , \4883 , \4886 );
and \U$2896 ( \4888 , \4882 , \4887 );
and \U$2897 ( \4889 , \4881 , \4888 );
and \U$2898 ( \4890 , \4880 , \4889 );
and \U$2899 ( \4891 , \4879 , \4890 );
and \U$2900 ( \4892 , \4878 , \4891 );
and \U$2901 ( \4893 , \4877 , \4892 );
and \U$2902 ( \4894 , \4876 , \4893 );
xor \U$2903 ( \4895 , \4875 , \4894 );
buf \U$2904 ( \4896 , \4895 );
buf \U$2905 ( \4897 , \4896 );
buf \U$2906 ( \4898 , RI2b5e785ae9b8_600);
buf \U$2907 ( \4899 , RI2b5e785aeb98_596);
buf \U$2908 ( \4900 , RI2b5e785aec10_595);
buf \U$2909 ( \4901 , RI2b5e785aec88_594);
buf \U$2910 ( \4902 , RI2b5e785aed00_593);
buf \U$2911 ( \4903 , RI2b5e785aed78_592);
buf \U$2912 ( \4904 , RI2b5e785aedf0_591);
buf \U$2913 ( \4905 , RI2b5e785aee68_590);
buf \U$2914 ( \4906 , RI2b5e785aeee0_589);
buf \U$2915 ( \4907 , RI2b5e785aef58_588);
buf \U$2916 ( \4908 , RI2b5e785ae9b8_600);
buf \U$2917 ( \4909 , RI2b5e785aea30_599);
buf \U$2918 ( \4910 , RI2b5e785aeaa8_598);
buf \U$2919 ( \4911 , RI2b5e785aeb20_597);
and \U$2920 ( \4912 , \4908 , \4909 , \4910 , \4911 );
nor \U$2921 ( \4913 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4912 );
buf \U$2922 ( \4914 , \4913 );
buf \U$2923 ( \4915 , \4914 );
xor \U$2924 ( \4916 , \4898 , \4915 );
buf \U$2925 ( \4917 , \4916 );
buf \U$2926 ( \4918 , RI2b5e785aea30_599);
and \U$2927 ( \4919 , \4898 , \4915 );
xor \U$2928 ( \4920 , \4918 , \4919 );
buf \U$2929 ( \4921 , \4920 );
buf \U$2930 ( \4922 , RI2b5e785aeaa8_598);
and \U$2931 ( \4923 , \4918 , \4919 );
xor \U$2932 ( \4924 , \4922 , \4923 );
buf \U$2933 ( \4925 , \4924 );
buf \U$2934 ( \4926 , RI2b5e785aeb20_597);
and \U$2935 ( \4927 , \4922 , \4923 );
xor \U$2936 ( \4928 , \4926 , \4927 );
buf \U$2937 ( \4929 , \4928 );
buf \U$2938 ( \4930 , RI2b5e785aeb98_596);
and \U$2939 ( \4931 , \4926 , \4927 );
xor \U$2940 ( \4932 , \4930 , \4931 );
buf \U$2941 ( \4933 , \4932 );
not \U$2942 ( \4934 , \4933 );
nor \U$2943 ( \4935 , \4917 , \4921 , \4925 , \4929 , \4934 );
and \U$2944 ( \4936 , RI2b5e785daa40_28, \4935 );
and \U$2945 ( \4937 , \4917 , \4921 , \4925 , \4929 , \4934 );
and \U$2946 ( \4938 , RI2b5e78549540_41, \4937 );
not \U$2947 ( \4939 , \4917 );
and \U$2948 ( \4940 , \4939 , \4921 , \4925 , \4929 , \4934 );
and \U$2949 ( \4941 , RI2b5e785388a8_54, \4940 );
not \U$2950 ( \4942 , \4921 );
and \U$2951 ( \4943 , \4917 , \4942 , \4925 , \4929 , \4934 );
and \U$2952 ( \4944 , RI2b5e784a6330_67, \4943 );
and \U$2953 ( \4945 , \4939 , \4942 , \4925 , \4929 , \4934 );
and \U$2954 ( \4946 , RI2b5e78495698_80, \4945 );
not \U$2955 ( \4947 , \4925 );
and \U$2956 ( \4948 , \4917 , \4921 , \4947 , \4929 , \4934 );
and \U$2957 ( \4949 , RI2b5e78495080_93, \4948 );
and \U$2958 ( \4950 , \4939 , \4921 , \4947 , \4929 , \4934 );
and \U$2959 ( \4951 , RI2b5e78403b80_106, \4950 );
and \U$2960 ( \4952 , \4917 , \4942 , \4947 , \4929 , \4934 );
and \U$2961 ( \4953 , RI2b5e775b1e60_119, \4952 );
and \U$2962 ( \4954 , \4939 , \4942 , \4947 , \4929 , \4934 );
and \U$2963 ( \4955 , RI2b5e7750bdf8_132, \4954 );
nor \U$2964 ( \4956 , \4939 , \4942 , \4947 , \4929 , \4933 );
and \U$2965 ( \4957 , RI2b5e774ff5d0_145, \4956 );
nor \U$2966 ( \4958 , \4917 , \4942 , \4947 , \4929 , \4933 );
and \U$2967 ( \4959 , RI2b5e774f65e8_158, \4958 );
nor \U$2968 ( \4960 , \4939 , \4921 , \4947 , \4929 , \4933 );
and \U$2969 ( \4961 , RI2b5e774eabd0_171, \4960 );
nor \U$2970 ( \4962 , \4917 , \4921 , \4947 , \4929 , \4933 );
and \U$2971 ( \4963 , RI2b5e774de3a8_184, \4962 );
nor \U$2972 ( \4964 , \4939 , \4942 , \4925 , \4929 , \4933 );
and \U$2973 ( \4965 , RI2b5e774d53c0_197, \4964 );
nor \U$2974 ( \4966 , \4917 , \4942 , \4925 , \4929 , \4933 );
and \U$2975 ( \4967 , RI2b5e785f4300_210, \4966 );
nor \U$2976 ( \4968 , \4939 , \4921 , \4925 , \4929 , \4933 );
and \U$2977 ( \4969 , RI2b5e785f3ce8_223, \4968 );
nor \U$2978 ( \4970 , \4917 , \4921 , \4925 , \4929 , \4933 );
and \U$2979 ( \4971 , RI2b5e785eb0c0_236, \4970 );
or \U$2980 ( \4972 , \4936 , \4938 , \4941 , \4944 , \4946 , \4949 , \4951 , \4953 , \4955 , \4957 , \4959 , \4961 , \4963 , \4965 , \4967 , \4969 , \4971 );
buf \U$2981 ( \4973 , \4933 );
buf \U$2982 ( \4974 , \4917 );
buf \U$2983 ( \4975 , \4921 );
buf \U$2984 ( \4976 , \4925 );
buf \U$2985 ( \4977 , \4929 );
or \U$2986 ( \4978 , \4974 , \4975 , \4976 , \4977 );
and \U$2987 ( \4979 , \4973 , \4978 );
buf \U$2988 ( \4980 , \4979 );
_DC r20e2 ( \4981_nR20e2 , \4972 , \4980 );
buf \U$2989 ( \4982 , \4981_nR20e2 );
not \U$2990 ( \4983 , \4982 );
xor \U$2991 ( \4984 , \4897 , \4983 );
xor \U$2992 ( \4985 , \4876 , \4893 );
buf \U$2993 ( \4986 , \4985 );
buf \U$2994 ( \4987 , \4986 );
and \U$2995 ( \4988 , RI2b5e785da9c8_29, \4935 );
and \U$2996 ( \4989 , RI2b5e785494c8_42, \4937 );
and \U$2997 ( \4990 , RI2b5e78538830_55, \4940 );
and \U$2998 ( \4991 , RI2b5e784a62b8_68, \4943 );
and \U$2999 ( \4992 , RI2b5e78495620_81, \4945 );
and \U$3000 ( \4993 , RI2b5e78495008_94, \4948 );
and \U$3001 ( \4994 , RI2b5e78403b08_107, \4950 );
and \U$3002 ( \4995 , RI2b5e775b1de8_120, \4952 );
and \U$3003 ( \4996 , RI2b5e7750bd80_133, \4954 );
and \U$3004 ( \4997 , RI2b5e774ff558_146, \4956 );
and \U$3005 ( \4998 , RI2b5e774f6570_159, \4958 );
and \U$3006 ( \4999 , RI2b5e774eab58_172, \4960 );
and \U$3007 ( \5000 , RI2b5e774de330_185, \4962 );
and \U$3008 ( \5001 , RI2b5e774d5348_198, \4964 );
and \U$3009 ( \5002 , RI2b5e785f4288_211, \4966 );
and \U$3010 ( \5003 , RI2b5e785f3658_224, \4968 );
and \U$3011 ( \5004 , RI2b5e785eb048_237, \4970 );
or \U$3012 ( \5005 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 );
_DC r20be ( \5006_nR20be , \5005 , \4980 );
buf \U$3013 ( \5007 , \5006_nR20be );
not \U$3014 ( \5008 , \5007 );
and \U$3015 ( \5009 , \4987 , \5008 );
xor \U$3016 ( \5010 , \4877 , \4892 );
buf \U$3017 ( \5011 , \5010 );
buf \U$3018 ( \5012 , \5011 );
and \U$3019 ( \5013 , RI2b5e785da950_30, \4935 );
and \U$3020 ( \5014 , RI2b5e78549450_43, \4937 );
and \U$3021 ( \5015 , RI2b5e785387b8_56, \4940 );
and \U$3022 ( \5016 , RI2b5e784a6240_69, \4943 );
and \U$3023 ( \5017 , RI2b5e784955a8_82, \4945 );
and \U$3024 ( \5018 , RI2b5e78494f90_95, \4948 );
and \U$3025 ( \5019 , RI2b5e78403a90_108, \4950 );
and \U$3026 ( \5020 , RI2b5e775b1d70_121, \4952 );
and \U$3027 ( \5021 , RI2b5e7750bd08_134, \4954 );
and \U$3028 ( \5022 , RI2b5e774ff4e0_147, \4956 );
and \U$3029 ( \5023 , RI2b5e774f64f8_160, \4958 );
and \U$3030 ( \5024 , RI2b5e774eaae0_173, \4960 );
and \U$3031 ( \5025 , RI2b5e774de2b8_186, \4962 );
and \U$3032 ( \5026 , RI2b5e774d52d0_199, \4964 );
and \U$3033 ( \5027 , RI2b5e785f4210_212, \4966 );
and \U$3034 ( \5028 , RI2b5e785eb5e8_225, \4968 );
and \U$3035 ( \5029 , RI2b5e785e6c50_238, \4970 );
or \U$3036 ( \5030 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 );
_DC r1f2b ( \5031_nR1f2b , \5030 , \4980 );
buf \U$3037 ( \5032 , \5031_nR1f2b );
not \U$3038 ( \5033 , \5032 );
and \U$3039 ( \5034 , \5012 , \5033 );
xor \U$3040 ( \5035 , \4878 , \4891 );
buf \U$3041 ( \5036 , \5035 );
buf \U$3042 ( \5037 , \5036 );
and \U$3043 ( \5038 , RI2b5e785da8d8_31, \4935 );
and \U$3044 ( \5039 , RI2b5e785493d8_44, \4937 );
and \U$3045 ( \5040 , RI2b5e78538740_57, \4940 );
and \U$3046 ( \5041 , RI2b5e784a61c8_70, \4943 );
and \U$3047 ( \5042 , RI2b5e78495530_83, \4945 );
and \U$3048 ( \5043 , RI2b5e78494f18_96, \4948 );
and \U$3049 ( \5044 , RI2b5e78403a18_109, \4950 );
and \U$3050 ( \5045 , RI2b5e775b1cf8_122, \4952 );
and \U$3051 ( \5046 , RI2b5e7750bc90_135, \4954 );
and \U$3052 ( \5047 , RI2b5e774ff468_148, \4956 );
and \U$3053 ( \5048 , RI2b5e774f6480_161, \4958 );
and \U$3054 ( \5049 , RI2b5e774eaa68_174, \4960 );
and \U$3055 ( \5050 , RI2b5e774de240_187, \4962 );
and \U$3056 ( \5051 , RI2b5e774d5258_200, \4964 );
and \U$3057 ( \5052 , RI2b5e785f4198_213, \4966 );
and \U$3058 ( \5053 , RI2b5e785eb570_226, \4968 );
and \U$3059 ( \5054 , RI2b5e785e6bd8_239, \4970 );
or \U$3060 ( \5055 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 );
_DC r1f07 ( \5056_nR1f07 , \5055 , \4980 );
buf \U$3061 ( \5057 , \5056_nR1f07 );
not \U$3062 ( \5058 , \5057 );
and \U$3063 ( \5059 , \5037 , \5058 );
xor \U$3064 ( \5060 , \4879 , \4890 );
buf \U$3065 ( \5061 , \5060 );
buf \U$3066 ( \5062 , \5061 );
and \U$3067 ( \5063 , RI2b5e785da860_32, \4935 );
and \U$3068 ( \5064 , RI2b5e78549360_45, \4937 );
and \U$3069 ( \5065 , RI2b5e785386c8_58, \4940 );
and \U$3070 ( \5066 , RI2b5e784a6150_71, \4943 );
and \U$3071 ( \5067 , RI2b5e784954b8_84, \4945 );
and \U$3072 ( \5068 , RI2b5e78494ea0_97, \4948 );
and \U$3073 ( \5069 , RI2b5e784039a0_110, \4950 );
and \U$3074 ( \5070 , RI2b5e775b1c80_123, \4952 );
and \U$3075 ( \5071 , RI2b5e7750bc18_136, \4954 );
and \U$3076 ( \5072 , RI2b5e774ff3f0_149, \4956 );
and \U$3077 ( \5073 , RI2b5e774f6408_162, \4958 );
and \U$3078 ( \5074 , RI2b5e774ea9f0_175, \4960 );
and \U$3079 ( \5075 , RI2b5e774de1c8_188, \4962 );
and \U$3080 ( \5076 , RI2b5e774d51e0_201, \4964 );
and \U$3081 ( \5077 , RI2b5e785f4120_214, \4966 );
and \U$3082 ( \5078 , RI2b5e785eb4f8_227, \4968 );
and \U$3083 ( \5079 , RI2b5e785e64d0_240, \4970 );
or \U$3084 ( \5080 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 );
_DC r1d88 ( \5081_nR1d88 , \5080 , \4980 );
buf \U$3085 ( \5082 , \5081_nR1d88 );
not \U$3086 ( \5083 , \5082 );
and \U$3087 ( \5084 , \5062 , \5083 );
xor \U$3088 ( \5085 , \4880 , \4889 );
buf \U$3089 ( \5086 , \5085 );
buf \U$3090 ( \5087 , \5086 );
and \U$3091 ( \5088 , RI2b5e78549900_33, \4935 );
and \U$3092 ( \5089 , RI2b5e78538c68_46, \4937 );
and \U$3093 ( \5090 , RI2b5e78538650_59, \4940 );
and \U$3094 ( \5091 , RI2b5e784a60d8_72, \4943 );
and \U$3095 ( \5092 , RI2b5e78495440_85, \4945 );
and \U$3096 ( \5093 , RI2b5e78494e28_98, \4948 );
and \U$3097 ( \5094 , RI2b5e78403928_111, \4950 );
and \U$3098 ( \5095 , RI2b5e775b1c08_124, \4952 );
and \U$3099 ( \5096 , RI2b5e7750bba0_137, \4954 );
and \U$3100 ( \5097 , RI2b5e774ff378_150, \4956 );
and \U$3101 ( \5098 , RI2b5e774f6390_163, \4958 );
and \U$3102 ( \5099 , RI2b5e774ea978_176, \4960 );
and \U$3103 ( \5100 , RI2b5e774de150_189, \4962 );
and \U$3104 ( \5101 , RI2b5e774d5168_202, \4964 );
and \U$3105 ( \5102 , RI2b5e785f40a8_215, \4966 );
and \U$3106 ( \5103 , RI2b5e785eb480_228, \4968 );
and \U$3107 ( \5104 , RI2b5e785da608_241, \4970 );
or \U$3108 ( \5105 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 );
_DC r1d64 ( \5106_nR1d64 , \5105 , \4980 );
buf \U$3109 ( \5107 , \5106_nR1d64 );
not \U$3110 ( \5108 , \5107 );
and \U$3111 ( \5109 , \5087 , \5108 );
xor \U$3112 ( \5110 , \4881 , \4888 );
buf \U$3113 ( \5111 , \5110 );
buf \U$3114 ( \5112 , \5111 );
and \U$3115 ( \5113 , RI2b5e78549888_34, \4935 );
and \U$3116 ( \5114 , RI2b5e78538bf0_47, \4937 );
and \U$3117 ( \5115 , RI2b5e785385d8_60, \4940 );
and \U$3118 ( \5116 , RI2b5e784a6060_73, \4943 );
and \U$3119 ( \5117 , RI2b5e784953c8_86, \4945 );
and \U$3120 ( \5118 , RI2b5e78403ec8_99, \4948 );
and \U$3121 ( \5119 , RI2b5e775b21a8_112, \4950 );
and \U$3122 ( \5120 , RI2b5e775b1b90_125, \4952 );
and \U$3123 ( \5121 , RI2b5e7750bb28_138, \4954 );
and \U$3124 ( \5122 , RI2b5e774ff300_151, \4956 );
and \U$3125 ( \5123 , RI2b5e774f6318_164, \4958 );
and \U$3126 ( \5124 , RI2b5e774ea900_177, \4960 );
and \U$3127 ( \5125 , RI2b5e774de0d8_190, \4962 );
and \U$3128 ( \5126 , RI2b5e774d50f0_203, \4964 );
and \U$3129 ( \5127 , RI2b5e785f4030_216, \4966 );
and \U$3130 ( \5128 , RI2b5e785eb408_229, \4968 );
and \U$3131 ( \5129 , RI2b5e785da590_242, \4970 );
or \U$3132 ( \5130 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 );
_DC r1c19 ( \5131_nR1c19 , \5130 , \4980 );
buf \U$3133 ( \5132 , \5131_nR1c19 );
not \U$3134 ( \5133 , \5132 );
and \U$3135 ( \5134 , \5112 , \5133 );
xor \U$3136 ( \5135 , \4882 , \4887 );
buf \U$3137 ( \5136 , \5135 );
buf \U$3138 ( \5137 , \5136 );
and \U$3139 ( \5138 , RI2b5e78549810_35, \4935 );
and \U$3140 ( \5139 , RI2b5e78538b78_48, \4937 );
and \U$3141 ( \5140 , RI2b5e78538560_61, \4940 );
and \U$3142 ( \5141 , RI2b5e784a5fe8_74, \4943 );
and \U$3143 ( \5142 , RI2b5e78495350_87, \4945 );
and \U$3144 ( \5143 , RI2b5e78403e50_100, \4948 );
and \U$3145 ( \5144 , RI2b5e775b2130_113, \4950 );
and \U$3146 ( \5145 , RI2b5e775b1b18_126, \4952 );
and \U$3147 ( \5146 , RI2b5e7750bab0_139, \4954 );
and \U$3148 ( \5147 , RI2b5e774ff288_152, \4956 );
and \U$3149 ( \5148 , RI2b5e774f62a0_165, \4958 );
and \U$3150 ( \5149 , RI2b5e774ea888_178, \4960 );
and \U$3151 ( \5150 , RI2b5e774de060_191, \4962 );
and \U$3152 ( \5151 , RI2b5e774d5078_204, \4964 );
and \U$3153 ( \5152 , RI2b5e785f3fb8_217, \4966 );
and \U$3154 ( \5153 , RI2b5e785eb390_230, \4968 );
and \U$3155 ( \5154 , RI2b5e785da518_243, \4970 );
or \U$3156 ( \5155 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 );
_DC r1bf5 ( \5156_nR1bf5 , \5155 , \4980 );
buf \U$3157 ( \5157 , \5156_nR1bf5 );
not \U$3158 ( \5158 , \5157 );
and \U$3159 ( \5159 , \5137 , \5158 );
xor \U$3160 ( \5160 , \4883 , \4886 );
buf \U$3161 ( \5161 , \5160 );
buf \U$3162 ( \5162 , \5161 );
and \U$3163 ( \5163 , RI2b5e78549798_36, \4935 );
and \U$3164 ( \5164 , RI2b5e78538b00_49, \4937 );
and \U$3165 ( \5165 , RI2b5e785384e8_62, \4940 );
and \U$3166 ( \5166 , RI2b5e784a5f70_75, \4943 );
and \U$3167 ( \5167 , RI2b5e784952d8_88, \4945 );
and \U$3168 ( \5168 , RI2b5e78403dd8_101, \4948 );
and \U$3169 ( \5169 , RI2b5e775b20b8_114, \4950 );
and \U$3170 ( \5170 , RI2b5e775b1aa0_127, \4952 );
and \U$3171 ( \5171 , RI2b5e7750ba38_140, \4954 );
and \U$3172 ( \5172 , RI2b5e774ff210_153, \4956 );
and \U$3173 ( \5173 , RI2b5e774f6228_166, \4958 );
and \U$3174 ( \5174 , RI2b5e774ea810_179, \4960 );
and \U$3175 ( \5175 , RI2b5e774ddfe8_192, \4962 );
and \U$3176 ( \5176 , RI2b5e774d5000_205, \4964 );
and \U$3177 ( \5177 , RI2b5e785f3f40_218, \4966 );
and \U$3178 ( \5178 , RI2b5e785eb318_231, \4968 );
and \U$3179 ( \5179 , RI2b5e785da4a0_244, \4970 );
or \U$3180 ( \5180 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 );
_DC r1ada ( \5181_nR1ada , \5180 , \4980 );
buf \U$3181 ( \5182 , \5181_nR1ada );
not \U$3182 ( \5183 , \5182 );
and \U$3183 ( \5184 , \5162 , \5183 );
xor \U$3184 ( \5185 , \4884 , \4885 );
buf \U$3185 ( \5186 , \5185 );
buf \U$3186 ( \5187 , \5186 );
and \U$3187 ( \5188 , RI2b5e78549720_37, \4935 );
and \U$3188 ( \5189 , RI2b5e78538a88_50, \4937 );
and \U$3189 ( \5190 , RI2b5e78538470_63, \4940 );
and \U$3190 ( \5191 , RI2b5e784a5ef8_76, \4943 );
and \U$3191 ( \5192 , RI2b5e78495260_89, \4945 );
and \U$3192 ( \5193 , RI2b5e78403d60_102, \4948 );
and \U$3193 ( \5194 , RI2b5e775b2040_115, \4950 );
and \U$3194 ( \5195 , RI2b5e775b1a28_128, \4952 );
and \U$3195 ( \5196 , RI2b5e7750b9c0_141, \4954 );
and \U$3196 ( \5197 , RI2b5e774ff198_154, \4956 );
and \U$3197 ( \5198 , RI2b5e774f61b0_167, \4958 );
and \U$3198 ( \5199 , RI2b5e774ea798_180, \4960 );
and \U$3199 ( \5200 , RI2b5e774ddf70_193, \4962 );
and \U$3200 ( \5201 , RI2b5e774d4f88_206, \4964 );
and \U$3201 ( \5202 , RI2b5e785f3ec8_219, \4966 );
and \U$3202 ( \5203 , RI2b5e785eb2a0_232, \4968 );
and \U$3203 ( \5204 , RI2b5e785da428_245, \4970 );
or \U$3204 ( \5205 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 );
_DC r1af3 ( \5206_nR1af3 , \5205 , \4980 );
buf \U$3205 ( \5207 , \5206_nR1af3 );
not \U$3206 ( \5208 , \5207 );
and \U$3207 ( \5209 , \5187 , \5208 );
not \U$3208 ( \5210 , \4885 );
buf \U$3209 ( \5211 , \5210 );
buf \U$3210 ( \5212 , \5211 );
and \U$3211 ( \5213 , RI2b5e785496a8_38, \4935 );
and \U$3212 ( \5214 , RI2b5e78538a10_51, \4937 );
and \U$3213 ( \5215 , RI2b5e785383f8_64, \4940 );
and \U$3214 ( \5216 , RI2b5e784a5e80_77, \4943 );
and \U$3215 ( \5217 , RI2b5e784951e8_90, \4945 );
and \U$3216 ( \5218 , RI2b5e78403ce8_103, \4948 );
and \U$3217 ( \5219 , RI2b5e775b1fc8_116, \4950 );
and \U$3218 ( \5220 , RI2b5e775b19b0_129, \4952 );
and \U$3219 ( \5221 , RI2b5e7750b948_142, \4954 );
and \U$3220 ( \5222 , RI2b5e774ff120_155, \4956 );
and \U$3221 ( \5223 , RI2b5e774f6138_168, \4958 );
and \U$3222 ( \5224 , RI2b5e774ea720_181, \4960 );
and \U$3223 ( \5225 , RI2b5e774ddef8_194, \4962 );
and \U$3224 ( \5226 , RI2b5e774d4f10_207, \4964 );
and \U$3225 ( \5227 , RI2b5e785f3e50_220, \4966 );
and \U$3226 ( \5228 , RI2b5e785eb228_233, \4968 );
and \U$3227 ( \5229 , RI2b5e785da3b0_246, \4970 );
or \U$3228 ( \5230 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 );
_DC r19f0 ( \5231_nR19f0 , \5230 , \4980 );
buf \U$3229 ( \5232 , \5231_nR19f0 );
not \U$3230 ( \5233 , \5232 );
and \U$3231 ( \5234 , \5212 , \5233 );
buf \U$3232 ( \5235 , RI2b5e785db148_13);
buf \U$3235 ( \5236 , \5235 );
and \U$3236 ( \5237 , RI2b5e78549630_39, \4935 );
and \U$3237 ( \5238 , RI2b5e78538998_52, \4937 );
and \U$3238 ( \5239 , RI2b5e78538380_65, \4940 );
and \U$3239 ( \5240 , RI2b5e784a5e08_78, \4943 );
and \U$3240 ( \5241 , RI2b5e78495170_91, \4945 );
and \U$3241 ( \5242 , RI2b5e78403c70_104, \4948 );
and \U$3242 ( \5243 , RI2b5e775b1f50_117, \4950 );
and \U$3243 ( \5244 , RI2b5e775b1938_130, \4952 );
and \U$3244 ( \5245 , RI2b5e7750b8d0_143, \4954 );
and \U$3245 ( \5246 , RI2b5e774ff0a8_156, \4956 );
and \U$3246 ( \5247 , RI2b5e774f60c0_169, \4958 );
and \U$3247 ( \5248 , RI2b5e774ea6a8_182, \4960 );
and \U$3248 ( \5249 , RI2b5e774dde80_195, \4962 );
and \U$3249 ( \5250 , RI2b5e774d4e98_208, \4964 );
and \U$3250 ( \5251 , RI2b5e785f3dd8_221, \4966 );
and \U$3251 ( \5252 , RI2b5e785eb1b0_234, \4968 );
and \U$3252 ( \5253 , RI2b5e785da338_247, \4970 );
or \U$3253 ( \5254 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 );
_DC r19d4 ( \5255_nR19d4 , \5254 , \4980 );
buf \U$3254 ( \5256 , \5255_nR19d4 );
not \U$3255 ( \5257 , \5256 );
or \U$3256 ( \5258 , \5236 , \5257 );
and \U$3257 ( \5259 , \5233 , \5258 );
and \U$3258 ( \5260 , \5212 , \5258 );
or \U$3259 ( \5261 , \5234 , \5259 , \5260 );
and \U$3260 ( \5262 , \5208 , \5261 );
and \U$3261 ( \5263 , \5187 , \5261 );
or \U$3262 ( \5264 , \5209 , \5262 , \5263 );
and \U$3263 ( \5265 , \5183 , \5264 );
and \U$3264 ( \5266 , \5162 , \5264 );
or \U$3265 ( \5267 , \5184 , \5265 , \5266 );
and \U$3266 ( \5268 , \5158 , \5267 );
and \U$3267 ( \5269 , \5137 , \5267 );
or \U$3268 ( \5270 , \5159 , \5268 , \5269 );
and \U$3269 ( \5271 , \5133 , \5270 );
and \U$3270 ( \5272 , \5112 , \5270 );
or \U$3271 ( \5273 , \5134 , \5271 , \5272 );
and \U$3272 ( \5274 , \5108 , \5273 );
and \U$3273 ( \5275 , \5087 , \5273 );
or \U$3274 ( \5276 , \5109 , \5274 , \5275 );
and \U$3275 ( \5277 , \5083 , \5276 );
and \U$3276 ( \5278 , \5062 , \5276 );
or \U$3277 ( \5279 , \5084 , \5277 , \5278 );
and \U$3278 ( \5280 , \5058 , \5279 );
and \U$3279 ( \5281 , \5037 , \5279 );
or \U$3280 ( \5282 , \5059 , \5280 , \5281 );
and \U$3281 ( \5283 , \5033 , \5282 );
and \U$3282 ( \5284 , \5012 , \5282 );
or \U$3283 ( \5285 , \5034 , \5283 , \5284 );
and \U$3284 ( \5286 , \5008 , \5285 );
and \U$3285 ( \5287 , \4987 , \5285 );
or \U$3286 ( \5288 , \5009 , \5286 , \5287 );
xor \U$3287 ( \5289 , \4984 , \5288 );
buf \U$3288 ( \5290 , \5289 );
buf \U$3289 ( \5291 , \5290 );
xor \U$3290 ( \5292 , \4987 , \5008 );
xor \U$3291 ( \5293 , \5292 , \5285 );
buf \U$3292 ( \5294 , \5293 );
buf \U$3293 ( \5295 , \5294 );
xor \U$3294 ( \5296 , \5012 , \5033 );
xor \U$3295 ( \5297 , \5296 , \5282 );
buf \U$3296 ( \5298 , \5297 );
buf \U$3297 ( \5299 , \5298 );
and \U$3298 ( \5300 , \5295 , \5299 );
not \U$3299 ( \5301 , \5300 );
and \U$3300 ( \5302 , \5291 , \5301 );
not \U$3301 ( \5303 , \5302 );
buf \U$3302 ( \5304 , \4917 );
buf \U$3303 ( \5305 , RI2b5e785aec10_595);
and \U$3304 ( \5306 , \4930 , \4931 );
xor \U$3305 ( \5307 , \5305 , \5306 );
buf \U$3306 ( \5308 , \5307 );
buf \U$3307 ( \5309 , \5308 );
buf \U$3308 ( \5310 , RI2b5e785aec88_594);
and \U$3309 ( \5311 , \5305 , \5306 );
xor \U$3310 ( \5312 , \5310 , \5311 );
buf \U$3311 ( \5313 , \5312 );
buf \U$3312 ( \5314 , \5313 );
buf \U$3313 ( \5315 , RI2b5e785aed00_593);
and \U$3314 ( \5316 , \5310 , \5311 );
xor \U$3315 ( \5317 , \5315 , \5316 );
buf \U$3316 ( \5318 , \5317 );
buf \U$3317 ( \5319 , \5318 );
buf \U$3318 ( \5320 , RI2b5e785aed78_592);
and \U$3319 ( \5321 , \5315 , \5316 );
xor \U$3320 ( \5322 , \5320 , \5321 );
buf \U$3321 ( \5323 , \5322 );
buf \U$3322 ( \5324 , \5323 );
buf \U$3323 ( \5325 , RI2b5e785aedf0_591);
and \U$3324 ( \5326 , \5320 , \5321 );
xor \U$3325 ( \5327 , \5325 , \5326 );
buf \U$3326 ( \5328 , \5327 );
buf \U$3327 ( \5329 , \5328 );
buf \U$3328 ( \5330 , RI2b5e785aee68_590);
and \U$3329 ( \5331 , \5325 , \5326 );
xor \U$3330 ( \5332 , \5330 , \5331 );
buf \U$3331 ( \5333 , \5332 );
buf \U$3332 ( \5334 , \5333 );
buf \U$3333 ( \5335 , RI2b5e785aeee0_589);
and \U$3334 ( \5336 , \5330 , \5331 );
xor \U$3335 ( \5337 , \5335 , \5336 );
buf \U$3336 ( \5338 , \5337 );
buf \U$3337 ( \5339 , \5338 );
buf \U$3338 ( \5340 , RI2b5e785aef58_588);
and \U$3339 ( \5341 , \5335 , \5336 );
xor \U$3340 ( \5342 , \5340 , \5341 );
buf \U$3341 ( \5343 , \5342 );
buf \U$3342 ( \5344 , \5343 );
buf \U$3343 ( \5345 , \4933 );
nor \U$3344 ( \5346 , \5309 , \5314 , \5319 , \5324 , \5329 , \5334 , \5339 , \5344 , \5345 );
buf \U$3345 ( \5347 , \5346 );
buf \U$3346 ( \5348 , \5347 );
xor \U$3347 ( \5349 , \5304 , \5348 );
buf \U$3348 ( \5350 , \5349 );
buf \U$3349 ( \5351 , \4921 );
and \U$3350 ( \5352 , \5304 , \5348 );
xor \U$3351 ( \5353 , \5351 , \5352 );
buf \U$3352 ( \5354 , \5353 );
buf \U$3353 ( \5355 , \4925 );
and \U$3354 ( \5356 , \5351 , \5352 );
xor \U$3355 ( \5357 , \5355 , \5356 );
buf \U$3356 ( \5358 , \5357 );
buf \U$3357 ( \5359 , \4929 );
and \U$3358 ( \5360 , \5355 , \5356 );
xor \U$3359 ( \5361 , \5359 , \5360 );
buf \U$3360 ( \5362 , \5361 );
buf \U$3361 ( \5363 , \4933 );
and \U$3362 ( \5364 , \5359 , \5360 );
xor \U$3363 ( \5365 , \5363 , \5364 );
buf \U$3364 ( \5366 , \5365 );
not \U$3365 ( \5367 , \5366 );
nor \U$3366 ( \5368 , \5350 , \5354 , \5358 , \5362 , \5367 );
and \U$3367 ( \5369 , RI2b5e785da248_249, \5368 );
and \U$3368 ( \5370 , \5350 , \5354 , \5358 , \5362 , \5367 );
and \U$3369 ( \5371 , RI2b5e785be750_269, \5370 );
not \U$3370 ( \5372 , \5350 );
and \U$3371 ( \5373 , \5372 , \5354 , \5358 , \5362 , \5367 );
and \U$3372 ( \5374 , RI2b5e785bc4a0_289, \5373 );
not \U$3373 ( \5375 , \5354 );
and \U$3374 ( \5376 , \5350 , \5375 , \5358 , \5362 , \5367 );
and \U$3375 ( \5377 , RI2b5e785bbb40_309, \5376 );
and \U$3376 ( \5378 , \5372 , \5375 , \5358 , \5362 , \5367 );
and \U$3377 ( \5379 , RI2b5e785b9c50_329, \5378 );
not \U$3378 ( \5380 , \5358 );
and \U$3379 ( \5381 , \5350 , \5354 , \5380 , \5362 , \5367 );
and \U$3380 ( \5382 , RI2b5e785b8120_349, \5381 );
and \U$3381 ( \5383 , \5372 , \5354 , \5380 , \5362 , \5367 );
and \U$3382 ( \5384 , RI2b5e785b77c0_369, \5383 );
and \U$3383 ( \5385 , \5350 , \5375 , \5380 , \5362 , \5367 );
and \U$3384 ( \5386 , RI2b5e785b6e60_389, \5385 );
and \U$3385 ( \5387 , \5372 , \5375 , \5380 , \5362 , \5367 );
and \U$3386 ( \5388 , RI2b5e785b56f0_409, \5387 );
nor \U$3387 ( \5389 , \5372 , \5375 , \5380 , \5362 , \5366 );
and \U$3388 ( \5390 , RI2b5e785b4d90_429, \5389 );
nor \U$3389 ( \5391 , \5350 , \5375 , \5380 , \5362 , \5366 );
and \U$3390 ( \5392 , RI2b5e785b39e0_449, \5391 );
nor \U$3391 ( \5393 , \5372 , \5354 , \5380 , \5362 , \5366 );
and \U$3392 ( \5394 , RI2b5e785b3080_469, \5393 );
nor \U$3393 ( \5395 , \5350 , \5354 , \5380 , \5362 , \5366 );
and \U$3394 ( \5396 , RI2b5e785b2720_489, \5395 );
nor \U$3395 ( \5397 , \5372 , \5375 , \5358 , \5362 , \5366 );
and \U$3396 ( \5398 , RI2b5e785b1730_509, \5397 );
nor \U$3397 ( \5399 , \5350 , \5375 , \5358 , \5362 , \5366 );
and \U$3398 ( \5400 , RI2b5e785b0dd0_529, \5399 );
nor \U$3399 ( \5401 , \5372 , \5354 , \5358 , \5362 , \5366 );
and \U$3400 ( \5402 , RI2b5e785b0470_549, \5401 );
nor \U$3401 ( \5403 , \5350 , \5354 , \5358 , \5362 , \5366 );
and \U$3402 ( \5404 , RI2b5e785af840_569, \5403 );
or \U$3403 ( \5405 , \5369 , \5371 , \5374 , \5377 , \5379 , \5382 , \5384 , \5386 , \5388 , \5390 , \5392 , \5394 , \5396 , \5398 , \5400 , \5402 , \5404 );
buf \U$3404 ( \5406 , \5366 );
buf \U$3405 ( \5407 , \5350 );
buf \U$3406 ( \5408 , \5354 );
buf \U$3407 ( \5409 , \5358 );
buf \U$3408 ( \5410 , \5362 );
or \U$3409 ( \5411 , \5407 , \5408 , \5409 , \5410 );
and \U$3410 ( \5412 , \5406 , \5411 );
buf \U$3411 ( \5413 , \5412 );
_DC r27bc ( \5414_nR27bc , \5405 , \5413 );
buf \U$3412 ( \5415 , \5414_nR27bc );
buf \U$3413 ( \5416 , RI2b5e785ebd68_1);
and \U$3414 ( \5417 , \4875 , \4894 );
and \U$3415 ( \5418 , \5416 , \5417 );
buf \U$3416 ( \5419 , \5418 );
buf \U$3417 ( \5420 , \5419 );
xor \U$3418 ( \5421 , \5416 , \5417 );
buf \U$3419 ( \5422 , \5421 );
buf \U$3420 ( \5423 , \5422 );
and \U$3421 ( \5424 , RI2b5e785daab8_27, \4935 );
and \U$3422 ( \5425 , RI2b5e785495b8_40, \4937 );
and \U$3423 ( \5426 , RI2b5e78538920_53, \4940 );
and \U$3424 ( \5427 , RI2b5e784a63a8_66, \4943 );
and \U$3425 ( \5428 , RI2b5e78495710_79, \4945 );
and \U$3426 ( \5429 , RI2b5e784950f8_92, \4948 );
and \U$3427 ( \5430 , RI2b5e78403bf8_105, \4950 );
and \U$3428 ( \5431 , RI2b5e775b1ed8_118, \4952 );
and \U$3429 ( \5432 , RI2b5e775b18c0_131, \4954 );
and \U$3430 ( \5433 , RI2b5e7750b858_144, \4956 );
and \U$3431 ( \5434 , RI2b5e774ff030_157, \4958 );
and \U$3432 ( \5435 , RI2b5e774f6048_170, \4960 );
and \U$3433 ( \5436 , RI2b5e774ea630_183, \4962 );
and \U$3434 ( \5437 , RI2b5e774dde08_196, \4964 );
and \U$3435 ( \5438 , RI2b5e774d4e20_209, \4966 );
and \U$3436 ( \5439 , RI2b5e785f3d60_222, \4968 );
and \U$3437 ( \5440 , RI2b5e785eb138_235, \4970 );
or \U$3438 ( \5441 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 );
_DC r229d ( \5442_nR229d , \5441 , \4980 );
buf \U$3439 ( \5443 , \5442_nR229d );
not \U$3440 ( \5444 , \5443 );
and \U$3441 ( \5445 , \5423 , \5444 );
and \U$3442 ( \5446 , \4897 , \4983 );
and \U$3443 ( \5447 , \4983 , \5288 );
and \U$3444 ( \5448 , \4897 , \5288 );
or \U$3445 ( \5449 , \5446 , \5447 , \5448 );
and \U$3446 ( \5450 , \5444 , \5449 );
and \U$3447 ( \5451 , \5423 , \5449 );
or \U$3448 ( \5452 , \5445 , \5450 , \5451 );
xnor \U$3449 ( \5453 , \5420 , \5452 );
buf \U$3450 ( \5454 , \5453 );
buf \U$3451 ( \5455 , \5454 );
xor \U$3452 ( \5456 , \5423 , \5444 );
xor \U$3453 ( \5457 , \5456 , \5449 );
buf \U$3454 ( \5458 , \5457 );
buf \U$3455 ( \5459 , \5458 );
xor \U$3456 ( \5460 , \5455 , \5459 );
xor \U$3457 ( \5461 , \5459 , \5291 );
not \U$3458 ( \5462 , \5461 );
and \U$3459 ( \5463 , \5460 , \5462 );
and \U$3460 ( \5464 , \5415 , \5463 );
and \U$3461 ( \5465 , RI2b5e785da2c0_248, \5368 );
and \U$3462 ( \5466 , RI2b5e785be7c8_268, \5370 );
and \U$3463 ( \5467 , RI2b5e785bc518_288, \5373 );
and \U$3464 ( \5468 , RI2b5e785bbbb8_308, \5376 );
and \U$3465 ( \5469 , RI2b5e785b9cc8_328, \5378 );
and \U$3466 ( \5470 , RI2b5e785b9368_348, \5381 );
and \U$3467 ( \5471 , RI2b5e785b7838_368, \5383 );
and \U$3468 ( \5472 , RI2b5e785b6ed8_388, \5385 );
and \U$3469 ( \5473 , RI2b5e785b5768_408, \5387 );
and \U$3470 ( \5474 , RI2b5e785b4e08_428, \5389 );
and \U$3471 ( \5475 , RI2b5e785b3a58_448, \5391 );
and \U$3472 ( \5476 , RI2b5e785b30f8_468, \5393 );
and \U$3473 ( \5477 , RI2b5e785b2798_488, \5395 );
and \U$3474 ( \5478 , RI2b5e785b17a8_508, \5397 );
and \U$3475 ( \5479 , RI2b5e785b0e48_528, \5399 );
and \U$3476 ( \5480 , RI2b5e785b04e8_548, \5401 );
and \U$3477 ( \5481 , RI2b5e785afb88_568, \5403 );
or \U$3478 ( \5482 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 );
_DC r28b1 ( \5483_nR28b1 , \5482 , \5413 );
buf \U$3479 ( \5484 , \5483_nR28b1 );
and \U$3480 ( \5485 , \5484 , \5461 );
nor \U$3481 ( \5486 , \5464 , \5485 );
and \U$3482 ( \5487 , \5459 , \5291 );
not \U$3483 ( \5488 , \5487 );
and \U$3484 ( \5489 , \5455 , \5488 );
xnor \U$3485 ( \5490 , \5486 , \5489 );
xor \U$3486 ( \5491 , \5303 , \5490 );
and \U$3488 ( \5492 , RI2b5e785da1d0_250, \5368 );
and \U$3489 ( \5493 , RI2b5e785be6d8_270, \5370 );
and \U$3490 ( \5494 , RI2b5e785bc428_290, \5373 );
and \U$3491 ( \5495 , RI2b5e785bbac8_310, \5376 );
and \U$3492 ( \5496 , RI2b5e785b9bd8_330, \5378 );
and \U$3493 ( \5497 , RI2b5e785b80a8_350, \5381 );
and \U$3494 ( \5498 , RI2b5e785b7748_370, \5383 );
and \U$3495 ( \5499 , RI2b5e785b6de8_390, \5385 );
and \U$3496 ( \5500 , RI2b5e785b5678_410, \5387 );
and \U$3497 ( \5501 , RI2b5e785b4d18_430, \5389 );
and \U$3498 ( \5502 , RI2b5e785b3968_450, \5391 );
and \U$3499 ( \5503 , RI2b5e785b3008_470, \5393 );
and \U$3500 ( \5504 , RI2b5e785b26a8_490, \5395 );
and \U$3501 ( \5505 , RI2b5e785b16b8_510, \5397 );
and \U$3502 ( \5506 , RI2b5e785b0d58_530, \5399 );
and \U$3503 ( \5507 , RI2b5e785b03f8_550, \5401 );
and \U$3504 ( \5508 , RI2b5e785af7c8_570, \5403 );
or \U$3505 ( \5509 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 );
_DC r26f3 ( \5510_nR26f3 , \5509 , \5413 );
buf \U$3506 ( \5511 , \5510_nR26f3 );
or \U$3507 ( \5512 , \5420 , \5452 );
not \U$3508 ( \5513 , \5512 );
buf \U$3509 ( \5514 , \5513 );
buf \U$3510 ( \5515 , \5514 );
xor \U$3511 ( \5516 , \5515 , \5455 );
and \U$3512 ( \5517 , \5511 , \5516 );
nor \U$3513 ( \5518 , 1'b0 , \5517 );
xnor \U$3515 ( \5519 , \5518 , 1'b0 );
xor \U$3516 ( \5520 , \5491 , \5519 );
xor \U$3517 ( \5521 , 1'b0 , \5520 );
xor \U$3519 ( \5522 , \5291 , \5295 );
xor \U$3520 ( \5523 , \5295 , \5299 );
not \U$3521 ( \5524 , \5523 );
and \U$3522 ( \5525 , \5522 , \5524 );
and \U$3523 ( \5526 , \5484 , \5525 );
not \U$3524 ( \5527 , \5526 );
xnor \U$3525 ( \5528 , \5527 , \5302 );
and \U$3526 ( \5529 , \5511 , \5463 );
and \U$3527 ( \5530 , \5415 , \5461 );
nor \U$3528 ( \5531 , \5529 , \5530 );
xnor \U$3529 ( \5532 , \5531 , \5489 );
and \U$3530 ( \5533 , \5528 , \5532 );
or \U$3532 ( \5534 , 1'b0 , \5533 , 1'b0 );
xor \U$3534 ( \5535 , \5534 , 1'b0 );
xor \U$3536 ( \5536 , \5535 , 1'b0 );
and \U$3537 ( \5537 , \5521 , \5536 );
or \U$3538 ( \5538 , 1'b0 , 1'b0 , \5537 );
and \U$3541 ( \5539 , \5484 , \5463 );
not \U$3542 ( \5540 , \5539 );
xnor \U$3543 ( \5541 , \5540 , \5489 );
xor \U$3544 ( \5542 , 1'b0 , \5541 );
and \U$3546 ( \5543 , \5415 , \5516 );
nor \U$3547 ( \5544 , 1'b0 , \5543 );
xnor \U$3548 ( \5545 , \5544 , 1'b0 );
xor \U$3549 ( \5546 , \5542 , \5545 );
xor \U$3550 ( \5547 , 1'b0 , \5546 );
xor \U$3552 ( \5548 , \5547 , 1'b1 );
and \U$3553 ( \5549 , \5303 , \5490 );
and \U$3554 ( \5550 , \5490 , \5519 );
and \U$3555 ( \5551 , \5303 , \5519 );
or \U$3556 ( \5552 , \5549 , \5550 , \5551 );
xor \U$3558 ( \5553 , \5552 , 1'b0 );
xor \U$3560 ( \5554 , \5553 , 1'b0 );
xor \U$3561 ( \5555 , \5548 , \5554 );
and \U$3562 ( \5556 , \5538 , \5555 );
or \U$3564 ( \5557 , 1'b0 , \5556 , 1'b0 );
xor \U$3566 ( \5558 , \5557 , 1'b0 );
and \U$3568 ( \5559 , \5547 , 1'b1 );
and \U$3569 ( \5560 , 1'b1 , \5554 );
and \U$3570 ( \5561 , \5547 , \5554 );
or \U$3571 ( \5562 , \5559 , \5560 , \5561 );
xor \U$3572 ( \5563 , 1'b0 , \5562 );
not \U$3574 ( \5564 , \5489 );
and \U$3576 ( \5565 , \5484 , \5516 );
nor \U$3577 ( \5566 , 1'b0 , \5565 );
xnor \U$3578 ( \5567 , \5566 , 1'b0 );
xor \U$3579 ( \5568 , \5564 , \5567 );
xor \U$3581 ( \5569 , \5568 , 1'b0 );
xor \U$3582 ( \5570 , 1'b0 , \5569 );
xor \U$3584 ( \5571 , \5570 , 1'b0 );
and \U$3586 ( \5572 , \5541 , \5545 );
or \U$3588 ( \5573 , 1'b0 , \5572 , 1'b0 );
xor \U$3590 ( \5574 , \5573 , 1'b0 );
xor \U$3592 ( \5575 , \5574 , 1'b0 );
xor \U$3593 ( \5576 , \5571 , \5575 );
xor \U$3594 ( \5577 , \5563 , \5576 );
xor \U$3595 ( \5578 , \5558 , \5577 );
xor \U$3601 ( \5579 , \5037 , \5058 );
xor \U$3602 ( \5580 , \5579 , \5279 );
buf \U$3603 ( \5581 , \5580 );
buf \U$3604 ( \5582 , \5581 );
xor \U$3605 ( \5583 , \5299 , \5582 );
xor \U$3606 ( \5584 , \5062 , \5083 );
xor \U$3607 ( \5585 , \5584 , \5276 );
buf \U$3608 ( \5586 , \5585 );
buf \U$3609 ( \5587 , \5586 );
xor \U$3610 ( \5588 , \5582 , \5587 );
not \U$3611 ( \5589 , \5588 );
and \U$3612 ( \5590 , \5583 , \5589 );
and \U$3613 ( \5591 , \5484 , \5590 );
not \U$3614 ( \5592 , \5591 );
and \U$3615 ( \5593 , \5582 , \5587 );
not \U$3616 ( \5594 , \5593 );
and \U$3617 ( \5595 , \5299 , \5594 );
xnor \U$3618 ( \5596 , \5592 , \5595 );
and \U$3619 ( \5597 , \5511 , \5525 );
and \U$3620 ( \5598 , \5415 , \5523 );
nor \U$3621 ( \5599 , \5597 , \5598 );
xnor \U$3622 ( \5600 , \5599 , \5302 );
and \U$3623 ( \5601 , \5596 , \5600 );
or \U$3625 ( \5602 , 1'b0 , \5601 , 1'b0 );
and \U$3626 ( \5603 , RI2b5e785da0e0_252, \5368 );
and \U$3627 ( \5604 , RI2b5e785be5e8_272, \5370 );
and \U$3628 ( \5605 , RI2b5e785bc338_292, \5373 );
and \U$3629 ( \5606 , RI2b5e785bb9d8_312, \5376 );
and \U$3630 ( \5607 , RI2b5e785b9ae8_332, \5378 );
and \U$3631 ( \5608 , RI2b5e785b7fb8_352, \5381 );
and \U$3632 ( \5609 , RI2b5e785b7658_372, \5383 );
and \U$3633 ( \5610 , RI2b5e785b5ee8_392, \5385 );
and \U$3634 ( \5611 , RI2b5e785b5588_412, \5387 );
and \U$3635 ( \5612 , RI2b5e785b4c28_432, \5389 );
and \U$3636 ( \5613 , RI2b5e785b3878_452, \5391 );
and \U$3637 ( \5614 , RI2b5e785b2f18_472, \5393 );
and \U$3638 ( \5615 , RI2b5e785b25b8_492, \5395 );
and \U$3639 ( \5616 , RI2b5e785b15c8_512, \5397 );
and \U$3640 ( \5617 , RI2b5e785b0c68_532, \5399 );
and \U$3641 ( \5618 , RI2b5e785b0308_552, \5401 );
and \U$3642 ( \5619 , RI2b5e785af6d8_572, \5403 );
or \U$3643 ( \5620 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 );
_DC r2554 ( \5621_nR2554 , \5620 , \5413 );
buf \U$3644 ( \5622 , \5621_nR2554 );
and \U$3645 ( \5623 , \5622 , \5463 );
and \U$3646 ( \5624 , RI2b5e785da158_251, \5368 );
and \U$3647 ( \5625 , RI2b5e785be660_271, \5370 );
and \U$3648 ( \5626 , RI2b5e785bc3b0_291, \5373 );
and \U$3649 ( \5627 , RI2b5e785bba50_311, \5376 );
and \U$3650 ( \5628 , RI2b5e785b9b60_331, \5378 );
and \U$3651 ( \5629 , RI2b5e785b8030_351, \5381 );
and \U$3652 ( \5630 , RI2b5e785b76d0_371, \5383 );
and \U$3653 ( \5631 , RI2b5e785b6d70_391, \5385 );
and \U$3654 ( \5632 , RI2b5e785b5600_411, \5387 );
and \U$3655 ( \5633 , RI2b5e785b4ca0_431, \5389 );
and \U$3656 ( \5634 , RI2b5e785b38f0_451, \5391 );
and \U$3657 ( \5635 , RI2b5e785b2f90_471, \5393 );
and \U$3658 ( \5636 , RI2b5e785b2630_491, \5395 );
and \U$3659 ( \5637 , RI2b5e785b1640_511, \5397 );
and \U$3660 ( \5638 , RI2b5e785b0ce0_531, \5399 );
and \U$3661 ( \5639 , RI2b5e785b0380_551, \5401 );
and \U$3662 ( \5640 , RI2b5e785af750_571, \5403 );
or \U$3663 ( \5641 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 );
_DC r2632 ( \5642_nR2632 , \5641 , \5413 );
buf \U$3664 ( \5643 , \5642_nR2632 );
and \U$3665 ( \5644 , \5643 , \5461 );
nor \U$3666 ( \5645 , \5623 , \5644 );
xnor \U$3667 ( \5646 , \5645 , \5489 );
and \U$3669 ( \5647 , RI2b5e785da068_253, \5368 );
and \U$3670 ( \5648 , RI2b5e785be570_273, \5370 );
and \U$3671 ( \5649 , RI2b5e785bc2c0_293, \5373 );
and \U$3672 ( \5650 , RI2b5e785bb960_313, \5376 );
and \U$3673 ( \5651 , RI2b5e785b9a70_333, \5378 );
and \U$3674 ( \5652 , RI2b5e785b7f40_353, \5381 );
and \U$3675 ( \5653 , RI2b5e785b75e0_373, \5383 );
and \U$3676 ( \5654 , RI2b5e785b5e70_393, \5385 );
and \U$3677 ( \5655 , RI2b5e785b5510_413, \5387 );
and \U$3678 ( \5656 , RI2b5e785b4bb0_433, \5389 );
and \U$3679 ( \5657 , RI2b5e785b3800_453, \5391 );
and \U$3680 ( \5658 , RI2b5e785b2ea0_473, \5393 );
and \U$3681 ( \5659 , RI2b5e785b2540_493, \5395 );
and \U$3682 ( \5660 , RI2b5e785b1550_513, \5397 );
and \U$3683 ( \5661 , RI2b5e785b0bf0_533, \5399 );
and \U$3684 ( \5662 , RI2b5e785b0290_553, \5401 );
and \U$3685 ( \5663 , RI2b5e785af660_573, \5403 );
or \U$3686 ( \5664 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 );
_DC r246b ( \5665_nR246b , \5664 , \5413 );
buf \U$3687 ( \5666 , \5665_nR246b );
and \U$3688 ( \5667 , \5666 , \5516 );
nor \U$3689 ( \5668 , 1'b0 , \5667 );
xnor \U$3690 ( \5669 , \5668 , 1'b0 );
and \U$3691 ( \5670 , \5646 , \5669 );
or \U$3694 ( \5671 , \5670 , 1'b0 , 1'b0 );
and \U$3695 ( \5672 , \5602 , \5671 );
or \U$3698 ( \5673 , \5672 , 1'b0 , 1'b0 );
and \U$3701 ( \5674 , \5622 , \5516 );
nor \U$3702 ( \5675 , 1'b0 , \5674 );
xnor \U$3703 ( \5676 , \5675 , 1'b0 );
xor \U$3705 ( \5677 , \5676 , 1'b0 );
xor \U$3707 ( \5678 , \5677 , 1'b0 );
not \U$3708 ( \5679 , \5595 );
and \U$3709 ( \5680 , \5415 , \5525 );
and \U$3710 ( \5681 , \5484 , \5523 );
nor \U$3711 ( \5682 , \5680 , \5681 );
xnor \U$3712 ( \5683 , \5682 , \5302 );
xor \U$3713 ( \5684 , \5679 , \5683 );
and \U$3714 ( \5685 , \5643 , \5463 );
and \U$3715 ( \5686 , \5511 , \5461 );
nor \U$3716 ( \5687 , \5685 , \5686 );
xnor \U$3717 ( \5688 , \5687 , \5489 );
xor \U$3718 ( \5689 , \5684 , \5688 );
and \U$3719 ( \5690 , \5678 , \5689 );
or \U$3721 ( \5691 , 1'b0 , \5690 , 1'b0 );
and \U$3722 ( \5692 , \5673 , \5691 );
or \U$3723 ( \5693 , 1'b0 , 1'b0 , \5692 );
and \U$3725 ( \5694 , \5643 , \5516 );
nor \U$3726 ( \5695 , 1'b0 , \5694 );
xnor \U$3727 ( \5696 , \5695 , 1'b0 );
xor \U$3729 ( \5697 , \5696 , 1'b0 );
xor \U$3731 ( \5698 , \5697 , 1'b0 );
xor \U$3733 ( \5699 , 1'b0 , \5528 );
xor \U$3734 ( \5700 , \5699 , \5532 );
xor \U$3735 ( \5701 , \5698 , \5700 );
and \U$3737 ( \5702 , \5701 , 1'b1 );
and \U$3738 ( \5703 , \5679 , \5683 );
and \U$3739 ( \5704 , \5683 , \5688 );
and \U$3740 ( \5705 , \5679 , \5688 );
or \U$3741 ( \5706 , \5703 , \5704 , \5705 );
xor \U$3743 ( \5707 , \5706 , 1'b0 );
xor \U$3745 ( \5708 , \5707 , 1'b0 );
and \U$3746 ( \5709 , 1'b1 , \5708 );
and \U$3747 ( \5710 , \5701 , \5708 );
or \U$3748 ( \5711 , \5702 , \5709 , \5710 );
and \U$3749 ( \5712 , \5693 , \5711 );
xor \U$3751 ( \5713 , \5521 , 1'b0 );
xor \U$3752 ( \5714 , \5713 , \5536 );
and \U$3753 ( \5715 , \5711 , \5714 );
and \U$3754 ( \5716 , \5693 , \5714 );
or \U$3755 ( \5717 , \5712 , \5715 , \5716 );
xor \U$3757 ( \5718 , 1'b0 , \5538 );
xor \U$3758 ( \5719 , \5718 , \5555 );
and \U$3759 ( \5720 , \5717 , \5719 );
or \U$3760 ( \5721 , 1'b0 , 1'b0 , \5720 );
nand \U$3761 ( \5722 , \5578 , \5721 );
nor \U$3762 ( \5723 , \5578 , \5721 );
not \U$3763 ( \5724 , \5723 );
nand \U$3764 ( \5725 , \5722 , \5724 );
xor \U$3765 ( \5726 , \5212 , \5233 );
xor \U$3766 ( \5727 , \5726 , \5258 );
buf \U$3767 ( \5728 , \5727 );
buf \U$3768 ( \5729 , \5728 );
xor \U$3769 ( \5730 , \5236 , \5256 );
buf \U$3770 ( \5731 , \5730 );
buf \U$3771 ( \5732 , \5731 );
xor \U$3772 ( \5733 , \5729 , \5732 );
not \U$3773 ( \5734 , \5732 );
and \U$3774 ( \5735 , \5733 , \5734 );
and \U$3775 ( \5736 , \5666 , \5735 );
and \U$3776 ( \5737 , \5622 , \5732 );
nor \U$3777 ( \5738 , \5736 , \5737 );
xnor \U$3778 ( \5739 , \5738 , \5729 );
and \U$3779 ( \5740 , RI2b5e785c2bc0_255, \5368 );
and \U$3780 ( \5741 , RI2b5e785be480_275, \5370 );
and \U$3781 ( \5742 , RI2b5e785bc1d0_295, \5373 );
and \U$3782 ( \5743 , RI2b5e785ba2e0_315, \5376 );
and \U$3783 ( \5744 , RI2b5e785b9980_335, \5378 );
and \U$3784 ( \5745 , RI2b5e785b7e50_355, \5381 );
and \U$3785 ( \5746 , RI2b5e785b74f0_375, \5383 );
and \U$3786 ( \5747 , RI2b5e785b5d80_395, \5385 );
and \U$3787 ( \5748 , RI2b5e785b5420_415, \5387 );
and \U$3788 ( \5749 , RI2b5e785b4ac0_435, \5389 );
and \U$3789 ( \5750 , RI2b5e785b3710_455, \5391 );
and \U$3790 ( \5751 , RI2b5e785b2db0_475, \5393 );
and \U$3791 ( \5752 , RI2b5e785b2450_495, \5395 );
and \U$3792 ( \5753 , RI2b5e785b1460_515, \5397 );
and \U$3793 ( \5754 , RI2b5e785b0b00_535, \5399 );
and \U$3794 ( \5755 , RI2b5e785b01a0_555, \5401 );
and \U$3795 ( \5756 , RI2b5e785af570_575, \5403 );
or \U$3796 ( \5757 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 );
_DC r22da ( \5758_nR22da , \5757 , \5413 );
buf \U$3797 ( \5759 , \5758_nR22da );
xor \U$3798 ( \5760 , \5162 , \5183 );
xor \U$3799 ( \5761 , \5760 , \5264 );
buf \U$3800 ( \5762 , \5761 );
buf \U$3801 ( \5763 , \5762 );
xor \U$3802 ( \5764 , \5187 , \5208 );
xor \U$3803 ( \5765 , \5764 , \5261 );
buf \U$3804 ( \5766 , \5765 );
buf \U$3805 ( \5767 , \5766 );
xor \U$3806 ( \5768 , \5763 , \5767 );
xor \U$3807 ( \5769 , \5767 , \5729 );
not \U$3808 ( \5770 , \5769 );
and \U$3809 ( \5771 , \5768 , \5770 );
and \U$3810 ( \5772 , \5759 , \5771 );
and \U$3811 ( \5773 , RI2b5e785c2c38_254, \5368 );
and \U$3812 ( \5774 , RI2b5e785be4f8_274, \5370 );
and \U$3813 ( \5775 , RI2b5e785bc248_294, \5373 );
and \U$3814 ( \5776 , RI2b5e785ba358_314, \5376 );
and \U$3815 ( \5777 , RI2b5e785b99f8_334, \5378 );
and \U$3816 ( \5778 , RI2b5e785b7ec8_354, \5381 );
and \U$3817 ( \5779 , RI2b5e785b7568_374, \5383 );
and \U$3818 ( \5780 , RI2b5e785b5df8_394, \5385 );
and \U$3819 ( \5781 , RI2b5e785b5498_414, \5387 );
and \U$3820 ( \5782 , RI2b5e785b4b38_434, \5389 );
and \U$3821 ( \5783 , RI2b5e785b3788_454, \5391 );
and \U$3822 ( \5784 , RI2b5e785b2e28_474, \5393 );
and \U$3823 ( \5785 , RI2b5e785b24c8_494, \5395 );
and \U$3824 ( \5786 , RI2b5e785b14d8_514, \5397 );
and \U$3825 ( \5787 , RI2b5e785b0b78_534, \5399 );
and \U$3826 ( \5788 , RI2b5e785b0218_554, \5401 );
and \U$3827 ( \5789 , RI2b5e785af5e8_574, \5403 );
or \U$3828 ( \5790 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 );
_DC r2387 ( \5791_nR2387 , \5790 , \5413 );
buf \U$3829 ( \5792 , \5791_nR2387 );
and \U$3830 ( \5793 , \5792 , \5769 );
nor \U$3831 ( \5794 , \5772 , \5793 );
and \U$3832 ( \5795 , \5767 , \5729 );
not \U$3833 ( \5796 , \5795 );
and \U$3834 ( \5797 , \5763 , \5796 );
xnor \U$3835 ( \5798 , \5794 , \5797 );
and \U$3836 ( \5799 , \5739 , \5798 );
and \U$3837 ( \5800 , RI2b5e785c0a00_257, \5368 );
and \U$3838 ( \5801 , RI2b5e785be390_277, \5370 );
and \U$3839 ( \5802 , RI2b5e785bc0e0_297, \5373 );
and \U$3840 ( \5803 , RI2b5e785ba1f0_317, \5376 );
and \U$3841 ( \5804 , RI2b5e785b9890_337, \5378 );
and \U$3842 ( \5805 , RI2b5e785b7d60_357, \5381 );
and \U$3843 ( \5806 , RI2b5e785b7400_377, \5383 );
and \U$3844 ( \5807 , RI2b5e785b5c90_397, \5385 );
and \U$3845 ( \5808 , RI2b5e785b5330_417, \5387 );
and \U$3846 ( \5809 , RI2b5e785b49d0_437, \5389 );
and \U$3847 ( \5810 , RI2b5e785b3620_457, \5391 );
and \U$3848 ( \5811 , RI2b5e785b2cc0_477, \5393 );
and \U$3849 ( \5812 , RI2b5e785b2360_497, \5395 );
and \U$3850 ( \5813 , RI2b5e785b1370_517, \5397 );
and \U$3851 ( \5814 , RI2b5e785b0a10_537, \5399 );
and \U$3852 ( \5815 , RI2b5e785b00b0_557, \5401 );
and \U$3853 ( \5816 , RI2b5e785af480_577, \5403 );
or \U$3854 ( \5817 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 );
_DC r211a ( \5818_nR211a , \5817 , \5413 );
buf \U$3855 ( \5819 , \5818_nR211a );
xor \U$3856 ( \5820 , \5112 , \5133 );
xor \U$3857 ( \5821 , \5820 , \5270 );
buf \U$3858 ( \5822 , \5821 );
buf \U$3859 ( \5823 , \5822 );
xor \U$3860 ( \5824 , \5137 , \5158 );
xor \U$3861 ( \5825 , \5824 , \5267 );
buf \U$3862 ( \5826 , \5825 );
buf \U$3863 ( \5827 , \5826 );
xor \U$3864 ( \5828 , \5823 , \5827 );
xor \U$3865 ( \5829 , \5827 , \5763 );
not \U$3866 ( \5830 , \5829 );
and \U$3867 ( \5831 , \5828 , \5830 );
and \U$3868 ( \5832 , \5819 , \5831 );
and \U$3869 ( \5833 , RI2b5e785c2b48_256, \5368 );
and \U$3870 ( \5834 , RI2b5e785be408_276, \5370 );
and \U$3871 ( \5835 , RI2b5e785bc158_296, \5373 );
and \U$3872 ( \5836 , RI2b5e785ba268_316, \5376 );
and \U$3873 ( \5837 , RI2b5e785b9908_336, \5378 );
and \U$3874 ( \5838 , RI2b5e785b7dd8_356, \5381 );
and \U$3875 ( \5839 , RI2b5e785b7478_376, \5383 );
and \U$3876 ( \5840 , RI2b5e785b5d08_396, \5385 );
and \U$3877 ( \5841 , RI2b5e785b53a8_416, \5387 );
and \U$3878 ( \5842 , RI2b5e785b4a48_436, \5389 );
and \U$3879 ( \5843 , RI2b5e785b3698_456, \5391 );
and \U$3880 ( \5844 , RI2b5e785b2d38_476, \5393 );
and \U$3881 ( \5845 , RI2b5e785b23d8_496, \5395 );
and \U$3882 ( \5846 , RI2b5e785b13e8_516, \5397 );
and \U$3883 ( \5847 , RI2b5e785b0a88_536, \5399 );
and \U$3884 ( \5848 , RI2b5e785b0128_556, \5401 );
and \U$3885 ( \5849 , RI2b5e785af4f8_576, \5403 );
or \U$3886 ( \5850 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 );
_DC r21b2 ( \5851_nR21b2 , \5850 , \5413 );
buf \U$3887 ( \5852 , \5851_nR21b2 );
and \U$3888 ( \5853 , \5852 , \5829 );
nor \U$3889 ( \5854 , \5832 , \5853 );
and \U$3890 ( \5855 , \5827 , \5763 );
not \U$3891 ( \5856 , \5855 );
and \U$3892 ( \5857 , \5823 , \5856 );
xnor \U$3893 ( \5858 , \5854 , \5857 );
and \U$3894 ( \5859 , \5798 , \5858 );
and \U$3895 ( \5860 , \5739 , \5858 );
or \U$3896 ( \5861 , \5799 , \5859 , \5860 );
and \U$3897 ( \5862 , RI2b5e785c0910_259, \5368 );
and \U$3898 ( \5863 , RI2b5e785be2a0_279, \5370 );
and \U$3899 ( \5864 , RI2b5e785bbff0_299, \5373 );
and \U$3900 ( \5865 , RI2b5e785ba100_319, \5376 );
and \U$3901 ( \5866 , RI2b5e785b97a0_339, \5378 );
and \U$3902 ( \5867 , RI2b5e785b7c70_359, \5381 );
and \U$3903 ( \5868 , RI2b5e785b7310_379, \5383 );
and \U$3904 ( \5869 , RI2b5e785b5ba0_399, \5385 );
and \U$3905 ( \5870 , RI2b5e785b5240_419, \5387 );
and \U$3906 ( \5871 , RI2b5e785b48e0_439, \5389 );
and \U$3907 ( \5872 , RI2b5e785b3530_459, \5391 );
and \U$3908 ( \5873 , RI2b5e785b2bd0_479, \5393 );
and \U$3909 ( \5874 , RI2b5e785b2270_499, \5395 );
and \U$3910 ( \5875 , RI2b5e785b1280_519, \5397 );
and \U$3911 ( \5876 , RI2b5e785b0920_539, \5399 );
and \U$3912 ( \5877 , RI2b5e785affc0_559, \5401 );
and \U$3913 ( \5878 , RI2b5e785af390_579, \5403 );
or \U$3914 ( \5879 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 );
_DC r1f4f ( \5880_nR1f4f , \5879 , \5413 );
buf \U$3915 ( \5881 , \5880_nR1f4f );
xor \U$3916 ( \5882 , \5087 , \5108 );
xor \U$3917 ( \5883 , \5882 , \5273 );
buf \U$3918 ( \5884 , \5883 );
buf \U$3919 ( \5885 , \5884 );
xor \U$3920 ( \5886 , \5587 , \5885 );
xor \U$3921 ( \5887 , \5885 , \5823 );
not \U$3922 ( \5888 , \5887 );
and \U$3923 ( \5889 , \5886 , \5888 );
and \U$3924 ( \5890 , \5881 , \5889 );
and \U$3925 ( \5891 , RI2b5e785c0988_258, \5368 );
and \U$3926 ( \5892 , RI2b5e785be318_278, \5370 );
and \U$3927 ( \5893 , RI2b5e785bc068_298, \5373 );
and \U$3928 ( \5894 , RI2b5e785ba178_318, \5376 );
and \U$3929 ( \5895 , RI2b5e785b9818_338, \5378 );
and \U$3930 ( \5896 , RI2b5e785b7ce8_358, \5381 );
and \U$3931 ( \5897 , RI2b5e785b7388_378, \5383 );
and \U$3932 ( \5898 , RI2b5e785b5c18_398, \5385 );
and \U$3933 ( \5899 , RI2b5e785b52b8_418, \5387 );
and \U$3934 ( \5900 , RI2b5e785b4958_438, \5389 );
and \U$3935 ( \5901 , RI2b5e785b35a8_458, \5391 );
and \U$3936 ( \5902 , RI2b5e785b2c48_478, \5393 );
and \U$3937 ( \5903 , RI2b5e785b22e8_498, \5395 );
and \U$3938 ( \5904 , RI2b5e785b12f8_518, \5397 );
and \U$3939 ( \5905 , RI2b5e785b0998_538, \5399 );
and \U$3940 ( \5906 , RI2b5e785b0038_558, \5401 );
and \U$3941 ( \5907 , RI2b5e785af408_578, \5403 );
or \U$3942 ( \5908 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 );
_DC r1fd9 ( \5909_nR1fd9 , \5908 , \5413 );
buf \U$3943 ( \5910 , \5909_nR1fd9 );
and \U$3944 ( \5911 , \5910 , \5887 );
nor \U$3945 ( \5912 , \5890 , \5911 );
and \U$3946 ( \5913 , \5885 , \5823 );
not \U$3947 ( \5914 , \5913 );
and \U$3948 ( \5915 , \5587 , \5914 );
xnor \U$3949 ( \5916 , \5912 , \5915 );
and \U$3950 ( \5917 , RI2b5e785c0820_261, \5368 );
and \U$3951 ( \5918 , RI2b5e785be1b0_281, \5370 );
and \U$3952 ( \5919 , RI2b5e785bbf00_301, \5373 );
and \U$3953 ( \5920 , RI2b5e785ba010_321, \5376 );
and \U$3954 ( \5921 , RI2b5e785b96b0_341, \5378 );
and \U$3955 ( \5922 , RI2b5e785b7b80_361, \5381 );
and \U$3956 ( \5923 , RI2b5e785b7220_381, \5383 );
and \U$3957 ( \5924 , RI2b5e785b5ab0_401, \5385 );
and \U$3958 ( \5925 , RI2b5e785b5150_421, \5387 );
and \U$3959 ( \5926 , RI2b5e785b47f0_441, \5389 );
and \U$3960 ( \5927 , RI2b5e785b3440_461, \5391 );
and \U$3961 ( \5928 , RI2b5e785b2ae0_481, \5393 );
and \U$3962 ( \5929 , RI2b5e785b2180_501, \5395 );
and \U$3963 ( \5930 , RI2b5e785b1190_521, \5397 );
and \U$3964 ( \5931 , RI2b5e785b0830_541, \5399 );
and \U$3965 ( \5932 , RI2b5e785afed0_561, \5401 );
and \U$3966 ( \5933 , RI2b5e785af2a0_581, \5403 );
or \U$3967 ( \5934 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 );
_DC r1dac ( \5935_nR1dac , \5934 , \5413 );
buf \U$3968 ( \5936 , \5935_nR1dac );
and \U$3969 ( \5937 , \5936 , \5590 );
and \U$3970 ( \5938 , RI2b5e785c0898_260, \5368 );
and \U$3971 ( \5939 , RI2b5e785be228_280, \5370 );
and \U$3972 ( \5940 , RI2b5e785bbf78_300, \5373 );
and \U$3973 ( \5941 , RI2b5e785ba088_320, \5376 );
and \U$3974 ( \5942 , RI2b5e785b9728_340, \5378 );
and \U$3975 ( \5943 , RI2b5e785b7bf8_360, \5381 );
and \U$3976 ( \5944 , RI2b5e785b7298_380, \5383 );
and \U$3977 ( \5945 , RI2b5e785b5b28_400, \5385 );
and \U$3978 ( \5946 , RI2b5e785b51c8_420, \5387 );
and \U$3979 ( \5947 , RI2b5e785b4868_440, \5389 );
and \U$3980 ( \5948 , RI2b5e785b34b8_460, \5391 );
and \U$3981 ( \5949 , RI2b5e785b2b58_480, \5393 );
and \U$3982 ( \5950 , RI2b5e785b21f8_500, \5395 );
and \U$3983 ( \5951 , RI2b5e785b1208_520, \5397 );
and \U$3984 ( \5952 , RI2b5e785b08a8_540, \5399 );
and \U$3985 ( \5953 , RI2b5e785aff48_560, \5401 );
and \U$3986 ( \5954 , RI2b5e785af318_580, \5403 );
or \U$3987 ( \5955 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 );
_DC r1e20 ( \5956_nR1e20 , \5955 , \5413 );
buf \U$3988 ( \5957 , \5956_nR1e20 );
and \U$3989 ( \5958 , \5957 , \5588 );
nor \U$3990 ( \5959 , \5937 , \5958 );
xnor \U$3991 ( \5960 , \5959 , \5595 );
and \U$3992 ( \5961 , \5916 , \5960 );
and \U$3993 ( \5962 , RI2b5e785c0730_263, \5368 );
and \U$3994 ( \5963 , RI2b5e785be0c0_283, \5370 );
and \U$3995 ( \5964 , RI2b5e785bbe10_303, \5373 );
and \U$3996 ( \5965 , RI2b5e785b9f20_323, \5376 );
and \U$3997 ( \5966 , RI2b5e785b95c0_343, \5378 );
and \U$3998 ( \5967 , RI2b5e785b7a90_363, \5381 );
and \U$3999 ( \5968 , RI2b5e785b7130_383, \5383 );
and \U$4000 ( \5969 , RI2b5e785b59c0_403, \5385 );
and \U$4001 ( \5970 , RI2b5e785b5060_423, \5387 );
and \U$4002 ( \5971 , RI2b5e785b3cb0_443, \5389 );
and \U$4003 ( \5972 , RI2b5e785b3350_463, \5391 );
and \U$4004 ( \5973 , RI2b5e785b29f0_483, \5393 );
and \U$4005 ( \5974 , RI2b5e785b1a00_503, \5395 );
and \U$4006 ( \5975 , RI2b5e785b10a0_523, \5397 );
and \U$4007 ( \5976 , RI2b5e785b0740_543, \5399 );
and \U$4008 ( \5977 , RI2b5e785afde0_563, \5401 );
and \U$4009 ( \5978 , RI2b5e785af1b0_583, \5403 );
or \U$4010 ( \5979 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 );
_DC r1c3b ( \5980_nR1c3b , \5979 , \5413 );
buf \U$4011 ( \5981 , \5980_nR1c3b );
and \U$4012 ( \5982 , \5981 , \5525 );
and \U$4013 ( \5983 , RI2b5e785c07a8_262, \5368 );
and \U$4014 ( \5984 , RI2b5e785be138_282, \5370 );
and \U$4015 ( \5985 , RI2b5e785bbe88_302, \5373 );
and \U$4016 ( \5986 , RI2b5e785b9f98_322, \5376 );
and \U$4017 ( \5987 , RI2b5e785b9638_342, \5378 );
and \U$4018 ( \5988 , RI2b5e785b7b08_362, \5381 );
and \U$4019 ( \5989 , RI2b5e785b71a8_382, \5383 );
and \U$4020 ( \5990 , RI2b5e785b5a38_402, \5385 );
and \U$4021 ( \5991 , RI2b5e785b50d8_422, \5387 );
and \U$4022 ( \5992 , RI2b5e785b4778_442, \5389 );
and \U$4023 ( \5993 , RI2b5e785b33c8_462, \5391 );
and \U$4024 ( \5994 , RI2b5e785b2a68_482, \5393 );
and \U$4025 ( \5995 , RI2b5e785b1a78_502, \5395 );
and \U$4026 ( \5996 , RI2b5e785b1118_522, \5397 );
and \U$4027 ( \5997 , RI2b5e785b07b8_542, \5399 );
and \U$4028 ( \5998 , RI2b5e785afe58_562, \5401 );
and \U$4029 ( \5999 , RI2b5e785af228_582, \5403 );
or \U$4030 ( \6000 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 );
_DC r1ca2 ( \6001_nR1ca2 , \6000 , \5413 );
buf \U$4031 ( \6002 , \6001_nR1ca2 );
and \U$4032 ( \6003 , \6002 , \5523 );
nor \U$4033 ( \6004 , \5982 , \6003 );
xnor \U$4034 ( \6005 , \6004 , \5302 );
and \U$4035 ( \6006 , \5960 , \6005 );
and \U$4036 ( \6007 , \5916 , \6005 );
or \U$4037 ( \6008 , \5961 , \6006 , \6007 );
and \U$4038 ( \6009 , \5861 , \6008 );
and \U$4039 ( \6010 , RI2b5e785c0640_265, \5368 );
and \U$4040 ( \6011 , RI2b5e785bdfd0_285, \5370 );
and \U$4041 ( \6012 , RI2b5e785bbd20_305, \5373 );
and \U$4042 ( \6013 , RI2b5e785b9e30_325, \5376 );
and \U$4043 ( \6014 , RI2b5e785b94d0_345, \5378 );
and \U$4044 ( \6015 , RI2b5e785b79a0_365, \5381 );
and \U$4045 ( \6016 , RI2b5e785b7040_385, \5383 );
and \U$4046 ( \6017 , RI2b5e785b58d0_405, \5385 );
and \U$4047 ( \6018 , RI2b5e785b4f70_425, \5387 );
and \U$4048 ( \6019 , RI2b5e785b3bc0_445, \5389 );
and \U$4049 ( \6020 , RI2b5e785b3260_465, \5391 );
and \U$4050 ( \6021 , RI2b5e785b2900_485, \5393 );
and \U$4051 ( \6022 , RI2b5e785b1910_505, \5395 );
and \U$4052 ( \6023 , RI2b5e785b0fb0_525, \5397 );
and \U$4053 ( \6024 , RI2b5e785b0650_545, \5399 );
and \U$4054 ( \6025 , RI2b5e785afcf0_565, \5401 );
and \U$4055 ( \6026 , RI2b5e785af0c0_585, \5403 );
or \U$4056 ( \6027 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 );
_DC r1abd ( \6028_nR1abd , \6027 , \5413 );
buf \U$4057 ( \6029 , \6028_nR1abd );
and \U$4058 ( \6030 , \6029 , \5463 );
and \U$4059 ( \6031 , RI2b5e785c06b8_264, \5368 );
and \U$4060 ( \6032 , RI2b5e785be048_284, \5370 );
and \U$4061 ( \6033 , RI2b5e785bbd98_304, \5373 );
and \U$4062 ( \6034 , RI2b5e785b9ea8_324, \5376 );
and \U$4063 ( \6035 , RI2b5e785b9548_344, \5378 );
and \U$4064 ( \6036 , RI2b5e785b7a18_364, \5381 );
and \U$4065 ( \6037 , RI2b5e785b70b8_384, \5383 );
and \U$4066 ( \6038 , RI2b5e785b5948_404, \5385 );
and \U$4067 ( \6039 , RI2b5e785b4fe8_424, \5387 );
and \U$4068 ( \6040 , RI2b5e785b3c38_444, \5389 );
and \U$4069 ( \6041 , RI2b5e785b32d8_464, \5391 );
and \U$4070 ( \6042 , RI2b5e785b2978_484, \5393 );
and \U$4071 ( \6043 , RI2b5e785b1988_504, \5395 );
and \U$4072 ( \6044 , RI2b5e785b1028_524, \5397 );
and \U$4073 ( \6045 , RI2b5e785b06c8_544, \5399 );
and \U$4074 ( \6046 , RI2b5e785afd68_564, \5401 );
and \U$4075 ( \6047 , RI2b5e785af138_584, \5403 );
or \U$4076 ( \6048 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 );
_DC r1b50 ( \6049_nR1b50 , \6048 , \5413 );
buf \U$4077 ( \6050 , \6049_nR1b50 );
and \U$4078 ( \6051 , \6050 , \5461 );
nor \U$4079 ( \6052 , \6030 , \6051 );
xnor \U$4080 ( \6053 , \6052 , \5489 );
and \U$4082 ( \6054 , RI2b5e785c05c8_266, \5368 );
and \U$4083 ( \6055 , RI2b5e785bdf58_286, \5370 );
and \U$4084 ( \6056 , RI2b5e785bbca8_306, \5373 );
and \U$4085 ( \6057 , RI2b5e785b9db8_326, \5376 );
and \U$4086 ( \6058 , RI2b5e785b9458_346, \5378 );
and \U$4087 ( \6059 , RI2b5e785b7928_366, \5381 );
and \U$4088 ( \6060 , RI2b5e785b6fc8_386, \5383 );
and \U$4089 ( \6061 , RI2b5e785b5858_406, \5385 );
and \U$4090 ( \6062 , RI2b5e785b4ef8_426, \5387 );
and \U$4091 ( \6063 , RI2b5e785b3b48_446, \5389 );
and \U$4092 ( \6064 , RI2b5e785b31e8_466, \5391 );
and \U$4093 ( \6065 , RI2b5e785b2888_486, \5393 );
and \U$4094 ( \6066 , RI2b5e785b1898_506, \5395 );
and \U$4095 ( \6067 , RI2b5e785b0f38_526, \5397 );
and \U$4096 ( \6068 , RI2b5e785b05d8_546, \5399 );
and \U$4097 ( \6069 , RI2b5e785afc78_566, \5401 );
and \U$4098 ( \6070 , RI2b5e785af048_586, \5403 );
or \U$4099 ( \6071 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 );
_DC r1a35 ( \6072_nR1a35 , \6071 , \5413 );
buf \U$4100 ( \6073 , \6072_nR1a35 );
and \U$4101 ( \6074 , \6073 , \5516 );
nor \U$4102 ( \6075 , 1'b0 , \6074 );
xnor \U$4103 ( \6076 , \6075 , 1'b0 );
and \U$4104 ( \6077 , \6053 , \6076 );
and \U$4105 ( \6078 , \6008 , \6077 );
and \U$4106 ( \6079 , \5861 , \6077 );
or \U$4107 ( \6080 , \6009 , \6078 , \6079 );
and \U$4109 ( \6081 , \6002 , \5525 );
and \U$4110 ( \6082 , \5936 , \5523 );
nor \U$4111 ( \6083 , \6081 , \6082 );
xnor \U$4112 ( \6084 , \6083 , \5302 );
and \U$4113 ( \6085 , \6050 , \5463 );
and \U$4114 ( \6086 , \5981 , \5461 );
nor \U$4115 ( \6087 , \6085 , \6086 );
xnor \U$4116 ( \6088 , \6087 , \5489 );
xor \U$4117 ( \6089 , \6084 , \6088 );
and \U$4119 ( \6090 , \6029 , \5516 );
nor \U$4120 ( \6091 , 1'b0 , \6090 );
xnor \U$4121 ( \6092 , \6091 , 1'b0 );
xor \U$4122 ( \6093 , \6089 , \6092 );
and \U$4123 ( \6094 , \5852 , \5831 );
and \U$4124 ( \6095 , \5759 , \5829 );
nor \U$4125 ( \6096 , \6094 , \6095 );
xnor \U$4126 ( \6097 , \6096 , \5857 );
and \U$4127 ( \6098 , \5910 , \5889 );
and \U$4128 ( \6099 , \5819 , \5887 );
nor \U$4129 ( \6100 , \6098 , \6099 );
xnor \U$4130 ( \6101 , \6100 , \5915 );
xor \U$4131 ( \6102 , \6097 , \6101 );
and \U$4132 ( \6103 , \5957 , \5590 );
and \U$4133 ( \6104 , \5881 , \5588 );
nor \U$4134 ( \6105 , \6103 , \6104 );
xnor \U$4135 ( \6106 , \6105 , \5595 );
xor \U$4136 ( \6107 , \6102 , \6106 );
and \U$4137 ( \6108 , \6093 , \6107 );
or \U$4139 ( \6109 , 1'b0 , \6108 , 1'b0 );
xor \U$4140 ( \6110 , \6080 , \6109 );
and \U$4141 ( \6111 , \5981 , \5463 );
and \U$4142 ( \6112 , \6002 , \5461 );
nor \U$4143 ( \6113 , \6111 , \6112 );
xnor \U$4144 ( \6114 , \6113 , \5489 );
and \U$4146 ( \6115 , \6050 , \5516 );
nor \U$4147 ( \6116 , 1'b0 , \6115 );
xnor \U$4148 ( \6117 , \6116 , 1'b0 );
xor \U$4149 ( \6118 , \6114 , \6117 );
xor \U$4151 ( \6119 , \6118 , 1'b0 );
and \U$4152 ( \6120 , \5819 , \5889 );
and \U$4153 ( \6121 , \5852 , \5887 );
nor \U$4154 ( \6122 , \6120 , \6121 );
xnor \U$4155 ( \6123 , \6122 , \5915 );
and \U$4156 ( \6124 , \5881 , \5590 );
and \U$4157 ( \6125 , \5910 , \5588 );
nor \U$4158 ( \6126 , \6124 , \6125 );
xnor \U$4159 ( \6127 , \6126 , \5595 );
xor \U$4160 ( \6128 , \6123 , \6127 );
and \U$4161 ( \6129 , \5936 , \5525 );
and \U$4162 ( \6130 , \5957 , \5523 );
nor \U$4163 ( \6131 , \6129 , \6130 );
xnor \U$4164 ( \6132 , \6131 , \5302 );
xor \U$4165 ( \6133 , \6128 , \6132 );
xor \U$4166 ( \6134 , \6119 , \6133 );
and \U$4167 ( \6135 , \5643 , \5735 );
and \U$4168 ( \6136 , \5511 , \5732 );
nor \U$4169 ( \6137 , \6135 , \6136 );
xnor \U$4170 ( \6138 , \6137 , \5729 );
and \U$4171 ( \6139 , \5666 , \5771 );
and \U$4172 ( \6140 , \5622 , \5769 );
nor \U$4173 ( \6141 , \6139 , \6140 );
xnor \U$4174 ( \6142 , \6141 , \5797 );
xor \U$4175 ( \6143 , \6138 , \6142 );
and \U$4176 ( \6144 , \5759 , \5831 );
and \U$4177 ( \6145 , \5792 , \5829 );
nor \U$4178 ( \6146 , \6144 , \6145 );
xnor \U$4179 ( \6147 , \6146 , \5857 );
xor \U$4180 ( \6148 , \6143 , \6147 );
xor \U$4181 ( \6149 , \6134 , \6148 );
xor \U$4182 ( \6150 , \6110 , \6149 );
and \U$4184 ( \6151 , \5792 , \5735 );
and \U$4185 ( \6152 , \5666 , \5732 );
nor \U$4186 ( \6153 , \6151 , \6152 );
xnor \U$4187 ( \6154 , \6153 , \5729 );
and \U$4188 ( \6155 , \5852 , \5771 );
and \U$4189 ( \6156 , \5759 , \5769 );
nor \U$4190 ( \6157 , \6155 , \6156 );
xnor \U$4191 ( \6158 , \6157 , \5797 );
and \U$4192 ( \6159 , \6154 , \6158 );
or \U$4194 ( \6160 , 1'b0 , \6159 , 1'b0 );
and \U$4195 ( \6161 , \5910 , \5831 );
and \U$4196 ( \6162 , \5819 , \5829 );
nor \U$4197 ( \6163 , \6161 , \6162 );
xnor \U$4198 ( \6164 , \6163 , \5857 );
and \U$4199 ( \6165 , \5957 , \5889 );
and \U$4200 ( \6166 , \5881 , \5887 );
nor \U$4201 ( \6167 , \6165 , \6166 );
xnor \U$4202 ( \6168 , \6167 , \5915 );
and \U$4203 ( \6169 , \6164 , \6168 );
and \U$4204 ( \6170 , \6002 , \5590 );
and \U$4205 ( \6171 , \5936 , \5588 );
nor \U$4206 ( \6172 , \6170 , \6171 );
xnor \U$4207 ( \6173 , \6172 , \5595 );
and \U$4208 ( \6174 , \6168 , \6173 );
and \U$4209 ( \6175 , \6164 , \6173 );
or \U$4210 ( \6176 , \6169 , \6174 , \6175 );
and \U$4211 ( \6177 , \6160 , \6176 );
and \U$4212 ( \6178 , \6050 , \5525 );
and \U$4213 ( \6179 , \5981 , \5523 );
nor \U$4214 ( \6180 , \6178 , \6179 );
xnor \U$4215 ( \6181 , \6180 , \5302 );
and \U$4216 ( \6182 , \6073 , \5463 );
and \U$4217 ( \6183 , \6029 , \5461 );
nor \U$4218 ( \6184 , \6182 , \6183 );
xnor \U$4219 ( \6185 , \6184 , \5489 );
and \U$4220 ( \6186 , \6181 , \6185 );
and \U$4221 ( \6187 , RI2b5e785c0550_267, \5368 );
and \U$4222 ( \6188 , RI2b5e785bc590_287, \5370 );
and \U$4223 ( \6189 , RI2b5e785bbc30_307, \5373 );
and \U$4224 ( \6190 , RI2b5e785b9d40_327, \5376 );
and \U$4225 ( \6191 , RI2b5e785b93e0_347, \5378 );
and \U$4226 ( \6192 , RI2b5e785b78b0_367, \5381 );
and \U$4227 ( \6193 , RI2b5e785b6f50_387, \5383 );
and \U$4228 ( \6194 , RI2b5e785b57e0_407, \5385 );
and \U$4229 ( \6195 , RI2b5e785b4e80_427, \5387 );
and \U$4230 ( \6196 , RI2b5e785b3ad0_447, \5389 );
and \U$4231 ( \6197 , RI2b5e785b3170_467, \5391 );
and \U$4232 ( \6198 , RI2b5e785b2810_487, \5393 );
and \U$4233 ( \6199 , RI2b5e785b1820_507, \5395 );
and \U$4234 ( \6200 , RI2b5e785b0ec0_527, \5397 );
and \U$4235 ( \6201 , RI2b5e785b0560_547, \5399 );
and \U$4236 ( \6202 , RI2b5e785afc00_567, \5401 );
and \U$4237 ( \6203 , RI2b5e785aefd0_587, \5403 );
or \U$4238 ( \6204 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 );
_DC r19a3 ( \6205_nR19a3 , \6204 , \5413 );
buf \U$4239 ( \6206 , \6205_nR19a3 );
nand \U$4240 ( \6207 , \6206 , \5516 );
xnor \U$4241 ( \6208 , \6207 , 1'b0 );
and \U$4242 ( \6209 , \6185 , \6208 );
and \U$4243 ( \6210 , \6181 , \6208 );
or \U$4244 ( \6211 , \6186 , \6209 , \6210 );
and \U$4245 ( \6212 , \6176 , \6211 );
and \U$4246 ( \6213 , \6160 , \6211 );
or \U$4247 ( \6214 , \6177 , \6212 , \6213 );
xor \U$4248 ( \6215 , \6053 , \6076 );
xor \U$4249 ( \6216 , \5916 , \5960 );
xor \U$4250 ( \6217 , \6216 , \6005 );
and \U$4251 ( \6218 , \6215 , \6217 );
xor \U$4252 ( \6219 , \5739 , \5798 );
xor \U$4253 ( \6220 , \6219 , \5858 );
and \U$4254 ( \6221 , \6217 , \6220 );
and \U$4255 ( \6222 , \6215 , \6220 );
or \U$4256 ( \6223 , \6218 , \6221 , \6222 );
and \U$4257 ( \6224 , \6214 , \6223 );
and \U$4259 ( \6225 , \5622 , \5735 );
and \U$4260 ( \6226 , \5643 , \5732 );
nor \U$4261 ( \6227 , \6225 , \6226 );
xnor \U$4262 ( \6228 , \6227 , \5729 );
xor \U$4263 ( \6229 , 1'b0 , \6228 );
and \U$4264 ( \6230 , \5792 , \5771 );
and \U$4265 ( \6231 , \5666 , \5769 );
nor \U$4266 ( \6232 , \6230 , \6231 );
xnor \U$4267 ( \6233 , \6232 , \5797 );
xor \U$4268 ( \6234 , \6229 , \6233 );
and \U$4269 ( \6235 , \6223 , \6234 );
and \U$4270 ( \6236 , \6214 , \6234 );
or \U$4271 ( \6237 , \6224 , \6235 , \6236 );
xor \U$4273 ( \6238 , 1'b0 , \6093 );
xor \U$4274 ( \6239 , \6238 , \6107 );
xor \U$4275 ( \6240 , \5861 , \6008 );
xor \U$4276 ( \6241 , \6240 , \6077 );
and \U$4277 ( \6242 , \6239 , \6241 );
xor \U$4278 ( \6243 , \6237 , \6242 );
and \U$4280 ( \6244 , \6228 , \6233 );
or \U$4282 ( \6245 , 1'b0 , \6244 , 1'b0 );
and \U$4283 ( \6246 , \6097 , \6101 );
and \U$4284 ( \6247 , \6101 , \6106 );
and \U$4285 ( \6248 , \6097 , \6106 );
or \U$4286 ( \6249 , \6246 , \6247 , \6248 );
xor \U$4287 ( \6250 , \6245 , \6249 );
and \U$4288 ( \6251 , \6084 , \6088 );
and \U$4289 ( \6252 , \6088 , \6092 );
and \U$4290 ( \6253 , \6084 , \6092 );
or \U$4291 ( \6254 , \6251 , \6252 , \6253 );
xor \U$4292 ( \6255 , \6250 , \6254 );
xor \U$4293 ( \6256 , \6243 , \6255 );
xor \U$4294 ( \6257 , \6150 , \6256 );
and \U$4295 ( \6258 , \5759 , \5735 );
and \U$4296 ( \6259 , \5792 , \5732 );
nor \U$4297 ( \6260 , \6258 , \6259 );
xnor \U$4298 ( \6261 , \6260 , \5729 );
and \U$4299 ( \6262 , \5819 , \5771 );
and \U$4300 ( \6263 , \5852 , \5769 );
nor \U$4301 ( \6264 , \6262 , \6263 );
xnor \U$4302 ( \6265 , \6264 , \5797 );
and \U$4303 ( \6266 , \6261 , \6265 );
and \U$4304 ( \6267 , \5881 , \5831 );
and \U$4305 ( \6268 , \5910 , \5829 );
nor \U$4306 ( \6269 , \6267 , \6268 );
xnor \U$4307 ( \6270 , \6269 , \5857 );
and \U$4308 ( \6271 , \6265 , \6270 );
and \U$4309 ( \6272 , \6261 , \6270 );
or \U$4310 ( \6273 , \6266 , \6271 , \6272 );
and \U$4311 ( \6274 , \5936 , \5889 );
and \U$4312 ( \6275 , \5957 , \5887 );
nor \U$4313 ( \6276 , \6274 , \6275 );
xnor \U$4314 ( \6277 , \6276 , \5915 );
and \U$4315 ( \6278 , \5981 , \5590 );
and \U$4316 ( \6279 , \6002 , \5588 );
nor \U$4317 ( \6280 , \6278 , \6279 );
xnor \U$4318 ( \6281 , \6280 , \5595 );
and \U$4319 ( \6282 , \6277 , \6281 );
and \U$4320 ( \6283 , \6029 , \5525 );
and \U$4321 ( \6284 , \6050 , \5523 );
nor \U$4322 ( \6285 , \6283 , \6284 );
xnor \U$4323 ( \6286 , \6285 , \5302 );
and \U$4324 ( \6287 , \6281 , \6286 );
and \U$4325 ( \6288 , \6277 , \6286 );
or \U$4326 ( \6289 , \6282 , \6287 , \6288 );
and \U$4327 ( \6290 , \6273 , \6289 );
xor \U$4328 ( \6291 , \6181 , \6185 );
xor \U$4329 ( \6292 , \6291 , \6208 );
and \U$4330 ( \6293 , \6289 , \6292 );
and \U$4331 ( \6294 , \6273 , \6292 );
or \U$4332 ( \6295 , \6290 , \6293 , \6294 );
xor \U$4333 ( \6296 , \6164 , \6168 );
xor \U$4334 ( \6297 , \6296 , \6173 );
xor \U$4335 ( \6298 , 1'b0 , \6154 );
xor \U$4336 ( \6299 , \6298 , \6158 );
and \U$4337 ( \6300 , \6297 , \6299 );
and \U$4338 ( \6301 , \6295 , \6300 );
xor \U$4339 ( \6302 , \6215 , \6217 );
xor \U$4340 ( \6303 , \6302 , \6220 );
and \U$4341 ( \6304 , \6300 , \6303 );
and \U$4342 ( \6305 , \6295 , \6303 );
or \U$4343 ( \6306 , \6301 , \6304 , \6305 );
xor \U$4344 ( \6307 , \6239 , \6241 );
and \U$4345 ( \6308 , \6306 , \6307 );
xor \U$4346 ( \6309 , \6214 , \6223 );
xor \U$4347 ( \6310 , \6309 , \6234 );
and \U$4348 ( \6311 , \6307 , \6310 );
and \U$4349 ( \6312 , \6306 , \6310 );
or \U$4350 ( \6313 , \6308 , \6311 , \6312 );
nor \U$4351 ( \6314 , \6257 , \6313 );
and \U$4352 ( \6315 , \6237 , \6242 );
and \U$4353 ( \6316 , \6242 , \6255 );
and \U$4354 ( \6317 , \6237 , \6255 );
or \U$4355 ( \6318 , \6315 , \6316 , \6317 );
and \U$4356 ( \6319 , \6080 , \6109 );
and \U$4357 ( \6320 , \6109 , \6149 );
and \U$4358 ( \6321 , \6080 , \6149 );
or \U$4359 ( \6322 , \6319 , \6320 , \6321 );
and \U$4361 ( \6323 , \5511 , \5735 );
and \U$4362 ( \6324 , \5415 , \5732 );
nor \U$4363 ( \6325 , \6323 , \6324 );
xnor \U$4364 ( \6326 , \6325 , \5729 );
xor \U$4365 ( \6327 , 1'b0 , \6326 );
and \U$4366 ( \6328 , \5622 , \5771 );
and \U$4367 ( \6329 , \5643 , \5769 );
nor \U$4368 ( \6330 , \6328 , \6329 );
xnor \U$4369 ( \6331 , \6330 , \5797 );
xor \U$4370 ( \6332 , \6327 , \6331 );
and \U$4372 ( \6333 , \5957 , \5525 );
and \U$4373 ( \6334 , \5881 , \5523 );
nor \U$4374 ( \6335 , \6333 , \6334 );
xnor \U$4375 ( \6336 , \6335 , \5302 );
and \U$4376 ( \6337 , \6002 , \5463 );
and \U$4377 ( \6338 , \5936 , \5461 );
nor \U$4378 ( \6339 , \6337 , \6338 );
xnor \U$4379 ( \6340 , \6339 , \5489 );
xor \U$4380 ( \6341 , \6336 , \6340 );
and \U$4382 ( \6342 , \5981 , \5516 );
nor \U$4383 ( \6343 , 1'b0 , \6342 );
xnor \U$4384 ( \6344 , \6343 , 1'b0 );
xor \U$4385 ( \6345 , \6341 , \6344 );
xor \U$4386 ( \6346 , 1'b0 , \6345 );
xor \U$4387 ( \6347 , \6332 , \6346 );
and \U$4388 ( \6348 , \6138 , \6142 );
and \U$4389 ( \6349 , \6142 , \6147 );
and \U$4390 ( \6350 , \6138 , \6147 );
or \U$4391 ( \6351 , \6348 , \6349 , \6350 );
and \U$4392 ( \6352 , \6123 , \6127 );
and \U$4393 ( \6353 , \6127 , \6132 );
and \U$4394 ( \6354 , \6123 , \6132 );
or \U$4395 ( \6355 , \6352 , \6353 , \6354 );
xor \U$4396 ( \6356 , \6351 , \6355 );
and \U$4397 ( \6357 , \6114 , \6117 );
or \U$4400 ( \6358 , \6357 , 1'b0 , 1'b0 );
xor \U$4401 ( \6359 , \6356 , \6358 );
xor \U$4402 ( \6360 , \6347 , \6359 );
xor \U$4403 ( \6361 , \6322 , \6360 );
and \U$4404 ( \6362 , \6245 , \6249 );
and \U$4405 ( \6363 , \6249 , \6254 );
and \U$4406 ( \6364 , \6245 , \6254 );
or \U$4407 ( \6365 , \6362 , \6363 , \6364 );
and \U$4408 ( \6366 , \6119 , \6133 );
and \U$4409 ( \6367 , \6133 , \6148 );
and \U$4410 ( \6368 , \6119 , \6148 );
or \U$4411 ( \6369 , \6366 , \6367 , \6368 );
xor \U$4412 ( \6370 , \6365 , \6369 );
and \U$4413 ( \6371 , \5792 , \5831 );
and \U$4414 ( \6372 , \5666 , \5829 );
nor \U$4415 ( \6373 , \6371 , \6372 );
xnor \U$4416 ( \6374 , \6373 , \5857 );
and \U$4417 ( \6375 , \5852 , \5889 );
and \U$4418 ( \6376 , \5759 , \5887 );
nor \U$4419 ( \6377 , \6375 , \6376 );
xnor \U$4420 ( \6378 , \6377 , \5915 );
xor \U$4421 ( \6379 , \6374 , \6378 );
and \U$4422 ( \6380 , \5910 , \5590 );
and \U$4423 ( \6381 , \5819 , \5588 );
nor \U$4424 ( \6382 , \6380 , \6381 );
xnor \U$4425 ( \6383 , \6382 , \5595 );
xor \U$4426 ( \6384 , \6379 , \6383 );
xor \U$4427 ( \6385 , \6370 , \6384 );
xor \U$4428 ( \6386 , \6361 , \6385 );
xor \U$4429 ( \6387 , \6318 , \6386 );
and \U$4430 ( \6388 , \6150 , \6256 );
nor \U$4431 ( \6389 , \6387 , \6388 );
nor \U$4432 ( \6390 , \6314 , \6389 );
and \U$4433 ( \6391 , \6322 , \6360 );
and \U$4434 ( \6392 , \6360 , \6385 );
and \U$4435 ( \6393 , \6322 , \6385 );
or \U$4436 ( \6394 , \6391 , \6392 , \6393 );
and \U$4438 ( \6395 , \6326 , \6331 );
or \U$4440 ( \6396 , 1'b0 , \6395 , 1'b0 );
and \U$4441 ( \6397 , \6374 , \6378 );
and \U$4442 ( \6398 , \6378 , \6383 );
and \U$4443 ( \6399 , \6374 , \6383 );
or \U$4444 ( \6400 , \6397 , \6398 , \6399 );
xor \U$4445 ( \6401 , \6396 , \6400 );
and \U$4446 ( \6402 , \6336 , \6340 );
and \U$4447 ( \6403 , \6340 , \6344 );
and \U$4448 ( \6404 , \6336 , \6344 );
or \U$4449 ( \6405 , \6402 , \6403 , \6404 );
xor \U$4450 ( \6406 , \6401 , \6405 );
and \U$4451 ( \6407 , \6351 , \6355 );
and \U$4452 ( \6408 , \6355 , \6358 );
and \U$4453 ( \6409 , \6351 , \6358 );
or \U$4454 ( \6410 , \6407 , \6408 , \6409 );
xor \U$4456 ( \6411 , \6410 , 1'b0 );
and \U$4457 ( \6412 , \5415 , \5735 );
and \U$4458 ( \6413 , \5484 , \5732 );
nor \U$4459 ( \6414 , \6412 , \6413 );
xnor \U$4460 ( \6415 , \6414 , \5729 );
and \U$4461 ( \6416 , \5643 , \5771 );
and \U$4462 ( \6417 , \5511 , \5769 );
nor \U$4463 ( \6418 , \6416 , \6417 );
xnor \U$4464 ( \6419 , \6418 , \5797 );
xor \U$4465 ( \6420 , \6415 , \6419 );
and \U$4466 ( \6421 , \5666 , \5831 );
and \U$4467 ( \6422 , \5622 , \5829 );
nor \U$4468 ( \6423 , \6421 , \6422 );
xnor \U$4469 ( \6424 , \6423 , \5857 );
xor \U$4470 ( \6425 , \6420 , \6424 );
xor \U$4471 ( \6426 , \6411 , \6425 );
xor \U$4472 ( \6427 , \6406 , \6426 );
xor \U$4473 ( \6428 , \6394 , \6427 );
and \U$4474 ( \6429 , \6365 , \6369 );
and \U$4475 ( \6430 , \6369 , \6384 );
and \U$4476 ( \6431 , \6365 , \6384 );
or \U$4477 ( \6432 , \6429 , \6430 , \6431 );
and \U$4478 ( \6433 , \6332 , \6346 );
and \U$4479 ( \6434 , \6346 , \6359 );
and \U$4480 ( \6435 , \6332 , \6359 );
or \U$4481 ( \6436 , \6433 , \6434 , \6435 );
xor \U$4482 ( \6437 , \6432 , \6436 );
and \U$4484 ( \6438 , \5936 , \5463 );
and \U$4485 ( \6439 , \5957 , \5461 );
nor \U$4486 ( \6440 , \6438 , \6439 );
xnor \U$4487 ( \6441 , \6440 , \5489 );
and \U$4489 ( \6442 , \6002 , \5516 );
nor \U$4490 ( \6443 , 1'b0 , \6442 );
xnor \U$4491 ( \6444 , \6443 , 1'b0 );
xor \U$4492 ( \6445 , \6441 , \6444 );
xor \U$4494 ( \6446 , \6445 , 1'b0 );
xor \U$4495 ( \6447 , 1'b0 , \6446 );
and \U$4496 ( \6448 , \5759 , \5889 );
and \U$4497 ( \6449 , \5792 , \5887 );
nor \U$4498 ( \6450 , \6448 , \6449 );
xnor \U$4499 ( \6451 , \6450 , \5915 );
and \U$4500 ( \6452 , \5819 , \5590 );
and \U$4501 ( \6453 , \5852 , \5588 );
nor \U$4502 ( \6454 , \6452 , \6453 );
xnor \U$4503 ( \6455 , \6454 , \5595 );
xor \U$4504 ( \6456 , \6451 , \6455 );
and \U$4505 ( \6457 , \5881 , \5525 );
and \U$4506 ( \6458 , \5910 , \5523 );
nor \U$4507 ( \6459 , \6457 , \6458 );
xnor \U$4508 ( \6460 , \6459 , \5302 );
xor \U$4509 ( \6461 , \6456 , \6460 );
xor \U$4510 ( \6462 , \6447 , \6461 );
xor \U$4511 ( \6463 , \6437 , \6462 );
xor \U$4512 ( \6464 , \6428 , \6463 );
and \U$4513 ( \6465 , \6318 , \6386 );
nor \U$4514 ( \6466 , \6464 , \6465 );
and \U$4515 ( \6467 , \6432 , \6436 );
and \U$4516 ( \6468 , \6436 , \6462 );
and \U$4517 ( \6469 , \6432 , \6462 );
or \U$4518 ( \6470 , \6467 , \6468 , \6469 );
and \U$4519 ( \6471 , \6406 , \6426 );
xor \U$4520 ( \6472 , \6470 , \6471 );
and \U$4523 ( \6473 , \6410 , \6425 );
or \U$4524 ( \6474 , 1'b0 , 1'b0 , \6473 );
and \U$4526 ( \6475 , \5910 , \5525 );
and \U$4527 ( \6476 , \5819 , \5523 );
nor \U$4528 ( \6477 , \6475 , \6476 );
xnor \U$4529 ( \6478 , \6477 , \5302 );
and \U$4530 ( \6479 , \5957 , \5463 );
and \U$4531 ( \6480 , \5881 , \5461 );
nor \U$4532 ( \6481 , \6479 , \6480 );
xnor \U$4533 ( \6482 , \6481 , \5489 );
xor \U$4534 ( \6483 , \6478 , \6482 );
and \U$4536 ( \6484 , \5936 , \5516 );
nor \U$4537 ( \6485 , 1'b0 , \6484 );
xnor \U$4538 ( \6486 , \6485 , 1'b0 );
xor \U$4539 ( \6487 , \6483 , \6486 );
xor \U$4540 ( \6488 , 1'b0 , \6487 );
and \U$4541 ( \6489 , \5622 , \5831 );
and \U$4542 ( \6490 , \5643 , \5829 );
nor \U$4543 ( \6491 , \6489 , \6490 );
xnor \U$4544 ( \6492 , \6491 , \5857 );
and \U$4545 ( \6493 , \5792 , \5889 );
and \U$4546 ( \6494 , \5666 , \5887 );
nor \U$4547 ( \6495 , \6493 , \6494 );
xnor \U$4548 ( \6496 , \6495 , \5915 );
xor \U$4549 ( \6497 , \6492 , \6496 );
and \U$4550 ( \6498 , \5852 , \5590 );
and \U$4551 ( \6499 , \5759 , \5588 );
nor \U$4552 ( \6500 , \6498 , \6499 );
xnor \U$4553 ( \6501 , \6500 , \5595 );
xor \U$4554 ( \6502 , \6497 , \6501 );
xor \U$4555 ( \6503 , \6488 , \6502 );
and \U$4556 ( \6504 , \6415 , \6419 );
and \U$4557 ( \6505 , \6419 , \6424 );
and \U$4558 ( \6506 , \6415 , \6424 );
or \U$4559 ( \6507 , \6504 , \6505 , \6506 );
and \U$4560 ( \6508 , \6451 , \6455 );
and \U$4561 ( \6509 , \6455 , \6460 );
and \U$4562 ( \6510 , \6451 , \6460 );
or \U$4563 ( \6511 , \6508 , \6509 , \6510 );
xor \U$4564 ( \6512 , \6507 , \6511 );
and \U$4565 ( \6513 , \6441 , \6444 );
or \U$4568 ( \6514 , \6513 , 1'b0 , 1'b0 );
xor \U$4569 ( \6515 , \6512 , \6514 );
xor \U$4570 ( \6516 , \6503 , \6515 );
xor \U$4571 ( \6517 , \6474 , \6516 );
and \U$4572 ( \6518 , \6396 , \6400 );
and \U$4573 ( \6519 , \6400 , \6405 );
and \U$4574 ( \6520 , \6396 , \6405 );
or \U$4575 ( \6521 , \6518 , \6519 , \6520 );
and \U$4577 ( \6522 , \6446 , \6461 );
or \U$4579 ( \6523 , 1'b0 , \6522 , 1'b0 );
xor \U$4580 ( \6524 , \6521 , \6523 );
and \U$4582 ( \6525 , \5484 , \5735 );
not \U$4583 ( \6526 , \6525 );
xnor \U$4584 ( \6527 , \6526 , \5729 );
xor \U$4585 ( \6528 , 1'b0 , \6527 );
and \U$4586 ( \6529 , \5511 , \5771 );
and \U$4587 ( \6530 , \5415 , \5769 );
nor \U$4588 ( \6531 , \6529 , \6530 );
xnor \U$4589 ( \6532 , \6531 , \5797 );
xor \U$4590 ( \6533 , \6528 , \6532 );
xor \U$4591 ( \6534 , \6524 , \6533 );
xor \U$4592 ( \6535 , \6517 , \6534 );
xor \U$4593 ( \6536 , \6472 , \6535 );
and \U$4594 ( \6537 , \6394 , \6427 );
and \U$4595 ( \6538 , \6427 , \6463 );
and \U$4596 ( \6539 , \6394 , \6463 );
or \U$4597 ( \6540 , \6537 , \6538 , \6539 );
nor \U$4598 ( \6541 , \6536 , \6540 );
nor \U$4599 ( \6542 , \6466 , \6541 );
nand \U$4600 ( \6543 , \6390 , \6542 );
and \U$4601 ( \6544 , \6474 , \6516 );
and \U$4602 ( \6545 , \6516 , \6534 );
and \U$4603 ( \6546 , \6474 , \6534 );
or \U$4604 ( \6547 , \6544 , \6545 , \6546 );
and \U$4605 ( \6548 , \6507 , \6511 );
and \U$4606 ( \6549 , \6511 , \6514 );
and \U$4607 ( \6550 , \6507 , \6514 );
or \U$4608 ( \6551 , \6548 , \6549 , \6550 );
and \U$4610 ( \6552 , \6487 , \6502 );
or \U$4612 ( \6553 , 1'b0 , \6552 , 1'b0 );
xor \U$4613 ( \6554 , \6551 , \6553 );
and \U$4614 ( \6555 , \5666 , \5889 );
and \U$4615 ( \6556 , \5622 , \5887 );
nor \U$4616 ( \6557 , \6555 , \6556 );
xnor \U$4617 ( \6558 , \6557 , \5915 );
and \U$4618 ( \6559 , \5759 , \5590 );
and \U$4619 ( \6560 , \5792 , \5588 );
nor \U$4620 ( \6561 , \6559 , \6560 );
xnor \U$4621 ( \6562 , \6561 , \5595 );
xor \U$4622 ( \6563 , \6558 , \6562 );
and \U$4623 ( \6564 , \5819 , \5525 );
and \U$4624 ( \6565 , \5852 , \5523 );
nor \U$4625 ( \6566 , \6564 , \6565 );
xnor \U$4626 ( \6567 , \6566 , \5302 );
xor \U$4627 ( \6568 , \6563 , \6567 );
xor \U$4628 ( \6569 , \6554 , \6568 );
xor \U$4629 ( \6570 , \6547 , \6569 );
and \U$4630 ( \6571 , \6521 , \6523 );
and \U$4631 ( \6572 , \6523 , \6533 );
and \U$4632 ( \6573 , \6521 , \6533 );
or \U$4633 ( \6574 , \6571 , \6572 , \6573 );
and \U$4634 ( \6575 , \6503 , \6515 );
xor \U$4635 ( \6576 , \6574 , \6575 );
not \U$4636 ( \6577 , \5729 );
and \U$4637 ( \6578 , \5415 , \5771 );
and \U$4638 ( \6579 , \5484 , \5769 );
nor \U$4639 ( \6580 , \6578 , \6579 );
xnor \U$4640 ( \6581 , \6580 , \5797 );
xor \U$4641 ( \6582 , \6577 , \6581 );
and \U$4642 ( \6583 , \5643 , \5831 );
and \U$4643 ( \6584 , \5511 , \5829 );
nor \U$4644 ( \6585 , \6583 , \6584 );
xnor \U$4645 ( \6586 , \6585 , \5857 );
xor \U$4646 ( \6587 , \6582 , \6586 );
and \U$4648 ( \6588 , \5881 , \5463 );
and \U$4649 ( \6589 , \5910 , \5461 );
nor \U$4650 ( \6590 , \6588 , \6589 );
xnor \U$4651 ( \6591 , \6590 , \5489 );
and \U$4653 ( \6592 , \5957 , \5516 );
nor \U$4654 ( \6593 , 1'b0 , \6592 );
xnor \U$4655 ( \6594 , \6593 , 1'b0 );
xor \U$4656 ( \6595 , \6591 , \6594 );
xor \U$4658 ( \6596 , \6595 , 1'b0 );
xor \U$4659 ( \6597 , 1'b1 , \6596 );
xor \U$4660 ( \6598 , \6587 , \6597 );
and \U$4662 ( \6599 , \6527 , \6532 );
or \U$4664 ( \6600 , 1'b0 , \6599 , 1'b0 );
and \U$4665 ( \6601 , \6492 , \6496 );
and \U$4666 ( \6602 , \6496 , \6501 );
and \U$4667 ( \6603 , \6492 , \6501 );
or \U$4668 ( \6604 , \6601 , \6602 , \6603 );
xor \U$4669 ( \6605 , \6600 , \6604 );
and \U$4670 ( \6606 , \6478 , \6482 );
and \U$4671 ( \6607 , \6482 , \6486 );
and \U$4672 ( \6608 , \6478 , \6486 );
or \U$4673 ( \6609 , \6606 , \6607 , \6608 );
xor \U$4674 ( \6610 , \6605 , \6609 );
xor \U$4675 ( \6611 , \6598 , \6610 );
xor \U$4676 ( \6612 , \6576 , \6611 );
xor \U$4677 ( \6613 , \6570 , \6612 );
and \U$4678 ( \6614 , \6470 , \6471 );
and \U$4679 ( \6615 , \6471 , \6535 );
and \U$4680 ( \6616 , \6470 , \6535 );
or \U$4681 ( \6617 , \6614 , \6615 , \6616 );
nor \U$4682 ( \6618 , \6613 , \6617 );
and \U$4683 ( \6619 , \6574 , \6575 );
and \U$4684 ( \6620 , \6575 , \6611 );
and \U$4685 ( \6621 , \6574 , \6611 );
or \U$4686 ( \6622 , \6619 , \6620 , \6621 );
and \U$4687 ( \6623 , \6577 , \6581 );
and \U$4688 ( \6624 , \6581 , \6586 );
and \U$4689 ( \6625 , \6577 , \6586 );
or \U$4690 ( \6626 , \6623 , \6624 , \6625 );
and \U$4691 ( \6627 , \6558 , \6562 );
and \U$4692 ( \6628 , \6562 , \6567 );
and \U$4693 ( \6629 , \6558 , \6567 );
or \U$4694 ( \6630 , \6627 , \6628 , \6629 );
xor \U$4695 ( \6631 , \6626 , \6630 );
and \U$4696 ( \6632 , \6591 , \6594 );
or \U$4699 ( \6633 , \6632 , 1'b0 , 1'b0 );
xor \U$4700 ( \6634 , \6631 , \6633 );
and \U$4701 ( \6635 , \6600 , \6604 );
and \U$4702 ( \6636 , \6604 , \6609 );
and \U$4703 ( \6637 , \6600 , \6609 );
or \U$4704 ( \6638 , \6635 , \6636 , \6637 );
and \U$4707 ( \6639 , 1'b1 , \6596 );
or \U$4709 ( \6640 , 1'b0 , \6639 , 1'b0 );
xor \U$4710 ( \6641 , \6638 , \6640 );
and \U$4711 ( \6642 , \5910 , \5463 );
and \U$4712 ( \6643 , \5819 , \5461 );
nor \U$4713 ( \6644 , \6642 , \6643 );
xnor \U$4714 ( \6645 , \6644 , \5489 );
and \U$4716 ( \6646 , \5881 , \5516 );
nor \U$4717 ( \6647 , 1'b0 , \6646 );
xnor \U$4718 ( \6648 , \6647 , 1'b0 );
xor \U$4719 ( \6649 , \6645 , \6648 );
xor \U$4721 ( \6650 , \6649 , 1'b0 );
and \U$4722 ( \6651 , \5622 , \5889 );
and \U$4723 ( \6652 , \5643 , \5887 );
nor \U$4724 ( \6653 , \6651 , \6652 );
xnor \U$4725 ( \6654 , \6653 , \5915 );
and \U$4726 ( \6655 , \5792 , \5590 );
and \U$4727 ( \6656 , \5666 , \5588 );
nor \U$4728 ( \6657 , \6655 , \6656 );
xnor \U$4729 ( \6658 , \6657 , \5595 );
xor \U$4730 ( \6659 , \6654 , \6658 );
and \U$4731 ( \6660 , \5852 , \5525 );
and \U$4732 ( \6661 , \5759 , \5523 );
nor \U$4733 ( \6662 , \6660 , \6661 );
xnor \U$4734 ( \6663 , \6662 , \5302 );
xor \U$4735 ( \6664 , \6659 , \6663 );
xor \U$4736 ( \6665 , \6650 , \6664 );
and \U$4738 ( \6666 , \5484 , \5771 );
not \U$4739 ( \6667 , \6666 );
xnor \U$4740 ( \6668 , \6667 , \5797 );
xor \U$4741 ( \6669 , 1'b0 , \6668 );
and \U$4742 ( \6670 , \5511 , \5831 );
and \U$4743 ( \6671 , \5415 , \5829 );
nor \U$4744 ( \6672 , \6670 , \6671 );
xnor \U$4745 ( \6673 , \6672 , \5857 );
xor \U$4746 ( \6674 , \6669 , \6673 );
xor \U$4747 ( \6675 , \6665 , \6674 );
xor \U$4748 ( \6676 , \6641 , \6675 );
xor \U$4749 ( \6677 , \6634 , \6676 );
xor \U$4750 ( \6678 , \6622 , \6677 );
and \U$4751 ( \6679 , \6551 , \6553 );
and \U$4752 ( \6680 , \6553 , \6568 );
and \U$4753 ( \6681 , \6551 , \6568 );
or \U$4754 ( \6682 , \6679 , \6680 , \6681 );
and \U$4755 ( \6683 , \6587 , \6597 );
and \U$4756 ( \6684 , \6597 , \6610 );
and \U$4757 ( \6685 , \6587 , \6610 );
or \U$4758 ( \6686 , \6683 , \6684 , \6685 );
xor \U$4759 ( \6687 , \6682 , \6686 );
xor \U$4761 ( \6688 , \6687 , 1'b1 );
xor \U$4762 ( \6689 , \6678 , \6688 );
and \U$4763 ( \6690 , \6547 , \6569 );
and \U$4764 ( \6691 , \6569 , \6612 );
and \U$4765 ( \6692 , \6547 , \6612 );
or \U$4766 ( \6693 , \6690 , \6691 , \6692 );
nor \U$4767 ( \6694 , \6689 , \6693 );
nor \U$4768 ( \6695 , \6618 , \6694 );
and \U$4769 ( \6696 , \6682 , \6686 );
and \U$4770 ( \6697 , \6686 , 1'b1 );
and \U$4771 ( \6698 , \6682 , 1'b1 );
or \U$4772 ( \6699 , \6696 , \6697 , \6698 );
and \U$4773 ( \6700 , \6634 , \6676 );
xor \U$4774 ( \6701 , \6699 , \6700 );
and \U$4775 ( \6702 , \6638 , \6640 );
and \U$4776 ( \6703 , \6640 , \6675 );
and \U$4777 ( \6704 , \6638 , \6675 );
or \U$4778 ( \6705 , \6702 , \6703 , \6704 );
and \U$4780 ( \6706 , \5910 , \5516 );
nor \U$4781 ( \6707 , 1'b0 , \6706 );
xnor \U$4782 ( \6708 , \6707 , 1'b0 );
xor \U$4784 ( \6709 , \6708 , 1'b0 );
xor \U$4786 ( \6710 , \6709 , 1'b0 );
and \U$4787 ( \6711 , \5666 , \5590 );
and \U$4788 ( \6712 , \5622 , \5588 );
nor \U$4789 ( \6713 , \6711 , \6712 );
xnor \U$4790 ( \6714 , \6713 , \5595 );
and \U$4791 ( \6715 , \5759 , \5525 );
and \U$4792 ( \6716 , \5792 , \5523 );
nor \U$4793 ( \6717 , \6715 , \6716 );
xnor \U$4794 ( \6718 , \6717 , \5302 );
xor \U$4795 ( \6719 , \6714 , \6718 );
and \U$4796 ( \6720 , \5819 , \5463 );
and \U$4797 ( \6721 , \5852 , \5461 );
nor \U$4798 ( \6722 , \6720 , \6721 );
xnor \U$4799 ( \6723 , \6722 , \5489 );
xor \U$4800 ( \6724 , \6719 , \6723 );
xor \U$4801 ( \6725 , \6710 , \6724 );
not \U$4802 ( \6726 , \5797 );
and \U$4803 ( \6727 , \5415 , \5831 );
and \U$4804 ( \6728 , \5484 , \5829 );
nor \U$4805 ( \6729 , \6727 , \6728 );
xnor \U$4806 ( \6730 , \6729 , \5857 );
xor \U$4807 ( \6731 , \6726 , \6730 );
and \U$4808 ( \6732 , \5643 , \5889 );
and \U$4809 ( \6733 , \5511 , \5887 );
nor \U$4810 ( \6734 , \6732 , \6733 );
xnor \U$4811 ( \6735 , \6734 , \5915 );
xor \U$4812 ( \6736 , \6731 , \6735 );
xor \U$4813 ( \6737 , \6725 , \6736 );
xor \U$4815 ( \6738 , \6737 , 1'b0 );
and \U$4817 ( \6739 , \6668 , \6673 );
or \U$4819 ( \6740 , 1'b0 , \6739 , 1'b0 );
and \U$4820 ( \6741 , \6654 , \6658 );
and \U$4821 ( \6742 , \6658 , \6663 );
and \U$4822 ( \6743 , \6654 , \6663 );
or \U$4823 ( \6744 , \6741 , \6742 , \6743 );
xor \U$4824 ( \6745 , \6740 , \6744 );
and \U$4825 ( \6746 , \6645 , \6648 );
or \U$4828 ( \6747 , \6746 , 1'b0 , 1'b0 );
xor \U$4829 ( \6748 , \6745 , \6747 );
xor \U$4830 ( \6749 , \6738 , \6748 );
xor \U$4831 ( \6750 , \6705 , \6749 );
and \U$4832 ( \6751 , \6626 , \6630 );
and \U$4833 ( \6752 , \6630 , \6633 );
and \U$4834 ( \6753 , \6626 , \6633 );
or \U$4835 ( \6754 , \6751 , \6752 , \6753 );
xor \U$4837 ( \6755 , \6754 , 1'b0 );
and \U$4838 ( \6756 , \6650 , \6664 );
and \U$4839 ( \6757 , \6664 , \6674 );
and \U$4840 ( \6758 , \6650 , \6674 );
or \U$4841 ( \6759 , \6756 , \6757 , \6758 );
xor \U$4842 ( \6760 , \6755 , \6759 );
xor \U$4843 ( \6761 , \6750 , \6760 );
xor \U$4844 ( \6762 , \6701 , \6761 );
and \U$4845 ( \6763 , \6622 , \6677 );
and \U$4846 ( \6764 , \6677 , \6688 );
and \U$4847 ( \6765 , \6622 , \6688 );
or \U$4848 ( \6766 , \6763 , \6764 , \6765 );
nor \U$4849 ( \6767 , \6762 , \6766 );
and \U$4850 ( \6768 , \6705 , \6749 );
and \U$4851 ( \6769 , \6749 , \6760 );
and \U$4852 ( \6770 , \6705 , \6760 );
or \U$4853 ( \6771 , \6768 , \6769 , \6770 );
and \U$4854 ( \6772 , \6740 , \6744 );
and \U$4855 ( \6773 , \6744 , \6747 );
and \U$4856 ( \6774 , \6740 , \6747 );
or \U$4857 ( \6775 , \6772 , \6773 , \6774 );
xor \U$4859 ( \6776 , \6775 , 1'b0 );
and \U$4860 ( \6777 , \6710 , \6724 );
and \U$4861 ( \6778 , \6724 , \6736 );
and \U$4862 ( \6779 , \6710 , \6736 );
or \U$4863 ( \6780 , \6777 , \6778 , \6779 );
xor \U$4864 ( \6781 , \6776 , \6780 );
xor \U$4865 ( \6782 , \6771 , \6781 );
and \U$4868 ( \6783 , \6754 , \6759 );
or \U$4869 ( \6784 , 1'b0 , 1'b0 , \6783 );
and \U$4872 ( \6785 , \6737 , \6748 );
or \U$4873 ( \6786 , 1'b0 , 1'b0 , \6785 );
xor \U$4874 ( \6787 , \6784 , \6786 );
and \U$4875 ( \6788 , \5622 , \5590 );
and \U$4876 ( \6789 , \5643 , \5588 );
nor \U$4877 ( \6790 , \6788 , \6789 );
xnor \U$4878 ( \6791 , \6790 , \5595 );
and \U$4879 ( \6792 , \5792 , \5525 );
and \U$4880 ( \6793 , \5666 , \5523 );
nor \U$4881 ( \6794 , \6792 , \6793 );
xnor \U$4882 ( \6795 , \6794 , \5302 );
xor \U$4883 ( \6796 , \6791 , \6795 );
and \U$4884 ( \6797 , \5852 , \5463 );
and \U$4885 ( \6798 , \5759 , \5461 );
nor \U$4886 ( \6799 , \6797 , \6798 );
xnor \U$4887 ( \6800 , \6799 , \5489 );
xor \U$4888 ( \6801 , \6796 , \6800 );
and \U$4890 ( \6802 , \5484 , \5831 );
not \U$4891 ( \6803 , \6802 );
xnor \U$4892 ( \6804 , \6803 , \5857 );
xor \U$4893 ( \6805 , 1'b0 , \6804 );
and \U$4894 ( \6806 , \5511 , \5889 );
and \U$4895 ( \6807 , \5415 , \5887 );
nor \U$4896 ( \6808 , \6806 , \6807 );
xnor \U$4897 ( \6809 , \6808 , \5915 );
xor \U$4898 ( \6810 , \6805 , \6809 );
xor \U$4899 ( \6811 , \6801 , \6810 );
and \U$4902 ( \6812 , \5819 , \5516 );
nor \U$4903 ( \6813 , 1'b0 , \6812 );
xnor \U$4904 ( \6814 , \6813 , 1'b0 );
xor \U$4906 ( \6815 , \6814 , 1'b0 );
xor \U$4908 ( \6816 , \6815 , 1'b0 );
xnor \U$4909 ( \6817 , 1'b0 , \6816 );
xor \U$4910 ( \6818 , \6811 , \6817 );
and \U$4911 ( \6819 , \6726 , \6730 );
and \U$4912 ( \6820 , \6730 , \6735 );
and \U$4913 ( \6821 , \6726 , \6735 );
or \U$4914 ( \6822 , \6819 , \6820 , \6821 );
and \U$4915 ( \6823 , \6714 , \6718 );
and \U$4916 ( \6824 , \6718 , \6723 );
and \U$4917 ( \6825 , \6714 , \6723 );
or \U$4918 ( \6826 , \6823 , \6824 , \6825 );
xor \U$4919 ( \6827 , \6822 , \6826 );
xor \U$4921 ( \6828 , \6827 , 1'b0 );
xor \U$4922 ( \6829 , \6818 , \6828 );
xor \U$4923 ( \6830 , \6787 , \6829 );
xor \U$4924 ( \6831 , \6782 , \6830 );
and \U$4925 ( \6832 , \6699 , \6700 );
and \U$4926 ( \6833 , \6700 , \6761 );
and \U$4927 ( \6834 , \6699 , \6761 );
or \U$4928 ( \6835 , \6832 , \6833 , \6834 );
nor \U$4929 ( \6836 , \6831 , \6835 );
nor \U$4930 ( \6837 , \6767 , \6836 );
nand \U$4931 ( \6838 , \6695 , \6837 );
nor \U$4932 ( \6839 , \6543 , \6838 );
and \U$4933 ( \6840 , \6784 , \6786 );
and \U$4934 ( \6841 , \6786 , \6829 );
and \U$4935 ( \6842 , \6784 , \6829 );
or \U$4936 ( \6843 , \6840 , \6841 , \6842 );
and \U$4937 ( \6844 , \6822 , \6826 );
or \U$4940 ( \6845 , \6844 , 1'b0 , 1'b0 );
or \U$4941 ( \6846 , 1'b0 , \6816 );
xor \U$4942 ( \6847 , \6845 , \6846 );
and \U$4943 ( \6848 , \6801 , \6810 );
xor \U$4944 ( \6849 , \6847 , \6848 );
xor \U$4945 ( \6850 , \6843 , \6849 );
and \U$4948 ( \6851 , \6775 , \6780 );
or \U$4949 ( \6852 , 1'b0 , 1'b0 , \6851 );
and \U$4950 ( \6853 , \6811 , \6817 );
and \U$4951 ( \6854 , \6817 , \6828 );
and \U$4952 ( \6855 , \6811 , \6828 );
or \U$4953 ( \6856 , \6853 , \6854 , \6855 );
xor \U$4954 ( \6857 , \6852 , \6856 );
and \U$4956 ( \6858 , \5666 , \5525 );
and \U$4957 ( \6859 , \5622 , \5523 );
nor \U$4958 ( \6860 , \6858 , \6859 );
xnor \U$4959 ( \6861 , \6860 , \5302 );
and \U$4960 ( \6862 , \5759 , \5463 );
and \U$4961 ( \6863 , \5792 , \5461 );
nor \U$4962 ( \6864 , \6862 , \6863 );
xnor \U$4963 ( \6865 , \6864 , \5489 );
xor \U$4964 ( \6866 , \6861 , \6865 );
and \U$4966 ( \6867 , \5852 , \5516 );
nor \U$4967 ( \6868 , 1'b0 , \6867 );
xnor \U$4968 ( \6869 , \6868 , 1'b0 );
xor \U$4969 ( \6870 , \6866 , \6869 );
xor \U$4970 ( \6871 , 1'b0 , \6870 );
not \U$4971 ( \6872 , \5857 );
and \U$4972 ( \6873 , \5415 , \5889 );
and \U$4973 ( \6874 , \5484 , \5887 );
nor \U$4974 ( \6875 , \6873 , \6874 );
xnor \U$4975 ( \6876 , \6875 , \5915 );
xor \U$4976 ( \6877 , \6872 , \6876 );
and \U$4977 ( \6878 , \5643 , \5590 );
and \U$4978 ( \6879 , \5511 , \5588 );
nor \U$4979 ( \6880 , \6878 , \6879 );
xnor \U$4980 ( \6881 , \6880 , \5595 );
xor \U$4981 ( \6882 , \6877 , \6881 );
xor \U$4982 ( \6883 , \6871 , \6882 );
xor \U$4984 ( \6884 , \6883 , 1'b0 );
and \U$4986 ( \6885 , \6804 , \6809 );
or \U$4988 ( \6886 , 1'b0 , \6885 , 1'b0 );
and \U$4989 ( \6887 , \6791 , \6795 );
and \U$4990 ( \6888 , \6795 , \6800 );
and \U$4991 ( \6889 , \6791 , \6800 );
or \U$4992 ( \6890 , \6887 , \6888 , \6889 );
xor \U$4993 ( \6891 , \6886 , \6890 );
xor \U$4995 ( \6892 , \6891 , 1'b0 );
xor \U$4996 ( \6893 , \6884 , \6892 );
xor \U$4997 ( \6894 , \6857 , \6893 );
xor \U$4998 ( \6895 , \6850 , \6894 );
and \U$4999 ( \6896 , \6771 , \6781 );
and \U$5000 ( \6897 , \6781 , \6830 );
and \U$5001 ( \6898 , \6771 , \6830 );
or \U$5002 ( \6899 , \6896 , \6897 , \6898 );
nor \U$5003 ( \6900 , \6895 , \6899 );
and \U$5004 ( \6901 , \6852 , \6856 );
and \U$5005 ( \6902 , \6856 , \6893 );
and \U$5006 ( \6903 , \6852 , \6893 );
or \U$5007 ( \6904 , \6901 , \6902 , \6903 );
and \U$5008 ( \6905 , \6886 , \6890 );
or \U$5011 ( \6906 , \6905 , 1'b0 , 1'b0 );
xor \U$5013 ( \6907 , \6906 , 1'b0 );
and \U$5015 ( \6908 , \6870 , \6882 );
or \U$5017 ( \6909 , 1'b0 , \6908 , 1'b0 );
xor \U$5018 ( \6910 , \6907 , \6909 );
xor \U$5019 ( \6911 , \6904 , \6910 );
and \U$5020 ( \6912 , \6845 , \6846 );
and \U$5021 ( \6913 , \6846 , \6848 );
and \U$5022 ( \6914 , \6845 , \6848 );
or \U$5023 ( \6915 , \6912 , \6913 , \6914 );
and \U$5026 ( \6916 , \6883 , \6892 );
or \U$5027 ( \6917 , 1'b0 , 1'b0 , \6916 );
xor \U$5028 ( \6918 , \6915 , \6917 );
and \U$5029 ( \6919 , \5622 , \5525 );
and \U$5030 ( \6920 , \5643 , \5523 );
nor \U$5031 ( \6921 , \6919 , \6920 );
xnor \U$5032 ( \6922 , \6921 , \5302 );
and \U$5033 ( \6923 , \5792 , \5463 );
and \U$5034 ( \6924 , \5666 , \5461 );
nor \U$5035 ( \6925 , \6923 , \6924 );
xnor \U$5036 ( \6926 , \6925 , \5489 );
xor \U$5037 ( \6927 , \6922 , \6926 );
and \U$5039 ( \6928 , \5759 , \5516 );
nor \U$5040 ( \6929 , 1'b0 , \6928 );
xnor \U$5041 ( \6930 , \6929 , 1'b0 );
xor \U$5042 ( \6931 , \6927 , \6930 );
and \U$5044 ( \6932 , \5484 , \5889 );
not \U$5045 ( \6933 , \6932 );
xnor \U$5046 ( \6934 , \6933 , \5915 );
xor \U$5047 ( \6935 , 1'b0 , \6934 );
and \U$5048 ( \6936 , \5511 , \5590 );
and \U$5049 ( \6937 , \5415 , \5588 );
nor \U$5050 ( \6938 , \6936 , \6937 );
xnor \U$5051 ( \6939 , \6938 , \5595 );
xor \U$5052 ( \6940 , \6935 , \6939 );
xor \U$5053 ( \6941 , \6931 , \6940 );
xor \U$5055 ( \6942 , \6941 , 1'b1 );
and \U$5056 ( \6943 , \6872 , \6876 );
and \U$5057 ( \6944 , \6876 , \6881 );
and \U$5058 ( \6945 , \6872 , \6881 );
or \U$5059 ( \6946 , \6943 , \6944 , \6945 );
and \U$5060 ( \6947 , \6861 , \6865 );
and \U$5061 ( \6948 , \6865 , \6869 );
and \U$5062 ( \6949 , \6861 , \6869 );
or \U$5063 ( \6950 , \6947 , \6948 , \6949 );
xor \U$5064 ( \6951 , \6946 , \6950 );
xor \U$5066 ( \6952 , \6951 , 1'b0 );
xor \U$5067 ( \6953 , \6942 , \6952 );
xor \U$5068 ( \6954 , \6918 , \6953 );
xor \U$5069 ( \6955 , \6911 , \6954 );
and \U$5070 ( \6956 , \6843 , \6849 );
and \U$5071 ( \6957 , \6849 , \6894 );
and \U$5072 ( \6958 , \6843 , \6894 );
or \U$5073 ( \6959 , \6956 , \6957 , \6958 );
nor \U$5074 ( \6960 , \6955 , \6959 );
nor \U$5075 ( \6961 , \6900 , \6960 );
and \U$5076 ( \6962 , \6915 , \6917 );
and \U$5077 ( \6963 , \6917 , \6953 );
and \U$5078 ( \6964 , \6915 , \6953 );
or \U$5079 ( \6965 , \6962 , \6963 , \6964 );
and \U$5080 ( \6966 , \6946 , \6950 );
or \U$5083 ( \6967 , \6966 , 1'b0 , 1'b0 );
xor \U$5085 ( \6968 , \6967 , 1'b0 );
and \U$5086 ( \6969 , \6931 , \6940 );
xor \U$5087 ( \6970 , \6968 , \6969 );
xor \U$5088 ( \6971 , \6965 , \6970 );
and \U$5091 ( \6972 , \6906 , \6909 );
or \U$5092 ( \6973 , 1'b0 , 1'b0 , \6972 );
and \U$5093 ( \6974 , \6941 , 1'b1 );
and \U$5094 ( \6975 , 1'b1 , \6952 );
and \U$5095 ( \6976 , \6941 , \6952 );
or \U$5096 ( \6977 , \6974 , \6975 , \6976 );
xor \U$5097 ( \6978 , \6973 , \6977 );
and \U$5099 ( \6979 , \5666 , \5463 );
and \U$5100 ( \6980 , \5622 , \5461 );
nor \U$5101 ( \6981 , \6979 , \6980 );
xnor \U$5102 ( \6982 , \6981 , \5489 );
and \U$5104 ( \6983 , \5792 , \5516 );
nor \U$5105 ( \6984 , 1'b0 , \6983 );
xnor \U$5106 ( \6985 , \6984 , 1'b0 );
xor \U$5107 ( \6986 , \6982 , \6985 );
xor \U$5109 ( \6987 , \6986 , 1'b0 );
xor \U$5110 ( \6988 , 1'b0 , \6987 );
not \U$5111 ( \6989 , \5915 );
and \U$5112 ( \6990 , \5415 , \5590 );
and \U$5113 ( \6991 , \5484 , \5588 );
nor \U$5114 ( \6992 , \6990 , \6991 );
xnor \U$5115 ( \6993 , \6992 , \5595 );
xor \U$5116 ( \6994 , \6989 , \6993 );
and \U$5117 ( \6995 , \5643 , \5525 );
and \U$5118 ( \6996 , \5511 , \5523 );
nor \U$5119 ( \6997 , \6995 , \6996 );
xnor \U$5120 ( \6998 , \6997 , \5302 );
xor \U$5121 ( \6999 , \6994 , \6998 );
xor \U$5122 ( \7000 , \6988 , \6999 );
xor \U$5124 ( \7001 , \7000 , 1'b0 );
and \U$5126 ( \7002 , \6934 , \6939 );
or \U$5128 ( \7003 , 1'b0 , \7002 , 1'b0 );
and \U$5129 ( \7004 , \6922 , \6926 );
and \U$5130 ( \7005 , \6926 , \6930 );
and \U$5131 ( \7006 , \6922 , \6930 );
or \U$5132 ( \7007 , \7004 , \7005 , \7006 );
xor \U$5133 ( \7008 , \7003 , \7007 );
xor \U$5135 ( \7009 , \7008 , 1'b0 );
xor \U$5136 ( \7010 , \7001 , \7009 );
xor \U$5137 ( \7011 , \6978 , \7010 );
xor \U$5138 ( \7012 , \6971 , \7011 );
and \U$5139 ( \7013 , \6904 , \6910 );
and \U$5140 ( \7014 , \6910 , \6954 );
and \U$5141 ( \7015 , \6904 , \6954 );
or \U$5142 ( \7016 , \7013 , \7014 , \7015 );
nor \U$5143 ( \7017 , \7012 , \7016 );
and \U$5144 ( \7018 , \6973 , \6977 );
and \U$5145 ( \7019 , \6977 , \7010 );
and \U$5146 ( \7020 , \6973 , \7010 );
or \U$5147 ( \7021 , \7018 , \7019 , \7020 );
and \U$5148 ( \7022 , \7003 , \7007 );
or \U$5151 ( \7023 , \7022 , 1'b0 , 1'b0 );
xor \U$5153 ( \7024 , \7023 , 1'b0 );
and \U$5155 ( \7025 , \6987 , \6999 );
or \U$5157 ( \7026 , 1'b0 , \7025 , 1'b0 );
xor \U$5158 ( \7027 , \7024 , \7026 );
xor \U$5159 ( \7028 , \7021 , \7027 );
and \U$5162 ( \7029 , \6967 , \6969 );
or \U$5163 ( \7030 , 1'b0 , 1'b0 , \7029 );
and \U$5166 ( \7031 , \7000 , \7009 );
or \U$5167 ( \7032 , 1'b0 , 1'b0 , \7031 );
xor \U$5168 ( \7033 , \7030 , \7032 );
xor \U$5169 ( \7034 , \5646 , \5669 );
xor \U$5171 ( \7035 , \7034 , 1'b0 );
xor \U$5173 ( \7036 , 1'b0 , \5596 );
xor \U$5174 ( \7037 , \7036 , \5600 );
xor \U$5175 ( \7038 , \7035 , \7037 );
xor \U$5177 ( \7039 , \7038 , 1'b1 );
and \U$5178 ( \7040 , \6989 , \6993 );
and \U$5179 ( \7041 , \6993 , \6998 );
and \U$5180 ( \7042 , \6989 , \6998 );
or \U$5181 ( \7043 , \7040 , \7041 , \7042 );
and \U$5182 ( \7044 , \6982 , \6985 );
or \U$5185 ( \7045 , \7044 , 1'b0 , 1'b0 );
xor \U$5186 ( \7046 , \7043 , \7045 );
xor \U$5188 ( \7047 , \7046 , 1'b0 );
xor \U$5189 ( \7048 , \7039 , \7047 );
xor \U$5190 ( \7049 , \7033 , \7048 );
xor \U$5191 ( \7050 , \7028 , \7049 );
and \U$5192 ( \7051 , \6965 , \6970 );
and \U$5193 ( \7052 , \6970 , \7011 );
and \U$5194 ( \7053 , \6965 , \7011 );
or \U$5195 ( \7054 , \7051 , \7052 , \7053 );
nor \U$5196 ( \7055 , \7050 , \7054 );
nor \U$5197 ( \7056 , \7017 , \7055 );
nand \U$5198 ( \7057 , \6961 , \7056 );
and \U$5199 ( \7058 , \7030 , \7032 );
and \U$5200 ( \7059 , \7032 , \7048 );
and \U$5201 ( \7060 , \7030 , \7048 );
or \U$5202 ( \7061 , \7058 , \7059 , \7060 );
and \U$5203 ( \7062 , \7043 , \7045 );
or \U$5206 ( \7063 , \7062 , 1'b0 , 1'b0 );
xor \U$5208 ( \7064 , \7063 , 1'b0 );
and \U$5209 ( \7065 , \7035 , \7037 );
xor \U$5210 ( \7066 , \7064 , \7065 );
xor \U$5211 ( \7067 , \7061 , \7066 );
and \U$5214 ( \7068 , \7023 , \7026 );
or \U$5215 ( \7069 , 1'b0 , 1'b0 , \7068 );
and \U$5216 ( \7070 , \7038 , 1'b1 );
and \U$5217 ( \7071 , 1'b1 , \7047 );
and \U$5218 ( \7072 , \7038 , \7047 );
or \U$5219 ( \7073 , \7070 , \7071 , \7072 );
xor \U$5220 ( \7074 , \7069 , \7073 );
xor \U$5222 ( \7075 , 1'b0 , \5678 );
xor \U$5223 ( \7076 , \7075 , \5689 );
xor \U$5225 ( \7077 , \7076 , 1'b0 );
xor \U$5226 ( \7078 , \5602 , \5671 );
xor \U$5228 ( \7079 , \7078 , 1'b0 );
xor \U$5229 ( \7080 , \7077 , \7079 );
xor \U$5230 ( \7081 , \7074 , \7080 );
xor \U$5231 ( \7082 , \7067 , \7081 );
and \U$5232 ( \7083 , \7021 , \7027 );
and \U$5233 ( \7084 , \7027 , \7049 );
and \U$5234 ( \7085 , \7021 , \7049 );
or \U$5235 ( \7086 , \7083 , \7084 , \7085 );
nor \U$5236 ( \7087 , \7082 , \7086 );
and \U$5237 ( \7088 , \7069 , \7073 );
and \U$5238 ( \7089 , \7073 , \7080 );
and \U$5239 ( \7090 , \7069 , \7080 );
or \U$5240 ( \7091 , \7088 , \7089 , \7090 );
xor \U$5242 ( \7092 , \5673 , 1'b0 );
xor \U$5243 ( \7093 , \7092 , \5691 );
xor \U$5244 ( \7094 , \7091 , \7093 );
and \U$5247 ( \7095 , \7063 , \7065 );
or \U$5248 ( \7096 , 1'b0 , 1'b0 , \7095 );
and \U$5251 ( \7097 , \7076 , \7079 );
or \U$5252 ( \7098 , 1'b0 , 1'b0 , \7097 );
xor \U$5253 ( \7099 , \7096 , \7098 );
xor \U$5254 ( \7100 , \5701 , 1'b1 );
xor \U$5255 ( \7101 , \7100 , \5708 );
xor \U$5256 ( \7102 , \7099 , \7101 );
xor \U$5257 ( \7103 , \7094 , \7102 );
and \U$5258 ( \7104 , \7061 , \7066 );
and \U$5259 ( \7105 , \7066 , \7081 );
and \U$5260 ( \7106 , \7061 , \7081 );
or \U$5261 ( \7107 , \7104 , \7105 , \7106 );
nor \U$5262 ( \7108 , \7103 , \7107 );
nor \U$5263 ( \7109 , \7087 , \7108 );
and \U$5264 ( \7110 , \7096 , \7098 );
and \U$5265 ( \7111 , \7098 , \7101 );
and \U$5266 ( \7112 , \7096 , \7101 );
or \U$5267 ( \7113 , \7110 , \7111 , \7112 );
and \U$5269 ( \7114 , \5698 , \5700 );
xor \U$5270 ( \7115 , 1'b0 , \7114 );
xor \U$5271 ( \7116 , \7113 , \7115 );
xor \U$5272 ( \7117 , \5693 , \5711 );
xor \U$5273 ( \7118 , \7117 , \5714 );
xor \U$5274 ( \7119 , \7116 , \7118 );
and \U$5275 ( \7120 , \7091 , \7093 );
and \U$5276 ( \7121 , \7093 , \7102 );
and \U$5277 ( \7122 , \7091 , \7102 );
or \U$5278 ( \7123 , \7120 , \7121 , \7122 );
nor \U$5279 ( \7124 , \7119 , \7123 );
xor \U$5281 ( \7125 , \5717 , 1'b0 );
xor \U$5282 ( \7126 , \7125 , \5719 );
and \U$5283 ( \7127 , \7113 , \7115 );
and \U$5284 ( \7128 , \7115 , \7118 );
and \U$5285 ( \7129 , \7113 , \7118 );
or \U$5286 ( \7130 , \7127 , \7128 , \7129 );
nor \U$5287 ( \7131 , \7126 , \7130 );
nor \U$5288 ( \7132 , \7124 , \7131 );
nand \U$5289 ( \7133 , \7109 , \7132 );
nor \U$5290 ( \7134 , \7057 , \7133 );
nand \U$5291 ( \7135 , \6839 , \7134 );
and \U$5292 ( \7136 , \5936 , \5735 );
and \U$5293 ( \7137 , \5957 , \5732 );
nor \U$5294 ( \7138 , \7136 , \7137 );
xnor \U$5295 ( \7139 , \7138 , \5729 );
and \U$5296 ( \7140 , \5981 , \5771 );
and \U$5297 ( \7141 , \6002 , \5769 );
nor \U$5298 ( \7142 , \7140 , \7141 );
xnor \U$5299 ( \7143 , \7142 , \5797 );
and \U$5300 ( \7144 , \7139 , \7143 );
and \U$5301 ( \7145 , \6029 , \5831 );
and \U$5302 ( \7146 , \6050 , \5829 );
nor \U$5303 ( \7147 , \7145 , \7146 );
xnor \U$5304 ( \7148 , \7147 , \5857 );
and \U$5305 ( \7149 , \7143 , \7148 );
and \U$5306 ( \7150 , \7139 , \7148 );
or \U$5307 ( \7151 , \7144 , \7149 , \7150 );
and \U$5308 ( \7152 , \6050 , \5831 );
and \U$5309 ( \7153 , \5981 , \5829 );
nor \U$5310 ( \7154 , \7152 , \7153 );
xnor \U$5311 ( \7155 , \7154 , \5857 );
and \U$5312 ( \7156 , \6073 , \5889 );
and \U$5313 ( \7157 , \6029 , \5887 );
nor \U$5314 ( \7158 , \7156 , \7157 );
xnor \U$5315 ( \7159 , \7158 , \5915 );
xor \U$5316 ( \7160 , \7155 , \7159 );
nand \U$5317 ( \7161 , \6206 , \5588 );
xnor \U$5318 ( \7162 , \7161 , \5595 );
xor \U$5319 ( \7163 , \7160 , \7162 );
and \U$5320 ( \7164 , \7151 , \7163 );
and \U$5321 ( \7165 , \5957 , \5735 );
and \U$5322 ( \7166 , \5881 , \5732 );
nor \U$5323 ( \7167 , \7165 , \7166 );
xnor \U$5324 ( \7168 , \7167 , \5729 );
xor \U$5325 ( \7169 , \5595 , \7168 );
and \U$5326 ( \7170 , \6002 , \5771 );
and \U$5327 ( \7171 , \5936 , \5769 );
nor \U$5328 ( \7172 , \7170 , \7171 );
xnor \U$5329 ( \7173 , \7172 , \5797 );
xor \U$5330 ( \7174 , \7169 , \7173 );
and \U$5331 ( \7175 , \7163 , \7174 );
and \U$5332 ( \7176 , \7151 , \7174 );
or \U$5333 ( \7177 , \7164 , \7175 , \7176 );
and \U$5334 ( \7178 , \6206 , \5590 );
and \U$5335 ( \7179 , \6073 , \5588 );
nor \U$5336 ( \7180 , \7178 , \7179 );
xnor \U$5337 ( \7181 , \7180 , \5595 );
and \U$5338 ( \7182 , \5881 , \5735 );
and \U$5339 ( \7183 , \5910 , \5732 );
nor \U$5340 ( \7184 , \7182 , \7183 );
xnor \U$5341 ( \7185 , \7184 , \5729 );
and \U$5342 ( \7186 , \5936 , \5771 );
and \U$5343 ( \7187 , \5957 , \5769 );
nor \U$5344 ( \7188 , \7186 , \7187 );
xnor \U$5345 ( \7189 , \7188 , \5797 );
xor \U$5346 ( \7190 , \7185 , \7189 );
and \U$5347 ( \7191 , \5981 , \5831 );
and \U$5348 ( \7192 , \6002 , \5829 );
nor \U$5349 ( \7193 , \7191 , \7192 );
xnor \U$5350 ( \7194 , \7193 , \5857 );
xor \U$5351 ( \7195 , \7190 , \7194 );
xor \U$5352 ( \7196 , \7181 , \7195 );
xor \U$5353 ( \7197 , \7177 , \7196 );
and \U$5354 ( \7198 , \5595 , \7168 );
and \U$5355 ( \7199 , \7168 , \7173 );
and \U$5356 ( \7200 , \5595 , \7173 );
or \U$5357 ( \7201 , \7198 , \7199 , \7200 );
and \U$5358 ( \7202 , \7155 , \7159 );
and \U$5359 ( \7203 , \7159 , \7162 );
and \U$5360 ( \7204 , \7155 , \7162 );
or \U$5361 ( \7205 , \7202 , \7203 , \7204 );
xor \U$5362 ( \7206 , \7201 , \7205 );
and \U$5363 ( \7207 , \6029 , \5889 );
and \U$5364 ( \7208 , \6050 , \5887 );
nor \U$5365 ( \7209 , \7207 , \7208 );
xnor \U$5366 ( \7210 , \7209 , \5915 );
xor \U$5367 ( \7211 , \7206 , \7210 );
xor \U$5368 ( \7212 , \7197 , \7211 );
and \U$5369 ( \7213 , \6002 , \5735 );
and \U$5370 ( \7214 , \5936 , \5732 );
nor \U$5371 ( \7215 , \7213 , \7214 );
xnor \U$5372 ( \7216 , \7215 , \5729 );
and \U$5373 ( \7217 , \5915 , \7216 );
and \U$5374 ( \7218 , \6050 , \5771 );
and \U$5375 ( \7219 , \5981 , \5769 );
nor \U$5376 ( \7220 , \7218 , \7219 );
xnor \U$5377 ( \7221 , \7220 , \5797 );
and \U$5378 ( \7222 , \7216 , \7221 );
and \U$5379 ( \7223 , \5915 , \7221 );
or \U$5380 ( \7224 , \7217 , \7222 , \7223 );
and \U$5381 ( \7225 , \6073 , \5831 );
and \U$5382 ( \7226 , \6029 , \5829 );
nor \U$5383 ( \7227 , \7225 , \7226 );
xnor \U$5384 ( \7228 , \7227 , \5857 );
nand \U$5385 ( \7229 , \6206 , \5887 );
xnor \U$5386 ( \7230 , \7229 , \5915 );
and \U$5387 ( \7231 , \7228 , \7230 );
and \U$5388 ( \7232 , \7224 , \7231 );
and \U$5389 ( \7233 , \6206 , \5889 );
and \U$5390 ( \7234 , \6073 , \5887 );
nor \U$5391 ( \7235 , \7233 , \7234 );
xnor \U$5392 ( \7236 , \7235 , \5915 );
and \U$5393 ( \7237 , \7231 , \7236 );
and \U$5394 ( \7238 , \7224 , \7236 );
or \U$5395 ( \7239 , \7232 , \7237 , \7238 );
xor \U$5396 ( \7240 , \7151 , \7163 );
xor \U$5397 ( \7241 , \7240 , \7174 );
and \U$5398 ( \7242 , \7239 , \7241 );
nor \U$5399 ( \7243 , \7212 , \7242 );
and \U$5400 ( \7244 , \7185 , \7189 );
and \U$5401 ( \7245 , \7189 , \7194 );
and \U$5402 ( \7246 , \7185 , \7194 );
or \U$5403 ( \7247 , \7244 , \7245 , \7246 );
nand \U$5404 ( \7248 , \6206 , \5523 );
xnor \U$5405 ( \7249 , \7248 , \5302 );
xor \U$5406 ( \7250 , \7247 , \7249 );
and \U$5407 ( \7251 , \6002 , \5831 );
and \U$5408 ( \7252 , \5936 , \5829 );
nor \U$5409 ( \7253 , \7251 , \7252 );
xnor \U$5410 ( \7254 , \7253 , \5857 );
and \U$5411 ( \7255 , \6050 , \5889 );
and \U$5412 ( \7256 , \5981 , \5887 );
nor \U$5413 ( \7257 , \7255 , \7256 );
xnor \U$5414 ( \7258 , \7257 , \5915 );
xor \U$5415 ( \7259 , \7254 , \7258 );
and \U$5416 ( \7260 , \6073 , \5590 );
and \U$5417 ( \7261 , \6029 , \5588 );
nor \U$5418 ( \7262 , \7260 , \7261 );
xnor \U$5419 ( \7263 , \7262 , \5595 );
xor \U$5420 ( \7264 , \7259 , \7263 );
xor \U$5421 ( \7265 , \7250 , \7264 );
and \U$5422 ( \7266 , \7201 , \7205 );
and \U$5423 ( \7267 , \7205 , \7210 );
and \U$5424 ( \7268 , \7201 , \7210 );
or \U$5425 ( \7269 , \7266 , \7267 , \7268 );
and \U$5426 ( \7270 , \7181 , \7195 );
xor \U$5427 ( \7271 , \7269 , \7270 );
and \U$5428 ( \7272 , \5910 , \5735 );
and \U$5429 ( \7273 , \5819 , \5732 );
nor \U$5430 ( \7274 , \7272 , \7273 );
xnor \U$5431 ( \7275 , \7274 , \5729 );
xor \U$5432 ( \7276 , \5302 , \7275 );
and \U$5433 ( \7277 , \5957 , \5771 );
and \U$5434 ( \7278 , \5881 , \5769 );
nor \U$5435 ( \7279 , \7277 , \7278 );
xnor \U$5436 ( \7280 , \7279 , \5797 );
xor \U$5437 ( \7281 , \7276 , \7280 );
xor \U$5438 ( \7282 , \7271 , \7281 );
xor \U$5439 ( \7283 , \7265 , \7282 );
and \U$5440 ( \7284 , \7177 , \7196 );
and \U$5441 ( \7285 , \7196 , \7211 );
and \U$5442 ( \7286 , \7177 , \7211 );
or \U$5443 ( \7287 , \7284 , \7285 , \7286 );
nor \U$5444 ( \7288 , \7283 , \7287 );
nor \U$5445 ( \7289 , \7243 , \7288 );
and \U$5446 ( \7290 , \7269 , \7270 );
and \U$5447 ( \7291 , \7270 , \7281 );
and \U$5448 ( \7292 , \7269 , \7281 );
or \U$5449 ( \7293 , \7290 , \7291 , \7292 );
and \U$5450 ( \7294 , \7247 , \7249 );
and \U$5451 ( \7295 , \7249 , \7264 );
and \U$5452 ( \7296 , \7247 , \7264 );
or \U$5453 ( \7297 , \7294 , \7295 , \7296 );
and \U$5454 ( \7298 , \5819 , \5735 );
and \U$5455 ( \7299 , \5852 , \5732 );
nor \U$5456 ( \7300 , \7298 , \7299 );
xnor \U$5457 ( \7301 , \7300 , \5729 );
and \U$5458 ( \7302 , \5881 , \5771 );
and \U$5459 ( \7303 , \5910 , \5769 );
nor \U$5460 ( \7304 , \7302 , \7303 );
xnor \U$5461 ( \7305 , \7304 , \5797 );
xor \U$5462 ( \7306 , \7301 , \7305 );
and \U$5463 ( \7307 , \5936 , \5831 );
and \U$5464 ( \7308 , \5957 , \5829 );
nor \U$5465 ( \7309 , \7307 , \7308 );
xnor \U$5466 ( \7310 , \7309 , \5857 );
xor \U$5467 ( \7311 , \7306 , \7310 );
xor \U$5468 ( \7312 , \7297 , \7311 );
and \U$5469 ( \7313 , \5302 , \7275 );
and \U$5470 ( \7314 , \7275 , \7280 );
and \U$5471 ( \7315 , \5302 , \7280 );
or \U$5472 ( \7316 , \7313 , \7314 , \7315 );
and \U$5473 ( \7317 , \7254 , \7258 );
and \U$5474 ( \7318 , \7258 , \7263 );
and \U$5475 ( \7319 , \7254 , \7263 );
or \U$5476 ( \7320 , \7317 , \7318 , \7319 );
xor \U$5477 ( \7321 , \7316 , \7320 );
and \U$5478 ( \7322 , \5981 , \5889 );
and \U$5479 ( \7323 , \6002 , \5887 );
nor \U$5480 ( \7324 , \7322 , \7323 );
xnor \U$5481 ( \7325 , \7324 , \5915 );
and \U$5482 ( \7326 , \6029 , \5590 );
and \U$5483 ( \7327 , \6050 , \5588 );
nor \U$5484 ( \7328 , \7326 , \7327 );
xnor \U$5485 ( \7329 , \7328 , \5595 );
xor \U$5486 ( \7330 , \7325 , \7329 );
and \U$5487 ( \7331 , \6206 , \5525 );
and \U$5488 ( \7332 , \6073 , \5523 );
nor \U$5489 ( \7333 , \7331 , \7332 );
xnor \U$5490 ( \7334 , \7333 , \5302 );
xor \U$5491 ( \7335 , \7330 , \7334 );
xor \U$5492 ( \7336 , \7321 , \7335 );
xor \U$5493 ( \7337 , \7312 , \7336 );
xor \U$5494 ( \7338 , \7293 , \7337 );
and \U$5495 ( \7339 , \7265 , \7282 );
nor \U$5496 ( \7340 , \7338 , \7339 );
and \U$5497 ( \7341 , \7297 , \7311 );
and \U$5498 ( \7342 , \7311 , \7336 );
and \U$5499 ( \7343 , \7297 , \7336 );
or \U$5500 ( \7344 , \7341 , \7342 , \7343 );
and \U$5501 ( \7345 , \7316 , \7320 );
and \U$5502 ( \7346 , \7320 , \7335 );
and \U$5503 ( \7347 , \7316 , \7335 );
or \U$5504 ( \7348 , \7345 , \7346 , \7347 );
nand \U$5505 ( \7349 , \6206 , \5461 );
xnor \U$5506 ( \7350 , \7349 , \5489 );
and \U$5507 ( \7351 , \5957 , \5831 );
and \U$5508 ( \7352 , \5881 , \5829 );
nor \U$5509 ( \7353 , \7351 , \7352 );
xnor \U$5510 ( \7354 , \7353 , \5857 );
and \U$5511 ( \7355 , \6002 , \5889 );
and \U$5512 ( \7356 , \5936 , \5887 );
nor \U$5513 ( \7357 , \7355 , \7356 );
xnor \U$5514 ( \7358 , \7357 , \5915 );
xor \U$5515 ( \7359 , \7354 , \7358 );
and \U$5516 ( \7360 , \6050 , \5590 );
and \U$5517 ( \7361 , \5981 , \5588 );
nor \U$5518 ( \7362 , \7360 , \7361 );
xnor \U$5519 ( \7363 , \7362 , \5595 );
xor \U$5520 ( \7364 , \7359 , \7363 );
xor \U$5521 ( \7365 , \7350 , \7364 );
and \U$5522 ( \7366 , \5852 , \5735 );
and \U$5523 ( \7367 , \5759 , \5732 );
nor \U$5524 ( \7368 , \7366 , \7367 );
xnor \U$5525 ( \7369 , \7368 , \5729 );
xor \U$5526 ( \7370 , \5489 , \7369 );
and \U$5527 ( \7371 , \5910 , \5771 );
and \U$5528 ( \7372 , \5819 , \5769 );
nor \U$5529 ( \7373 , \7371 , \7372 );
xnor \U$5530 ( \7374 , \7373 , \5797 );
xor \U$5531 ( \7375 , \7370 , \7374 );
xor \U$5532 ( \7376 , \7365 , \7375 );
xor \U$5533 ( \7377 , \7348 , \7376 );
and \U$5534 ( \7378 , \7301 , \7305 );
and \U$5535 ( \7379 , \7305 , \7310 );
and \U$5536 ( \7380 , \7301 , \7310 );
or \U$5537 ( \7381 , \7378 , \7379 , \7380 );
and \U$5538 ( \7382 , \7325 , \7329 );
and \U$5539 ( \7383 , \7329 , \7334 );
and \U$5540 ( \7384 , \7325 , \7334 );
or \U$5541 ( \7385 , \7382 , \7383 , \7384 );
xor \U$5542 ( \7386 , \7381 , \7385 );
and \U$5543 ( \7387 , \6073 , \5525 );
and \U$5544 ( \7388 , \6029 , \5523 );
nor \U$5545 ( \7389 , \7387 , \7388 );
xnor \U$5546 ( \7390 , \7389 , \5302 );
xor \U$5547 ( \7391 , \7386 , \7390 );
xor \U$5548 ( \7392 , \7377 , \7391 );
xor \U$5549 ( \7393 , \7344 , \7392 );
and \U$5550 ( \7394 , \7293 , \7337 );
nor \U$5551 ( \7395 , \7393 , \7394 );
nor \U$5552 ( \7396 , \7340 , \7395 );
nand \U$5553 ( \7397 , \7289 , \7396 );
and \U$5554 ( \7398 , \7348 , \7376 );
and \U$5555 ( \7399 , \7376 , \7391 );
and \U$5556 ( \7400 , \7348 , \7391 );
or \U$5557 ( \7401 , \7398 , \7399 , \7400 );
xor \U$5558 ( \7402 , \6261 , \6265 );
xor \U$5559 ( \7403 , \7402 , \6270 );
and \U$5560 ( \7404 , \5489 , \7369 );
and \U$5561 ( \7405 , \7369 , \7374 );
and \U$5562 ( \7406 , \5489 , \7374 );
or \U$5563 ( \7407 , \7404 , \7405 , \7406 );
and \U$5564 ( \7408 , \7354 , \7358 );
and \U$5565 ( \7409 , \7358 , \7363 );
and \U$5566 ( \7410 , \7354 , \7363 );
or \U$5567 ( \7411 , \7408 , \7409 , \7410 );
xor \U$5568 ( \7412 , \7407 , \7411 );
and \U$5569 ( \7413 , \6206 , \5463 );
and \U$5570 ( \7414 , \6073 , \5461 );
nor \U$5571 ( \7415 , \7413 , \7414 );
xnor \U$5572 ( \7416 , \7415 , \5489 );
xor \U$5573 ( \7417 , \7412 , \7416 );
xor \U$5574 ( \7418 , \7403 , \7417 );
xor \U$5575 ( \7419 , \7401 , \7418 );
and \U$5576 ( \7420 , \7381 , \7385 );
and \U$5577 ( \7421 , \7385 , \7390 );
and \U$5578 ( \7422 , \7381 , \7390 );
or \U$5579 ( \7423 , \7420 , \7421 , \7422 );
and \U$5580 ( \7424 , \7350 , \7364 );
and \U$5581 ( \7425 , \7364 , \7375 );
and \U$5582 ( \7426 , \7350 , \7375 );
or \U$5583 ( \7427 , \7424 , \7425 , \7426 );
xor \U$5584 ( \7428 , \7423 , \7427 );
xor \U$5585 ( \7429 , \6277 , \6281 );
xor \U$5586 ( \7430 , \7429 , \6286 );
xor \U$5587 ( \7431 , \7428 , \7430 );
xor \U$5588 ( \7432 , \7419 , \7431 );
and \U$5589 ( \7433 , \7344 , \7392 );
nor \U$5590 ( \7434 , \7432 , \7433 );
and \U$5591 ( \7435 , \7423 , \7427 );
and \U$5592 ( \7436 , \7427 , \7430 );
and \U$5593 ( \7437 , \7423 , \7430 );
or \U$5594 ( \7438 , \7435 , \7436 , \7437 );
and \U$5595 ( \7439 , \7403 , \7417 );
xor \U$5596 ( \7440 , \7438 , \7439 );
and \U$5597 ( \7441 , \7407 , \7411 );
and \U$5598 ( \7442 , \7411 , \7416 );
and \U$5599 ( \7443 , \7407 , \7416 );
or \U$5600 ( \7444 , \7441 , \7442 , \7443 );
xor \U$5601 ( \7445 , \6297 , \6299 );
xor \U$5602 ( \7446 , \7444 , \7445 );
xor \U$5603 ( \7447 , \6273 , \6289 );
xor \U$5604 ( \7448 , \7447 , \6292 );
xor \U$5605 ( \7449 , \7446 , \7448 );
xor \U$5606 ( \7450 , \7440 , \7449 );
and \U$5607 ( \7451 , \7401 , \7418 );
and \U$5608 ( \7452 , \7418 , \7431 );
and \U$5609 ( \7453 , \7401 , \7431 );
or \U$5610 ( \7454 , \7451 , \7452 , \7453 );
nor \U$5611 ( \7455 , \7450 , \7454 );
nor \U$5612 ( \7456 , \7434 , \7455 );
and \U$5613 ( \7457 , \7444 , \7445 );
and \U$5614 ( \7458 , \7445 , \7448 );
and \U$5615 ( \7459 , \7444 , \7448 );
or \U$5616 ( \7460 , \7457 , \7458 , \7459 );
xor \U$5617 ( \7461 , \6160 , \6176 );
xor \U$5618 ( \7462 , \7461 , \6211 );
xor \U$5619 ( \7463 , \7460 , \7462 );
xor \U$5620 ( \7464 , \6295 , \6300 );
xor \U$5621 ( \7465 , \7464 , \6303 );
xor \U$5622 ( \7466 , \7463 , \7465 );
and \U$5623 ( \7467 , \7438 , \7439 );
and \U$5624 ( \7468 , \7439 , \7449 );
and \U$5625 ( \7469 , \7438 , \7449 );
or \U$5626 ( \7470 , \7467 , \7468 , \7469 );
nor \U$5627 ( \7471 , \7466 , \7470 );
xor \U$5628 ( \7472 , \6306 , \6307 );
xor \U$5629 ( \7473 , \7472 , \6310 );
and \U$5630 ( \7474 , \7460 , \7462 );
and \U$5631 ( \7475 , \7462 , \7465 );
and \U$5632 ( \7476 , \7460 , \7465 );
or \U$5633 ( \7477 , \7474 , \7475 , \7476 );
nor \U$5634 ( \7478 , \7473 , \7477 );
nor \U$5635 ( \7479 , \7471 , \7478 );
nand \U$5636 ( \7480 , \7456 , \7479 );
nor \U$5637 ( \7481 , \7397 , \7480 );
and \U$5638 ( \7482 , \6050 , \5735 );
and \U$5639 ( \7483 , \5981 , \5732 );
nor \U$5640 ( \7484 , \7482 , \7483 );
xnor \U$5641 ( \7485 , \7484 , \5729 );
and \U$5642 ( \7486 , \5857 , \7485 );
and \U$5643 ( \7487 , \6073 , \5771 );
and \U$5644 ( \7488 , \6029 , \5769 );
nor \U$5645 ( \7489 , \7487 , \7488 );
xnor \U$5646 ( \7490 , \7489 , \5797 );
and \U$5647 ( \7491 , \7485 , \7490 );
and \U$5648 ( \7492 , \5857 , \7490 );
or \U$5649 ( \7493 , \7486 , \7491 , \7492 );
and \U$5650 ( \7494 , \5981 , \5735 );
and \U$5651 ( \7495 , \6002 , \5732 );
nor \U$5652 ( \7496 , \7494 , \7495 );
xnor \U$5653 ( \7497 , \7496 , \5729 );
and \U$5654 ( \7498 , \6029 , \5771 );
and \U$5655 ( \7499 , \6050 , \5769 );
nor \U$5656 ( \7500 , \7498 , \7499 );
xnor \U$5657 ( \7501 , \7500 , \5797 );
xor \U$5658 ( \7502 , \7497 , \7501 );
and \U$5659 ( \7503 , \6206 , \5831 );
and \U$5660 ( \7504 , \6073 , \5829 );
nor \U$5661 ( \7505 , \7503 , \7504 );
xnor \U$5662 ( \7506 , \7505 , \5857 );
xor \U$5663 ( \7507 , \7502 , \7506 );
xor \U$5664 ( \7508 , \7493 , \7507 );
nand \U$5665 ( \7509 , \6206 , \5829 );
xnor \U$5666 ( \7510 , \7509 , \5857 );
xor \U$5667 ( \7511 , \5857 , \7485 );
xor \U$5668 ( \7512 , \7511 , \7490 );
and \U$5669 ( \7513 , \7510 , \7512 );
nor \U$5670 ( \7514 , \7508 , \7513 );
and \U$5671 ( \7515 , \7497 , \7501 );
and \U$5672 ( \7516 , \7501 , \7506 );
and \U$5673 ( \7517 , \7497 , \7506 );
or \U$5674 ( \7518 , \7515 , \7516 , \7517 );
xor \U$5675 ( \7519 , \7228 , \7230 );
xor \U$5676 ( \7520 , \7518 , \7519 );
xor \U$5677 ( \7521 , \5915 , \7216 );
xor \U$5678 ( \7522 , \7521 , \7221 );
xor \U$5679 ( \7523 , \7520 , \7522 );
and \U$5680 ( \7524 , \7493 , \7507 );
nor \U$5681 ( \7525 , \7523 , \7524 );
nor \U$5682 ( \7526 , \7514 , \7525 );
xor \U$5683 ( \7527 , \7139 , \7143 );
xor \U$5684 ( \7528 , \7527 , \7148 );
xor \U$5685 ( \7529 , \7224 , \7231 );
xor \U$5686 ( \7530 , \7529 , \7236 );
xor \U$5687 ( \7531 , \7528 , \7530 );
and \U$5688 ( \7532 , \7518 , \7519 );
and \U$5689 ( \7533 , \7519 , \7522 );
and \U$5690 ( \7534 , \7518 , \7522 );
or \U$5691 ( \7535 , \7532 , \7533 , \7534 );
nor \U$5692 ( \7536 , \7531 , \7535 );
xor \U$5693 ( \7537 , \7239 , \7241 );
and \U$5694 ( \7538 , \7528 , \7530 );
nor \U$5695 ( \7539 , \7537 , \7538 );
nor \U$5696 ( \7540 , \7536 , \7539 );
nand \U$5697 ( \7541 , \7526 , \7540 );
and \U$5698 ( \7542 , \6029 , \5735 );
and \U$5699 ( \7543 , \6050 , \5732 );
nor \U$5700 ( \7544 , \7542 , \7543 );
xnor \U$5701 ( \7545 , \7544 , \5729 );
and \U$5702 ( \7546 , \6206 , \5771 );
and \U$5703 ( \7547 , \6073 , \5769 );
nor \U$5704 ( \7548 , \7546 , \7547 );
xnor \U$5705 ( \7549 , \7548 , \5797 );
xor \U$5706 ( \7550 , \7545 , \7549 );
and \U$5707 ( \7551 , \6073 , \5735 );
and \U$5708 ( \7552 , \6029 , \5732 );
nor \U$5709 ( \7553 , \7551 , \7552 );
xnor \U$5710 ( \7554 , \7553 , \5729 );
and \U$5711 ( \7555 , \7554 , \5797 );
nor \U$5712 ( \7556 , \7550 , \7555 );
xor \U$5713 ( \7557 , \7510 , \7512 );
and \U$5714 ( \7558 , \7545 , \7549 );
nor \U$5715 ( \7559 , \7557 , \7558 );
nor \U$5716 ( \7560 , \7556 , \7559 );
xor \U$5717 ( \7561 , \7554 , \5797 );
nand \U$5718 ( \7562 , \6206 , \5769 );
xnor \U$5719 ( \7563 , \7562 , \5797 );
nor \U$5720 ( \7564 , \7561 , \7563 );
and \U$5721 ( \7565 , \6206 , \5735 );
and \U$5722 ( \7566 , \6073 , \5732 );
nor \U$5723 ( \7567 , \7565 , \7566 );
xnor \U$5724 ( \7568 , \7567 , \5729 );
nand \U$5725 ( \7569 , \6206 , \5732 );
xnor \U$5726 ( \7570 , \7569 , \5729 );
and \U$5727 ( \7571 , \7570 , \5729 );
nand \U$5728 ( \7572 , \7568 , \7571 );
or \U$5729 ( \7573 , \7564 , \7572 );
nand \U$5730 ( \7574 , \7561 , \7563 );
nand \U$5731 ( \7575 , \7573 , \7574 );
and \U$5732 ( \7576 , \7560 , \7575 );
nand \U$5733 ( \7577 , \7550 , \7555 );
or \U$5734 ( \7578 , \7559 , \7577 );
nand \U$5735 ( \7579 , \7557 , \7558 );
nand \U$5736 ( \7580 , \7578 , \7579 );
nor \U$5737 ( \7581 , \7576 , \7580 );
or \U$5738 ( \7582 , \7541 , \7581 );
nand \U$5739 ( \7583 , \7508 , \7513 );
or \U$5740 ( \7584 , \7525 , \7583 );
nand \U$5741 ( \7585 , \7523 , \7524 );
nand \U$5742 ( \7586 , \7584 , \7585 );
and \U$5743 ( \7587 , \7540 , \7586 );
nand \U$5744 ( \7588 , \7531 , \7535 );
or \U$5745 ( \7589 , \7539 , \7588 );
nand \U$5746 ( \7590 , \7537 , \7538 );
nand \U$5747 ( \7591 , \7589 , \7590 );
nor \U$5748 ( \7592 , \7587 , \7591 );
nand \U$5749 ( \7593 , \7582 , \7592 );
and \U$5750 ( \7594 , \7481 , \7593 );
nand \U$5751 ( \7595 , \7212 , \7242 );
or \U$5752 ( \7596 , \7288 , \7595 );
nand \U$5753 ( \7597 , \7283 , \7287 );
nand \U$5754 ( \7598 , \7596 , \7597 );
and \U$5755 ( \7599 , \7396 , \7598 );
nand \U$5756 ( \7600 , \7338 , \7339 );
or \U$5757 ( \7601 , \7395 , \7600 );
nand \U$5758 ( \7602 , \7393 , \7394 );
nand \U$5759 ( \7603 , \7601 , \7602 );
nor \U$5760 ( \7604 , \7599 , \7603 );
or \U$5761 ( \7605 , \7480 , \7604 );
nand \U$5762 ( \7606 , \7432 , \7433 );
or \U$5763 ( \7607 , \7455 , \7606 );
nand \U$5764 ( \7608 , \7450 , \7454 );
nand \U$5765 ( \7609 , \7607 , \7608 );
and \U$5766 ( \7610 , \7479 , \7609 );
nand \U$5767 ( \7611 , \7466 , \7470 );
or \U$5768 ( \7612 , \7478 , \7611 );
nand \U$5769 ( \7613 , \7473 , \7477 );
nand \U$5770 ( \7614 , \7612 , \7613 );
nor \U$5771 ( \7615 , \7610 , \7614 );
nand \U$5772 ( \7616 , \7605 , \7615 );
nor \U$5773 ( \7617 , \7594 , \7616 );
or \U$5774 ( \7618 , \7135 , \7617 );
nand \U$5775 ( \7619 , \6257 , \6313 );
or \U$5776 ( \7620 , \6389 , \7619 );
nand \U$5777 ( \7621 , \6387 , \6388 );
nand \U$5778 ( \7622 , \7620 , \7621 );
and \U$5779 ( \7623 , \6542 , \7622 );
nand \U$5780 ( \7624 , \6464 , \6465 );
or \U$5781 ( \7625 , \6541 , \7624 );
nand \U$5782 ( \7626 , \6536 , \6540 );
nand \U$5783 ( \7627 , \7625 , \7626 );
nor \U$5784 ( \7628 , \7623 , \7627 );
or \U$5785 ( \7629 , \6838 , \7628 );
nand \U$5786 ( \7630 , \6613 , \6617 );
or \U$5787 ( \7631 , \6694 , \7630 );
nand \U$5788 ( \7632 , \6689 , \6693 );
nand \U$5789 ( \7633 , \7631 , \7632 );
and \U$5790 ( \7634 , \6837 , \7633 );
nand \U$5791 ( \7635 , \6762 , \6766 );
or \U$5792 ( \7636 , \6836 , \7635 );
nand \U$5793 ( \7637 , \6831 , \6835 );
nand \U$5794 ( \7638 , \7636 , \7637 );
nor \U$5795 ( \7639 , \7634 , \7638 );
nand \U$5796 ( \7640 , \7629 , \7639 );
and \U$5797 ( \7641 , \7134 , \7640 );
nand \U$5798 ( \7642 , \6895 , \6899 );
or \U$5799 ( \7643 , \6960 , \7642 );
nand \U$5800 ( \7644 , \6955 , \6959 );
nand \U$5801 ( \7645 , \7643 , \7644 );
and \U$5802 ( \7646 , \7056 , \7645 );
nand \U$5803 ( \7647 , \7012 , \7016 );
or \U$5804 ( \7648 , \7055 , \7647 );
nand \U$5805 ( \7649 , \7050 , \7054 );
nand \U$5806 ( \7650 , \7648 , \7649 );
nor \U$5807 ( \7651 , \7646 , \7650 );
or \U$5808 ( \7652 , \7133 , \7651 );
nand \U$5809 ( \7653 , \7082 , \7086 );
or \U$5810 ( \7654 , \7108 , \7653 );
nand \U$5811 ( \7655 , \7103 , \7107 );
nand \U$5812 ( \7656 , \7654 , \7655 );
and \U$5813 ( \7657 , \7132 , \7656 );
nand \U$5814 ( \7658 , \7119 , \7123 );
or \U$5815 ( \7659 , \7131 , \7658 );
nand \U$5816 ( \7660 , \7126 , \7130 );
nand \U$5817 ( \7661 , \7659 , \7660 );
nor \U$5818 ( \7662 , \7657 , \7661 );
nand \U$5819 ( \7663 , \7652 , \7662 );
nor \U$5820 ( \7664 , \7641 , \7663 );
nand \U$5821 ( \7665 , \7618 , \7664 );
not \U$5822 ( \7666 , \7665 );
xor \U$5823 ( \7667 , \5725 , \7666 );
buf \U$5824 ( \7668 , \7667 );
buf \U$5825 ( \7669 , RI2b5e785ebd68_1);
buf \U$5826 ( \7670 , RI2b5e785ebcf0_2);
buf \U$5827 ( \7671 , RI2b5e785ebc78_3);
buf \U$5828 ( \7672 , RI2b5e785ebc00_4);
buf \U$5829 ( \7673 , RI2b5e785ebb88_5);
buf \U$5830 ( \7674 , RI2b5e785ebb10_6);
buf \U$5831 ( \7675 , RI2b5e785eba98_7);
buf \U$5832 ( \7676 , RI2b5e785eba20_8);
buf \U$5833 ( \7677 , RI2b5e785eb9a8_9);
buf \U$5834 ( \7678 , RI2b5e785eb930_10);
buf \U$5835 ( \7679 , RI2b5e785eb8b8_11);
buf \U$5836 ( \7680 , RI2b5e785eb840_12);
not \U$5837 ( \7681 , RI2b5e785ae328_614);
buf \U$5838 ( \7682 , \7681 );
and \U$5839 ( \7683 , \7680 , \7682 );
and \U$5840 ( \7684 , \7679 , \7683 );
and \U$5841 ( \7685 , \7678 , \7684 );
and \U$5842 ( \7686 , \7677 , \7685 );
and \U$5843 ( \7687 , \7676 , \7686 );
and \U$5844 ( \7688 , \7675 , \7687 );
and \U$5845 ( \7689 , \7674 , \7688 );
and \U$5846 ( \7690 , \7673 , \7689 );
and \U$5847 ( \7691 , \7672 , \7690 );
and \U$5848 ( \7692 , \7671 , \7691 );
and \U$5849 ( \7693 , \7670 , \7692 );
xor \U$5850 ( \7694 , \7669 , \7693 );
buf \U$5851 ( \7695 , \7694 );
buf \U$5852 ( \7696 , \7695 );
not \U$5853 ( \7697 , \7696 );
nor \U$5854 ( \7698 , \4917 , \4921 , \4925 , \4929 , \4934 );
and \U$5855 ( \7699 , RI2b5e785daab8_27, \7698 );
and \U$5856 ( \7700 , \4917 , \4921 , \4925 , \4929 , \4934 );
and \U$5857 ( \7701 , RI2b5e785495b8_40, \7700 );
and \U$5858 ( \7702 , \4939 , \4921 , \4925 , \4929 , \4934 );
and \U$5859 ( \7703 , RI2b5e78538920_53, \7702 );
and \U$5860 ( \7704 , \4917 , \4942 , \4925 , \4929 , \4934 );
and \U$5861 ( \7705 , RI2b5e784a63a8_66, \7704 );
and \U$5862 ( \7706 , \4939 , \4942 , \4925 , \4929 , \4934 );
and \U$5863 ( \7707 , RI2b5e78495710_79, \7706 );
and \U$5864 ( \7708 , \4917 , \4921 , \4947 , \4929 , \4934 );
and \U$5865 ( \7709 , RI2b5e784950f8_92, \7708 );
and \U$5866 ( \7710 , \4939 , \4921 , \4947 , \4929 , \4934 );
and \U$5867 ( \7711 , RI2b5e78403bf8_105, \7710 );
and \U$5868 ( \7712 , \4917 , \4942 , \4947 , \4929 , \4934 );
and \U$5869 ( \7713 , RI2b5e775b1ed8_118, \7712 );
and \U$5870 ( \7714 , \4939 , \4942 , \4947 , \4929 , \4934 );
and \U$5871 ( \7715 , RI2b5e775b18c0_131, \7714 );
nor \U$5872 ( \7716 , \4939 , \4942 , \4947 , \4929 , \4933 );
and \U$5873 ( \7717 , RI2b5e7750b858_144, \7716 );
nor \U$5874 ( \7718 , \4917 , \4942 , \4947 , \4929 , \4933 );
and \U$5875 ( \7719 , RI2b5e774ff030_157, \7718 );
nor \U$5876 ( \7720 , \4939 , \4921 , \4947 , \4929 , \4933 );
and \U$5877 ( \7721 , RI2b5e774f6048_170, \7720 );
nor \U$5878 ( \7722 , \4917 , \4921 , \4947 , \4929 , \4933 );
and \U$5879 ( \7723 , RI2b5e774ea630_183, \7722 );
nor \U$5880 ( \7724 , \4939 , \4942 , \4925 , \4929 , \4933 );
and \U$5881 ( \7725 , RI2b5e774dde08_196, \7724 );
nor \U$5882 ( \7726 , \4917 , \4942 , \4925 , \4929 , \4933 );
and \U$5883 ( \7727 , RI2b5e774d4e20_209, \7726 );
nor \U$5884 ( \7728 , \4939 , \4921 , \4925 , \4929 , \4933 );
and \U$5885 ( \7729 , RI2b5e785f3d60_222, \7728 );
nor \U$5886 ( \7730 , \4917 , \4921 , \4925 , \4929 , \4933 );
and \U$5887 ( \7731 , RI2b5e785eb138_235, \7730 );
or \U$5888 ( \7732 , \7699 , \7701 , \7703 , \7705 , \7707 , \7709 , \7711 , \7713 , \7715 , \7717 , \7719 , \7721 , \7723 , \7725 , \7727 , \7729 , \7731 );
buf \U$5889 ( \7733 , \4933 );
buf \U$5890 ( \7734 , \4917 );
buf \U$5891 ( \7735 , \4921 );
buf \U$5892 ( \7736 , \4925 );
buf \U$5893 ( \7737 , \4929 );
or \U$5894 ( \7738 , \7734 , \7735 , \7736 , \7737 );
and \U$5895 ( \7739 , \7733 , \7738 );
buf \U$5896 ( \7740 , \7739 );
_DC rfe6 ( \7741_nRfe6 , \7732 , \7740 );
buf \U$5897 ( \7742 , \7741_nRfe6 );
and \U$5898 ( \7743 , \7697 , \7742 );
xor \U$5899 ( \7744 , \7670 , \7692 );
buf \U$5900 ( \7745 , \7744 );
buf \U$5901 ( \7746 , \7745 );
not \U$5902 ( \7747 , \7746 );
and \U$5903 ( \7748 , RI2b5e785daa40_28, \7698 );
and \U$5904 ( \7749 , RI2b5e78549540_41, \7700 );
and \U$5905 ( \7750 , RI2b5e785388a8_54, \7702 );
and \U$5906 ( \7751 , RI2b5e784a6330_67, \7704 );
and \U$5907 ( \7752 , RI2b5e78495698_80, \7706 );
and \U$5908 ( \7753 , RI2b5e78495080_93, \7708 );
and \U$5909 ( \7754 , RI2b5e78403b80_106, \7710 );
and \U$5910 ( \7755 , RI2b5e775b1e60_119, \7712 );
and \U$5911 ( \7756 , RI2b5e7750bdf8_132, \7714 );
and \U$5912 ( \7757 , RI2b5e774ff5d0_145, \7716 );
and \U$5913 ( \7758 , RI2b5e774f65e8_158, \7718 );
and \U$5914 ( \7759 , RI2b5e774eabd0_171, \7720 );
and \U$5915 ( \7760 , RI2b5e774de3a8_184, \7722 );
and \U$5916 ( \7761 , RI2b5e774d53c0_197, \7724 );
and \U$5917 ( \7762 , RI2b5e785f4300_210, \7726 );
and \U$5918 ( \7763 , RI2b5e785f3ce8_223, \7728 );
and \U$5919 ( \7764 , RI2b5e785eb0c0_236, \7730 );
or \U$5920 ( \7765 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 );
_DC rfff ( \7766_nRfff , \7765 , \7740 );
buf \U$5921 ( \7767 , \7766_nRfff );
and \U$5922 ( \7768 , \7747 , \7767 );
xor \U$5923 ( \7769 , \7671 , \7691 );
buf \U$5924 ( \7770 , \7769 );
buf \U$5925 ( \7771 , \7770 );
not \U$5926 ( \7772 , \7771 );
and \U$5927 ( \7773 , RI2b5e785da9c8_29, \7698 );
and \U$5928 ( \7774 , RI2b5e785494c8_42, \7700 );
and \U$5929 ( \7775 , RI2b5e78538830_55, \7702 );
and \U$5930 ( \7776 , RI2b5e784a62b8_68, \7704 );
and \U$5931 ( \7777 , RI2b5e78495620_81, \7706 );
and \U$5932 ( \7778 , RI2b5e78495008_94, \7708 );
and \U$5933 ( \7779 , RI2b5e78403b08_107, \7710 );
and \U$5934 ( \7780 , RI2b5e775b1de8_120, \7712 );
and \U$5935 ( \7781 , RI2b5e7750bd80_133, \7714 );
and \U$5936 ( \7782 , RI2b5e774ff558_146, \7716 );
and \U$5937 ( \7783 , RI2b5e774f6570_159, \7718 );
and \U$5938 ( \7784 , RI2b5e774eab58_172, \7720 );
and \U$5939 ( \7785 , RI2b5e774de330_185, \7722 );
and \U$5940 ( \7786 , RI2b5e774d5348_198, \7724 );
and \U$5941 ( \7787 , RI2b5e785f4288_211, \7726 );
and \U$5942 ( \7788 , RI2b5e785f3658_224, \7728 );
and \U$5943 ( \7789 , RI2b5e785eb048_237, \7730 );
or \U$5944 ( \7790 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 );
_DC r1018 ( \7791_nR1018 , \7790 , \7740 );
buf \U$5945 ( \7792 , \7791_nR1018 );
and \U$5946 ( \7793 , \7772 , \7792 );
xor \U$5947 ( \7794 , \7672 , \7690 );
buf \U$5948 ( \7795 , \7794 );
buf \U$5949 ( \7796 , \7795 );
not \U$5950 ( \7797 , \7796 );
and \U$5951 ( \7798 , RI2b5e785da950_30, \7698 );
and \U$5952 ( \7799 , RI2b5e78549450_43, \7700 );
and \U$5953 ( \7800 , RI2b5e785387b8_56, \7702 );
and \U$5954 ( \7801 , RI2b5e784a6240_69, \7704 );
and \U$5955 ( \7802 , RI2b5e784955a8_82, \7706 );
and \U$5956 ( \7803 , RI2b5e78494f90_95, \7708 );
and \U$5957 ( \7804 , RI2b5e78403a90_108, \7710 );
and \U$5958 ( \7805 , RI2b5e775b1d70_121, \7712 );
and \U$5959 ( \7806 , RI2b5e7750bd08_134, \7714 );
and \U$5960 ( \7807 , RI2b5e774ff4e0_147, \7716 );
and \U$5961 ( \7808 , RI2b5e774f64f8_160, \7718 );
and \U$5962 ( \7809 , RI2b5e774eaae0_173, \7720 );
and \U$5963 ( \7810 , RI2b5e774de2b8_186, \7722 );
and \U$5964 ( \7811 , RI2b5e774d52d0_199, \7724 );
and \U$5965 ( \7812 , RI2b5e785f4210_212, \7726 );
and \U$5966 ( \7813 , RI2b5e785eb5e8_225, \7728 );
and \U$5967 ( \7814 , RI2b5e785e6c50_238, \7730 );
or \U$5968 ( \7815 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 );
_DC r1031 ( \7816_nR1031 , \7815 , \7740 );
buf \U$5969 ( \7817 , \7816_nR1031 );
and \U$5970 ( \7818 , \7797 , \7817 );
xor \U$5971 ( \7819 , \7673 , \7689 );
buf \U$5972 ( \7820 , \7819 );
buf \U$5973 ( \7821 , \7820 );
not \U$5974 ( \7822 , \7821 );
and \U$5975 ( \7823 , RI2b5e785da8d8_31, \7698 );
and \U$5976 ( \7824 , RI2b5e785493d8_44, \7700 );
and \U$5977 ( \7825 , RI2b5e78538740_57, \7702 );
and \U$5978 ( \7826 , RI2b5e784a61c8_70, \7704 );
and \U$5979 ( \7827 , RI2b5e78495530_83, \7706 );
and \U$5980 ( \7828 , RI2b5e78494f18_96, \7708 );
and \U$5981 ( \7829 , RI2b5e78403a18_109, \7710 );
and \U$5982 ( \7830 , RI2b5e775b1cf8_122, \7712 );
and \U$5983 ( \7831 , RI2b5e7750bc90_135, \7714 );
and \U$5984 ( \7832 , RI2b5e774ff468_148, \7716 );
and \U$5985 ( \7833 , RI2b5e774f6480_161, \7718 );
and \U$5986 ( \7834 , RI2b5e774eaa68_174, \7720 );
and \U$5987 ( \7835 , RI2b5e774de240_187, \7722 );
and \U$5988 ( \7836 , RI2b5e774d5258_200, \7724 );
and \U$5989 ( \7837 , RI2b5e785f4198_213, \7726 );
and \U$5990 ( \7838 , RI2b5e785eb570_226, \7728 );
and \U$5991 ( \7839 , RI2b5e785e6bd8_239, \7730 );
or \U$5992 ( \7840 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 );
_DC r104a ( \7841_nR104a , \7840 , \7740 );
buf \U$5993 ( \7842 , \7841_nR104a );
and \U$5994 ( \7843 , \7822 , \7842 );
xor \U$5995 ( \7844 , \7674 , \7688 );
buf \U$5996 ( \7845 , \7844 );
buf \U$5997 ( \7846 , \7845 );
not \U$5998 ( \7847 , \7846 );
and \U$5999 ( \7848 , RI2b5e785da860_32, \7698 );
and \U$6000 ( \7849 , RI2b5e78549360_45, \7700 );
and \U$6001 ( \7850 , RI2b5e785386c8_58, \7702 );
and \U$6002 ( \7851 , RI2b5e784a6150_71, \7704 );
and \U$6003 ( \7852 , RI2b5e784954b8_84, \7706 );
and \U$6004 ( \7853 , RI2b5e78494ea0_97, \7708 );
and \U$6005 ( \7854 , RI2b5e784039a0_110, \7710 );
and \U$6006 ( \7855 , RI2b5e775b1c80_123, \7712 );
and \U$6007 ( \7856 , RI2b5e7750bc18_136, \7714 );
and \U$6008 ( \7857 , RI2b5e774ff3f0_149, \7716 );
and \U$6009 ( \7858 , RI2b5e774f6408_162, \7718 );
and \U$6010 ( \7859 , RI2b5e774ea9f0_175, \7720 );
and \U$6011 ( \7860 , RI2b5e774de1c8_188, \7722 );
and \U$6012 ( \7861 , RI2b5e774d51e0_201, \7724 );
and \U$6013 ( \7862 , RI2b5e785f4120_214, \7726 );
and \U$6014 ( \7863 , RI2b5e785eb4f8_227, \7728 );
and \U$6015 ( \7864 , RI2b5e785e64d0_240, \7730 );
or \U$6016 ( \7865 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 );
_DC r1063 ( \7866_nR1063 , \7865 , \7740 );
buf \U$6017 ( \7867 , \7866_nR1063 );
and \U$6018 ( \7868 , \7847 , \7867 );
xor \U$6019 ( \7869 , \7675 , \7687 );
buf \U$6020 ( \7870 , \7869 );
buf \U$6021 ( \7871 , \7870 );
not \U$6022 ( \7872 , \7871 );
and \U$6023 ( \7873 , RI2b5e78549900_33, \7698 );
and \U$6024 ( \7874 , RI2b5e78538c68_46, \7700 );
and \U$6025 ( \7875 , RI2b5e78538650_59, \7702 );
and \U$6026 ( \7876 , RI2b5e784a60d8_72, \7704 );
and \U$6027 ( \7877 , RI2b5e78495440_85, \7706 );
and \U$6028 ( \7878 , RI2b5e78494e28_98, \7708 );
and \U$6029 ( \7879 , RI2b5e78403928_111, \7710 );
and \U$6030 ( \7880 , RI2b5e775b1c08_124, \7712 );
and \U$6031 ( \7881 , RI2b5e7750bba0_137, \7714 );
and \U$6032 ( \7882 , RI2b5e774ff378_150, \7716 );
and \U$6033 ( \7883 , RI2b5e774f6390_163, \7718 );
and \U$6034 ( \7884 , RI2b5e774ea978_176, \7720 );
and \U$6035 ( \7885 , RI2b5e774de150_189, \7722 );
and \U$6036 ( \7886 , RI2b5e774d5168_202, \7724 );
and \U$6037 ( \7887 , RI2b5e785f40a8_215, \7726 );
and \U$6038 ( \7888 , RI2b5e785eb480_228, \7728 );
and \U$6039 ( \7889 , RI2b5e785da608_241, \7730 );
or \U$6040 ( \7890 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 );
_DC r107c ( \7891_nR107c , \7890 , \7740 );
buf \U$6041 ( \7892 , \7891_nR107c );
and \U$6042 ( \7893 , \7872 , \7892 );
xor \U$6043 ( \7894 , \7676 , \7686 );
buf \U$6044 ( \7895 , \7894 );
buf \U$6045 ( \7896 , \7895 );
not \U$6046 ( \7897 , \7896 );
and \U$6047 ( \7898 , RI2b5e78549888_34, \7698 );
and \U$6048 ( \7899 , RI2b5e78538bf0_47, \7700 );
and \U$6049 ( \7900 , RI2b5e785385d8_60, \7702 );
and \U$6050 ( \7901 , RI2b5e784a6060_73, \7704 );
and \U$6051 ( \7902 , RI2b5e784953c8_86, \7706 );
and \U$6052 ( \7903 , RI2b5e78403ec8_99, \7708 );
and \U$6053 ( \7904 , RI2b5e775b21a8_112, \7710 );
and \U$6054 ( \7905 , RI2b5e775b1b90_125, \7712 );
and \U$6055 ( \7906 , RI2b5e7750bb28_138, \7714 );
and \U$6056 ( \7907 , RI2b5e774ff300_151, \7716 );
and \U$6057 ( \7908 , RI2b5e774f6318_164, \7718 );
and \U$6058 ( \7909 , RI2b5e774ea900_177, \7720 );
and \U$6059 ( \7910 , RI2b5e774de0d8_190, \7722 );
and \U$6060 ( \7911 , RI2b5e774d50f0_203, \7724 );
and \U$6061 ( \7912 , RI2b5e785f4030_216, \7726 );
and \U$6062 ( \7913 , RI2b5e785eb408_229, \7728 );
and \U$6063 ( \7914 , RI2b5e785da590_242, \7730 );
or \U$6064 ( \7915 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 );
_DC r1095 ( \7916_nR1095 , \7915 , \7740 );
buf \U$6065 ( \7917 , \7916_nR1095 );
and \U$6066 ( \7918 , \7897 , \7917 );
xor \U$6067 ( \7919 , \7677 , \7685 );
buf \U$6068 ( \7920 , \7919 );
buf \U$6069 ( \7921 , \7920 );
not \U$6070 ( \7922 , \7921 );
and \U$6071 ( \7923 , RI2b5e78549810_35, \7698 );
and \U$6072 ( \7924 , RI2b5e78538b78_48, \7700 );
and \U$6073 ( \7925 , RI2b5e78538560_61, \7702 );
and \U$6074 ( \7926 , RI2b5e784a5fe8_74, \7704 );
and \U$6075 ( \7927 , RI2b5e78495350_87, \7706 );
and \U$6076 ( \7928 , RI2b5e78403e50_100, \7708 );
and \U$6077 ( \7929 , RI2b5e775b2130_113, \7710 );
and \U$6078 ( \7930 , RI2b5e775b1b18_126, \7712 );
and \U$6079 ( \7931 , RI2b5e7750bab0_139, \7714 );
and \U$6080 ( \7932 , RI2b5e774ff288_152, \7716 );
and \U$6081 ( \7933 , RI2b5e774f62a0_165, \7718 );
and \U$6082 ( \7934 , RI2b5e774ea888_178, \7720 );
and \U$6083 ( \7935 , RI2b5e774de060_191, \7722 );
and \U$6084 ( \7936 , RI2b5e774d5078_204, \7724 );
and \U$6085 ( \7937 , RI2b5e785f3fb8_217, \7726 );
and \U$6086 ( \7938 , RI2b5e785eb390_230, \7728 );
and \U$6087 ( \7939 , RI2b5e785da518_243, \7730 );
or \U$6088 ( \7940 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 );
_DC r10ae ( \7941_nR10ae , \7940 , \7740 );
buf \U$6089 ( \7942 , \7941_nR10ae );
and \U$6090 ( \7943 , \7922 , \7942 );
xor \U$6091 ( \7944 , \7678 , \7684 );
buf \U$6092 ( \7945 , \7944 );
buf \U$6093 ( \7946 , \7945 );
not \U$6094 ( \7947 , \7946 );
and \U$6095 ( \7948 , RI2b5e78549798_36, \7698 );
and \U$6096 ( \7949 , RI2b5e78538b00_49, \7700 );
and \U$6097 ( \7950 , RI2b5e785384e8_62, \7702 );
and \U$6098 ( \7951 , RI2b5e784a5f70_75, \7704 );
and \U$6099 ( \7952 , RI2b5e784952d8_88, \7706 );
and \U$6100 ( \7953 , RI2b5e78403dd8_101, \7708 );
and \U$6101 ( \7954 , RI2b5e775b20b8_114, \7710 );
and \U$6102 ( \7955 , RI2b5e775b1aa0_127, \7712 );
and \U$6103 ( \7956 , RI2b5e7750ba38_140, \7714 );
and \U$6104 ( \7957 , RI2b5e774ff210_153, \7716 );
and \U$6105 ( \7958 , RI2b5e774f6228_166, \7718 );
and \U$6106 ( \7959 , RI2b5e774ea810_179, \7720 );
and \U$6107 ( \7960 , RI2b5e774ddfe8_192, \7722 );
and \U$6108 ( \7961 , RI2b5e774d5000_205, \7724 );
and \U$6109 ( \7962 , RI2b5e785f3f40_218, \7726 );
and \U$6110 ( \7963 , RI2b5e785eb318_231, \7728 );
and \U$6111 ( \7964 , RI2b5e785da4a0_244, \7730 );
or \U$6112 ( \7965 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 );
_DC r10c7 ( \7966_nR10c7 , \7965 , \7740 );
buf \U$6113 ( \7967 , \7966_nR10c7 );
and \U$6114 ( \7968 , \7947 , \7967 );
xor \U$6115 ( \7969 , \7679 , \7683 );
buf \U$6116 ( \7970 , \7969 );
buf \U$6117 ( \7971 , \7970 );
not \U$6118 ( \7972 , \7971 );
and \U$6119 ( \7973 , RI2b5e78549720_37, \7698 );
and \U$6120 ( \7974 , RI2b5e78538a88_50, \7700 );
and \U$6121 ( \7975 , RI2b5e78538470_63, \7702 );
and \U$6122 ( \7976 , RI2b5e784a5ef8_76, \7704 );
and \U$6123 ( \7977 , RI2b5e78495260_89, \7706 );
and \U$6124 ( \7978 , RI2b5e78403d60_102, \7708 );
and \U$6125 ( \7979 , RI2b5e775b2040_115, \7710 );
and \U$6126 ( \7980 , RI2b5e775b1a28_128, \7712 );
and \U$6127 ( \7981 , RI2b5e7750b9c0_141, \7714 );
and \U$6128 ( \7982 , RI2b5e774ff198_154, \7716 );
and \U$6129 ( \7983 , RI2b5e774f61b0_167, \7718 );
and \U$6130 ( \7984 , RI2b5e774ea798_180, \7720 );
and \U$6131 ( \7985 , RI2b5e774ddf70_193, \7722 );
and \U$6132 ( \7986 , RI2b5e774d4f88_206, \7724 );
and \U$6133 ( \7987 , RI2b5e785f3ec8_219, \7726 );
and \U$6134 ( \7988 , RI2b5e785eb2a0_232, \7728 );
and \U$6135 ( \7989 , RI2b5e785da428_245, \7730 );
or \U$6136 ( \7990 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 );
_DC r10e0 ( \7991_nR10e0 , \7990 , \7740 );
buf \U$6137 ( \7992 , \7991_nR10e0 );
and \U$6138 ( \7993 , \7972 , \7992 );
xor \U$6139 ( \7994 , \7680 , \7682 );
buf \U$6140 ( \7995 , \7994 );
buf \U$6141 ( \7996 , \7995 );
not \U$6142 ( \7997 , \7996 );
and \U$6143 ( \7998 , RI2b5e785496a8_38, \7698 );
and \U$6144 ( \7999 , RI2b5e78538a10_51, \7700 );
and \U$6145 ( \8000 , RI2b5e785383f8_64, \7702 );
and \U$6146 ( \8001 , RI2b5e784a5e80_77, \7704 );
and \U$6147 ( \8002 , RI2b5e784951e8_90, \7706 );
and \U$6148 ( \8003 , RI2b5e78403ce8_103, \7708 );
and \U$6149 ( \8004 , RI2b5e775b1fc8_116, \7710 );
and \U$6150 ( \8005 , RI2b5e775b19b0_129, \7712 );
and \U$6151 ( \8006 , RI2b5e7750b948_142, \7714 );
and \U$6152 ( \8007 , RI2b5e774ff120_155, \7716 );
and \U$6153 ( \8008 , RI2b5e774f6138_168, \7718 );
and \U$6154 ( \8009 , RI2b5e774ea720_181, \7720 );
and \U$6155 ( \8010 , RI2b5e774ddef8_194, \7722 );
and \U$6156 ( \8011 , RI2b5e774d4f10_207, \7724 );
and \U$6157 ( \8012 , RI2b5e785f3e50_220, \7726 );
and \U$6158 ( \8013 , RI2b5e785eb228_233, \7728 );
and \U$6159 ( \8014 , RI2b5e785da3b0_246, \7730 );
or \U$6160 ( \8015 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 );
_DC r10f9 ( \8016_nR10f9 , \8015 , \7740 );
buf \U$6161 ( \8017 , \8016_nR10f9 );
and \U$6162 ( \8018 , \7997 , \8017 );
buf \U$6163 ( \8019 , RI2b5e785db148_13);
buf \U$6166 ( \8020 , \8019 );
not \U$6167 ( \8021 , \8020 );
and \U$6168 ( \8022 , RI2b5e78549630_39, \7698 );
and \U$6169 ( \8023 , RI2b5e78538998_52, \7700 );
and \U$6170 ( \8024 , RI2b5e78538380_65, \7702 );
and \U$6171 ( \8025 , RI2b5e784a5e08_78, \7704 );
and \U$6172 ( \8026 , RI2b5e78495170_91, \7706 );
and \U$6173 ( \8027 , RI2b5e78403c70_104, \7708 );
and \U$6174 ( \8028 , RI2b5e775b1f50_117, \7710 );
and \U$6175 ( \8029 , RI2b5e775b1938_130, \7712 );
and \U$6176 ( \8030 , RI2b5e7750b8d0_143, \7714 );
and \U$6177 ( \8031 , RI2b5e774ff0a8_156, \7716 );
and \U$6178 ( \8032 , RI2b5e774f60c0_169, \7718 );
and \U$6179 ( \8033 , RI2b5e774ea6a8_182, \7720 );
and \U$6180 ( \8034 , RI2b5e774dde80_195, \7722 );
and \U$6181 ( \8035 , RI2b5e774d4e98_208, \7724 );
and \U$6182 ( \8036 , RI2b5e785f3dd8_221, \7726 );
and \U$6183 ( \8037 , RI2b5e785eb1b0_234, \7728 );
and \U$6184 ( \8038 , RI2b5e785da338_247, \7730 );
or \U$6185 ( \8039 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 );
_DC r1113 ( \8040_nR1113 , \8039 , \7740 );
buf \U$6186 ( \8041 , \8040_nR1113 );
and \U$6187 ( \8042 , \8021 , \8041 );
xnor \U$6188 ( \8043 , \7996 , \8017 );
and \U$6189 ( \8044 , \8042 , \8043 );
or \U$6190 ( \8045 , \8018 , \8044 );
xnor \U$6191 ( \8046 , \7971 , \7992 );
and \U$6192 ( \8047 , \8045 , \8046 );
or \U$6193 ( \8048 , \7993 , \8047 );
xnor \U$6194 ( \8049 , \7946 , \7967 );
and \U$6195 ( \8050 , \8048 , \8049 );
or \U$6196 ( \8051 , \7968 , \8050 );
xnor \U$6197 ( \8052 , \7921 , \7942 );
and \U$6198 ( \8053 , \8051 , \8052 );
or \U$6199 ( \8054 , \7943 , \8053 );
xnor \U$6200 ( \8055 , \7896 , \7917 );
and \U$6201 ( \8056 , \8054 , \8055 );
or \U$6202 ( \8057 , \7918 , \8056 );
xnor \U$6203 ( \8058 , \7871 , \7892 );
and \U$6204 ( \8059 , \8057 , \8058 );
or \U$6205 ( \8060 , \7893 , \8059 );
xnor \U$6206 ( \8061 , \7846 , \7867 );
and \U$6207 ( \8062 , \8060 , \8061 );
or \U$6208 ( \8063 , \7868 , \8062 );
xnor \U$6209 ( \8064 , \7821 , \7842 );
and \U$6210 ( \8065 , \8063 , \8064 );
or \U$6211 ( \8066 , \7843 , \8065 );
xnor \U$6212 ( \8067 , \7796 , \7817 );
and \U$6213 ( \8068 , \8066 , \8067 );
or \U$6214 ( \8069 , \7818 , \8068 );
xnor \U$6215 ( \8070 , \7771 , \7792 );
and \U$6216 ( \8071 , \8069 , \8070 );
or \U$6217 ( \8072 , \7793 , \8071 );
xnor \U$6218 ( \8073 , \7746 , \7767 );
and \U$6219 ( \8074 , \8072 , \8073 );
or \U$6220 ( \8075 , \7768 , \8074 );
xnor \U$6221 ( \8076 , \7696 , \7742 );
and \U$6222 ( \8077 , \8075 , \8076 );
or \U$6223 ( \8078 , \7743 , \8077 );
not \U$6224 ( \8079 , \8078 );
buf \U$6225 ( \8080 , \8079 );
buf \U$6226 ( \8081 , RI2b5e785aeb98_596);
buf \U$6227 ( \8082 , RI2b5e785aec10_595);
buf \U$6228 ( \8083 , RI2b5e785aec88_594);
buf \U$6229 ( \8084 , RI2b5e785aed00_593);
buf \U$6230 ( \8085 , RI2b5e785aed78_592);
buf \U$6231 ( \8086 , RI2b5e785aedf0_591);
buf \U$6232 ( \8087 , RI2b5e785aee68_590);
buf \U$6233 ( \8088 , RI2b5e785aeee0_589);
buf \U$6234 ( \8089 , RI2b5e785aef58_588);
buf \U$6235 ( \8090 , RI2b5e785ae9b8_600);
buf \U$6236 ( \8091 , RI2b5e785aea30_599);
buf \U$6237 ( \8092 , RI2b5e785aeaa8_598);
buf \U$6238 ( \8093 , RI2b5e785aeb20_597);
and \U$6239 ( \8094 , \8090 , \8091 , \8092 , \8093 );
nor \U$6240 ( \8095 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8094 );
buf \U$6241 ( \8096 , \8095 );
and \U$6242 ( \8097 , \8080 , \8096 );
nor \U$6243 ( \8098 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$6244 ( \8099 , RI2b5e785daab8_27, \8098 );
and \U$6245 ( \8100 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$6246 ( \8101 , RI2b5e785495b8_40, \8100 );
and \U$6247 ( \8102 , \2177 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$6248 ( \8103 , RI2b5e78538920_53, \8102 );
and \U$6249 ( \8104 , RI2b5e785ae9b8_600, \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$6250 ( \8105 , RI2b5e784a63a8_66, \8104 );
and \U$6251 ( \8106 , \2177 , \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, \2172 );
and \U$6252 ( \8107 , RI2b5e78495710_79, \8106 );
and \U$6253 ( \8108 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, \2172 );
and \U$6254 ( \8109 , RI2b5e784950f8_92, \8108 );
and \U$6255 ( \8110 , \2177 , RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, \2172 );
and \U$6256 ( \8111 , RI2b5e78403bf8_105, \8110 );
and \U$6257 ( \8112 , RI2b5e785ae9b8_600, \2180 , \2185 , RI2b5e785aeb20_597, \2172 );
and \U$6258 ( \8113 , RI2b5e775b1ed8_118, \8112 );
and \U$6259 ( \8114 , \2177 , \2180 , \2185 , RI2b5e785aeb20_597, \2172 );
and \U$6260 ( \8115 , RI2b5e775b18c0_131, \8114 );
nor \U$6261 ( \8116 , \2177 , \2180 , \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6262 ( \8117 , RI2b5e7750b858_144, \8116 );
nor \U$6263 ( \8118 , RI2b5e785ae9b8_600, \2180 , \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6264 ( \8119 , RI2b5e774ff030_157, \8118 );
nor \U$6265 ( \8120 , \2177 , RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6266 ( \8121 , RI2b5e774f6048_170, \8120 );
nor \U$6267 ( \8122 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, \2185 , RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6268 ( \8123 , RI2b5e774ea630_183, \8122 );
nor \U$6269 ( \8124 , \2177 , \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6270 ( \8125 , RI2b5e774dde08_196, \8124 );
nor \U$6271 ( \8126 , RI2b5e785ae9b8_600, \2180 , RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6272 ( \8127 , RI2b5e774d4e20_209, \8126 );
nor \U$6273 ( \8128 , \2177 , RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6274 ( \8129 , RI2b5e785f3d60_222, \8128 );
nor \U$6275 ( \8130 , RI2b5e785ae9b8_600, RI2b5e785aea30_599, RI2b5e785aeaa8_598, RI2b5e785aeb20_597, RI2b5e785aeb98_596);
and \U$6276 ( \8131 , RI2b5e785eb138_235, \8130 );
or \U$6277 ( \8132 , \8099 , \8101 , \8103 , \8105 , \8107 , \8109 , \8111 , \8113 , \8115 , \8117 , \8119 , \8121 , \8123 , \8125 , \8127 , \8129 , \8131 );
buf \U$6278 ( \8133 , RI2b5e785aeb98_596);
buf \U$6279 ( \8134 , RI2b5e785ae9b8_600);
buf \U$6280 ( \8135 , RI2b5e785aea30_599);
buf \U$6281 ( \8136 , RI2b5e785aeaa8_598);
buf \U$6282 ( \8137 , RI2b5e785aeb20_597);
or \U$6283 ( \8138 , \8134 , \8135 , \8136 , \8137 );
and \U$6284 ( \8139 , \8133 , \8138 );
buf \U$6285 ( \8140 , \8139 );
_DC r117c ( \8141_nR117c , \8132 , \8140 );
buf \U$6286 ( \8142 , \8141_nR117c );
not \U$6287 ( \8143 , \8142 );
nor \U$6288 ( \8144 , \4917 , \4921 , \4925 , \4929 , \4934 );
and \U$6289 ( \8145 , RI2b5e785daab8_27, \8144 );
and \U$6290 ( \8146 , \4917 , \4921 , \4925 , \4929 , \4934 );
and \U$6291 ( \8147 , RI2b5e785495b8_40, \8146 );
and \U$6292 ( \8148 , \4939 , \4921 , \4925 , \4929 , \4934 );
and \U$6293 ( \8149 , RI2b5e78538920_53, \8148 );
and \U$6294 ( \8150 , \4917 , \4942 , \4925 , \4929 , \4934 );
and \U$6295 ( \8151 , RI2b5e784a63a8_66, \8150 );
and \U$6296 ( \8152 , \4939 , \4942 , \4925 , \4929 , \4934 );
and \U$6297 ( \8153 , RI2b5e78495710_79, \8152 );
and \U$6298 ( \8154 , \4917 , \4921 , \4947 , \4929 , \4934 );
and \U$6299 ( \8155 , RI2b5e784950f8_92, \8154 );
and \U$6300 ( \8156 , \4939 , \4921 , \4947 , \4929 , \4934 );
and \U$6301 ( \8157 , RI2b5e78403bf8_105, \8156 );
and \U$6302 ( \8158 , \4917 , \4942 , \4947 , \4929 , \4934 );
and \U$6303 ( \8159 , RI2b5e775b1ed8_118, \8158 );
and \U$6304 ( \8160 , \4939 , \4942 , \4947 , \4929 , \4934 );
and \U$6305 ( \8161 , RI2b5e775b18c0_131, \8160 );
nor \U$6306 ( \8162 , \4939 , \4942 , \4947 , \4929 , \4933 );
and \U$6307 ( \8163 , RI2b5e7750b858_144, \8162 );
nor \U$6308 ( \8164 , \4917 , \4942 , \4947 , \4929 , \4933 );
and \U$6309 ( \8165 , RI2b5e774ff030_157, \8164 );
nor \U$6310 ( \8166 , \4939 , \4921 , \4947 , \4929 , \4933 );
and \U$6311 ( \8167 , RI2b5e774f6048_170, \8166 );
nor \U$6312 ( \8168 , \4917 , \4921 , \4947 , \4929 , \4933 );
and \U$6313 ( \8169 , RI2b5e774ea630_183, \8168 );
nor \U$6314 ( \8170 , \4939 , \4942 , \4925 , \4929 , \4933 );
and \U$6315 ( \8171 , RI2b5e774dde08_196, \8170 );
nor \U$6316 ( \8172 , \4917 , \4942 , \4925 , \4929 , \4933 );
and \U$6317 ( \8173 , RI2b5e774d4e20_209, \8172 );
nor \U$6318 ( \8174 , \4939 , \4921 , \4925 , \4929 , \4933 );
and \U$6319 ( \8175 , RI2b5e785f3d60_222, \8174 );
nor \U$6320 ( \8176 , \4917 , \4921 , \4925 , \4929 , \4933 );
and \U$6321 ( \8177 , RI2b5e785eb138_235, \8176 );
or \U$6322 ( \8178 , \8145 , \8147 , \8149 , \8151 , \8153 , \8155 , \8157 , \8159 , \8161 , \8163 , \8165 , \8167 , \8169 , \8171 , \8173 , \8175 , \8177 );
buf \U$6323 ( \8179 , \4933 );
buf \U$6324 ( \8180 , \4917 );
buf \U$6325 ( \8181 , \4921 );
buf \U$6326 ( \8182 , \4925 );
buf \U$6327 ( \8183 , \4929 );
or \U$6328 ( \8184 , \8180 , \8181 , \8182 , \8183 );
and \U$6329 ( \8185 , \8179 , \8184 );
buf \U$6330 ( \8186 , \8185 );
_DC r11aa ( \8187_nR11aa , \8178 , \8186 );
buf \U$6331 ( \8188 , \8187_nR11aa );
and \U$6332 ( \8189 , \8143 , \8188 );
and \U$6333 ( \8190 , RI2b5e785daa40_28, \8098 );
and \U$6334 ( \8191 , RI2b5e78549540_41, \8100 );
and \U$6335 ( \8192 , RI2b5e785388a8_54, \8102 );
and \U$6336 ( \8193 , RI2b5e784a6330_67, \8104 );
and \U$6337 ( \8194 , RI2b5e78495698_80, \8106 );
and \U$6338 ( \8195 , RI2b5e78495080_93, \8108 );
and \U$6339 ( \8196 , RI2b5e78403b80_106, \8110 );
and \U$6340 ( \8197 , RI2b5e775b1e60_119, \8112 );
and \U$6341 ( \8198 , RI2b5e7750bdf8_132, \8114 );
and \U$6342 ( \8199 , RI2b5e774ff5d0_145, \8116 );
and \U$6343 ( \8200 , RI2b5e774f65e8_158, \8118 );
and \U$6344 ( \8201 , RI2b5e774eabd0_171, \8120 );
and \U$6345 ( \8202 , RI2b5e774de3a8_184, \8122 );
and \U$6346 ( \8203 , RI2b5e774d53c0_197, \8124 );
and \U$6347 ( \8204 , RI2b5e785f4300_210, \8126 );
and \U$6348 ( \8205 , RI2b5e785f3ce8_223, \8128 );
and \U$6349 ( \8206 , RI2b5e785eb0c0_236, \8130 );
or \U$6350 ( \8207 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 );
_DC r11bf ( \8208_nR11bf , \8207 , \8140 );
buf \U$6351 ( \8209 , \8208_nR11bf );
not \U$6352 ( \8210 , \8209 );
and \U$6353 ( \8211 , RI2b5e785daa40_28, \8144 );
and \U$6354 ( \8212 , RI2b5e78549540_41, \8146 );
and \U$6355 ( \8213 , RI2b5e785388a8_54, \8148 );
and \U$6356 ( \8214 , RI2b5e784a6330_67, \8150 );
and \U$6357 ( \8215 , RI2b5e78495698_80, \8152 );
and \U$6358 ( \8216 , RI2b5e78495080_93, \8154 );
and \U$6359 ( \8217 , RI2b5e78403b80_106, \8156 );
and \U$6360 ( \8218 , RI2b5e775b1e60_119, \8158 );
and \U$6361 ( \8219 , RI2b5e7750bdf8_132, \8160 );
and \U$6362 ( \8220 , RI2b5e774ff5d0_145, \8162 );
and \U$6363 ( \8221 , RI2b5e774f65e8_158, \8164 );
and \U$6364 ( \8222 , RI2b5e774eabd0_171, \8166 );
and \U$6365 ( \8223 , RI2b5e774de3a8_184, \8168 );
and \U$6366 ( \8224 , RI2b5e774d53c0_197, \8170 );
and \U$6367 ( \8225 , RI2b5e785f4300_210, \8172 );
and \U$6368 ( \8226 , RI2b5e785f3ce8_223, \8174 );
and \U$6369 ( \8227 , RI2b5e785eb0c0_236, \8176 );
or \U$6370 ( \8228 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 );
_DC r11d4 ( \8229_nR11d4 , \8228 , \8186 );
buf \U$6371 ( \8230 , \8229_nR11d4 );
and \U$6372 ( \8231 , \8210 , \8230 );
and \U$6373 ( \8232 , RI2b5e785da9c8_29, \8098 );
and \U$6374 ( \8233 , RI2b5e785494c8_42, \8100 );
and \U$6375 ( \8234 , RI2b5e78538830_55, \8102 );
and \U$6376 ( \8235 , RI2b5e784a62b8_68, \8104 );
and \U$6377 ( \8236 , RI2b5e78495620_81, \8106 );
and \U$6378 ( \8237 , RI2b5e78495008_94, \8108 );
and \U$6379 ( \8238 , RI2b5e78403b08_107, \8110 );
and \U$6380 ( \8239 , RI2b5e775b1de8_120, \8112 );
and \U$6381 ( \8240 , RI2b5e7750bd80_133, \8114 );
and \U$6382 ( \8241 , RI2b5e774ff558_146, \8116 );
and \U$6383 ( \8242 , RI2b5e774f6570_159, \8118 );
and \U$6384 ( \8243 , RI2b5e774eab58_172, \8120 );
and \U$6385 ( \8244 , RI2b5e774de330_185, \8122 );
and \U$6386 ( \8245 , RI2b5e774d5348_198, \8124 );
and \U$6387 ( \8246 , RI2b5e785f4288_211, \8126 );
and \U$6388 ( \8247 , RI2b5e785f3658_224, \8128 );
and \U$6389 ( \8248 , RI2b5e785eb048_237, \8130 );
or \U$6390 ( \8249 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 );
_DC r11e9 ( \8250_nR11e9 , \8249 , \8140 );
buf \U$6391 ( \8251 , \8250_nR11e9 );
not \U$6392 ( \8252 , \8251 );
and \U$6393 ( \8253 , RI2b5e785da9c8_29, \8144 );
and \U$6394 ( \8254 , RI2b5e785494c8_42, \8146 );
and \U$6395 ( \8255 , RI2b5e78538830_55, \8148 );
and \U$6396 ( \8256 , RI2b5e784a62b8_68, \8150 );
and \U$6397 ( \8257 , RI2b5e78495620_81, \8152 );
and \U$6398 ( \8258 , RI2b5e78495008_94, \8154 );
and \U$6399 ( \8259 , RI2b5e78403b08_107, \8156 );
and \U$6400 ( \8260 , RI2b5e775b1de8_120, \8158 );
and \U$6401 ( \8261 , RI2b5e7750bd80_133, \8160 );
and \U$6402 ( \8262 , RI2b5e774ff558_146, \8162 );
and \U$6403 ( \8263 , RI2b5e774f6570_159, \8164 );
and \U$6404 ( \8264 , RI2b5e774eab58_172, \8166 );
and \U$6405 ( \8265 , RI2b5e774de330_185, \8168 );
and \U$6406 ( \8266 , RI2b5e774d5348_198, \8170 );
and \U$6407 ( \8267 , RI2b5e785f4288_211, \8172 );
and \U$6408 ( \8268 , RI2b5e785f3658_224, \8174 );
and \U$6409 ( \8269 , RI2b5e785eb048_237, \8176 );
or \U$6410 ( \8270 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 );
_DC r11fe ( \8271_nR11fe , \8270 , \8186 );
buf \U$6411 ( \8272 , \8271_nR11fe );
and \U$6412 ( \8273 , \8252 , \8272 );
and \U$6413 ( \8274 , RI2b5e785da950_30, \8098 );
and \U$6414 ( \8275 , RI2b5e78549450_43, \8100 );
and \U$6415 ( \8276 , RI2b5e785387b8_56, \8102 );
and \U$6416 ( \8277 , RI2b5e784a6240_69, \8104 );
and \U$6417 ( \8278 , RI2b5e784955a8_82, \8106 );
and \U$6418 ( \8279 , RI2b5e78494f90_95, \8108 );
and \U$6419 ( \8280 , RI2b5e78403a90_108, \8110 );
and \U$6420 ( \8281 , RI2b5e775b1d70_121, \8112 );
and \U$6421 ( \8282 , RI2b5e7750bd08_134, \8114 );
and \U$6422 ( \8283 , RI2b5e774ff4e0_147, \8116 );
and \U$6423 ( \8284 , RI2b5e774f64f8_160, \8118 );
and \U$6424 ( \8285 , RI2b5e774eaae0_173, \8120 );
and \U$6425 ( \8286 , RI2b5e774de2b8_186, \8122 );
and \U$6426 ( \8287 , RI2b5e774d52d0_199, \8124 );
and \U$6427 ( \8288 , RI2b5e785f4210_212, \8126 );
and \U$6428 ( \8289 , RI2b5e785eb5e8_225, \8128 );
and \U$6429 ( \8290 , RI2b5e785e6c50_238, \8130 );
or \U$6430 ( \8291 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 );
_DC r1213 ( \8292_nR1213 , \8291 , \8140 );
buf \U$6431 ( \8293 , \8292_nR1213 );
not \U$6432 ( \8294 , \8293 );
and \U$6433 ( \8295 , RI2b5e785da950_30, \8144 );
and \U$6434 ( \8296 , RI2b5e78549450_43, \8146 );
and \U$6435 ( \8297 , RI2b5e785387b8_56, \8148 );
and \U$6436 ( \8298 , RI2b5e784a6240_69, \8150 );
and \U$6437 ( \8299 , RI2b5e784955a8_82, \8152 );
and \U$6438 ( \8300 , RI2b5e78494f90_95, \8154 );
and \U$6439 ( \8301 , RI2b5e78403a90_108, \8156 );
and \U$6440 ( \8302 , RI2b5e775b1d70_121, \8158 );
and \U$6441 ( \8303 , RI2b5e7750bd08_134, \8160 );
and \U$6442 ( \8304 , RI2b5e774ff4e0_147, \8162 );
and \U$6443 ( \8305 , RI2b5e774f64f8_160, \8164 );
and \U$6444 ( \8306 , RI2b5e774eaae0_173, \8166 );
and \U$6445 ( \8307 , RI2b5e774de2b8_186, \8168 );
and \U$6446 ( \8308 , RI2b5e774d52d0_199, \8170 );
and \U$6447 ( \8309 , RI2b5e785f4210_212, \8172 );
and \U$6448 ( \8310 , RI2b5e785eb5e8_225, \8174 );
and \U$6449 ( \8311 , RI2b5e785e6c50_238, \8176 );
or \U$6450 ( \8312 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 );
_DC r1228 ( \8313_nR1228 , \8312 , \8186 );
buf \U$6451 ( \8314 , \8313_nR1228 );
and \U$6452 ( \8315 , \8294 , \8314 );
and \U$6453 ( \8316 , RI2b5e785da8d8_31, \8098 );
and \U$6454 ( \8317 , RI2b5e785493d8_44, \8100 );
and \U$6455 ( \8318 , RI2b5e78538740_57, \8102 );
and \U$6456 ( \8319 , RI2b5e784a61c8_70, \8104 );
and \U$6457 ( \8320 , RI2b5e78495530_83, \8106 );
and \U$6458 ( \8321 , RI2b5e78494f18_96, \8108 );
and \U$6459 ( \8322 , RI2b5e78403a18_109, \8110 );
and \U$6460 ( \8323 , RI2b5e775b1cf8_122, \8112 );
and \U$6461 ( \8324 , RI2b5e7750bc90_135, \8114 );
and \U$6462 ( \8325 , RI2b5e774ff468_148, \8116 );
and \U$6463 ( \8326 , RI2b5e774f6480_161, \8118 );
and \U$6464 ( \8327 , RI2b5e774eaa68_174, \8120 );
and \U$6465 ( \8328 , RI2b5e774de240_187, \8122 );
and \U$6466 ( \8329 , RI2b5e774d5258_200, \8124 );
and \U$6467 ( \8330 , RI2b5e785f4198_213, \8126 );
and \U$6468 ( \8331 , RI2b5e785eb570_226, \8128 );
and \U$6469 ( \8332 , RI2b5e785e6bd8_239, \8130 );
or \U$6470 ( \8333 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 );
_DC r123d ( \8334_nR123d , \8333 , \8140 );
buf \U$6471 ( \8335 , \8334_nR123d );
not \U$6472 ( \8336 , \8335 );
and \U$6473 ( \8337 , RI2b5e785da8d8_31, \8144 );
and \U$6474 ( \8338 , RI2b5e785493d8_44, \8146 );
and \U$6475 ( \8339 , RI2b5e78538740_57, \8148 );
and \U$6476 ( \8340 , RI2b5e784a61c8_70, \8150 );
and \U$6477 ( \8341 , RI2b5e78495530_83, \8152 );
and \U$6478 ( \8342 , RI2b5e78494f18_96, \8154 );
and \U$6479 ( \8343 , RI2b5e78403a18_109, \8156 );
and \U$6480 ( \8344 , RI2b5e775b1cf8_122, \8158 );
and \U$6481 ( \8345 , RI2b5e7750bc90_135, \8160 );
and \U$6482 ( \8346 , RI2b5e774ff468_148, \8162 );
and \U$6483 ( \8347 , RI2b5e774f6480_161, \8164 );
and \U$6484 ( \8348 , RI2b5e774eaa68_174, \8166 );
and \U$6485 ( \8349 , RI2b5e774de240_187, \8168 );
and \U$6486 ( \8350 , RI2b5e774d5258_200, \8170 );
and \U$6487 ( \8351 , RI2b5e785f4198_213, \8172 );
and \U$6488 ( \8352 , RI2b5e785eb570_226, \8174 );
and \U$6489 ( \8353 , RI2b5e785e6bd8_239, \8176 );
or \U$6490 ( \8354 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 );
_DC r1252 ( \8355_nR1252 , \8354 , \8186 );
buf \U$6491 ( \8356 , \8355_nR1252 );
and \U$6492 ( \8357 , \8336 , \8356 );
and \U$6493 ( \8358 , RI2b5e785da860_32, \8098 );
and \U$6494 ( \8359 , RI2b5e78549360_45, \8100 );
and \U$6495 ( \8360 , RI2b5e785386c8_58, \8102 );
and \U$6496 ( \8361 , RI2b5e784a6150_71, \8104 );
and \U$6497 ( \8362 , RI2b5e784954b8_84, \8106 );
and \U$6498 ( \8363 , RI2b5e78494ea0_97, \8108 );
and \U$6499 ( \8364 , RI2b5e784039a0_110, \8110 );
and \U$6500 ( \8365 , RI2b5e775b1c80_123, \8112 );
and \U$6501 ( \8366 , RI2b5e7750bc18_136, \8114 );
and \U$6502 ( \8367 , RI2b5e774ff3f0_149, \8116 );
and \U$6503 ( \8368 , RI2b5e774f6408_162, \8118 );
and \U$6504 ( \8369 , RI2b5e774ea9f0_175, \8120 );
and \U$6505 ( \8370 , RI2b5e774de1c8_188, \8122 );
and \U$6506 ( \8371 , RI2b5e774d51e0_201, \8124 );
and \U$6507 ( \8372 , RI2b5e785f4120_214, \8126 );
and \U$6508 ( \8373 , RI2b5e785eb4f8_227, \8128 );
and \U$6509 ( \8374 , RI2b5e785e64d0_240, \8130 );
or \U$6510 ( \8375 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 );
_DC r1267 ( \8376_nR1267 , \8375 , \8140 );
buf \U$6511 ( \8377 , \8376_nR1267 );
not \U$6512 ( \8378 , \8377 );
and \U$6513 ( \8379 , RI2b5e785da860_32, \8144 );
and \U$6514 ( \8380 , RI2b5e78549360_45, \8146 );
and \U$6515 ( \8381 , RI2b5e785386c8_58, \8148 );
and \U$6516 ( \8382 , RI2b5e784a6150_71, \8150 );
and \U$6517 ( \8383 , RI2b5e784954b8_84, \8152 );
and \U$6518 ( \8384 , RI2b5e78494ea0_97, \8154 );
and \U$6519 ( \8385 , RI2b5e784039a0_110, \8156 );
and \U$6520 ( \8386 , RI2b5e775b1c80_123, \8158 );
and \U$6521 ( \8387 , RI2b5e7750bc18_136, \8160 );
and \U$6522 ( \8388 , RI2b5e774ff3f0_149, \8162 );
and \U$6523 ( \8389 , RI2b5e774f6408_162, \8164 );
and \U$6524 ( \8390 , RI2b5e774ea9f0_175, \8166 );
and \U$6525 ( \8391 , RI2b5e774de1c8_188, \8168 );
and \U$6526 ( \8392 , RI2b5e774d51e0_201, \8170 );
and \U$6527 ( \8393 , RI2b5e785f4120_214, \8172 );
and \U$6528 ( \8394 , RI2b5e785eb4f8_227, \8174 );
and \U$6529 ( \8395 , RI2b5e785e64d0_240, \8176 );
or \U$6530 ( \8396 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 );
_DC r127c ( \8397_nR127c , \8396 , \8186 );
buf \U$6531 ( \8398 , \8397_nR127c );
and \U$6532 ( \8399 , \8378 , \8398 );
and \U$6533 ( \8400 , RI2b5e78549900_33, \8098 );
and \U$6534 ( \8401 , RI2b5e78538c68_46, \8100 );
and \U$6535 ( \8402 , RI2b5e78538650_59, \8102 );
and \U$6536 ( \8403 , RI2b5e784a60d8_72, \8104 );
and \U$6537 ( \8404 , RI2b5e78495440_85, \8106 );
and \U$6538 ( \8405 , RI2b5e78494e28_98, \8108 );
and \U$6539 ( \8406 , RI2b5e78403928_111, \8110 );
and \U$6540 ( \8407 , RI2b5e775b1c08_124, \8112 );
and \U$6541 ( \8408 , RI2b5e7750bba0_137, \8114 );
and \U$6542 ( \8409 , RI2b5e774ff378_150, \8116 );
and \U$6543 ( \8410 , RI2b5e774f6390_163, \8118 );
and \U$6544 ( \8411 , RI2b5e774ea978_176, \8120 );
and \U$6545 ( \8412 , RI2b5e774de150_189, \8122 );
and \U$6546 ( \8413 , RI2b5e774d5168_202, \8124 );
and \U$6547 ( \8414 , RI2b5e785f40a8_215, \8126 );
and \U$6548 ( \8415 , RI2b5e785eb480_228, \8128 );
and \U$6549 ( \8416 , RI2b5e785da608_241, \8130 );
or \U$6550 ( \8417 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 );
_DC r1291 ( \8418_nR1291 , \8417 , \8140 );
buf \U$6551 ( \8419 , \8418_nR1291 );
not \U$6552 ( \8420 , \8419 );
and \U$6553 ( \8421 , RI2b5e78549900_33, \8144 );
and \U$6554 ( \8422 , RI2b5e78538c68_46, \8146 );
and \U$6555 ( \8423 , RI2b5e78538650_59, \8148 );
and \U$6556 ( \8424 , RI2b5e784a60d8_72, \8150 );
and \U$6557 ( \8425 , RI2b5e78495440_85, \8152 );
and \U$6558 ( \8426 , RI2b5e78494e28_98, \8154 );
and \U$6559 ( \8427 , RI2b5e78403928_111, \8156 );
and \U$6560 ( \8428 , RI2b5e775b1c08_124, \8158 );
and \U$6561 ( \8429 , RI2b5e7750bba0_137, \8160 );
and \U$6562 ( \8430 , RI2b5e774ff378_150, \8162 );
and \U$6563 ( \8431 , RI2b5e774f6390_163, \8164 );
and \U$6564 ( \8432 , RI2b5e774ea978_176, \8166 );
and \U$6565 ( \8433 , RI2b5e774de150_189, \8168 );
and \U$6566 ( \8434 , RI2b5e774d5168_202, \8170 );
and \U$6567 ( \8435 , RI2b5e785f40a8_215, \8172 );
and \U$6568 ( \8436 , RI2b5e785eb480_228, \8174 );
and \U$6569 ( \8437 , RI2b5e785da608_241, \8176 );
or \U$6570 ( \8438 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 );
_DC r12a6 ( \8439_nR12a6 , \8438 , \8186 );
buf \U$6571 ( \8440 , \8439_nR12a6 );
and \U$6572 ( \8441 , \8420 , \8440 );
and \U$6573 ( \8442 , RI2b5e78549888_34, \8098 );
and \U$6574 ( \8443 , RI2b5e78538bf0_47, \8100 );
and \U$6575 ( \8444 , RI2b5e785385d8_60, \8102 );
and \U$6576 ( \8445 , RI2b5e784a6060_73, \8104 );
and \U$6577 ( \8446 , RI2b5e784953c8_86, \8106 );
and \U$6578 ( \8447 , RI2b5e78403ec8_99, \8108 );
and \U$6579 ( \8448 , RI2b5e775b21a8_112, \8110 );
and \U$6580 ( \8449 , RI2b5e775b1b90_125, \8112 );
and \U$6581 ( \8450 , RI2b5e7750bb28_138, \8114 );
and \U$6582 ( \8451 , RI2b5e774ff300_151, \8116 );
and \U$6583 ( \8452 , RI2b5e774f6318_164, \8118 );
and \U$6584 ( \8453 , RI2b5e774ea900_177, \8120 );
and \U$6585 ( \8454 , RI2b5e774de0d8_190, \8122 );
and \U$6586 ( \8455 , RI2b5e774d50f0_203, \8124 );
and \U$6587 ( \8456 , RI2b5e785f4030_216, \8126 );
and \U$6588 ( \8457 , RI2b5e785eb408_229, \8128 );
and \U$6589 ( \8458 , RI2b5e785da590_242, \8130 );
or \U$6590 ( \8459 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 );
_DC r12bb ( \8460_nR12bb , \8459 , \8140 );
buf \U$6591 ( \8461 , \8460_nR12bb );
not \U$6592 ( \8462 , \8461 );
and \U$6593 ( \8463 , RI2b5e78549888_34, \8144 );
and \U$6594 ( \8464 , RI2b5e78538bf0_47, \8146 );
and \U$6595 ( \8465 , RI2b5e785385d8_60, \8148 );
and \U$6596 ( \8466 , RI2b5e784a6060_73, \8150 );
and \U$6597 ( \8467 , RI2b5e784953c8_86, \8152 );
and \U$6598 ( \8468 , RI2b5e78403ec8_99, \8154 );
and \U$6599 ( \8469 , RI2b5e775b21a8_112, \8156 );
and \U$6600 ( \8470 , RI2b5e775b1b90_125, \8158 );
and \U$6601 ( \8471 , RI2b5e7750bb28_138, \8160 );
and \U$6602 ( \8472 , RI2b5e774ff300_151, \8162 );
and \U$6603 ( \8473 , RI2b5e774f6318_164, \8164 );
and \U$6604 ( \8474 , RI2b5e774ea900_177, \8166 );
and \U$6605 ( \8475 , RI2b5e774de0d8_190, \8168 );
and \U$6606 ( \8476 , RI2b5e774d50f0_203, \8170 );
and \U$6607 ( \8477 , RI2b5e785f4030_216, \8172 );
and \U$6608 ( \8478 , RI2b5e785eb408_229, \8174 );
and \U$6609 ( \8479 , RI2b5e785da590_242, \8176 );
or \U$6610 ( \8480 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 );
_DC r12d0 ( \8481_nR12d0 , \8480 , \8186 );
buf \U$6611 ( \8482 , \8481_nR12d0 );
and \U$6612 ( \8483 , \8462 , \8482 );
and \U$6613 ( \8484 , RI2b5e78549810_35, \8098 );
and \U$6614 ( \8485 , RI2b5e78538b78_48, \8100 );
and \U$6615 ( \8486 , RI2b5e78538560_61, \8102 );
and \U$6616 ( \8487 , RI2b5e784a5fe8_74, \8104 );
and \U$6617 ( \8488 , RI2b5e78495350_87, \8106 );
and \U$6618 ( \8489 , RI2b5e78403e50_100, \8108 );
and \U$6619 ( \8490 , RI2b5e775b2130_113, \8110 );
and \U$6620 ( \8491 , RI2b5e775b1b18_126, \8112 );
and \U$6621 ( \8492 , RI2b5e7750bab0_139, \8114 );
and \U$6622 ( \8493 , RI2b5e774ff288_152, \8116 );
and \U$6623 ( \8494 , RI2b5e774f62a0_165, \8118 );
and \U$6624 ( \8495 , RI2b5e774ea888_178, \8120 );
and \U$6625 ( \8496 , RI2b5e774de060_191, \8122 );
and \U$6626 ( \8497 , RI2b5e774d5078_204, \8124 );
and \U$6627 ( \8498 , RI2b5e785f3fb8_217, \8126 );
and \U$6628 ( \8499 , RI2b5e785eb390_230, \8128 );
and \U$6629 ( \8500 , RI2b5e785da518_243, \8130 );
or \U$6630 ( \8501 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 );
_DC r12e5 ( \8502_nR12e5 , \8501 , \8140 );
buf \U$6631 ( \8503 , \8502_nR12e5 );
not \U$6632 ( \8504 , \8503 );
and \U$6633 ( \8505 , RI2b5e78549810_35, \8144 );
and \U$6634 ( \8506 , RI2b5e78538b78_48, \8146 );
and \U$6635 ( \8507 , RI2b5e78538560_61, \8148 );
and \U$6636 ( \8508 , RI2b5e784a5fe8_74, \8150 );
and \U$6637 ( \8509 , RI2b5e78495350_87, \8152 );
and \U$6638 ( \8510 , RI2b5e78403e50_100, \8154 );
and \U$6639 ( \8511 , RI2b5e775b2130_113, \8156 );
and \U$6640 ( \8512 , RI2b5e775b1b18_126, \8158 );
and \U$6641 ( \8513 , RI2b5e7750bab0_139, \8160 );
and \U$6642 ( \8514 , RI2b5e774ff288_152, \8162 );
and \U$6643 ( \8515 , RI2b5e774f62a0_165, \8164 );
and \U$6644 ( \8516 , RI2b5e774ea888_178, \8166 );
and \U$6645 ( \8517 , RI2b5e774de060_191, \8168 );
and \U$6646 ( \8518 , RI2b5e774d5078_204, \8170 );
and \U$6647 ( \8519 , RI2b5e785f3fb8_217, \8172 );
and \U$6648 ( \8520 , RI2b5e785eb390_230, \8174 );
and \U$6649 ( \8521 , RI2b5e785da518_243, \8176 );
or \U$6650 ( \8522 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 );
_DC r12fa ( \8523_nR12fa , \8522 , \8186 );
buf \U$6651 ( \8524 , \8523_nR12fa );
and \U$6652 ( \8525 , \8504 , \8524 );
and \U$6653 ( \8526 , RI2b5e78549798_36, \8098 );
and \U$6654 ( \8527 , RI2b5e78538b00_49, \8100 );
and \U$6655 ( \8528 , RI2b5e785384e8_62, \8102 );
and \U$6656 ( \8529 , RI2b5e784a5f70_75, \8104 );
and \U$6657 ( \8530 , RI2b5e784952d8_88, \8106 );
and \U$6658 ( \8531 , RI2b5e78403dd8_101, \8108 );
and \U$6659 ( \8532 , RI2b5e775b20b8_114, \8110 );
and \U$6660 ( \8533 , RI2b5e775b1aa0_127, \8112 );
and \U$6661 ( \8534 , RI2b5e7750ba38_140, \8114 );
and \U$6662 ( \8535 , RI2b5e774ff210_153, \8116 );
and \U$6663 ( \8536 , RI2b5e774f6228_166, \8118 );
and \U$6664 ( \8537 , RI2b5e774ea810_179, \8120 );
and \U$6665 ( \8538 , RI2b5e774ddfe8_192, \8122 );
and \U$6666 ( \8539 , RI2b5e774d5000_205, \8124 );
and \U$6667 ( \8540 , RI2b5e785f3f40_218, \8126 );
and \U$6668 ( \8541 , RI2b5e785eb318_231, \8128 );
and \U$6669 ( \8542 , RI2b5e785da4a0_244, \8130 );
or \U$6670 ( \8543 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 );
_DC r130f ( \8544_nR130f , \8543 , \8140 );
buf \U$6671 ( \8545 , \8544_nR130f );
not \U$6672 ( \8546 , \8545 );
and \U$6673 ( \8547 , RI2b5e78549798_36, \8144 );
and \U$6674 ( \8548 , RI2b5e78538b00_49, \8146 );
and \U$6675 ( \8549 , RI2b5e785384e8_62, \8148 );
and \U$6676 ( \8550 , RI2b5e784a5f70_75, \8150 );
and \U$6677 ( \8551 , RI2b5e784952d8_88, \8152 );
and \U$6678 ( \8552 , RI2b5e78403dd8_101, \8154 );
and \U$6679 ( \8553 , RI2b5e775b20b8_114, \8156 );
and \U$6680 ( \8554 , RI2b5e775b1aa0_127, \8158 );
and \U$6681 ( \8555 , RI2b5e7750ba38_140, \8160 );
and \U$6682 ( \8556 , RI2b5e774ff210_153, \8162 );
and \U$6683 ( \8557 , RI2b5e774f6228_166, \8164 );
and \U$6684 ( \8558 , RI2b5e774ea810_179, \8166 );
and \U$6685 ( \8559 , RI2b5e774ddfe8_192, \8168 );
and \U$6686 ( \8560 , RI2b5e774d5000_205, \8170 );
and \U$6687 ( \8561 , RI2b5e785f3f40_218, \8172 );
and \U$6688 ( \8562 , RI2b5e785eb318_231, \8174 );
and \U$6689 ( \8563 , RI2b5e785da4a0_244, \8176 );
or \U$6690 ( \8564 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 );
_DC r1324 ( \8565_nR1324 , \8564 , \8186 );
buf \U$6691 ( \8566 , \8565_nR1324 );
and \U$6692 ( \8567 , \8546 , \8566 );
and \U$6693 ( \8568 , RI2b5e78549720_37, \8098 );
and \U$6694 ( \8569 , RI2b5e78538a88_50, \8100 );
and \U$6695 ( \8570 , RI2b5e78538470_63, \8102 );
and \U$6696 ( \8571 , RI2b5e784a5ef8_76, \8104 );
and \U$6697 ( \8572 , RI2b5e78495260_89, \8106 );
and \U$6698 ( \8573 , RI2b5e78403d60_102, \8108 );
and \U$6699 ( \8574 , RI2b5e775b2040_115, \8110 );
and \U$6700 ( \8575 , RI2b5e775b1a28_128, \8112 );
and \U$6701 ( \8576 , RI2b5e7750b9c0_141, \8114 );
and \U$6702 ( \8577 , RI2b5e774ff198_154, \8116 );
and \U$6703 ( \8578 , RI2b5e774f61b0_167, \8118 );
and \U$6704 ( \8579 , RI2b5e774ea798_180, \8120 );
and \U$6705 ( \8580 , RI2b5e774ddf70_193, \8122 );
and \U$6706 ( \8581 , RI2b5e774d4f88_206, \8124 );
and \U$6707 ( \8582 , RI2b5e785f3ec8_219, \8126 );
and \U$6708 ( \8583 , RI2b5e785eb2a0_232, \8128 );
and \U$6709 ( \8584 , RI2b5e785da428_245, \8130 );
or \U$6710 ( \8585 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 );
_DC r1339 ( \8586_nR1339 , \8585 , \8140 );
buf \U$6711 ( \8587 , \8586_nR1339 );
not \U$6712 ( \8588 , \8587 );
and \U$6713 ( \8589 , RI2b5e78549720_37, \8144 );
and \U$6714 ( \8590 , RI2b5e78538a88_50, \8146 );
and \U$6715 ( \8591 , RI2b5e78538470_63, \8148 );
and \U$6716 ( \8592 , RI2b5e784a5ef8_76, \8150 );
and \U$6717 ( \8593 , RI2b5e78495260_89, \8152 );
and \U$6718 ( \8594 , RI2b5e78403d60_102, \8154 );
and \U$6719 ( \8595 , RI2b5e775b2040_115, \8156 );
and \U$6720 ( \8596 , RI2b5e775b1a28_128, \8158 );
and \U$6721 ( \8597 , RI2b5e7750b9c0_141, \8160 );
and \U$6722 ( \8598 , RI2b5e774ff198_154, \8162 );
and \U$6723 ( \8599 , RI2b5e774f61b0_167, \8164 );
and \U$6724 ( \8600 , RI2b5e774ea798_180, \8166 );
and \U$6725 ( \8601 , RI2b5e774ddf70_193, \8168 );
and \U$6726 ( \8602 , RI2b5e774d4f88_206, \8170 );
and \U$6727 ( \8603 , RI2b5e785f3ec8_219, \8172 );
and \U$6728 ( \8604 , RI2b5e785eb2a0_232, \8174 );
and \U$6729 ( \8605 , RI2b5e785da428_245, \8176 );
or \U$6730 ( \8606 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 );
_DC r134e ( \8607_nR134e , \8606 , \8186 );
buf \U$6731 ( \8608 , \8607_nR134e );
and \U$6732 ( \8609 , \8588 , \8608 );
and \U$6733 ( \8610 , RI2b5e785496a8_38, \8098 );
and \U$6734 ( \8611 , RI2b5e78538a10_51, \8100 );
and \U$6735 ( \8612 , RI2b5e785383f8_64, \8102 );
and \U$6736 ( \8613 , RI2b5e784a5e80_77, \8104 );
and \U$6737 ( \8614 , RI2b5e784951e8_90, \8106 );
and \U$6738 ( \8615 , RI2b5e78403ce8_103, \8108 );
and \U$6739 ( \8616 , RI2b5e775b1fc8_116, \8110 );
and \U$6740 ( \8617 , RI2b5e775b19b0_129, \8112 );
and \U$6741 ( \8618 , RI2b5e7750b948_142, \8114 );
and \U$6742 ( \8619 , RI2b5e774ff120_155, \8116 );
and \U$6743 ( \8620 , RI2b5e774f6138_168, \8118 );
and \U$6744 ( \8621 , RI2b5e774ea720_181, \8120 );
and \U$6745 ( \8622 , RI2b5e774ddef8_194, \8122 );
and \U$6746 ( \8623 , RI2b5e774d4f10_207, \8124 );
and \U$6747 ( \8624 , RI2b5e785f3e50_220, \8126 );
and \U$6748 ( \8625 , RI2b5e785eb228_233, \8128 );
and \U$6749 ( \8626 , RI2b5e785da3b0_246, \8130 );
or \U$6750 ( \8627 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 );
_DC r1363 ( \8628_nR1363 , \8627 , \8140 );
buf \U$6751 ( \8629 , \8628_nR1363 );
not \U$6752 ( \8630 , \8629 );
and \U$6753 ( \8631 , RI2b5e785496a8_38, \8144 );
and \U$6754 ( \8632 , RI2b5e78538a10_51, \8146 );
and \U$6755 ( \8633 , RI2b5e785383f8_64, \8148 );
and \U$6756 ( \8634 , RI2b5e784a5e80_77, \8150 );
and \U$6757 ( \8635 , RI2b5e784951e8_90, \8152 );
and \U$6758 ( \8636 , RI2b5e78403ce8_103, \8154 );
and \U$6759 ( \8637 , RI2b5e775b1fc8_116, \8156 );
and \U$6760 ( \8638 , RI2b5e775b19b0_129, \8158 );
and \U$6761 ( \8639 , RI2b5e7750b948_142, \8160 );
and \U$6762 ( \8640 , RI2b5e774ff120_155, \8162 );
and \U$6763 ( \8641 , RI2b5e774f6138_168, \8164 );
and \U$6764 ( \8642 , RI2b5e774ea720_181, \8166 );
and \U$6765 ( \8643 , RI2b5e774ddef8_194, \8168 );
and \U$6766 ( \8644 , RI2b5e774d4f10_207, \8170 );
and \U$6767 ( \8645 , RI2b5e785f3e50_220, \8172 );
and \U$6768 ( \8646 , RI2b5e785eb228_233, \8174 );
and \U$6769 ( \8647 , RI2b5e785da3b0_246, \8176 );
or \U$6770 ( \8648 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 );
_DC r1378 ( \8649_nR1378 , \8648 , \8186 );
buf \U$6771 ( \8650 , \8649_nR1378 );
and \U$6772 ( \8651 , \8630 , \8650 );
and \U$6773 ( \8652 , RI2b5e78549630_39, \8098 );
and \U$6774 ( \8653 , RI2b5e78538998_52, \8100 );
and \U$6775 ( \8654 , RI2b5e78538380_65, \8102 );
and \U$6776 ( \8655 , RI2b5e784a5e08_78, \8104 );
and \U$6777 ( \8656 , RI2b5e78495170_91, \8106 );
and \U$6778 ( \8657 , RI2b5e78403c70_104, \8108 );
and \U$6779 ( \8658 , RI2b5e775b1f50_117, \8110 );
and \U$6780 ( \8659 , RI2b5e775b1938_130, \8112 );
and \U$6781 ( \8660 , RI2b5e7750b8d0_143, \8114 );
and \U$6782 ( \8661 , RI2b5e774ff0a8_156, \8116 );
and \U$6783 ( \8662 , RI2b5e774f60c0_169, \8118 );
and \U$6784 ( \8663 , RI2b5e774ea6a8_182, \8120 );
and \U$6785 ( \8664 , RI2b5e774dde80_195, \8122 );
and \U$6786 ( \8665 , RI2b5e774d4e98_208, \8124 );
and \U$6787 ( \8666 , RI2b5e785f3dd8_221, \8126 );
and \U$6788 ( \8667 , RI2b5e785eb1b0_234, \8128 );
and \U$6789 ( \8668 , RI2b5e785da338_247, \8130 );
or \U$6790 ( \8669 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 );
_DC r138d ( \8670_nR138d , \8669 , \8140 );
buf \U$6791 ( \8671 , \8670_nR138d );
not \U$6792 ( \8672 , \8671 );
and \U$6793 ( \8673 , RI2b5e78549630_39, \8144 );
and \U$6794 ( \8674 , RI2b5e78538998_52, \8146 );
and \U$6795 ( \8675 , RI2b5e78538380_65, \8148 );
and \U$6796 ( \8676 , RI2b5e784a5e08_78, \8150 );
and \U$6797 ( \8677 , RI2b5e78495170_91, \8152 );
and \U$6798 ( \8678 , RI2b5e78403c70_104, \8154 );
and \U$6799 ( \8679 , RI2b5e775b1f50_117, \8156 );
and \U$6800 ( \8680 , RI2b5e775b1938_130, \8158 );
and \U$6801 ( \8681 , RI2b5e7750b8d0_143, \8160 );
and \U$6802 ( \8682 , RI2b5e774ff0a8_156, \8162 );
and \U$6803 ( \8683 , RI2b5e774f60c0_169, \8164 );
and \U$6804 ( \8684 , RI2b5e774ea6a8_182, \8166 );
and \U$6805 ( \8685 , RI2b5e774dde80_195, \8168 );
and \U$6806 ( \8686 , RI2b5e774d4e98_208, \8170 );
and \U$6807 ( \8687 , RI2b5e785f3dd8_221, \8172 );
and \U$6808 ( \8688 , RI2b5e785eb1b0_234, \8174 );
and \U$6809 ( \8689 , RI2b5e785da338_247, \8176 );
or \U$6810 ( \8690 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 );
_DC r13a2 ( \8691_nR13a2 , \8690 , \8186 );
buf \U$6811 ( \8692 , \8691_nR13a2 );
and \U$6812 ( \8693 , \8672 , \8692 );
xnor \U$6813 ( \8694 , \8650 , \8629 );
and \U$6814 ( \8695 , \8693 , \8694 );
or \U$6815 ( \8696 , \8651 , \8695 );
xnor \U$6816 ( \8697 , \8608 , \8587 );
and \U$6817 ( \8698 , \8696 , \8697 );
or \U$6818 ( \8699 , \8609 , \8698 );
xnor \U$6819 ( \8700 , \8566 , \8545 );
and \U$6820 ( \8701 , \8699 , \8700 );
or \U$6821 ( \8702 , \8567 , \8701 );
xnor \U$6822 ( \8703 , \8524 , \8503 );
and \U$6823 ( \8704 , \8702 , \8703 );
or \U$6824 ( \8705 , \8525 , \8704 );
xnor \U$6825 ( \8706 , \8482 , \8461 );
and \U$6826 ( \8707 , \8705 , \8706 );
or \U$6827 ( \8708 , \8483 , \8707 );
xnor \U$6828 ( \8709 , \8440 , \8419 );
and \U$6829 ( \8710 , \8708 , \8709 );
or \U$6830 ( \8711 , \8441 , \8710 );
xnor \U$6831 ( \8712 , \8398 , \8377 );
and \U$6832 ( \8713 , \8711 , \8712 );
or \U$6833 ( \8714 , \8399 , \8713 );
xnor \U$6834 ( \8715 , \8356 , \8335 );
and \U$6835 ( \8716 , \8714 , \8715 );
or \U$6836 ( \8717 , \8357 , \8716 );
xnor \U$6837 ( \8718 , \8314 , \8293 );
and \U$6838 ( \8719 , \8717 , \8718 );
or \U$6839 ( \8720 , \8315 , \8719 );
xnor \U$6840 ( \8721 , \8272 , \8251 );
and \U$6841 ( \8722 , \8720 , \8721 );
or \U$6842 ( \8723 , \8273 , \8722 );
xnor \U$6843 ( \8724 , \8230 , \8209 );
and \U$6844 ( \8725 , \8723 , \8724 );
or \U$6845 ( \8726 , \8231 , \8725 );
xnor \U$6846 ( \8727 , \8188 , \8142 );
and \U$6847 ( \8728 , \8726 , \8727 );
or \U$6848 ( \8729 , \8189 , \8728 );
buf \U$6849 ( \8730 , \8729 );
and \U$6850 ( \8731 , \8097 , \8730 );
_HMUX r3163 ( \8732_nR3163 , \4874 , \7668 , \8731 );
buf \U$6851 ( \8733 , \8732_nR3163 );
not \U$6852 ( \8734 , \4337 );
nand \U$6853 ( \8735 , \4866 , \8734 );
nor \U$6854 ( \8736 , \4684 , \3520 );
nor \U$6855 ( \8737 , \3595 , \3672 );
nand \U$6856 ( \8738 , \8736 , \8737 );
nor \U$6857 ( \8739 , \3747 , \3824 );
nor \U$6858 ( \8740 , \3900 , \3973 );
nand \U$6859 ( \8741 , \8739 , \8740 );
nor \U$6860 ( \8742 , \8738 , \8741 );
nor \U$6861 ( \8743 , \4042 , \4106 );
nor \U$6862 ( \8744 , \4166 , \4223 );
nand \U$6863 ( \8745 , \8743 , \8744 );
nor \U$6864 ( \8746 , \4261 , \4293 );
nor \U$6865 ( \8747 , \4314 , \4330 );
nand \U$6866 ( \8748 , \8746 , \8747 );
nor \U$6867 ( \8749 , \8745 , \8748 );
nand \U$6868 ( \8750 , \8742 , \8749 );
nor \U$6869 ( \8751 , \4745 , \4449 );
nor \U$6870 ( \8752 , \4494 , \4546 );
nand \U$6871 ( \8753 , \8751 , \8752 );
nor \U$6872 ( \8754 , \4601 , \4640 );
nor \U$6873 ( \8755 , \4661 , \4677 );
nand \U$6874 ( \8756 , \8754 , \8755 );
nor \U$6875 ( \8757 , \8753 , \8756 );
nor \U$6876 ( \8758 , \4765 , \4720 );
nor \U$6877 ( \8759 , \4731 , \4742 );
nand \U$6878 ( \8760 , \8758 , \8759 );
nor \U$6879 ( \8761 , \4770 , \4762 );
not \U$6880 ( \8762 , \4778 );
and \U$6881 ( \8763 , \8761 , \8762 );
or \U$6882 ( \8764 , \4762 , \4780 );
nand \U$6883 ( \8765 , \8764 , \4783 );
nor \U$6884 ( \8766 , \8763 , \8765 );
or \U$6885 ( \8767 , \8760 , \8766 );
or \U$6886 ( \8768 , \4720 , \4785 );
nand \U$6887 ( \8769 , \8768 , \4789 );
and \U$6888 ( \8770 , \8759 , \8769 );
or \U$6889 ( \8771 , \4742 , \4791 );
nand \U$6890 ( \8772 , \8771 , \4794 );
nor \U$6891 ( \8773 , \8770 , \8772 );
nand \U$6892 ( \8774 , \8767 , \8773 );
and \U$6893 ( \8775 , \8757 , \8774 );
or \U$6894 ( \8776 , \4449 , \4796 );
nand \U$6895 ( \8777 , \8776 , \4801 );
and \U$6896 ( \8778 , \8752 , \8777 );
or \U$6897 ( \8779 , \4546 , \4803 );
nand \U$6898 ( \8780 , \8779 , \4806 );
nor \U$6899 ( \8781 , \8778 , \8780 );
or \U$6900 ( \8782 , \8756 , \8781 );
or \U$6901 ( \8783 , \4640 , \4808 );
nand \U$6902 ( \8784 , \8783 , \4812 );
and \U$6903 ( \8785 , \8755 , \8784 );
or \U$6904 ( \8786 , \4677 , \4814 );
nand \U$6905 ( \8787 , \8786 , \4817 );
nor \U$6906 ( \8788 , \8785 , \8787 );
nand \U$6907 ( \8789 , \8782 , \8788 );
nor \U$6908 ( \8790 , \8775 , \8789 );
or \U$6909 ( \8791 , \8750 , \8790 );
or \U$6910 ( \8792 , \3520 , \4819 );
nand \U$6911 ( \8793 , \8792 , \4825 );
and \U$6912 ( \8794 , \8737 , \8793 );
or \U$6913 ( \8795 , \3672 , \4827 );
nand \U$6914 ( \8796 , \8795 , \4830 );
nor \U$6915 ( \8797 , \8794 , \8796 );
or \U$6916 ( \8798 , \8741 , \8797 );
or \U$6917 ( \8799 , \3824 , \4832 );
nand \U$6918 ( \8800 , \8799 , \4836 );
and \U$6919 ( \8801 , \8740 , \8800 );
or \U$6920 ( \8802 , \3973 , \4838 );
nand \U$6921 ( \8803 , \8802 , \4841 );
nor \U$6922 ( \8804 , \8801 , \8803 );
nand \U$6923 ( \8805 , \8798 , \8804 );
and \U$6924 ( \8806 , \8749 , \8805 );
or \U$6925 ( \8807 , \4106 , \4843 );
nand \U$6926 ( \8808 , \8807 , \4848 );
and \U$6927 ( \8809 , \8744 , \8808 );
or \U$6928 ( \8810 , \4223 , \4850 );
nand \U$6929 ( \8811 , \8810 , \4853 );
nor \U$6930 ( \8812 , \8809 , \8811 );
or \U$6931 ( \8813 , \8748 , \8812 );
or \U$6932 ( \8814 , \4293 , \4855 );
nand \U$6933 ( \8815 , \8814 , \4859 );
and \U$6934 ( \8816 , \8747 , \8815 );
or \U$6935 ( \8817 , \4330 , \4861 );
nand \U$6936 ( \8818 , \8817 , \4864 );
nor \U$6937 ( \8819 , \8816 , \8818 );
nand \U$6938 ( \8820 , \8813 , \8819 );
nor \U$6939 ( \8821 , \8806 , \8820 );
nand \U$6940 ( \8822 , \8791 , \8821 );
not \U$6941 ( \8823 , \8822 );
xor \U$6942 ( \8824 , \8735 , \8823 );
buf \U$6943 ( \8825 , \8824 );
not \U$6944 ( \8826 , \7131 );
nand \U$6945 ( \8827 , \7660 , \8826 );
nor \U$6946 ( \8828 , \7478 , \6314 );
nor \U$6947 ( \8829 , \6389 , \6466 );
nand \U$6948 ( \8830 , \8828 , \8829 );
nor \U$6949 ( \8831 , \6541 , \6618 );
nor \U$6950 ( \8832 , \6694 , \6767 );
nand \U$6951 ( \8833 , \8831 , \8832 );
nor \U$6952 ( \8834 , \8830 , \8833 );
nor \U$6953 ( \8835 , \6836 , \6900 );
nor \U$6954 ( \8836 , \6960 , \7017 );
nand \U$6955 ( \8837 , \8835 , \8836 );
nor \U$6956 ( \8838 , \7055 , \7087 );
nor \U$6957 ( \8839 , \7108 , \7124 );
nand \U$6958 ( \8840 , \8838 , \8839 );
nor \U$6959 ( \8841 , \8837 , \8840 );
nand \U$6960 ( \8842 , \8834 , \8841 );
nor \U$6961 ( \8843 , \7539 , \7243 );
nor \U$6962 ( \8844 , \7288 , \7340 );
nand \U$6963 ( \8845 , \8843 , \8844 );
nor \U$6964 ( \8846 , \7395 , \7434 );
nor \U$6965 ( \8847 , \7455 , \7471 );
nand \U$6966 ( \8848 , \8846 , \8847 );
nor \U$6967 ( \8849 , \8845 , \8848 );
nor \U$6968 ( \8850 , \7559 , \7514 );
nor \U$6969 ( \8851 , \7525 , \7536 );
nand \U$6970 ( \8852 , \8850 , \8851 );
nor \U$6971 ( \8853 , \7564 , \7556 );
not \U$6972 ( \8854 , \7572 );
and \U$6973 ( \8855 , \8853 , \8854 );
or \U$6974 ( \8856 , \7556 , \7574 );
nand \U$6975 ( \8857 , \8856 , \7577 );
nor \U$6976 ( \8858 , \8855 , \8857 );
or \U$6977 ( \8859 , \8852 , \8858 );
or \U$6978 ( \8860 , \7514 , \7579 );
nand \U$6979 ( \8861 , \8860 , \7583 );
and \U$6980 ( \8862 , \8851 , \8861 );
or \U$6981 ( \8863 , \7536 , \7585 );
nand \U$6982 ( \8864 , \8863 , \7588 );
nor \U$6983 ( \8865 , \8862 , \8864 );
nand \U$6984 ( \8866 , \8859 , \8865 );
and \U$6985 ( \8867 , \8849 , \8866 );
or \U$6986 ( \8868 , \7243 , \7590 );
nand \U$6987 ( \8869 , \8868 , \7595 );
and \U$6988 ( \8870 , \8844 , \8869 );
or \U$6989 ( \8871 , \7340 , \7597 );
nand \U$6990 ( \8872 , \8871 , \7600 );
nor \U$6991 ( \8873 , \8870 , \8872 );
or \U$6992 ( \8874 , \8848 , \8873 );
or \U$6993 ( \8875 , \7434 , \7602 );
nand \U$6994 ( \8876 , \8875 , \7606 );
and \U$6995 ( \8877 , \8847 , \8876 );
or \U$6996 ( \8878 , \7471 , \7608 );
nand \U$6997 ( \8879 , \8878 , \7611 );
nor \U$6998 ( \8880 , \8877 , \8879 );
nand \U$6999 ( \8881 , \8874 , \8880 );
nor \U$7000 ( \8882 , \8867 , \8881 );
or \U$7001 ( \8883 , \8842 , \8882 );
or \U$7002 ( \8884 , \6314 , \7613 );
nand \U$7003 ( \8885 , \8884 , \7619 );
and \U$7004 ( \8886 , \8829 , \8885 );
or \U$7005 ( \8887 , \6466 , \7621 );
nand \U$7006 ( \8888 , \8887 , \7624 );
nor \U$7007 ( \8889 , \8886 , \8888 );
or \U$7008 ( \8890 , \8833 , \8889 );
or \U$7009 ( \8891 , \6618 , \7626 );
nand \U$7010 ( \8892 , \8891 , \7630 );
and \U$7011 ( \8893 , \8832 , \8892 );
or \U$7012 ( \8894 , \6767 , \7632 );
nand \U$7013 ( \8895 , \8894 , \7635 );
nor \U$7014 ( \8896 , \8893 , \8895 );
nand \U$7015 ( \8897 , \8890 , \8896 );
and \U$7016 ( \8898 , \8841 , \8897 );
or \U$7017 ( \8899 , \6900 , \7637 );
nand \U$7018 ( \8900 , \8899 , \7642 );
and \U$7019 ( \8901 , \8836 , \8900 );
or \U$7020 ( \8902 , \7017 , \7644 );
nand \U$7021 ( \8903 , \8902 , \7647 );
nor \U$7022 ( \8904 , \8901 , \8903 );
or \U$7023 ( \8905 , \8840 , \8904 );
or \U$7024 ( \8906 , \7087 , \7649 );
nand \U$7025 ( \8907 , \8906 , \7653 );
and \U$7026 ( \8908 , \8839 , \8907 );
or \U$7027 ( \8909 , \7124 , \7655 );
nand \U$7028 ( \8910 , \8909 , \7658 );
nor \U$7029 ( \8911 , \8908 , \8910 );
nand \U$7030 ( \8912 , \8905 , \8911 );
nor \U$7031 ( \8913 , \8898 , \8912 );
nand \U$7032 ( \8914 , \8883 , \8913 );
not \U$7033 ( \8915 , \8914 );
xor \U$7034 ( \8916 , \8827 , \8915 );
buf \U$7035 ( \8917 , \8916 );
_HMUX r3106 ( \8918_nR3106 , \8825 , \8917 , \8731 );
buf \U$7036 ( \8919 , \8918_nR3106 );
not \U$7037 ( \8920 , \4330 );
nand \U$7038 ( \8921 , \4864 , \8920 );
nand \U$7039 ( \8922 , \4685 , \3596 );
nand \U$7040 ( \8923 , \3748 , \3901 );
nor \U$7041 ( \8924 , \8922 , \8923 );
nand \U$7042 ( \8925 , \4043 , \4167 );
nand \U$7043 ( \8926 , \4262 , \4315 );
nor \U$7044 ( \8927 , \8925 , \8926 );
nand \U$7045 ( \8928 , \8924 , \8927 );
nand \U$7046 ( \8929 , \4746 , \4495 );
nand \U$7047 ( \8930 , \4602 , \4662 );
nor \U$7048 ( \8931 , \8929 , \8930 );
nand \U$7049 ( \8932 , \4766 , \4732 );
not \U$7050 ( \8933 , \4781 );
or \U$7051 ( \8934 , \8932 , \8933 );
and \U$7052 ( \8935 , \4732 , \4786 );
nor \U$7053 ( \8936 , \8935 , \4792 );
nand \U$7054 ( \8937 , \8934 , \8936 );
and \U$7055 ( \8938 , \8931 , \8937 );
and \U$7056 ( \8939 , \4495 , \4797 );
nor \U$7057 ( \8940 , \8939 , \4804 );
or \U$7058 ( \8941 , \8930 , \8940 );
and \U$7059 ( \8942 , \4662 , \4809 );
nor \U$7060 ( \8943 , \8942 , \4815 );
nand \U$7061 ( \8944 , \8941 , \8943 );
nor \U$7062 ( \8945 , \8938 , \8944 );
or \U$7063 ( \8946 , \8928 , \8945 );
and \U$7064 ( \8947 , \3596 , \4820 );
nor \U$7065 ( \8948 , \8947 , \4828 );
or \U$7066 ( \8949 , \8923 , \8948 );
and \U$7067 ( \8950 , \3901 , \4833 );
nor \U$7068 ( \8951 , \8950 , \4839 );
nand \U$7069 ( \8952 , \8949 , \8951 );
and \U$7070 ( \8953 , \8927 , \8952 );
and \U$7071 ( \8954 , \4167 , \4844 );
nor \U$7072 ( \8955 , \8954 , \4851 );
or \U$7073 ( \8956 , \8926 , \8955 );
and \U$7074 ( \8957 , \4315 , \4856 );
nor \U$7075 ( \8958 , \8957 , \4862 );
nand \U$7076 ( \8959 , \8956 , \8958 );
nor \U$7077 ( \8960 , \8953 , \8959 );
nand \U$7078 ( \8961 , \8946 , \8960 );
not \U$7079 ( \8962 , \8961 );
xor \U$7080 ( \8963 , \8921 , \8962 );
buf \U$7081 ( \8964 , \8963 );
not \U$7082 ( \8965 , \7124 );
nand \U$7083 ( \8966 , \7658 , \8965 );
nand \U$7084 ( \8967 , \7479 , \6390 );
nand \U$7085 ( \8968 , \6542 , \6695 );
nor \U$7086 ( \8969 , \8967 , \8968 );
nand \U$7087 ( \8970 , \6837 , \6961 );
nand \U$7088 ( \8971 , \7056 , \7109 );
nor \U$7089 ( \8972 , \8970 , \8971 );
nand \U$7090 ( \8973 , \8969 , \8972 );
nand \U$7091 ( \8974 , \7540 , \7289 );
nand \U$7092 ( \8975 , \7396 , \7456 );
nor \U$7093 ( \8976 , \8974 , \8975 );
nand \U$7094 ( \8977 , \7560 , \7526 );
not \U$7095 ( \8978 , \7575 );
or \U$7096 ( \8979 , \8977 , \8978 );
and \U$7097 ( \8980 , \7526 , \7580 );
nor \U$7098 ( \8981 , \8980 , \7586 );
nand \U$7099 ( \8982 , \8979 , \8981 );
and \U$7100 ( \8983 , \8976 , \8982 );
and \U$7101 ( \8984 , \7289 , \7591 );
nor \U$7102 ( \8985 , \8984 , \7598 );
or \U$7103 ( \8986 , \8975 , \8985 );
and \U$7104 ( \8987 , \7456 , \7603 );
nor \U$7105 ( \8988 , \8987 , \7609 );
nand \U$7106 ( \8989 , \8986 , \8988 );
nor \U$7107 ( \8990 , \8983 , \8989 );
or \U$7108 ( \8991 , \8973 , \8990 );
and \U$7109 ( \8992 , \6390 , \7614 );
nor \U$7110 ( \8993 , \8992 , \7622 );
or \U$7111 ( \8994 , \8968 , \8993 );
and \U$7112 ( \8995 , \6695 , \7627 );
nor \U$7113 ( \8996 , \8995 , \7633 );
nand \U$7114 ( \8997 , \8994 , \8996 );
and \U$7115 ( \8998 , \8972 , \8997 );
and \U$7116 ( \8999 , \6961 , \7638 );
nor \U$7117 ( \9000 , \8999 , \7645 );
or \U$7118 ( \9001 , \8971 , \9000 );
and \U$7119 ( \9002 , \7109 , \7650 );
nor \U$7120 ( \9003 , \9002 , \7656 );
nand \U$7121 ( \9004 , \9001 , \9003 );
nor \U$7122 ( \9005 , \8998 , \9004 );
nand \U$7123 ( \9006 , \8991 , \9005 );
not \U$7124 ( \9007 , \9006 );
xor \U$7125 ( \9008 , \8966 , \9007 );
buf \U$7126 ( \9009 , \9008 );
_HMUX r309d ( \9010_nR309d , \8964 , \9009 , \8731 );
buf \U$7127 ( \9011 , \9010_nR309d );
not \U$7128 ( \9012 , \4314 );
nand \U$7129 ( \9013 , \4861 , \9012 );
nand \U$7130 ( \9014 , \8755 , \8736 );
nand \U$7131 ( \9015 , \8737 , \8739 );
nor \U$7132 ( \9016 , \9014 , \9015 );
nand \U$7133 ( \9017 , \8740 , \8743 );
nand \U$7134 ( \9018 , \8744 , \8746 );
nor \U$7135 ( \9019 , \9017 , \9018 );
nand \U$7136 ( \9020 , \9016 , \9019 );
nand \U$7137 ( \9021 , \8759 , \8751 );
nand \U$7138 ( \9022 , \8752 , \8754 );
nor \U$7139 ( \9023 , \9021 , \9022 );
nand \U$7140 ( \9024 , \8761 , \8758 );
or \U$7141 ( \9025 , \9024 , \4778 );
and \U$7142 ( \9026 , \8758 , \8765 );
nor \U$7143 ( \9027 , \9026 , \8769 );
nand \U$7144 ( \9028 , \9025 , \9027 );
and \U$7145 ( \9029 , \9023 , \9028 );
and \U$7146 ( \9030 , \8751 , \8772 );
nor \U$7147 ( \9031 , \9030 , \8777 );
or \U$7148 ( \9032 , \9022 , \9031 );
and \U$7149 ( \9033 , \8754 , \8780 );
nor \U$7150 ( \9034 , \9033 , \8784 );
nand \U$7151 ( \9035 , \9032 , \9034 );
nor \U$7152 ( \9036 , \9029 , \9035 );
or \U$7153 ( \9037 , \9020 , \9036 );
and \U$7154 ( \9038 , \8736 , \8787 );
nor \U$7155 ( \9039 , \9038 , \8793 );
or \U$7156 ( \9040 , \9015 , \9039 );
and \U$7157 ( \9041 , \8739 , \8796 );
nor \U$7158 ( \9042 , \9041 , \8800 );
nand \U$7159 ( \9043 , \9040 , \9042 );
and \U$7160 ( \9044 , \9019 , \9043 );
and \U$7161 ( \9045 , \8743 , \8803 );
nor \U$7162 ( \9046 , \9045 , \8808 );
or \U$7163 ( \9047 , \9018 , \9046 );
and \U$7164 ( \9048 , \8746 , \8811 );
nor \U$7165 ( \9049 , \9048 , \8815 );
nand \U$7166 ( \9050 , \9047 , \9049 );
nor \U$7167 ( \9051 , \9044 , \9050 );
nand \U$7168 ( \9052 , \9037 , \9051 );
not \U$7169 ( \9053 , \9052 );
xor \U$7170 ( \9054 , \9013 , \9053 );
buf \U$7171 ( \9055 , \9054 );
not \U$7172 ( \9056 , \7108 );
nand \U$7173 ( \9057 , \7655 , \9056 );
nand \U$7174 ( \9058 , \8847 , \8828 );
nand \U$7175 ( \9059 , \8829 , \8831 );
nor \U$7176 ( \9060 , \9058 , \9059 );
nand \U$7177 ( \9061 , \8832 , \8835 );
nand \U$7178 ( \9062 , \8836 , \8838 );
nor \U$7179 ( \9063 , \9061 , \9062 );
nand \U$7180 ( \9064 , \9060 , \9063 );
nand \U$7181 ( \9065 , \8851 , \8843 );
nand \U$7182 ( \9066 , \8844 , \8846 );
nor \U$7183 ( \9067 , \9065 , \9066 );
nand \U$7184 ( \9068 , \8853 , \8850 );
or \U$7185 ( \9069 , \9068 , \7572 );
and \U$7186 ( \9070 , \8850 , \8857 );
nor \U$7187 ( \9071 , \9070 , \8861 );
nand \U$7188 ( \9072 , \9069 , \9071 );
and \U$7189 ( \9073 , \9067 , \9072 );
and \U$7190 ( \9074 , \8843 , \8864 );
nor \U$7191 ( \9075 , \9074 , \8869 );
or \U$7192 ( \9076 , \9066 , \9075 );
and \U$7193 ( \9077 , \8846 , \8872 );
nor \U$7194 ( \9078 , \9077 , \8876 );
nand \U$7195 ( \9079 , \9076 , \9078 );
nor \U$7196 ( \9080 , \9073 , \9079 );
or \U$7197 ( \9081 , \9064 , \9080 );
and \U$7198 ( \9082 , \8828 , \8879 );
nor \U$7199 ( \9083 , \9082 , \8885 );
or \U$7200 ( \9084 , \9059 , \9083 );
and \U$7201 ( \9085 , \8831 , \8888 );
nor \U$7202 ( \9086 , \9085 , \8892 );
nand \U$7203 ( \9087 , \9084 , \9086 );
and \U$7204 ( \9088 , \9063 , \9087 );
and \U$7205 ( \9089 , \8835 , \8895 );
nor \U$7206 ( \9090 , \9089 , \8900 );
or \U$7207 ( \9091 , \9062 , \9090 );
and \U$7208 ( \9092 , \8838 , \8903 );
nor \U$7209 ( \9093 , \9092 , \8907 );
nand \U$7210 ( \9094 , \9091 , \9093 );
nor \U$7211 ( \9095 , \9088 , \9094 );
nand \U$7212 ( \9096 , \9081 , \9095 );
not \U$7213 ( \9097 , \9096 );
xor \U$7214 ( \9098 , \9057 , \9097 );
buf \U$7215 ( \9099 , \9098 );
_HMUX r3028 ( \9100_nR3028 , \9055 , \9099 , \8731 );
buf \U$7216 ( \9101 , \9100_nR3028 );
not \U$7217 ( \9102 , \4293 );
nand \U$7218 ( \9103 , \4859 , \9102 );
nor \U$7219 ( \9104 , \4686 , \3749 );
nor \U$7220 ( \9105 , \4044 , \4263 );
nand \U$7221 ( \9106 , \9104 , \9105 );
nor \U$7222 ( \9107 , \4747 , \4603 );
not \U$7223 ( \9108 , \4787 );
and \U$7224 ( \9109 , \9107 , \9108 );
or \U$7225 ( \9110 , \4603 , \4798 );
nand \U$7226 ( \9111 , \9110 , \4810 );
nor \U$7227 ( \9112 , \9109 , \9111 );
or \U$7228 ( \9113 , \9106 , \9112 );
or \U$7229 ( \9114 , \3749 , \4821 );
nand \U$7230 ( \9115 , \9114 , \4834 );
and \U$7231 ( \9116 , \9105 , \9115 );
or \U$7232 ( \9117 , \4263 , \4845 );
nand \U$7233 ( \9118 , \9117 , \4857 );
nor \U$7234 ( \9119 , \9116 , \9118 );
nand \U$7235 ( \9120 , \9113 , \9119 );
not \U$7236 ( \9121 , \9120 );
xor \U$7237 ( \9122 , \9103 , \9121 );
buf \U$7238 ( \9123 , \9122 );
not \U$7239 ( \9124 , \7087 );
nand \U$7240 ( \9125 , \7653 , \9124 );
nor \U$7241 ( \9126 , \7480 , \6543 );
nor \U$7242 ( \9127 , \6838 , \7057 );
nand \U$7243 ( \9128 , \9126 , \9127 );
nor \U$7244 ( \9129 , \7541 , \7397 );
not \U$7245 ( \9130 , \7581 );
and \U$7246 ( \9131 , \9129 , \9130 );
or \U$7247 ( \9132 , \7397 , \7592 );
nand \U$7248 ( \9133 , \9132 , \7604 );
nor \U$7249 ( \9134 , \9131 , \9133 );
or \U$7250 ( \9135 , \9128 , \9134 );
or \U$7251 ( \9136 , \6543 , \7615 );
nand \U$7252 ( \9137 , \9136 , \7628 );
and \U$7253 ( \9138 , \9127 , \9137 );
or \U$7254 ( \9139 , \7057 , \7639 );
nand \U$7255 ( \9140 , \9139 , \7651 );
nor \U$7256 ( \9141 , \9138 , \9140 );
nand \U$7257 ( \9142 , \9135 , \9141 );
not \U$7258 ( \9143 , \9142 );
xor \U$7259 ( \9144 , \9125 , \9143 );
buf \U$7260 ( \9145 , \9144 );
_HMUX r2fa3 ( \9146_nR2fa3 , \9123 , \9145 , \8731 );
buf \U$7261 ( \9147 , \9146_nR2fa3 );
not \U$7262 ( \9148 , \4261 );
nand \U$7263 ( \9149 , \4855 , \9148 );
nor \U$7264 ( \9150 , \8756 , \8738 );
nor \U$7265 ( \9151 , \8741 , \8745 );
nand \U$7266 ( \9152 , \9150 , \9151 );
nor \U$7267 ( \9153 , \8760 , \8753 );
not \U$7268 ( \9154 , \8766 );
and \U$7269 ( \9155 , \9153 , \9154 );
or \U$7270 ( \9156 , \8753 , \8773 );
nand \U$7271 ( \9157 , \9156 , \8781 );
nor \U$7272 ( \9158 , \9155 , \9157 );
or \U$7273 ( \9159 , \9152 , \9158 );
or \U$7274 ( \9160 , \8738 , \8788 );
nand \U$7275 ( \9161 , \9160 , \8797 );
and \U$7276 ( \9162 , \9151 , \9161 );
or \U$7277 ( \9163 , \8745 , \8804 );
nand \U$7278 ( \9164 , \9163 , \8812 );
nor \U$7279 ( \9165 , \9162 , \9164 );
nand \U$7280 ( \9166 , \9159 , \9165 );
not \U$7281 ( \9167 , \9166 );
xor \U$7282 ( \9168 , \9149 , \9167 );
buf \U$7283 ( \9169 , \9168 );
not \U$7284 ( \9170 , \7055 );
nand \U$7285 ( \9171 , \7649 , \9170 );
nor \U$7286 ( \9172 , \8848 , \8830 );
nor \U$7287 ( \9173 , \8833 , \8837 );
nand \U$7288 ( \9174 , \9172 , \9173 );
nor \U$7289 ( \9175 , \8852 , \8845 );
not \U$7290 ( \9176 , \8858 );
and \U$7291 ( \9177 , \9175 , \9176 );
or \U$7292 ( \9178 , \8845 , \8865 );
nand \U$7293 ( \9179 , \9178 , \8873 );
nor \U$7294 ( \9180 , \9177 , \9179 );
or \U$7295 ( \9181 , \9174 , \9180 );
or \U$7296 ( \9182 , \8830 , \8880 );
nand \U$7297 ( \9183 , \9182 , \8889 );
and \U$7298 ( \9184 , \9173 , \9183 );
or \U$7299 ( \9185 , \8837 , \8896 );
nand \U$7300 ( \9186 , \9185 , \8904 );
nor \U$7301 ( \9187 , \9184 , \9186 );
nand \U$7302 ( \9188 , \9181 , \9187 );
not \U$7303 ( \9189 , \9188 );
xor \U$7304 ( \9190 , \9171 , \9189 );
buf \U$7305 ( \9191 , \9190 );
_HMUX r2f16 ( \9192_nR2f16 , \9169 , \9191 , \8731 );
buf \U$7306 ( \9193 , \9192_nR2f16 );
not \U$7307 ( \9194 , \4223 );
nand \U$7308 ( \9195 , \4853 , \9194 );
nor \U$7309 ( \9196 , \8930 , \8922 );
nor \U$7310 ( \9197 , \8923 , \8925 );
nand \U$7311 ( \9198 , \9196 , \9197 );
nor \U$7312 ( \9199 , \8932 , \8929 );
and \U$7313 ( \9200 , \9199 , \4781 );
or \U$7314 ( \9201 , \8929 , \8936 );
nand \U$7315 ( \9202 , \9201 , \8940 );
nor \U$7316 ( \9203 , \9200 , \9202 );
or \U$7317 ( \9204 , \9198 , \9203 );
or \U$7318 ( \9205 , \8922 , \8943 );
nand \U$7319 ( \9206 , \9205 , \8948 );
and \U$7320 ( \9207 , \9197 , \9206 );
or \U$7321 ( \9208 , \8925 , \8951 );
nand \U$7322 ( \9209 , \9208 , \8955 );
nor \U$7323 ( \9210 , \9207 , \9209 );
nand \U$7324 ( \9211 , \9204 , \9210 );
not \U$7325 ( \9212 , \9211 );
xor \U$7326 ( \9213 , \9195 , \9212 );
buf \U$7327 ( \9214 , \9213 );
not \U$7328 ( \9215 , \7017 );
nand \U$7329 ( \9216 , \7647 , \9215 );
nor \U$7330 ( \9217 , \8975 , \8967 );
nor \U$7331 ( \9218 , \8968 , \8970 );
nand \U$7332 ( \9219 , \9217 , \9218 );
nor \U$7333 ( \9220 , \8977 , \8974 );
and \U$7334 ( \9221 , \9220 , \7575 );
or \U$7335 ( \9222 , \8974 , \8981 );
nand \U$7336 ( \9223 , \9222 , \8985 );
nor \U$7337 ( \9224 , \9221 , \9223 );
or \U$7338 ( \9225 , \9219 , \9224 );
or \U$7339 ( \9226 , \8967 , \8988 );
nand \U$7340 ( \9227 , \9226 , \8993 );
and \U$7341 ( \9228 , \9218 , \9227 );
or \U$7342 ( \9229 , \8970 , \8996 );
nand \U$7343 ( \9230 , \9229 , \9000 );
nor \U$7344 ( \9231 , \9228 , \9230 );
nand \U$7345 ( \9232 , \9225 , \9231 );
not \U$7346 ( \9233 , \9232 );
xor \U$7347 ( \9234 , \9216 , \9233 );
buf \U$7348 ( \9235 , \9234 );
_HMUX r2e85 ( \9236_nR2e85 , \9214 , \9235 , \8731 );
buf \U$7349 ( \9237 , \9236_nR2e85 );
not \U$7350 ( \9238 , \4166 );
nand \U$7351 ( \9239 , \4850 , \9238 );
nor \U$7352 ( \9240 , \9022 , \9014 );
nor \U$7353 ( \9241 , \9015 , \9017 );
nand \U$7354 ( \9242 , \9240 , \9241 );
nor \U$7355 ( \9243 , \9024 , \9021 );
and \U$7356 ( \9244 , \9243 , \8762 );
or \U$7357 ( \9245 , \9021 , \9027 );
nand \U$7358 ( \9246 , \9245 , \9031 );
nor \U$7359 ( \9247 , \9244 , \9246 );
or \U$7360 ( \9248 , \9242 , \9247 );
or \U$7361 ( \9249 , \9014 , \9034 );
nand \U$7362 ( \9250 , \9249 , \9039 );
and \U$7363 ( \9251 , \9241 , \9250 );
or \U$7364 ( \9252 , \9017 , \9042 );
nand \U$7365 ( \9253 , \9252 , \9046 );
nor \U$7366 ( \9254 , \9251 , \9253 );
nand \U$7367 ( \9255 , \9248 , \9254 );
not \U$7368 ( \9256 , \9255 );
xor \U$7369 ( \9257 , \9239 , \9256 );
buf \U$7370 ( \9258 , \9257 );
not \U$7371 ( \9259 , \6960 );
nand \U$7372 ( \9260 , \7644 , \9259 );
nor \U$7373 ( \9261 , \9066 , \9058 );
nor \U$7374 ( \9262 , \9059 , \9061 );
nand \U$7375 ( \9263 , \9261 , \9262 );
nor \U$7376 ( \9264 , \9068 , \9065 );
and \U$7377 ( \9265 , \9264 , \8854 );
or \U$7378 ( \9266 , \9065 , \9071 );
nand \U$7379 ( \9267 , \9266 , \9075 );
nor \U$7380 ( \9268 , \9265 , \9267 );
or \U$7381 ( \9269 , \9263 , \9268 );
or \U$7382 ( \9270 , \9058 , \9078 );
nand \U$7383 ( \9271 , \9270 , \9083 );
and \U$7384 ( \9272 , \9262 , \9271 );
or \U$7385 ( \9273 , \9061 , \9086 );
nand \U$7386 ( \9274 , \9273 , \9090 );
nor \U$7387 ( \9275 , \9272 , \9274 );
nand \U$7388 ( \9276 , \9269 , \9275 );
not \U$7389 ( \9277 , \9276 );
xor \U$7390 ( \9278 , \9260 , \9277 );
buf \U$7391 ( \9279 , \9278 );
_HMUX r2dec ( \9280_nR2dec , \9258 , \9279 , \8731 );
buf \U$7392 ( \9281 , \9280_nR2dec );
not \U$7393 ( \9282 , \4106 );
nand \U$7394 ( \9283 , \4848 , \9282 );
nand \U$7395 ( \9284 , \4687 , \4045 );
not \U$7396 ( \9285 , \4799 );
or \U$7397 ( \9286 , \9284 , \9285 );
and \U$7398 ( \9287 , \4045 , \4822 );
nor \U$7399 ( \9288 , \9287 , \4846 );
nand \U$7400 ( \9289 , \9286 , \9288 );
not \U$7401 ( \9290 , \9289 );
xor \U$7402 ( \9291 , \9283 , \9290 );
buf \U$7403 ( \9292 , \9291 );
not \U$7404 ( \9293 , \6900 );
nand \U$7405 ( \9294 , \7642 , \9293 );
nand \U$7406 ( \9295 , \7481 , \6839 );
not \U$7407 ( \9296 , \7593 );
or \U$7408 ( \9297 , \9295 , \9296 );
and \U$7409 ( \9298 , \6839 , \7616 );
nor \U$7410 ( \9299 , \9298 , \7640 );
nand \U$7411 ( \9300 , \9297 , \9299 );
not \U$7412 ( \9301 , \9300 );
xor \U$7413 ( \9302 , \9294 , \9301 );
buf \U$7414 ( \9303 , \9302 );
_HMUX r2d4b ( \9304_nR2d4b , \9292 , \9303 , \8731 );
buf \U$7415 ( \9305 , \9304_nR2d4b );
not \U$7416 ( \9306 , \4042 );
nand \U$7417 ( \9307 , \4843 , \9306 );
nand \U$7418 ( \9308 , \8757 , \8742 );
not \U$7419 ( \9309 , \8774 );
or \U$7420 ( \9310 , \9308 , \9309 );
and \U$7421 ( \9311 , \8742 , \8789 );
nor \U$7422 ( \9312 , \9311 , \8805 );
nand \U$7423 ( \9313 , \9310 , \9312 );
not \U$7424 ( \9314 , \9313 );
xor \U$7425 ( \9315 , \9307 , \9314 );
buf \U$7426 ( \9316 , \9315 );
not \U$7427 ( \9317 , \6836 );
nand \U$7428 ( \9318 , \7637 , \9317 );
nand \U$7429 ( \9319 , \8849 , \8834 );
not \U$7430 ( \9320 , \8866 );
or \U$7431 ( \9321 , \9319 , \9320 );
and \U$7432 ( \9322 , \8834 , \8881 );
nor \U$7433 ( \9323 , \9322 , \8897 );
nand \U$7434 ( \9324 , \9321 , \9323 );
not \U$7435 ( \9325 , \9324 );
xor \U$7436 ( \9326 , \9318 , \9325 );
buf \U$7437 ( \9327 , \9326 );
_HMUX r2ca8 ( \9328_nR2ca8 , \9316 , \9327 , \8731 );
buf \U$7438 ( \9329 , \9328_nR2ca8 );
not \U$7439 ( \9330 , \3973 );
nand \U$7440 ( \9331 , \4841 , \9330 );
nand \U$7441 ( \9332 , \8931 , \8924 );
not \U$7442 ( \9333 , \8937 );
or \U$7443 ( \9334 , \9332 , \9333 );
and \U$7444 ( \9335 , \8924 , \8944 );
nor \U$7445 ( \9336 , \9335 , \8952 );
nand \U$7446 ( \9337 , \9334 , \9336 );
not \U$7447 ( \9338 , \9337 );
xor \U$7448 ( \9339 , \9331 , \9338 );
buf \U$7449 ( \9340 , \9339 );
not \U$7450 ( \9341 , \6767 );
nand \U$7451 ( \9342 , \7635 , \9341 );
nand \U$7452 ( \9343 , \8976 , \8969 );
not \U$7453 ( \9344 , \8982 );
or \U$7454 ( \9345 , \9343 , \9344 );
and \U$7455 ( \9346 , \8969 , \8989 );
nor \U$7456 ( \9347 , \9346 , \8997 );
nand \U$7457 ( \9348 , \9345 , \9347 );
not \U$7458 ( \9349 , \9348 );
xor \U$7459 ( \9350 , \9342 , \9349 );
buf \U$7460 ( \9351 , \9350 );
_HMUX r2bf5 ( \9352_nR2bf5 , \9340 , \9351 , \8731 );
buf \U$7461 ( \9353 , \9352_nR2bf5 );
not \U$7462 ( \9354 , \3900 );
nand \U$7463 ( \9355 , \4838 , \9354 );
nand \U$7464 ( \9356 , \9023 , \9016 );
not \U$7465 ( \9357 , \9028 );
or \U$7466 ( \9358 , \9356 , \9357 );
and \U$7467 ( \9359 , \9016 , \9035 );
nor \U$7468 ( \9360 , \9359 , \9043 );
nand \U$7469 ( \9361 , \9358 , \9360 );
not \U$7470 ( \9362 , \9361 );
xor \U$7471 ( \9363 , \9355 , \9362 );
buf \U$7472 ( \9364 , \9363 );
not \U$7473 ( \9365 , \6694 );
nand \U$7474 ( \9366 , \7632 , \9365 );
nand \U$7475 ( \9367 , \9067 , \9060 );
not \U$7476 ( \9368 , \9072 );
or \U$7477 ( \9369 , \9367 , \9368 );
and \U$7478 ( \9370 , \9060 , \9079 );
nor \U$7479 ( \9371 , \9370 , \9087 );
nand \U$7480 ( \9372 , \9369 , \9371 );
not \U$7481 ( \9373 , \9372 );
xor \U$7482 ( \9374 , \9366 , \9373 );
buf \U$7483 ( \9375 , \9374 );
_HMUX r2b3c ( \9376_nR2b3c , \9364 , \9375 , \8731 );
buf \U$7484 ( \9377 , \9376_nR2b3c );
not \U$7485 ( \9378 , \3824 );
nand \U$7486 ( \9379 , \4836 , \9378 );
nand \U$7487 ( \9380 , \9107 , \9104 );
or \U$7488 ( \9381 , \9380 , \4787 );
and \U$7489 ( \9382 , \9104 , \9111 );
nor \U$7490 ( \9383 , \9382 , \9115 );
nand \U$7491 ( \9384 , \9381 , \9383 );
not \U$7492 ( \9385 , \9384 );
xor \U$7493 ( \9386 , \9379 , \9385 );
buf \U$7494 ( \9387 , \9386 );
not \U$7495 ( \9388 , \6618 );
nand \U$7496 ( \9389 , \7630 , \9388 );
nand \U$7497 ( \9390 , \9129 , \9126 );
or \U$7498 ( \9391 , \9390 , \7581 );
and \U$7499 ( \9392 , \9126 , \9133 );
nor \U$7500 ( \9393 , \9392 , \9137 );
nand \U$7501 ( \9394 , \9391 , \9393 );
not \U$7502 ( \9395 , \9394 );
xor \U$7503 ( \9396 , \9389 , \9395 );
buf \U$7504 ( \9397 , \9396 );
_HMUX r2a7b ( \9398_nR2a7b , \9387 , \9397 , \8731 );
buf \U$7505 ( \9399 , \9398_nR2a7b );
not \U$7506 ( \9400 , \3747 );
nand \U$7507 ( \9401 , \4832 , \9400 );
nand \U$7508 ( \9402 , \9153 , \9150 );
or \U$7509 ( \9403 , \9402 , \8766 );
and \U$7510 ( \9404 , \9150 , \9157 );
nor \U$7511 ( \9405 , \9404 , \9161 );
nand \U$7512 ( \9406 , \9403 , \9405 );
not \U$7513 ( \9407 , \9406 );
xor \U$7514 ( \9408 , \9401 , \9407 );
buf \U$7515 ( \9409 , \9408 );
not \U$7516 ( \9410 , \6541 );
nand \U$7517 ( \9411 , \7626 , \9410 );
nand \U$7518 ( \9412 , \9175 , \9172 );
or \U$7519 ( \9413 , \9412 , \8858 );
and \U$7520 ( \9414 , \9172 , \9179 );
nor \U$7521 ( \9415 , \9414 , \9183 );
nand \U$7522 ( \9416 , \9413 , \9415 );
not \U$7523 ( \9417 , \9416 );
xor \U$7524 ( \9418 , \9411 , \9417 );
buf \U$7525 ( \9419 , \9418 );
_HMUX r29bc ( \9420_nR29bc , \9409 , \9419 , \8731 );
buf \U$7526 ( \9421 , \9420_nR29bc );
not \U$7527 ( \9422 , \3672 );
nand \U$7528 ( \9423 , \4830 , \9422 );
nand \U$7529 ( \9424 , \9199 , \9196 );
or \U$7530 ( \9425 , \9424 , \8933 );
and \U$7531 ( \9426 , \9196 , \9202 );
nor \U$7532 ( \9427 , \9426 , \9206 );
nand \U$7533 ( \9428 , \9425 , \9427 );
not \U$7534 ( \9429 , \9428 );
xor \U$7535 ( \9430 , \9423 , \9429 );
buf \U$7536 ( \9431 , \9430 );
not \U$7537 ( \9432 , \6466 );
nand \U$7538 ( \9433 , \7624 , \9432 );
nand \U$7539 ( \9434 , \9220 , \9217 );
or \U$7540 ( \9435 , \9434 , \8978 );
and \U$7541 ( \9436 , \9217 , \9223 );
nor \U$7542 ( \9437 , \9436 , \9227 );
nand \U$7543 ( \9438 , \9435 , \9437 );
not \U$7544 ( \9439 , \9438 );
xor \U$7545 ( \9440 , \9433 , \9439 );
buf \U$7546 ( \9441 , \9440 );
_HMUX r28fd ( \9442_nR28fd , \9431 , \9441 , \8731 );
buf \U$7547 ( \9443 , \9442_nR28fd );
not \U$7548 ( \9444 , \3595 );
nand \U$7549 ( \9445 , \4827 , \9444 );
nand \U$7550 ( \9446 , \9243 , \9240 );
or \U$7551 ( \9447 , \9446 , \4778 );
and \U$7552 ( \9448 , \9240 , \9246 );
nor \U$7553 ( \9449 , \9448 , \9250 );
nand \U$7554 ( \9450 , \9447 , \9449 );
not \U$7555 ( \9451 , \9450 );
xor \U$7556 ( \9452 , \9445 , \9451 );
buf \U$7557 ( \9453 , \9452 );
not \U$7558 ( \9454 , \6389 );
nand \U$7559 ( \9455 , \7621 , \9454 );
nand \U$7560 ( \9456 , \9264 , \9261 );
or \U$7561 ( \9457 , \9456 , \7572 );
and \U$7562 ( \9458 , \9261 , \9267 );
nor \U$7563 ( \9459 , \9458 , \9271 );
nand \U$7564 ( \9460 , \9457 , \9459 );
not \U$7565 ( \9461 , \9460 );
xor \U$7566 ( \9462 , \9455 , \9461 );
buf \U$7567 ( \9463 , \9462 );
_HMUX r2814 ( \9464_nR2814 , \9453 , \9463 , \8731 );
buf \U$7568 ( \9465 , \9464_nR2814 );
not \U$7569 ( \9466 , \3520 );
nand \U$7570 ( \9467 , \4825 , \9466 );
xor \U$7571 ( \9468 , \9467 , \4823 );
buf \U$7572 ( \9469 , \9468 );
not \U$7573 ( \9470 , \6314 );
nand \U$7574 ( \9471 , \7619 , \9470 );
xor \U$7575 ( \9472 , \9471 , \7617 );
buf \U$7576 ( \9473 , \9472 );
_HMUX r272d ( \9474_nR272d , \9469 , \9473 , \8731 );
buf \U$7577 ( \9475 , \9474_nR272d );
not \U$7578 ( \9476 , \4684 );
nand \U$7579 ( \9477 , \4819 , \9476 );
xor \U$7580 ( \9478 , \9477 , \8790 );
buf \U$7581 ( \9479 , \9478 );
not \U$7582 ( \9480 , \7478 );
nand \U$7583 ( \9481 , \7613 , \9480 );
xor \U$7584 ( \9482 , \9481 , \8882 );
buf \U$7585 ( \9483 , \9482 );
_HMUX r2654 ( \9484_nR2654 , \9479 , \9483 , \8731 );
buf \U$7586 ( \9485 , \9484_nR2654 );
not \U$7587 ( \9486 , \4677 );
nand \U$7588 ( \9487 , \4817 , \9486 );
xor \U$7589 ( \9488 , \9487 , \8945 );
buf \U$7590 ( \9489 , \9488 );
not \U$7591 ( \9490 , \7471 );
nand \U$7592 ( \9491 , \7611 , \9490 );
xor \U$7593 ( \9492 , \9491 , \8990 );
buf \U$7594 ( \9493 , \9492 );
_HMUX r257b ( \9494_nR257b , \9489 , \9493 , \8731 );
buf \U$7595 ( \9495 , \9494_nR257b );
not \U$7596 ( \9496 , \4661 );
nand \U$7597 ( \9497 , \4814 , \9496 );
xor \U$7598 ( \9498 , \9497 , \9036 );
buf \U$7599 ( \9499 , \9498 );
not \U$7600 ( \9500 , \7455 );
nand \U$7601 ( \9501 , \7608 , \9500 );
xor \U$7602 ( \9502 , \9501 , \9080 );
buf \U$7603 ( \9503 , \9502 );
_HMUX r24aa ( \9504_nR24aa , \9499 , \9503 , \8731 );
buf \U$7604 ( \9505 , \9504_nR24aa );
not \U$7605 ( \9506 , \4640 );
nand \U$7606 ( \9507 , \4812 , \9506 );
xor \U$7607 ( \9508 , \9507 , \9112 );
buf \U$7608 ( \9509 , \9508 );
not \U$7609 ( \9510 , \7434 );
nand \U$7610 ( \9511 , \7606 , \9510 );
xor \U$7611 ( \9512 , \9511 , \9134 );
buf \U$7612 ( \9513 , \9512 );
_HMUX r23d5 ( \9514_nR23d5 , \9509 , \9513 , \8731 );
buf \U$7613 ( \9515 , \9514_nR23d5 );
not \U$7614 ( \9516 , \4601 );
nand \U$7615 ( \9517 , \4808 , \9516 );
xor \U$7616 ( \9518 , \9517 , \9158 );
buf \U$7617 ( \9519 , \9518 );
not \U$7618 ( \9520 , \7395 );
nand \U$7619 ( \9521 , \7602 , \9520 );
xor \U$7620 ( \9522 , \9521 , \9180 );
buf \U$7621 ( \9523 , \9522 );
_HMUX r230a ( \9524_nR230a , \9519 , \9523 , \8731 );
buf \U$7622 ( \9525 , \9524_nR230a );
not \U$7623 ( \9526 , \4546 );
nand \U$7624 ( \9527 , \4806 , \9526 );
xor \U$7625 ( \9528 , \9527 , \9203 );
buf \U$7626 ( \9529 , \9528 );
not \U$7627 ( \9530 , \7340 );
nand \U$7628 ( \9531 , \7600 , \9530 );
xor \U$7629 ( \9532 , \9531 , \9224 );
buf \U$7630 ( \9533 , \9532 );
_HMUX r21f1 ( \9534_nR21f1 , \9529 , \9533 , \8731 );
buf \U$7631 ( \9535 , \9534_nR21f1 );
not \U$7632 ( \9536 , \4494 );
nand \U$7633 ( \9537 , \4803 , \9536 );
xor \U$7634 ( \9538 , \9537 , \9247 );
buf \U$7635 ( \9539 , \9538 );
not \U$7636 ( \9540 , \7288 );
nand \U$7637 ( \9541 , \7597 , \9540 );
xor \U$7638 ( \9542 , \9541 , \9268 );
buf \U$7639 ( \9543 , \9542 );
_HMUX r213c ( \9544_nR213c , \9539 , \9543 , \8731 );
buf \U$7640 ( \9545 , \9544_nR213c );
not \U$7641 ( \9546 , \4449 );
nand \U$7642 ( \9547 , \4801 , \9546 );
xor \U$7643 ( \9548 , \9547 , \9285 );
buf \U$7644 ( \9549 , \9548 );
not \U$7645 ( \9550 , \7243 );
nand \U$7646 ( \9551 , \7595 , \9550 );
xor \U$7647 ( \9552 , \9551 , \9296 );
buf \U$7648 ( \9553 , \9552 );
_HMUX r2009 ( \9554_nR2009 , \9549 , \9553 , \8731 );
buf \U$7649 ( \9555 , \9554_nR2009 );
not \U$7650 ( \9556 , \4745 );
nand \U$7651 ( \9557 , \4796 , \9556 );
xor \U$7652 ( \9558 , \9557 , \9309 );
buf \U$7653 ( \9559 , \9558 );
not \U$7654 ( \9560 , \7539 );
nand \U$7655 ( \9561 , \7590 , \9560 );
xor \U$7656 ( \9562 , \9561 , \9320 );
buf \U$7657 ( \9563 , \9562 );
_HMUX r1f6c ( \9564_nR1f6c , \9559 , \9563 , \8731 );
buf \U$7658 ( \9565 , \9564_nR1f6c );
not \U$7659 ( \9566 , \4742 );
nand \U$7660 ( \9567 , \4794 , \9566 );
xor \U$7661 ( \9568 , \9567 , \9333 );
buf \U$7662 ( \9569 , \9568 );
not \U$7663 ( \9570 , \7536 );
nand \U$7664 ( \9571 , \7588 , \9570 );
xor \U$7665 ( \9572 , \9571 , \9344 );
buf \U$7666 ( \9573 , \9572 );
_HMUX r1e51 ( \9574_nR1e51 , \9569 , \9573 , \8731 );
buf \U$7667 ( \9575 , \9574_nR1e51 );
not \U$7668 ( \9576 , \4731 );
nand \U$7669 ( \9577 , \4791 , \9576 );
xor \U$7670 ( \9578 , \9577 , \9357 );
buf \U$7671 ( \9579 , \9578 );
not \U$7672 ( \9580 , \7525 );
nand \U$7673 ( \9581 , \7585 , \9580 );
xor \U$7674 ( \9582 , \9581 , \9368 );
buf \U$7675 ( \9583 , \9582 );
_HMUX r1dc8 ( \9584_nR1dc8 , \9579 , \9583 , \8731 );
buf \U$7676 ( \9585 , \9584_nR1dc8 );
not \U$7677 ( \9586 , \4720 );
nand \U$7678 ( \9587 , \4789 , \9586 );
xor \U$7679 ( \9588 , \9587 , \4787 );
buf \U$7680 ( \9589 , \9588 );
not \U$7681 ( \9590 , \7514 );
nand \U$7682 ( \9591 , \7583 , \9590 );
xor \U$7683 ( \9592 , \9591 , \7581 );
buf \U$7684 ( \9593 , \9592 );
_HMUX r1cc1 ( \9594_nR1cc1 , \9589 , \9593 , \8731 );
buf \U$7685 ( \9595 , \9594_nR1cc1 );
not \U$7686 ( \9596 , \4765 );
nand \U$7687 ( \9597 , \4785 , \9596 );
xor \U$7688 ( \9598 , \9597 , \8766 );
buf \U$7689 ( \9599 , \9598 );
not \U$7690 ( \9600 , \7559 );
nand \U$7691 ( \9601 , \7579 , \9600 );
xor \U$7692 ( \9602 , \9601 , \8858 );
buf \U$7693 ( \9603 , \9602 );
_HMUX r1c54 ( \9604_nR1c54 , \9599 , \9603 , \8731 );
buf \U$7694 ( \9605 , \9604_nR1c54 );
not \U$7695 ( \9606 , \4762 );
nand \U$7696 ( \9607 , \4783 , \9606 );
xor \U$7697 ( \9608 , \9607 , \8933 );
buf \U$7698 ( \9609 , \9608 );
not \U$7699 ( \9610 , \7556 );
nand \U$7700 ( \9611 , \7577 , \9610 );
xor \U$7701 ( \9612 , \9611 , \8978 );
buf \U$7702 ( \9613 , \9612 );
_HMUX r1b67 ( \9614_nR1b67 , \9609 , \9613 , \8731 );
buf \U$7703 ( \9615 , \9614_nR1b67 );
not \U$7704 ( \9616 , \4770 );
nand \U$7705 ( \9617 , \4780 , \9616 );
xor \U$7706 ( \9618 , \9617 , \4778 );
buf \U$7707 ( \9619 , \9618 );
not \U$7708 ( \9620 , \7564 );
nand \U$7709 ( \9621 , \7574 , \9620 );
xor \U$7710 ( \9622 , \9621 , \7572 );
buf \U$7711 ( \9623 , \9622 );
_HMUX r1b12 ( \9624_nR1b12 , \9619 , \9623 , \8731 );
buf \U$7712 ( \9625 , \9624_nR1b12 );
nor \U$7713 ( \9626 , \4774 , \4777 );
not \U$7714 ( \9627 , \9626 );
nand \U$7715 ( \9628 , \4778 , \9627 );
not \U$7716 ( \9629 , \9628 );
buf \U$7717 ( \9630 , \9629 );
nor \U$7718 ( \9631 , \7568 , \7571 );
not \U$7719 ( \9632 , \9631 );
nand \U$7720 ( \9633 , \7572 , \9632 );
not \U$7721 ( \9634 , \9633 );
buf \U$7722 ( \9635 , \9634 );
_HMUX r1a41 ( \9636_nR1a41 , \9630 , \9635 , \8731 );
buf \U$7723 ( \9637 , \9636_nR1a41 );
xor \U$7724 ( \9638 , \4776 , \2935 );
buf \U$7725 ( \9639 , \9638 );
xor \U$7726 ( \9640 , \7570 , \5729 );
buf \U$7727 ( \9641 , \9640 );
_HMUX r19fc ( \9642_nR19fc , \9639 , \9641 , \8731 );
buf \U$7728 ( \9643 , \9642_nR19fc );
buf \U$7733 ( \9644 , RI2b5e785db058_15);
buf \U$7734 ( \9645 , RI2b5e785dafe0_16);
buf \U$7735 ( \9646 , RI2b5e785daf68_17);
buf \U$7736 ( \9647 , RI2b5e785daef0_18);
buf \U$7737 ( \9648 , RI2b5e785dae78_19);
buf \U$7738 ( \9649 , RI2b5e785dae00_20);
buf \U$7739 ( \9650 , RI2b5e785dad88_21);
buf \U$7740 ( \9651 , RI2b5e785dad10_22);
buf \U$7741 ( \9652 , RI2b5e785dac98_23);
buf \U$7742 ( \9653 , RI2b5e785dac20_24);
buf \U$7743 ( \9654 , RI2b5e785daba8_25);
and \U$7744 ( \9655 , \9653 , \9654 );
and \U$7745 ( \9656 , \9652 , \9655 );
and \U$7746 ( \9657 , \9651 , \9656 );
and \U$7747 ( \9658 , \9650 , \9657 );
and \U$7748 ( \9659 , \9649 , \9658 );
and \U$7749 ( \9660 , \9648 , \9659 );
and \U$7750 ( \9661 , \9647 , \9660 );
and \U$7751 ( \9662 , \9646 , \9661 );
and \U$7752 ( \9663 , \9645 , \9662 );
xor \U$7753 ( \9664 , \9644 , \9663 );
buf \U$7754 ( \9665 , \9664 );
buf \U$7755 ( \9666 , \9665 );
not \U$7756 ( \9667 , RI2b5e785ae580_609);
nor \U$7757 ( \9668 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$7758 ( \9669 , RI2b5e785daa40_28, \9668 );
and \U$7759 ( \9670 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$7760 ( \9671 , RI2b5e78549540_41, \9670 );
not \U$7761 ( \9672 , RI2b5e785ae3a0_613);
and \U$7762 ( \9673 , \9672 , RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$7763 ( \9674 , RI2b5e785388a8_54, \9673 );
not \U$7764 ( \9675 , RI2b5e785ae418_612);
and \U$7765 ( \9676 , RI2b5e785ae3a0_613, \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$7766 ( \9677 , RI2b5e784a6330_67, \9676 );
and \U$7767 ( \9678 , \9672 , \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$7768 ( \9679 , RI2b5e78495698_80, \9678 );
not \U$7769 ( \9680 , RI2b5e785ae490_611);
and \U$7770 ( \9681 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, \9667 );
and \U$7771 ( \9682 , RI2b5e78495080_93, \9681 );
and \U$7772 ( \9683 , \9672 , RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, \9667 );
and \U$7773 ( \9684 , RI2b5e78403b80_106, \9683 );
and \U$7774 ( \9685 , RI2b5e785ae3a0_613, \9675 , \9680 , RI2b5e785ae508_610, \9667 );
and \U$7775 ( \9686 , RI2b5e775b1e60_119, \9685 );
and \U$7776 ( \9687 , \9672 , \9675 , \9680 , RI2b5e785ae508_610, \9667 );
and \U$7777 ( \9688 , RI2b5e7750bdf8_132, \9687 );
nor \U$7778 ( \9689 , \9672 , \9675 , \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7779 ( \9690 , RI2b5e774ff5d0_145, \9689 );
nor \U$7780 ( \9691 , RI2b5e785ae3a0_613, \9675 , \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7781 ( \9692 , RI2b5e774f65e8_158, \9691 );
nor \U$7782 ( \9693 , \9672 , RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7783 ( \9694 , RI2b5e774eabd0_171, \9693 );
nor \U$7784 ( \9695 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7785 ( \9696 , RI2b5e774de3a8_184, \9695 );
nor \U$7786 ( \9697 , \9672 , \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7787 ( \9698 , RI2b5e774d53c0_197, \9697 );
nor \U$7788 ( \9699 , RI2b5e785ae3a0_613, \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7789 ( \9700 , RI2b5e785f4300_210, \9699 );
nor \U$7790 ( \9701 , \9672 , RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7791 ( \9702 , RI2b5e785f3ce8_223, \9701 );
nor \U$7792 ( \9703 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$7793 ( \9704 , RI2b5e785eb0c0_236, \9703 );
or \U$7794 ( \9705 , \9669 , \9671 , \9674 , \9677 , \9679 , \9682 , \9684 , \9686 , \9688 , \9690 , \9692 , \9694 , \9696 , \9698 , \9700 , \9702 , \9704 );
buf \U$7795 ( \9706 , RI2b5e785ae580_609);
buf \U$7796 ( \9707 , RI2b5e785ae3a0_613);
buf \U$7797 ( \9708 , RI2b5e785ae418_612);
buf \U$7798 ( \9709 , RI2b5e785ae490_611);
buf \U$7799 ( \9710 , RI2b5e785ae508_610);
or \U$7800 ( \9711 , \9707 , \9708 , \9709 , \9710 );
and \U$7801 ( \9712 , \9706 , \9711 );
buf \U$7802 ( \9713 , \9712 );
_DC r3911 ( \9714_nR3911 , \9705 , \9713 );
buf \U$7803 ( \9715 , \9714_nR3911 );
not \U$7804 ( \9716 , \9715 );
xor \U$7805 ( \9717 , \9666 , \9716 );
xor \U$7806 ( \9718 , \9645 , \9662 );
buf \U$7807 ( \9719 , \9718 );
buf \U$7808 ( \9720 , \9719 );
and \U$7809 ( \9721 , RI2b5e785da9c8_29, \9668 );
and \U$7810 ( \9722 , RI2b5e785494c8_42, \9670 );
and \U$7811 ( \9723 , RI2b5e78538830_55, \9673 );
and \U$7812 ( \9724 , RI2b5e784a62b8_68, \9676 );
and \U$7813 ( \9725 , RI2b5e78495620_81, \9678 );
and \U$7814 ( \9726 , RI2b5e78495008_94, \9681 );
and \U$7815 ( \9727 , RI2b5e78403b08_107, \9683 );
and \U$7816 ( \9728 , RI2b5e775b1de8_120, \9685 );
and \U$7817 ( \9729 , RI2b5e7750bd80_133, \9687 );
and \U$7818 ( \9730 , RI2b5e774ff558_146, \9689 );
and \U$7819 ( \9731 , RI2b5e774f6570_159, \9691 );
and \U$7820 ( \9732 , RI2b5e774eab58_172, \9693 );
and \U$7821 ( \9733 , RI2b5e774de330_185, \9695 );
and \U$7822 ( \9734 , RI2b5e774d5348_198, \9697 );
and \U$7823 ( \9735 , RI2b5e785f4288_211, \9699 );
and \U$7824 ( \9736 , RI2b5e785f3658_224, \9701 );
and \U$7825 ( \9737 , RI2b5e785eb048_237, \9703 );
or \U$7826 ( \9738 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 );
_DC r38ed ( \9739_nR38ed , \9738 , \9713 );
buf \U$7827 ( \9740 , \9739_nR38ed );
not \U$7828 ( \9741 , \9740 );
and \U$7829 ( \9742 , \9720 , \9741 );
xor \U$7830 ( \9743 , \9646 , \9661 );
buf \U$7831 ( \9744 , \9743 );
buf \U$7832 ( \9745 , \9744 );
and \U$7833 ( \9746 , RI2b5e785da950_30, \9668 );
and \U$7834 ( \9747 , RI2b5e78549450_43, \9670 );
and \U$7835 ( \9748 , RI2b5e785387b8_56, \9673 );
and \U$7836 ( \9749 , RI2b5e784a6240_69, \9676 );
and \U$7837 ( \9750 , RI2b5e784955a8_82, \9678 );
and \U$7838 ( \9751 , RI2b5e78494f90_95, \9681 );
and \U$7839 ( \9752 , RI2b5e78403a90_108, \9683 );
and \U$7840 ( \9753 , RI2b5e775b1d70_121, \9685 );
and \U$7841 ( \9754 , RI2b5e7750bd08_134, \9687 );
and \U$7842 ( \9755 , RI2b5e774ff4e0_147, \9689 );
and \U$7843 ( \9756 , RI2b5e774f64f8_160, \9691 );
and \U$7844 ( \9757 , RI2b5e774eaae0_173, \9693 );
and \U$7845 ( \9758 , RI2b5e774de2b8_186, \9695 );
and \U$7846 ( \9759 , RI2b5e774d52d0_199, \9697 );
and \U$7847 ( \9760 , RI2b5e785f4210_212, \9699 );
and \U$7848 ( \9761 , RI2b5e785eb5e8_225, \9701 );
and \U$7849 ( \9762 , RI2b5e785e6c50_238, \9703 );
or \U$7850 ( \9763 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 );
_DC r3766 ( \9764_nR3766 , \9763 , \9713 );
buf \U$7851 ( \9765 , \9764_nR3766 );
not \U$7852 ( \9766 , \9765 );
and \U$7853 ( \9767 , \9745 , \9766 );
xor \U$7854 ( \9768 , \9647 , \9660 );
buf \U$7855 ( \9769 , \9768 );
buf \U$7856 ( \9770 , \9769 );
and \U$7857 ( \9771 , RI2b5e785da8d8_31, \9668 );
and \U$7858 ( \9772 , RI2b5e785493d8_44, \9670 );
and \U$7859 ( \9773 , RI2b5e78538740_57, \9673 );
and \U$7860 ( \9774 , RI2b5e784a61c8_70, \9676 );
and \U$7861 ( \9775 , RI2b5e78495530_83, \9678 );
and \U$7862 ( \9776 , RI2b5e78494f18_96, \9681 );
and \U$7863 ( \9777 , RI2b5e78403a18_109, \9683 );
and \U$7864 ( \9778 , RI2b5e775b1cf8_122, \9685 );
and \U$7865 ( \9779 , RI2b5e7750bc90_135, \9687 );
and \U$7866 ( \9780 , RI2b5e774ff468_148, \9689 );
and \U$7867 ( \9781 , RI2b5e774f6480_161, \9691 );
and \U$7868 ( \9782 , RI2b5e774eaa68_174, \9693 );
and \U$7869 ( \9783 , RI2b5e774de240_187, \9695 );
and \U$7870 ( \9784 , RI2b5e774d5258_200, \9697 );
and \U$7871 ( \9785 , RI2b5e785f4198_213, \9699 );
and \U$7872 ( \9786 , RI2b5e785eb570_226, \9701 );
and \U$7873 ( \9787 , RI2b5e785e6bd8_239, \9703 );
or \U$7874 ( \9788 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 );
_DC r3742 ( \9789_nR3742 , \9788 , \9713 );
buf \U$7875 ( \9790 , \9789_nR3742 );
not \U$7876 ( \9791 , \9790 );
and \U$7877 ( \9792 , \9770 , \9791 );
xor \U$7878 ( \9793 , \9648 , \9659 );
buf \U$7879 ( \9794 , \9793 );
buf \U$7880 ( \9795 , \9794 );
and \U$7881 ( \9796 , RI2b5e785da860_32, \9668 );
and \U$7882 ( \9797 , RI2b5e78549360_45, \9670 );
and \U$7883 ( \9798 , RI2b5e785386c8_58, \9673 );
and \U$7884 ( \9799 , RI2b5e784a6150_71, \9676 );
and \U$7885 ( \9800 , RI2b5e784954b8_84, \9678 );
and \U$7886 ( \9801 , RI2b5e78494ea0_97, \9681 );
and \U$7887 ( \9802 , RI2b5e784039a0_110, \9683 );
and \U$7888 ( \9803 , RI2b5e775b1c80_123, \9685 );
and \U$7889 ( \9804 , RI2b5e7750bc18_136, \9687 );
and \U$7890 ( \9805 , RI2b5e774ff3f0_149, \9689 );
and \U$7891 ( \9806 , RI2b5e774f6408_162, \9691 );
and \U$7892 ( \9807 , RI2b5e774ea9f0_175, \9693 );
and \U$7893 ( \9808 , RI2b5e774de1c8_188, \9695 );
and \U$7894 ( \9809 , RI2b5e774d51e0_201, \9697 );
and \U$7895 ( \9810 , RI2b5e785f4120_214, \9699 );
and \U$7896 ( \9811 , RI2b5e785eb4f8_227, \9701 );
and \U$7897 ( \9812 , RI2b5e785e64d0_240, \9703 );
or \U$7898 ( \9813 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 );
_DC r35cd ( \9814_nR35cd , \9813 , \9713 );
buf \U$7899 ( \9815 , \9814_nR35cd );
not \U$7900 ( \9816 , \9815 );
and \U$7901 ( \9817 , \9795 , \9816 );
xor \U$7902 ( \9818 , \9649 , \9658 );
buf \U$7903 ( \9819 , \9818 );
buf \U$7904 ( \9820 , \9819 );
and \U$7905 ( \9821 , RI2b5e78549900_33, \9668 );
and \U$7906 ( \9822 , RI2b5e78538c68_46, \9670 );
and \U$7907 ( \9823 , RI2b5e78538650_59, \9673 );
and \U$7908 ( \9824 , RI2b5e784a60d8_72, \9676 );
and \U$7909 ( \9825 , RI2b5e78495440_85, \9678 );
and \U$7910 ( \9826 , RI2b5e78494e28_98, \9681 );
and \U$7911 ( \9827 , RI2b5e78403928_111, \9683 );
and \U$7912 ( \9828 , RI2b5e775b1c08_124, \9685 );
and \U$7913 ( \9829 , RI2b5e7750bba0_137, \9687 );
and \U$7914 ( \9830 , RI2b5e774ff378_150, \9689 );
and \U$7915 ( \9831 , RI2b5e774f6390_163, \9691 );
and \U$7916 ( \9832 , RI2b5e774ea978_176, \9693 );
and \U$7917 ( \9833 , RI2b5e774de150_189, \9695 );
and \U$7918 ( \9834 , RI2b5e774d5168_202, \9697 );
and \U$7919 ( \9835 , RI2b5e785f40a8_215, \9699 );
and \U$7920 ( \9836 , RI2b5e785eb480_228, \9701 );
and \U$7921 ( \9837 , RI2b5e785da608_241, \9703 );
or \U$7922 ( \9838 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 );
_DC r35a9 ( \9839_nR35a9 , \9838 , \9713 );
buf \U$7923 ( \9840 , \9839_nR35a9 );
not \U$7924 ( \9841 , \9840 );
and \U$7925 ( \9842 , \9820 , \9841 );
xor \U$7926 ( \9843 , \9650 , \9657 );
buf \U$7927 ( \9844 , \9843 );
buf \U$7928 ( \9845 , \9844 );
and \U$7929 ( \9846 , RI2b5e78549888_34, \9668 );
and \U$7930 ( \9847 , RI2b5e78538bf0_47, \9670 );
and \U$7931 ( \9848 , RI2b5e785385d8_60, \9673 );
and \U$7932 ( \9849 , RI2b5e784a6060_73, \9676 );
and \U$7933 ( \9850 , RI2b5e784953c8_86, \9678 );
and \U$7934 ( \9851 , RI2b5e78403ec8_99, \9681 );
and \U$7935 ( \9852 , RI2b5e775b21a8_112, \9683 );
and \U$7936 ( \9853 , RI2b5e775b1b90_125, \9685 );
and \U$7937 ( \9854 , RI2b5e7750bb28_138, \9687 );
and \U$7938 ( \9855 , RI2b5e774ff300_151, \9689 );
and \U$7939 ( \9856 , RI2b5e774f6318_164, \9691 );
and \U$7940 ( \9857 , RI2b5e774ea900_177, \9693 );
and \U$7941 ( \9858 , RI2b5e774de0d8_190, \9695 );
and \U$7942 ( \9859 , RI2b5e774d50f0_203, \9697 );
and \U$7943 ( \9860 , RI2b5e785f4030_216, \9699 );
and \U$7944 ( \9861 , RI2b5e785eb408_229, \9701 );
and \U$7945 ( \9862 , RI2b5e785da590_242, \9703 );
or \U$7946 ( \9863 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 );
_DC r346b ( \9864_nR346b , \9863 , \9713 );
buf \U$7947 ( \9865 , \9864_nR346b );
not \U$7948 ( \9866 , \9865 );
and \U$7949 ( \9867 , \9845 , \9866 );
xor \U$7950 ( \9868 , \9651 , \9656 );
buf \U$7951 ( \9869 , \9868 );
buf \U$7952 ( \9870 , \9869 );
and \U$7953 ( \9871 , RI2b5e78549810_35, \9668 );
and \U$7954 ( \9872 , RI2b5e78538b78_48, \9670 );
and \U$7955 ( \9873 , RI2b5e78538560_61, \9673 );
and \U$7956 ( \9874 , RI2b5e784a5fe8_74, \9676 );
and \U$7957 ( \9875 , RI2b5e78495350_87, \9678 );
and \U$7958 ( \9876 , RI2b5e78403e50_100, \9681 );
and \U$7959 ( \9877 , RI2b5e775b2130_113, \9683 );
and \U$7960 ( \9878 , RI2b5e775b1b18_126, \9685 );
and \U$7961 ( \9879 , RI2b5e7750bab0_139, \9687 );
and \U$7962 ( \9880 , RI2b5e774ff288_152, \9689 );
and \U$7963 ( \9881 , RI2b5e774f62a0_165, \9691 );
and \U$7964 ( \9882 , RI2b5e774ea888_178, \9693 );
and \U$7965 ( \9883 , RI2b5e774de060_191, \9695 );
and \U$7966 ( \9884 , RI2b5e774d5078_204, \9697 );
and \U$7967 ( \9885 , RI2b5e785f3fb8_217, \9699 );
and \U$7968 ( \9886 , RI2b5e785eb390_230, \9701 );
and \U$7969 ( \9887 , RI2b5e785da518_243, \9703 );
or \U$7970 ( \9888 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 );
_DC r3447 ( \9889_nR3447 , \9888 , \9713 );
buf \U$7971 ( \9890 , \9889_nR3447 );
not \U$7972 ( \9891 , \9890 );
and \U$7973 ( \9892 , \9870 , \9891 );
xor \U$7974 ( \9893 , \9652 , \9655 );
buf \U$7975 ( \9894 , \9893 );
buf \U$7976 ( \9895 , \9894 );
and \U$7977 ( \9896 , RI2b5e78549798_36, \9668 );
and \U$7978 ( \9897 , RI2b5e78538b00_49, \9670 );
and \U$7979 ( \9898 , RI2b5e785384e8_62, \9673 );
and \U$7980 ( \9899 , RI2b5e784a5f70_75, \9676 );
and \U$7981 ( \9900 , RI2b5e784952d8_88, \9678 );
and \U$7982 ( \9901 , RI2b5e78403dd8_101, \9681 );
and \U$7983 ( \9902 , RI2b5e775b20b8_114, \9683 );
and \U$7984 ( \9903 , RI2b5e775b1aa0_127, \9685 );
and \U$7985 ( \9904 , RI2b5e7750ba38_140, \9687 );
and \U$7986 ( \9905 , RI2b5e774ff210_153, \9689 );
and \U$7987 ( \9906 , RI2b5e774f6228_166, \9691 );
and \U$7988 ( \9907 , RI2b5e774ea810_179, \9693 );
and \U$7989 ( \9908 , RI2b5e774ddfe8_192, \9695 );
and \U$7990 ( \9909 , RI2b5e774d5000_205, \9697 );
and \U$7991 ( \9910 , RI2b5e785f3f40_218, \9699 );
and \U$7992 ( \9911 , RI2b5e785eb318_231, \9701 );
and \U$7993 ( \9912 , RI2b5e785da4a0_244, \9703 );
or \U$7994 ( \9913 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 );
_DC r333a ( \9914_nR333a , \9913 , \9713 );
buf \U$7995 ( \9915 , \9914_nR333a );
not \U$7996 ( \9916 , \9915 );
and \U$7997 ( \9917 , \9895 , \9916 );
xor \U$7998 ( \9918 , \9653 , \9654 );
buf \U$7999 ( \9919 , \9918 );
buf \U$8000 ( \9920 , \9919 );
and \U$8001 ( \9921 , RI2b5e78549720_37, \9668 );
and \U$8002 ( \9922 , RI2b5e78538a88_50, \9670 );
and \U$8003 ( \9923 , RI2b5e78538470_63, \9673 );
and \U$8004 ( \9924 , RI2b5e784a5ef8_76, \9676 );
and \U$8005 ( \9925 , RI2b5e78495260_89, \9678 );
and \U$8006 ( \9926 , RI2b5e78403d60_102, \9681 );
and \U$8007 ( \9927 , RI2b5e775b2040_115, \9683 );
and \U$8008 ( \9928 , RI2b5e775b1a28_128, \9685 );
and \U$8009 ( \9929 , RI2b5e7750b9c0_141, \9687 );
and \U$8010 ( \9930 , RI2b5e774ff198_154, \9689 );
and \U$8011 ( \9931 , RI2b5e774f61b0_167, \9691 );
and \U$8012 ( \9932 , RI2b5e774ea798_180, \9693 );
and \U$8013 ( \9933 , RI2b5e774ddf70_193, \9695 );
and \U$8014 ( \9934 , RI2b5e774d4f88_206, \9697 );
and \U$8015 ( \9935 , RI2b5e785f3ec8_219, \9699 );
and \U$8016 ( \9936 , RI2b5e785eb2a0_232, \9701 );
and \U$8017 ( \9937 , RI2b5e785da428_245, \9703 );
or \U$8018 ( \9938 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 );
_DC r3353 ( \9939_nR3353 , \9938 , \9713 );
buf \U$8019 ( \9940 , \9939_nR3353 );
not \U$8020 ( \9941 , \9940 );
and \U$8021 ( \9942 , \9920 , \9941 );
not \U$8022 ( \9943 , \9654 );
buf \U$8023 ( \9944 , \9943 );
buf \U$8024 ( \9945 , \9944 );
and \U$8025 ( \9946 , RI2b5e785496a8_38, \9668 );
and \U$8026 ( \9947 , RI2b5e78538a10_51, \9670 );
and \U$8027 ( \9948 , RI2b5e785383f8_64, \9673 );
and \U$8028 ( \9949 , RI2b5e784a5e80_77, \9676 );
and \U$8029 ( \9950 , RI2b5e784951e8_90, \9678 );
and \U$8030 ( \9951 , RI2b5e78403ce8_103, \9681 );
and \U$8031 ( \9952 , RI2b5e775b1fc8_116, \9683 );
and \U$8032 ( \9953 , RI2b5e775b19b0_129, \9685 );
and \U$8033 ( \9954 , RI2b5e7750b948_142, \9687 );
and \U$8034 ( \9955 , RI2b5e774ff120_155, \9689 );
and \U$8035 ( \9956 , RI2b5e774f6138_168, \9691 );
and \U$8036 ( \9957 , RI2b5e774ea720_181, \9693 );
and \U$8037 ( \9958 , RI2b5e774ddef8_194, \9695 );
and \U$8038 ( \9959 , RI2b5e774d4f10_207, \9697 );
and \U$8039 ( \9960 , RI2b5e785f3e50_220, \9699 );
and \U$8040 ( \9961 , RI2b5e785eb228_233, \9701 );
and \U$8041 ( \9962 , RI2b5e785da3b0_246, \9703 );
or \U$8042 ( \9963 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 );
_DC r3230 ( \9964_nR3230 , \9963 , \9713 );
buf \U$8043 ( \9965 , \9964_nR3230 );
not \U$8044 ( \9966 , \9965 );
and \U$8045 ( \9967 , \9945 , \9966 );
buf \U$8046 ( \9968 , RI2b5e785dab30_26);
buf \U$8049 ( \9969 , \9968 );
and \U$8050 ( \9970 , RI2b5e78549630_39, \9668 );
and \U$8051 ( \9971 , RI2b5e78538998_52, \9670 );
and \U$8052 ( \9972 , RI2b5e78538380_65, \9673 );
and \U$8053 ( \9973 , RI2b5e784a5e08_78, \9676 );
and \U$8054 ( \9974 , RI2b5e78495170_91, \9678 );
and \U$8055 ( \9975 , RI2b5e78403c70_104, \9681 );
and \U$8056 ( \9976 , RI2b5e775b1f50_117, \9683 );
and \U$8057 ( \9977 , RI2b5e775b1938_130, \9685 );
and \U$8058 ( \9978 , RI2b5e7750b8d0_143, \9687 );
and \U$8059 ( \9979 , RI2b5e774ff0a8_156, \9689 );
and \U$8060 ( \9980 , RI2b5e774f60c0_169, \9691 );
and \U$8061 ( \9981 , RI2b5e774ea6a8_182, \9693 );
and \U$8062 ( \9982 , RI2b5e774dde80_195, \9695 );
and \U$8063 ( \9983 , RI2b5e774d4e98_208, \9697 );
and \U$8064 ( \9984 , RI2b5e785f3dd8_221, \9699 );
and \U$8065 ( \9985 , RI2b5e785eb1b0_234, \9701 );
and \U$8066 ( \9986 , RI2b5e785da338_247, \9703 );
or \U$8067 ( \9987 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 );
_DC r3214 ( \9988_nR3214 , \9987 , \9713 );
buf \U$8068 ( \9989 , \9988_nR3214 );
not \U$8069 ( \9990 , \9989 );
or \U$8070 ( \9991 , \9969 , \9990 );
and \U$8071 ( \9992 , \9966 , \9991 );
and \U$8072 ( \9993 , \9945 , \9991 );
or \U$8073 ( \9994 , \9967 , \9992 , \9993 );
and \U$8074 ( \9995 , \9941 , \9994 );
and \U$8075 ( \9996 , \9920 , \9994 );
or \U$8076 ( \9997 , \9942 , \9995 , \9996 );
and \U$8077 ( \9998 , \9916 , \9997 );
and \U$8078 ( \9999 , \9895 , \9997 );
or \U$8079 ( \10000 , \9917 , \9998 , \9999 );
and \U$8080 ( \10001 , \9891 , \10000 );
and \U$8081 ( \10002 , \9870 , \10000 );
or \U$8082 ( \10003 , \9892 , \10001 , \10002 );
and \U$8083 ( \10004 , \9866 , \10003 );
and \U$8084 ( \10005 , \9845 , \10003 );
or \U$8085 ( \10006 , \9867 , \10004 , \10005 );
and \U$8086 ( \10007 , \9841 , \10006 );
and \U$8087 ( \10008 , \9820 , \10006 );
or \U$8088 ( \10009 , \9842 , \10007 , \10008 );
and \U$8089 ( \10010 , \9816 , \10009 );
and \U$8090 ( \10011 , \9795 , \10009 );
or \U$8091 ( \10012 , \9817 , \10010 , \10011 );
and \U$8092 ( \10013 , \9791 , \10012 );
and \U$8093 ( \10014 , \9770 , \10012 );
or \U$8094 ( \10015 , \9792 , \10013 , \10014 );
and \U$8095 ( \10016 , \9766 , \10015 );
and \U$8096 ( \10017 , \9745 , \10015 );
or \U$8097 ( \10018 , \9767 , \10016 , \10017 );
and \U$8098 ( \10019 , \9741 , \10018 );
and \U$8099 ( \10020 , \9720 , \10018 );
or \U$8100 ( \10021 , \9742 , \10019 , \10020 );
xor \U$8101 ( \10022 , \9717 , \10021 );
buf \U$8102 ( \10023 , \10022 );
buf \U$8103 ( \10024 , \10023 );
xor \U$8104 ( \10025 , \9720 , \9741 );
xor \U$8105 ( \10026 , \10025 , \10018 );
buf \U$8106 ( \10027 , \10026 );
buf \U$8107 ( \10028 , \10027 );
xor \U$8108 ( \10029 , \9745 , \9766 );
xor \U$8109 ( \10030 , \10029 , \10015 );
buf \U$8110 ( \10031 , \10030 );
buf \U$8111 ( \10032 , \10031 );
and \U$8112 ( \10033 , \10028 , \10032 );
not \U$8113 ( \10034 , \10033 );
and \U$8114 ( \10035 , \10024 , \10034 );
not \U$8115 ( \10036 , \10035 );
buf \U$8116 ( \10037 , RI2b5e785ae3a0_613);
buf \U$8117 ( \10038 , RI2b5e785ae5f8_608);
buf \U$8118 ( \10039 , RI2b5e785ae670_607);
buf \U$8119 ( \10040 , RI2b5e785ae6e8_606);
buf \U$8120 ( \10041 , RI2b5e785ae760_605);
buf \U$8121 ( \10042 , RI2b5e785ae7d8_604);
buf \U$8122 ( \10043 , RI2b5e785ae850_603);
buf \U$8123 ( \10044 , RI2b5e785ae8c8_602);
buf \U$8124 ( \10045 , RI2b5e785ae940_601);
buf \U$8125 ( \10046 , RI2b5e785ae580_609);
nor \U$8126 ( \10047 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 );
buf \U$8127 ( \10048 , \10047 );
buf \U$8128 ( \10049 , \10048 );
xor \U$8129 ( \10050 , \10037 , \10049 );
buf \U$8130 ( \10051 , \10050 );
buf \U$8131 ( \10052 , RI2b5e785ae418_612);
and \U$8132 ( \10053 , \10037 , \10049 );
xor \U$8133 ( \10054 , \10052 , \10053 );
buf \U$8134 ( \10055 , \10054 );
buf \U$8135 ( \10056 , RI2b5e785ae490_611);
and \U$8136 ( \10057 , \10052 , \10053 );
xor \U$8137 ( \10058 , \10056 , \10057 );
buf \U$8138 ( \10059 , \10058 );
buf \U$8139 ( \10060 , RI2b5e785ae508_610);
and \U$8140 ( \10061 , \10056 , \10057 );
xor \U$8141 ( \10062 , \10060 , \10061 );
buf \U$8142 ( \10063 , \10062 );
buf \U$8143 ( \10064 , RI2b5e785ae580_609);
and \U$8144 ( \10065 , \10060 , \10061 );
xor \U$8145 ( \10066 , \10064 , \10065 );
buf \U$8146 ( \10067 , \10066 );
not \U$8147 ( \10068 , \10067 );
nor \U$8148 ( \10069 , \10051 , \10055 , \10059 , \10063 , \10068 );
and \U$8149 ( \10070 , RI2b5e785da248_249, \10069 );
and \U$8150 ( \10071 , \10051 , \10055 , \10059 , \10063 , \10068 );
and \U$8151 ( \10072 , RI2b5e785be750_269, \10071 );
not \U$8152 ( \10073 , \10051 );
and \U$8153 ( \10074 , \10073 , \10055 , \10059 , \10063 , \10068 );
and \U$8154 ( \10075 , RI2b5e785bc4a0_289, \10074 );
not \U$8155 ( \10076 , \10055 );
and \U$8156 ( \10077 , \10051 , \10076 , \10059 , \10063 , \10068 );
and \U$8157 ( \10078 , RI2b5e785bbb40_309, \10077 );
and \U$8158 ( \10079 , \10073 , \10076 , \10059 , \10063 , \10068 );
and \U$8159 ( \10080 , RI2b5e785b9c50_329, \10079 );
not \U$8160 ( \10081 , \10059 );
and \U$8161 ( \10082 , \10051 , \10055 , \10081 , \10063 , \10068 );
and \U$8162 ( \10083 , RI2b5e785b8120_349, \10082 );
and \U$8163 ( \10084 , \10073 , \10055 , \10081 , \10063 , \10068 );
and \U$8164 ( \10085 , RI2b5e785b77c0_369, \10084 );
and \U$8165 ( \10086 , \10051 , \10076 , \10081 , \10063 , \10068 );
and \U$8166 ( \10087 , RI2b5e785b6e60_389, \10086 );
and \U$8167 ( \10088 , \10073 , \10076 , \10081 , \10063 , \10068 );
and \U$8168 ( \10089 , RI2b5e785b56f0_409, \10088 );
nor \U$8169 ( \10090 , \10073 , \10076 , \10081 , \10063 , \10067 );
and \U$8170 ( \10091 , RI2b5e785b4d90_429, \10090 );
nor \U$8171 ( \10092 , \10051 , \10076 , \10081 , \10063 , \10067 );
and \U$8172 ( \10093 , RI2b5e785b39e0_449, \10092 );
nor \U$8173 ( \10094 , \10073 , \10055 , \10081 , \10063 , \10067 );
and \U$8174 ( \10095 , RI2b5e785b3080_469, \10094 );
nor \U$8175 ( \10096 , \10051 , \10055 , \10081 , \10063 , \10067 );
and \U$8176 ( \10097 , RI2b5e785b2720_489, \10096 );
nor \U$8177 ( \10098 , \10073 , \10076 , \10059 , \10063 , \10067 );
and \U$8178 ( \10099 , RI2b5e785b1730_509, \10098 );
nor \U$8179 ( \10100 , \10051 , \10076 , \10059 , \10063 , \10067 );
and \U$8180 ( \10101 , RI2b5e785b0dd0_529, \10100 );
nor \U$8181 ( \10102 , \10073 , \10055 , \10059 , \10063 , \10067 );
and \U$8182 ( \10103 , RI2b5e785b0470_549, \10102 );
nor \U$8183 ( \10104 , \10051 , \10055 , \10059 , \10063 , \10067 );
and \U$8184 ( \10105 , RI2b5e785af840_569, \10104 );
or \U$8185 ( \10106 , \10070 , \10072 , \10075 , \10078 , \10080 , \10083 , \10085 , \10087 , \10089 , \10091 , \10093 , \10095 , \10097 , \10099 , \10101 , \10103 , \10105 );
buf \U$8186 ( \10107 , \10067 );
buf \U$8187 ( \10108 , \10051 );
buf \U$8188 ( \10109 , \10055 );
buf \U$8189 ( \10110 , \10059 );
buf \U$8190 ( \10111 , \10063 );
or \U$8191 ( \10112 , \10108 , \10109 , \10110 , \10111 );
and \U$8192 ( \10113 , \10107 , \10112 );
buf \U$8193 ( \10114 , \10113 );
_DC r4011 ( \10115_nR4011 , \10106 , \10114 );
buf \U$8194 ( \10116 , \10115_nR4011 );
buf \U$8195 ( \10117 , RI2b5e785db0d0_14);
and \U$8196 ( \10118 , \9644 , \9663 );
and \U$8197 ( \10119 , \10117 , \10118 );
buf \U$8198 ( \10120 , \10119 );
buf \U$8199 ( \10121 , \10120 );
xor \U$8200 ( \10122 , \10117 , \10118 );
buf \U$8201 ( \10123 , \10122 );
buf \U$8202 ( \10124 , \10123 );
and \U$8203 ( \10125 , RI2b5e785daab8_27, \9668 );
and \U$8204 ( \10126 , RI2b5e785495b8_40, \9670 );
and \U$8205 ( \10127 , RI2b5e78538920_53, \9673 );
and \U$8206 ( \10128 , RI2b5e784a63a8_66, \9676 );
and \U$8207 ( \10129 , RI2b5e78495710_79, \9678 );
and \U$8208 ( \10130 , RI2b5e784950f8_92, \9681 );
and \U$8209 ( \10131 , RI2b5e78403bf8_105, \9683 );
and \U$8210 ( \10132 , RI2b5e775b1ed8_118, \9685 );
and \U$8211 ( \10133 , RI2b5e775b18c0_131, \9687 );
and \U$8212 ( \10134 , RI2b5e7750b858_144, \9689 );
and \U$8213 ( \10135 , RI2b5e774ff030_157, \9691 );
and \U$8214 ( \10136 , RI2b5e774f6048_170, \9693 );
and \U$8215 ( \10137 , RI2b5e774ea630_183, \9695 );
and \U$8216 ( \10138 , RI2b5e774dde08_196, \9697 );
and \U$8217 ( \10139 , RI2b5e774d4e20_209, \9699 );
and \U$8218 ( \10140 , RI2b5e785f3d60_222, \9701 );
and \U$8219 ( \10141 , RI2b5e785eb138_235, \9703 );
or \U$8220 ( \10142 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 );
_DC r3ad9 ( \10143_nR3ad9 , \10142 , \9713 );
buf \U$8221 ( \10144 , \10143_nR3ad9 );
not \U$8222 ( \10145 , \10144 );
and \U$8223 ( \10146 , \10124 , \10145 );
and \U$8224 ( \10147 , \9666 , \9716 );
and \U$8225 ( \10148 , \9716 , \10021 );
and \U$8226 ( \10149 , \9666 , \10021 );
or \U$8227 ( \10150 , \10147 , \10148 , \10149 );
and \U$8228 ( \10151 , \10145 , \10150 );
and \U$8229 ( \10152 , \10124 , \10150 );
or \U$8230 ( \10153 , \10146 , \10151 , \10152 );
xnor \U$8231 ( \10154 , \10121 , \10153 );
buf \U$8232 ( \10155 , \10154 );
buf \U$8233 ( \10156 , \10155 );
xor \U$8234 ( \10157 , \10124 , \10145 );
xor \U$8235 ( \10158 , \10157 , \10150 );
buf \U$8236 ( \10159 , \10158 );
buf \U$8237 ( \10160 , \10159 );
xor \U$8238 ( \10161 , \10156 , \10160 );
xor \U$8239 ( \10162 , \10160 , \10024 );
not \U$8240 ( \10163 , \10162 );
and \U$8241 ( \10164 , \10161 , \10163 );
and \U$8242 ( \10165 , \10116 , \10164 );
and \U$8243 ( \10166 , RI2b5e785da2c0_248, \10069 );
and \U$8244 ( \10167 , RI2b5e785be7c8_268, \10071 );
and \U$8245 ( \10168 , RI2b5e785bc518_288, \10074 );
and \U$8246 ( \10169 , RI2b5e785bbbb8_308, \10077 );
and \U$8247 ( \10170 , RI2b5e785b9cc8_328, \10079 );
and \U$8248 ( \10171 , RI2b5e785b9368_348, \10082 );
and \U$8249 ( \10172 , RI2b5e785b7838_368, \10084 );
and \U$8250 ( \10173 , RI2b5e785b6ed8_388, \10086 );
and \U$8251 ( \10174 , RI2b5e785b5768_408, \10088 );
and \U$8252 ( \10175 , RI2b5e785b4e08_428, \10090 );
and \U$8253 ( \10176 , RI2b5e785b3a58_448, \10092 );
and \U$8254 ( \10177 , RI2b5e785b30f8_468, \10094 );
and \U$8255 ( \10178 , RI2b5e785b2798_488, \10096 );
and \U$8256 ( \10179 , RI2b5e785b17a8_508, \10098 );
and \U$8257 ( \10180 , RI2b5e785b0e48_528, \10100 );
and \U$8258 ( \10181 , RI2b5e785b04e8_548, \10102 );
and \U$8259 ( \10182 , RI2b5e785afb88_568, \10104 );
or \U$8260 ( \10183 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 );
_DC r4105 ( \10184_nR4105 , \10183 , \10114 );
buf \U$8261 ( \10185 , \10184_nR4105 );
and \U$8262 ( \10186 , \10185 , \10162 );
nor \U$8263 ( \10187 , \10165 , \10186 );
and \U$8264 ( \10188 , \10160 , \10024 );
not \U$8265 ( \10189 , \10188 );
and \U$8266 ( \10190 , \10156 , \10189 );
xnor \U$8267 ( \10191 , \10187 , \10190 );
xor \U$8268 ( \10192 , \10036 , \10191 );
and \U$8270 ( \10193 , RI2b5e785da1d0_250, \10069 );
and \U$8271 ( \10194 , RI2b5e785be6d8_270, \10071 );
and \U$8272 ( \10195 , RI2b5e785bc428_290, \10074 );
and \U$8273 ( \10196 , RI2b5e785bbac8_310, \10077 );
and \U$8274 ( \10197 , RI2b5e785b9bd8_330, \10079 );
and \U$8275 ( \10198 , RI2b5e785b80a8_350, \10082 );
and \U$8276 ( \10199 , RI2b5e785b7748_370, \10084 );
and \U$8277 ( \10200 , RI2b5e785b6de8_390, \10086 );
and \U$8278 ( \10201 , RI2b5e785b5678_410, \10088 );
and \U$8279 ( \10202 , RI2b5e785b4d18_430, \10090 );
and \U$8280 ( \10203 , RI2b5e785b3968_450, \10092 );
and \U$8281 ( \10204 , RI2b5e785b3008_470, \10094 );
and \U$8282 ( \10205 , RI2b5e785b26a8_490, \10096 );
and \U$8283 ( \10206 , RI2b5e785b16b8_510, \10098 );
and \U$8284 ( \10207 , RI2b5e785b0d58_530, \10100 );
and \U$8285 ( \10208 , RI2b5e785b03f8_550, \10102 );
and \U$8286 ( \10209 , RI2b5e785af7c8_570, \10104 );
or \U$8287 ( \10210 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 );
_DC r3f4f ( \10211_nR3f4f , \10210 , \10114 );
buf \U$8288 ( \10212 , \10211_nR3f4f );
or \U$8289 ( \10213 , \10121 , \10153 );
not \U$8290 ( \10214 , \10213 );
buf \U$8291 ( \10215 , \10214 );
buf \U$8292 ( \10216 , \10215 );
xor \U$8293 ( \10217 , \10216 , \10156 );
and \U$8294 ( \10218 , \10212 , \10217 );
nor \U$8295 ( \10219 , 1'b0 , \10218 );
xnor \U$8297 ( \10220 , \10219 , 1'b0 );
xor \U$8298 ( \10221 , \10192 , \10220 );
xor \U$8299 ( \10222 , 1'b0 , \10221 );
xor \U$8301 ( \10223 , \10024 , \10028 );
xor \U$8302 ( \10224 , \10028 , \10032 );
not \U$8303 ( \10225 , \10224 );
and \U$8304 ( \10226 , \10223 , \10225 );
and \U$8305 ( \10227 , \10185 , \10226 );
not \U$8306 ( \10228 , \10227 );
xnor \U$8307 ( \10229 , \10228 , \10035 );
and \U$8308 ( \10230 , \10212 , \10164 );
and \U$8309 ( \10231 , \10116 , \10162 );
nor \U$8310 ( \10232 , \10230 , \10231 );
xnor \U$8311 ( \10233 , \10232 , \10190 );
and \U$8312 ( \10234 , \10229 , \10233 );
or \U$8314 ( \10235 , 1'b0 , \10234 , 1'b0 );
xor \U$8316 ( \10236 , \10235 , 1'b0 );
xor \U$8318 ( \10237 , \10236 , 1'b0 );
and \U$8319 ( \10238 , \10222 , \10237 );
or \U$8320 ( \10239 , 1'b0 , 1'b0 , \10238 );
and \U$8323 ( \10240 , \10185 , \10164 );
not \U$8324 ( \10241 , \10240 );
xnor \U$8325 ( \10242 , \10241 , \10190 );
xor \U$8326 ( \10243 , 1'b0 , \10242 );
and \U$8328 ( \10244 , \10116 , \10217 );
nor \U$8329 ( \10245 , 1'b0 , \10244 );
xnor \U$8330 ( \10246 , \10245 , 1'b0 );
xor \U$8331 ( \10247 , \10243 , \10246 );
xor \U$8332 ( \10248 , 1'b0 , \10247 );
xor \U$8334 ( \10249 , \10248 , 1'b1 );
and \U$8335 ( \10250 , \10036 , \10191 );
and \U$8336 ( \10251 , \10191 , \10220 );
and \U$8337 ( \10252 , \10036 , \10220 );
or \U$8338 ( \10253 , \10250 , \10251 , \10252 );
xor \U$8340 ( \10254 , \10253 , 1'b0 );
xor \U$8342 ( \10255 , \10254 , 1'b0 );
xor \U$8343 ( \10256 , \10249 , \10255 );
and \U$8344 ( \10257 , \10239 , \10256 );
or \U$8346 ( \10258 , 1'b0 , \10257 , 1'b0 );
xor \U$8348 ( \10259 , \10258 , 1'b0 );
and \U$8350 ( \10260 , \10248 , 1'b1 );
and \U$8351 ( \10261 , 1'b1 , \10255 );
and \U$8352 ( \10262 , \10248 , \10255 );
or \U$8353 ( \10263 , \10260 , \10261 , \10262 );
xor \U$8354 ( \10264 , 1'b0 , \10263 );
not \U$8356 ( \10265 , \10190 );
and \U$8358 ( \10266 , \10185 , \10217 );
nor \U$8359 ( \10267 , 1'b0 , \10266 );
xnor \U$8360 ( \10268 , \10267 , 1'b0 );
xor \U$8361 ( \10269 , \10265 , \10268 );
xor \U$8363 ( \10270 , \10269 , 1'b0 );
xor \U$8364 ( \10271 , 1'b0 , \10270 );
xor \U$8366 ( \10272 , \10271 , 1'b0 );
and \U$8368 ( \10273 , \10242 , \10246 );
or \U$8370 ( \10274 , 1'b0 , \10273 , 1'b0 );
xor \U$8372 ( \10275 , \10274 , 1'b0 );
xor \U$8374 ( \10276 , \10275 , 1'b0 );
xor \U$8375 ( \10277 , \10272 , \10276 );
xor \U$8376 ( \10278 , \10264 , \10277 );
xor \U$8377 ( \10279 , \10259 , \10278 );
xor \U$8383 ( \10280 , \9770 , \9791 );
xor \U$8384 ( \10281 , \10280 , \10012 );
buf \U$8385 ( \10282 , \10281 );
buf \U$8386 ( \10283 , \10282 );
xor \U$8387 ( \10284 , \10032 , \10283 );
xor \U$8388 ( \10285 , \9795 , \9816 );
xor \U$8389 ( \10286 , \10285 , \10009 );
buf \U$8390 ( \10287 , \10286 );
buf \U$8391 ( \10288 , \10287 );
xor \U$8392 ( \10289 , \10283 , \10288 );
not \U$8393 ( \10290 , \10289 );
and \U$8394 ( \10291 , \10284 , \10290 );
and \U$8395 ( \10292 , \10185 , \10291 );
not \U$8396 ( \10293 , \10292 );
and \U$8397 ( \10294 , \10283 , \10288 );
not \U$8398 ( \10295 , \10294 );
and \U$8399 ( \10296 , \10032 , \10295 );
xnor \U$8400 ( \10297 , \10293 , \10296 );
and \U$8401 ( \10298 , \10212 , \10226 );
and \U$8402 ( \10299 , \10116 , \10224 );
nor \U$8403 ( \10300 , \10298 , \10299 );
xnor \U$8404 ( \10301 , \10300 , \10035 );
and \U$8405 ( \10302 , \10297 , \10301 );
or \U$8407 ( \10303 , 1'b0 , \10302 , 1'b0 );
and \U$8408 ( \10304 , RI2b5e785da0e0_252, \10069 );
and \U$8409 ( \10305 , RI2b5e785be5e8_272, \10071 );
and \U$8410 ( \10306 , RI2b5e785bc338_292, \10074 );
and \U$8411 ( \10307 , RI2b5e785bb9d8_312, \10077 );
and \U$8412 ( \10308 , RI2b5e785b9ae8_332, \10079 );
and \U$8413 ( \10309 , RI2b5e785b7fb8_352, \10082 );
and \U$8414 ( \10310 , RI2b5e785b7658_372, \10084 );
and \U$8415 ( \10311 , RI2b5e785b5ee8_392, \10086 );
and \U$8416 ( \10312 , RI2b5e785b5588_412, \10088 );
and \U$8417 ( \10313 , RI2b5e785b4c28_432, \10090 );
and \U$8418 ( \10314 , RI2b5e785b3878_452, \10092 );
and \U$8419 ( \10315 , RI2b5e785b2f18_472, \10094 );
and \U$8420 ( \10316 , RI2b5e785b25b8_492, \10096 );
and \U$8421 ( \10317 , RI2b5e785b15c8_512, \10098 );
and \U$8422 ( \10318 , RI2b5e785b0c68_532, \10100 );
and \U$8423 ( \10319 , RI2b5e785b0308_552, \10102 );
and \U$8424 ( \10320 , RI2b5e785af6d8_572, \10104 );
or \U$8425 ( \10321 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 );
_DC r3db4 ( \10322_nR3db4 , \10321 , \10114 );
buf \U$8426 ( \10323 , \10322_nR3db4 );
and \U$8427 ( \10324 , \10323 , \10164 );
and \U$8428 ( \10325 , RI2b5e785da158_251, \10069 );
and \U$8429 ( \10326 , RI2b5e785be660_271, \10071 );
and \U$8430 ( \10327 , RI2b5e785bc3b0_291, \10074 );
and \U$8431 ( \10328 , RI2b5e785bba50_311, \10077 );
and \U$8432 ( \10329 , RI2b5e785b9b60_331, \10079 );
and \U$8433 ( \10330 , RI2b5e785b8030_351, \10082 );
and \U$8434 ( \10331 , RI2b5e785b76d0_371, \10084 );
and \U$8435 ( \10332 , RI2b5e785b6d70_391, \10086 );
and \U$8436 ( \10333 , RI2b5e785b5600_411, \10088 );
and \U$8437 ( \10334 , RI2b5e785b4ca0_431, \10090 );
and \U$8438 ( \10335 , RI2b5e785b38f0_451, \10092 );
and \U$8439 ( \10336 , RI2b5e785b2f90_471, \10094 );
and \U$8440 ( \10337 , RI2b5e785b2630_491, \10096 );
and \U$8441 ( \10338 , RI2b5e785b1640_511, \10098 );
and \U$8442 ( \10339 , RI2b5e785b0ce0_531, \10100 );
and \U$8443 ( \10340 , RI2b5e785b0380_551, \10102 );
and \U$8444 ( \10341 , RI2b5e785af750_571, \10104 );
or \U$8445 ( \10342 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 );
_DC r3e8e ( \10343_nR3e8e , \10342 , \10114 );
buf \U$8446 ( \10344 , \10343_nR3e8e );
and \U$8447 ( \10345 , \10344 , \10162 );
nor \U$8448 ( \10346 , \10324 , \10345 );
xnor \U$8449 ( \10347 , \10346 , \10190 );
and \U$8451 ( \10348 , RI2b5e785da068_253, \10069 );
and \U$8452 ( \10349 , RI2b5e785be570_273, \10071 );
and \U$8453 ( \10350 , RI2b5e785bc2c0_293, \10074 );
and \U$8454 ( \10351 , RI2b5e785bb960_313, \10077 );
and \U$8455 ( \10352 , RI2b5e785b9a70_333, \10079 );
and \U$8456 ( \10353 , RI2b5e785b7f40_353, \10082 );
and \U$8457 ( \10354 , RI2b5e785b75e0_373, \10084 );
and \U$8458 ( \10355 , RI2b5e785b5e70_393, \10086 );
and \U$8459 ( \10356 , RI2b5e785b5510_413, \10088 );
and \U$8460 ( \10357 , RI2b5e785b4bb0_433, \10090 );
and \U$8461 ( \10358 , RI2b5e785b3800_453, \10092 );
and \U$8462 ( \10359 , RI2b5e785b2ea0_473, \10094 );
and \U$8463 ( \10360 , RI2b5e785b2540_493, \10096 );
and \U$8464 ( \10361 , RI2b5e785b1550_513, \10098 );
and \U$8465 ( \10362 , RI2b5e785b0bf0_533, \10100 );
and \U$8466 ( \10363 , RI2b5e785b0290_553, \10102 );
and \U$8467 ( \10364 , RI2b5e785af660_573, \10104 );
or \U$8468 ( \10365 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 );
_DC r3cc9 ( \10366_nR3cc9 , \10365 , \10114 );
buf \U$8469 ( \10367 , \10366_nR3cc9 );
and \U$8470 ( \10368 , \10367 , \10217 );
nor \U$8471 ( \10369 , 1'b0 , \10368 );
xnor \U$8472 ( \10370 , \10369 , 1'b0 );
and \U$8473 ( \10371 , \10347 , \10370 );
or \U$8476 ( \10372 , \10371 , 1'b0 , 1'b0 );
and \U$8477 ( \10373 , \10303 , \10372 );
or \U$8480 ( \10374 , \10373 , 1'b0 , 1'b0 );
and \U$8483 ( \10375 , \10323 , \10217 );
nor \U$8484 ( \10376 , 1'b0 , \10375 );
xnor \U$8485 ( \10377 , \10376 , 1'b0 );
xor \U$8487 ( \10378 , \10377 , 1'b0 );
xor \U$8489 ( \10379 , \10378 , 1'b0 );
not \U$8490 ( \10380 , \10296 );
and \U$8491 ( \10381 , \10116 , \10226 );
and \U$8492 ( \10382 , \10185 , \10224 );
nor \U$8493 ( \10383 , \10381 , \10382 );
xnor \U$8494 ( \10384 , \10383 , \10035 );
xor \U$8495 ( \10385 , \10380 , \10384 );
and \U$8496 ( \10386 , \10344 , \10164 );
and \U$8497 ( \10387 , \10212 , \10162 );
nor \U$8498 ( \10388 , \10386 , \10387 );
xnor \U$8499 ( \10389 , \10388 , \10190 );
xor \U$8500 ( \10390 , \10385 , \10389 );
and \U$8501 ( \10391 , \10379 , \10390 );
or \U$8503 ( \10392 , 1'b0 , \10391 , 1'b0 );
and \U$8504 ( \10393 , \10374 , \10392 );
or \U$8505 ( \10394 , 1'b0 , 1'b0 , \10393 );
and \U$8507 ( \10395 , \10344 , \10217 );
nor \U$8508 ( \10396 , 1'b0 , \10395 );
xnor \U$8509 ( \10397 , \10396 , 1'b0 );
xor \U$8511 ( \10398 , \10397 , 1'b0 );
xor \U$8513 ( \10399 , \10398 , 1'b0 );
xor \U$8515 ( \10400 , 1'b0 , \10229 );
xor \U$8516 ( \10401 , \10400 , \10233 );
xor \U$8517 ( \10402 , \10399 , \10401 );
and \U$8519 ( \10403 , \10402 , 1'b1 );
and \U$8520 ( \10404 , \10380 , \10384 );
and \U$8521 ( \10405 , \10384 , \10389 );
and \U$8522 ( \10406 , \10380 , \10389 );
or \U$8523 ( \10407 , \10404 , \10405 , \10406 );
xor \U$8525 ( \10408 , \10407 , 1'b0 );
xor \U$8527 ( \10409 , \10408 , 1'b0 );
and \U$8528 ( \10410 , 1'b1 , \10409 );
and \U$8529 ( \10411 , \10402 , \10409 );
or \U$8530 ( \10412 , \10403 , \10410 , \10411 );
and \U$8531 ( \10413 , \10394 , \10412 );
xor \U$8533 ( \10414 , \10222 , 1'b0 );
xor \U$8534 ( \10415 , \10414 , \10237 );
and \U$8535 ( \10416 , \10412 , \10415 );
and \U$8536 ( \10417 , \10394 , \10415 );
or \U$8537 ( \10418 , \10413 , \10416 , \10417 );
xor \U$8539 ( \10419 , 1'b0 , \10239 );
xor \U$8540 ( \10420 , \10419 , \10256 );
and \U$8541 ( \10421 , \10418 , \10420 );
or \U$8542 ( \10422 , 1'b0 , 1'b0 , \10421 );
nand \U$8543 ( \10423 , \10279 , \10422 );
nor \U$8544 ( \10424 , \10279 , \10422 );
not \U$8545 ( \10425 , \10424 );
nand \U$8546 ( \10426 , \10423 , \10425 );
xor \U$8547 ( \10427 , \9945 , \9966 );
xor \U$8548 ( \10428 , \10427 , \9991 );
buf \U$8549 ( \10429 , \10428 );
buf \U$8550 ( \10430 , \10429 );
xor \U$8551 ( \10431 , \9969 , \9989 );
buf \U$8552 ( \10432 , \10431 );
buf \U$8553 ( \10433 , \10432 );
xor \U$8554 ( \10434 , \10430 , \10433 );
not \U$8555 ( \10435 , \10433 );
and \U$8556 ( \10436 , \10434 , \10435 );
and \U$8557 ( \10437 , \10367 , \10436 );
and \U$8558 ( \10438 , \10323 , \10433 );
nor \U$8559 ( \10439 , \10437 , \10438 );
xnor \U$8560 ( \10440 , \10439 , \10430 );
and \U$8561 ( \10441 , RI2b5e785c2bc0_255, \10069 );
and \U$8562 ( \10442 , RI2b5e785be480_275, \10071 );
and \U$8563 ( \10443 , RI2b5e785bc1d0_295, \10074 );
and \U$8564 ( \10444 , RI2b5e785ba2e0_315, \10077 );
and \U$8565 ( \10445 , RI2b5e785b9980_335, \10079 );
and \U$8566 ( \10446 , RI2b5e785b7e50_355, \10082 );
and \U$8567 ( \10447 , RI2b5e785b74f0_375, \10084 );
and \U$8568 ( \10448 , RI2b5e785b5d80_395, \10086 );
and \U$8569 ( \10449 , RI2b5e785b5420_415, \10088 );
and \U$8570 ( \10450 , RI2b5e785b4ac0_435, \10090 );
and \U$8571 ( \10451 , RI2b5e785b3710_455, \10092 );
and \U$8572 ( \10452 , RI2b5e785b2db0_475, \10094 );
and \U$8573 ( \10453 , RI2b5e785b2450_495, \10096 );
and \U$8574 ( \10454 , RI2b5e785b1460_515, \10098 );
and \U$8575 ( \10455 , RI2b5e785b0b00_535, \10100 );
and \U$8576 ( \10456 , RI2b5e785b01a0_555, \10102 );
and \U$8577 ( \10457 , RI2b5e785af570_575, \10104 );
or \U$8578 ( \10458 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 );
_DC r3b16 ( \10459_nR3b16 , \10458 , \10114 );
buf \U$8579 ( \10460 , \10459_nR3b16 );
xor \U$8580 ( \10461 , \9895 , \9916 );
xor \U$8581 ( \10462 , \10461 , \9997 );
buf \U$8582 ( \10463 , \10462 );
buf \U$8583 ( \10464 , \10463 );
xor \U$8584 ( \10465 , \9920 , \9941 );
xor \U$8585 ( \10466 , \10465 , \9994 );
buf \U$8586 ( \10467 , \10466 );
buf \U$8587 ( \10468 , \10467 );
xor \U$8588 ( \10469 , \10464 , \10468 );
xor \U$8589 ( \10470 , \10468 , \10430 );
not \U$8590 ( \10471 , \10470 );
and \U$8591 ( \10472 , \10469 , \10471 );
and \U$8592 ( \10473 , \10460 , \10472 );
and \U$8593 ( \10474 , RI2b5e785c2c38_254, \10069 );
and \U$8594 ( \10475 , RI2b5e785be4f8_274, \10071 );
and \U$8595 ( \10476 , RI2b5e785bc248_294, \10074 );
and \U$8596 ( \10477 , RI2b5e785ba358_314, \10077 );
and \U$8597 ( \10478 , RI2b5e785b99f8_334, \10079 );
and \U$8598 ( \10479 , RI2b5e785b7ec8_354, \10082 );
and \U$8599 ( \10480 , RI2b5e785b7568_374, \10084 );
and \U$8600 ( \10481 , RI2b5e785b5df8_394, \10086 );
and \U$8601 ( \10482 , RI2b5e785b5498_414, \10088 );
and \U$8602 ( \10483 , RI2b5e785b4b38_434, \10090 );
and \U$8603 ( \10484 , RI2b5e785b3788_454, \10092 );
and \U$8604 ( \10485 , RI2b5e785b2e28_474, \10094 );
and \U$8605 ( \10486 , RI2b5e785b24c8_494, \10096 );
and \U$8606 ( \10487 , RI2b5e785b14d8_514, \10098 );
and \U$8607 ( \10488 , RI2b5e785b0b78_534, \10100 );
and \U$8608 ( \10489 , RI2b5e785b0218_554, \10102 );
and \U$8609 ( \10490 , RI2b5e785af5e8_574, \10104 );
or \U$8610 ( \10491 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 );
_DC r3bea ( \10492_nR3bea , \10491 , \10114 );
buf \U$8611 ( \10493 , \10492_nR3bea );
and \U$8612 ( \10494 , \10493 , \10470 );
nor \U$8613 ( \10495 , \10473 , \10494 );
and \U$8614 ( \10496 , \10468 , \10430 );
not \U$8615 ( \10497 , \10496 );
and \U$8616 ( \10498 , \10464 , \10497 );
xnor \U$8617 ( \10499 , \10495 , \10498 );
and \U$8618 ( \10500 , \10440 , \10499 );
and \U$8619 ( \10501 , RI2b5e785c0a00_257, \10069 );
and \U$8620 ( \10502 , RI2b5e785be390_277, \10071 );
and \U$8621 ( \10503 , RI2b5e785bc0e0_297, \10074 );
and \U$8622 ( \10504 , RI2b5e785ba1f0_317, \10077 );
and \U$8623 ( \10505 , RI2b5e785b9890_337, \10079 );
and \U$8624 ( \10506 , RI2b5e785b7d60_357, \10082 );
and \U$8625 ( \10507 , RI2b5e785b7400_377, \10084 );
and \U$8626 ( \10508 , RI2b5e785b5c90_397, \10086 );
and \U$8627 ( \10509 , RI2b5e785b5330_417, \10088 );
and \U$8628 ( \10510 , RI2b5e785b49d0_437, \10090 );
and \U$8629 ( \10511 , RI2b5e785b3620_457, \10092 );
and \U$8630 ( \10512 , RI2b5e785b2cc0_477, \10094 );
and \U$8631 ( \10513 , RI2b5e785b2360_497, \10096 );
and \U$8632 ( \10514 , RI2b5e785b1370_517, \10098 );
and \U$8633 ( \10515 , RI2b5e785b0a10_537, \10100 );
and \U$8634 ( \10516 , RI2b5e785b00b0_557, \10102 );
and \U$8635 ( \10517 , RI2b5e785af480_577, \10104 );
or \U$8636 ( \10518 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 );
_DC r3949 ( \10519_nR3949 , \10518 , \10114 );
buf \U$8637 ( \10520 , \10519_nR3949 );
xor \U$8638 ( \10521 , \9845 , \9866 );
xor \U$8639 ( \10522 , \10521 , \10003 );
buf \U$8640 ( \10523 , \10522 );
buf \U$8641 ( \10524 , \10523 );
xor \U$8642 ( \10525 , \9870 , \9891 );
xor \U$8643 ( \10526 , \10525 , \10000 );
buf \U$8644 ( \10527 , \10526 );
buf \U$8645 ( \10528 , \10527 );
xor \U$8646 ( \10529 , \10524 , \10528 );
xor \U$8647 ( \10530 , \10528 , \10464 );
not \U$8648 ( \10531 , \10530 );
and \U$8649 ( \10532 , \10529 , \10531 );
and \U$8650 ( \10533 , \10520 , \10532 );
and \U$8651 ( \10534 , RI2b5e785c2b48_256, \10069 );
and \U$8652 ( \10535 , RI2b5e785be408_276, \10071 );
and \U$8653 ( \10536 , RI2b5e785bc158_296, \10074 );
and \U$8654 ( \10537 , RI2b5e785ba268_316, \10077 );
and \U$8655 ( \10538 , RI2b5e785b9908_336, \10079 );
and \U$8656 ( \10539 , RI2b5e785b7dd8_356, \10082 );
and \U$8657 ( \10540 , RI2b5e785b7478_376, \10084 );
and \U$8658 ( \10541 , RI2b5e785b5d08_396, \10086 );
and \U$8659 ( \10542 , RI2b5e785b53a8_416, \10088 );
and \U$8660 ( \10543 , RI2b5e785b4a48_436, \10090 );
and \U$8661 ( \10544 , RI2b5e785b3698_456, \10092 );
and \U$8662 ( \10545 , RI2b5e785b2d38_476, \10094 );
and \U$8663 ( \10546 , RI2b5e785b23d8_496, \10096 );
and \U$8664 ( \10547 , RI2b5e785b13e8_516, \10098 );
and \U$8665 ( \10548 , RI2b5e785b0a88_536, \10100 );
and \U$8666 ( \10549 , RI2b5e785b0128_556, \10102 );
and \U$8667 ( \10550 , RI2b5e785af4f8_576, \10104 );
or \U$8668 ( \10551 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 );
_DC r3a20 ( \10552_nR3a20 , \10551 , \10114 );
buf \U$8669 ( \10553 , \10552_nR3a20 );
and \U$8670 ( \10554 , \10553 , \10530 );
nor \U$8671 ( \10555 , \10533 , \10554 );
and \U$8672 ( \10556 , \10528 , \10464 );
not \U$8673 ( \10557 , \10556 );
and \U$8674 ( \10558 , \10524 , \10557 );
xnor \U$8675 ( \10559 , \10555 , \10558 );
and \U$8676 ( \10560 , \10499 , \10559 );
and \U$8677 ( \10561 , \10440 , \10559 );
or \U$8678 ( \10562 , \10500 , \10560 , \10561 );
and \U$8679 ( \10563 , RI2b5e785c0910_259, \10069 );
and \U$8680 ( \10564 , RI2b5e785be2a0_279, \10071 );
and \U$8681 ( \10565 , RI2b5e785bbff0_299, \10074 );
and \U$8682 ( \10566 , RI2b5e785ba100_319, \10077 );
and \U$8683 ( \10567 , RI2b5e785b97a0_339, \10079 );
and \U$8684 ( \10568 , RI2b5e785b7c70_359, \10082 );
and \U$8685 ( \10569 , RI2b5e785b7310_379, \10084 );
and \U$8686 ( \10570 , RI2b5e785b5ba0_399, \10086 );
and \U$8687 ( \10571 , RI2b5e785b5240_419, \10088 );
and \U$8688 ( \10572 , RI2b5e785b48e0_439, \10090 );
and \U$8689 ( \10573 , RI2b5e785b3530_459, \10092 );
and \U$8690 ( \10574 , RI2b5e785b2bd0_479, \10094 );
and \U$8691 ( \10575 , RI2b5e785b2270_499, \10096 );
and \U$8692 ( \10576 , RI2b5e785b1280_519, \10098 );
and \U$8693 ( \10577 , RI2b5e785b0920_539, \10100 );
and \U$8694 ( \10578 , RI2b5e785affc0_559, \10102 );
and \U$8695 ( \10579 , RI2b5e785af390_579, \10104 );
or \U$8696 ( \10580 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 );
_DC r378a ( \10581_nR378a , \10580 , \10114 );
buf \U$8697 ( \10582 , \10581_nR378a );
xor \U$8698 ( \10583 , \9820 , \9841 );
xor \U$8699 ( \10584 , \10583 , \10006 );
buf \U$8700 ( \10585 , \10584 );
buf \U$8701 ( \10586 , \10585 );
xor \U$8702 ( \10587 , \10288 , \10586 );
xor \U$8703 ( \10588 , \10586 , \10524 );
not \U$8704 ( \10589 , \10588 );
and \U$8705 ( \10590 , \10587 , \10589 );
and \U$8706 ( \10591 , \10582 , \10590 );
and \U$8707 ( \10592 , RI2b5e785c0988_258, \10069 );
and \U$8708 ( \10593 , RI2b5e785be318_278, \10071 );
and \U$8709 ( \10594 , RI2b5e785bc068_298, \10074 );
and \U$8710 ( \10595 , RI2b5e785ba178_318, \10077 );
and \U$8711 ( \10596 , RI2b5e785b9818_338, \10079 );
and \U$8712 ( \10597 , RI2b5e785b7ce8_358, \10082 );
and \U$8713 ( \10598 , RI2b5e785b7388_378, \10084 );
and \U$8714 ( \10599 , RI2b5e785b5c18_398, \10086 );
and \U$8715 ( \10600 , RI2b5e785b52b8_418, \10088 );
and \U$8716 ( \10601 , RI2b5e785b4958_438, \10090 );
and \U$8717 ( \10602 , RI2b5e785b35a8_458, \10092 );
and \U$8718 ( \10603 , RI2b5e785b2c48_478, \10094 );
and \U$8719 ( \10604 , RI2b5e785b22e8_498, \10096 );
and \U$8720 ( \10605 , RI2b5e785b12f8_518, \10098 );
and \U$8721 ( \10606 , RI2b5e785b0998_538, \10100 );
and \U$8722 ( \10607 , RI2b5e785b0038_558, \10102 );
and \U$8723 ( \10608 , RI2b5e785af408_578, \10104 );
or \U$8724 ( \10609 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 );
_DC r3853 ( \10610_nR3853 , \10609 , \10114 );
buf \U$8725 ( \10611 , \10610_nR3853 );
and \U$8726 ( \10612 , \10611 , \10588 );
nor \U$8727 ( \10613 , \10591 , \10612 );
and \U$8728 ( \10614 , \10586 , \10524 );
not \U$8729 ( \10615 , \10614 );
and \U$8730 ( \10616 , \10288 , \10615 );
xnor \U$8731 ( \10617 , \10613 , \10616 );
and \U$8732 ( \10618 , RI2b5e785c0820_261, \10069 );
and \U$8733 ( \10619 , RI2b5e785be1b0_281, \10071 );
and \U$8734 ( \10620 , RI2b5e785bbf00_301, \10074 );
and \U$8735 ( \10621 , RI2b5e785ba010_321, \10077 );
and \U$8736 ( \10622 , RI2b5e785b96b0_341, \10079 );
and \U$8737 ( \10623 , RI2b5e785b7b80_361, \10082 );
and \U$8738 ( \10624 , RI2b5e785b7220_381, \10084 );
and \U$8739 ( \10625 , RI2b5e785b5ab0_401, \10086 );
and \U$8740 ( \10626 , RI2b5e785b5150_421, \10088 );
and \U$8741 ( \10627 , RI2b5e785b47f0_441, \10090 );
and \U$8742 ( \10628 , RI2b5e785b3440_461, \10092 );
and \U$8743 ( \10629 , RI2b5e785b2ae0_481, \10094 );
and \U$8744 ( \10630 , RI2b5e785b2180_501, \10096 );
and \U$8745 ( \10631 , RI2b5e785b1190_521, \10098 );
and \U$8746 ( \10632 , RI2b5e785b0830_541, \10100 );
and \U$8747 ( \10633 , RI2b5e785afed0_561, \10102 );
and \U$8748 ( \10634 , RI2b5e785af2a0_581, \10104 );
or \U$8749 ( \10635 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 );
_DC r35f1 ( \10636_nR35f1 , \10635 , \10114 );
buf \U$8750 ( \10637 , \10636_nR35f1 );
and \U$8751 ( \10638 , \10637 , \10291 );
and \U$8752 ( \10639 , RI2b5e785c0898_260, \10069 );
and \U$8753 ( \10640 , RI2b5e785be228_280, \10071 );
and \U$8754 ( \10641 , RI2b5e785bbf78_300, \10074 );
and \U$8755 ( \10642 , RI2b5e785ba088_320, \10077 );
and \U$8756 ( \10643 , RI2b5e785b9728_340, \10079 );
and \U$8757 ( \10644 , RI2b5e785b7bf8_360, \10082 );
and \U$8758 ( \10645 , RI2b5e785b7298_380, \10084 );
and \U$8759 ( \10646 , RI2b5e785b5b28_400, \10086 );
and \U$8760 ( \10647 , RI2b5e785b51c8_420, \10088 );
and \U$8761 ( \10648 , RI2b5e785b4868_440, \10090 );
and \U$8762 ( \10649 , RI2b5e785b34b8_460, \10092 );
and \U$8763 ( \10650 , RI2b5e785b2b58_480, \10094 );
and \U$8764 ( \10651 , RI2b5e785b21f8_500, \10096 );
and \U$8765 ( \10652 , RI2b5e785b1208_520, \10098 );
and \U$8766 ( \10653 , RI2b5e785b08a8_540, \10100 );
and \U$8767 ( \10654 , RI2b5e785aff48_560, \10102 );
and \U$8768 ( \10655 , RI2b5e785af318_580, \10104 );
or \U$8769 ( \10656 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 );
_DC r36a4 ( \10657_nR36a4 , \10656 , \10114 );
buf \U$8770 ( \10658 , \10657_nR36a4 );
and \U$8771 ( \10659 , \10658 , \10289 );
nor \U$8772 ( \10660 , \10638 , \10659 );
xnor \U$8773 ( \10661 , \10660 , \10296 );
and \U$8774 ( \10662 , \10617 , \10661 );
and \U$8775 ( \10663 , RI2b5e785c0730_263, \10069 );
and \U$8776 ( \10664 , RI2b5e785be0c0_283, \10071 );
and \U$8777 ( \10665 , RI2b5e785bbe10_303, \10074 );
and \U$8778 ( \10666 , RI2b5e785b9f20_323, \10077 );
and \U$8779 ( \10667 , RI2b5e785b95c0_343, \10079 );
and \U$8780 ( \10668 , RI2b5e785b7a90_363, \10082 );
and \U$8781 ( \10669 , RI2b5e785b7130_383, \10084 );
and \U$8782 ( \10670 , RI2b5e785b59c0_403, \10086 );
and \U$8783 ( \10671 , RI2b5e785b5060_423, \10088 );
and \U$8784 ( \10672 , RI2b5e785b3cb0_443, \10090 );
and \U$8785 ( \10673 , RI2b5e785b3350_463, \10092 );
and \U$8786 ( \10674 , RI2b5e785b29f0_483, \10094 );
and \U$8787 ( \10675 , RI2b5e785b1a00_503, \10096 );
and \U$8788 ( \10676 , RI2b5e785b10a0_523, \10098 );
and \U$8789 ( \10677 , RI2b5e785b0740_543, \10100 );
and \U$8790 ( \10678 , RI2b5e785afde0_563, \10102 );
and \U$8791 ( \10679 , RI2b5e785af1b0_583, \10104 );
or \U$8792 ( \10680 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 );
_DC r348d ( \10681_nR348d , \10680 , \10114 );
buf \U$8793 ( \10682 , \10681_nR348d );
and \U$8794 ( \10683 , \10682 , \10226 );
and \U$8795 ( \10684 , RI2b5e785c07a8_262, \10069 );
and \U$8796 ( \10685 , RI2b5e785be138_282, \10071 );
and \U$8797 ( \10686 , RI2b5e785bbe88_302, \10074 );
and \U$8798 ( \10687 , RI2b5e785b9f98_322, \10077 );
and \U$8799 ( \10688 , RI2b5e785b9638_342, \10079 );
and \U$8800 ( \10689 , RI2b5e785b7b08_362, \10082 );
and \U$8801 ( \10690 , RI2b5e785b71a8_382, \10084 );
and \U$8802 ( \10691 , RI2b5e785b5a38_402, \10086 );
and \U$8803 ( \10692 , RI2b5e785b50d8_422, \10088 );
and \U$8804 ( \10693 , RI2b5e785b4778_442, \10090 );
and \U$8805 ( \10694 , RI2b5e785b33c8_462, \10092 );
and \U$8806 ( \10695 , RI2b5e785b2a68_482, \10094 );
and \U$8807 ( \10696 , RI2b5e785b1a78_502, \10096 );
and \U$8808 ( \10697 , RI2b5e785b1118_522, \10098 );
and \U$8809 ( \10698 , RI2b5e785b07b8_542, \10100 );
and \U$8810 ( \10699 , RI2b5e785afe58_562, \10102 );
and \U$8811 ( \10700 , RI2b5e785af228_582, \10104 );
or \U$8812 ( \10701 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 );
_DC r3534 ( \10702_nR3534 , \10701 , \10114 );
buf \U$8813 ( \10703 , \10702_nR3534 );
and \U$8814 ( \10704 , \10703 , \10224 );
nor \U$8815 ( \10705 , \10683 , \10704 );
xnor \U$8816 ( \10706 , \10705 , \10035 );
and \U$8817 ( \10707 , \10661 , \10706 );
and \U$8818 ( \10708 , \10617 , \10706 );
or \U$8819 ( \10709 , \10662 , \10707 , \10708 );
and \U$8820 ( \10710 , \10562 , \10709 );
and \U$8821 ( \10711 , RI2b5e785c0640_265, \10069 );
and \U$8822 ( \10712 , RI2b5e785bdfd0_285, \10071 );
and \U$8823 ( \10713 , RI2b5e785bbd20_305, \10074 );
and \U$8824 ( \10714 , RI2b5e785b9e30_325, \10077 );
and \U$8825 ( \10715 , RI2b5e785b94d0_345, \10079 );
and \U$8826 ( \10716 , RI2b5e785b79a0_365, \10082 );
and \U$8827 ( \10717 , RI2b5e785b7040_385, \10084 );
and \U$8828 ( \10718 , RI2b5e785b58d0_405, \10086 );
and \U$8829 ( \10719 , RI2b5e785b4f70_425, \10088 );
and \U$8830 ( \10720 , RI2b5e785b3bc0_445, \10090 );
and \U$8831 ( \10721 , RI2b5e785b3260_465, \10092 );
and \U$8832 ( \10722 , RI2b5e785b2900_485, \10094 );
and \U$8833 ( \10723 , RI2b5e785b1910_505, \10096 );
and \U$8834 ( \10724 , RI2b5e785b0fb0_525, \10098 );
and \U$8835 ( \10725 , RI2b5e785b0650_545, \10100 );
and \U$8836 ( \10726 , RI2b5e785afcf0_565, \10102 );
and \U$8837 ( \10727 , RI2b5e785af0c0_585, \10104 );
or \U$8838 ( \10728 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 );
_DC r331d ( \10729_nR331d , \10728 , \10114 );
buf \U$8839 ( \10730 , \10729_nR331d );
and \U$8840 ( \10731 , \10730 , \10164 );
and \U$8841 ( \10732 , RI2b5e785c06b8_264, \10069 );
and \U$8842 ( \10733 , RI2b5e785be048_284, \10071 );
and \U$8843 ( \10734 , RI2b5e785bbd98_304, \10074 );
and \U$8844 ( \10735 , RI2b5e785b9ea8_324, \10077 );
and \U$8845 ( \10736 , RI2b5e785b9548_344, \10079 );
and \U$8846 ( \10737 , RI2b5e785b7a18_364, \10082 );
and \U$8847 ( \10738 , RI2b5e785b70b8_384, \10084 );
and \U$8848 ( \10739 , RI2b5e785b5948_404, \10086 );
and \U$8849 ( \10740 , RI2b5e785b4fe8_424, \10088 );
and \U$8850 ( \10741 , RI2b5e785b3c38_444, \10090 );
and \U$8851 ( \10742 , RI2b5e785b32d8_464, \10092 );
and \U$8852 ( \10743 , RI2b5e785b2978_484, \10094 );
and \U$8853 ( \10744 , RI2b5e785b1988_504, \10096 );
and \U$8854 ( \10745 , RI2b5e785b1028_524, \10098 );
and \U$8855 ( \10746 , RI2b5e785b06c8_544, \10100 );
and \U$8856 ( \10747 , RI2b5e785afd68_564, \10102 );
and \U$8857 ( \10748 , RI2b5e785af138_584, \10104 );
or \U$8858 ( \10749 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 );
_DC r33ee ( \10750_nR33ee , \10749 , \10114 );
buf \U$8859 ( \10751 , \10750_nR33ee );
and \U$8860 ( \10752 , \10751 , \10162 );
nor \U$8861 ( \10753 , \10731 , \10752 );
xnor \U$8862 ( \10754 , \10753 , \10190 );
and \U$8864 ( \10755 , RI2b5e785c05c8_266, \10069 );
and \U$8865 ( \10756 , RI2b5e785bdf58_286, \10071 );
and \U$8866 ( \10757 , RI2b5e785bbca8_306, \10074 );
and \U$8867 ( \10758 , RI2b5e785b9db8_326, \10077 );
and \U$8868 ( \10759 , RI2b5e785b9458_346, \10079 );
and \U$8869 ( \10760 , RI2b5e785b7928_366, \10082 );
and \U$8870 ( \10761 , RI2b5e785b6fc8_386, \10084 );
and \U$8871 ( \10762 , RI2b5e785b5858_406, \10086 );
and \U$8872 ( \10763 , RI2b5e785b4ef8_426, \10088 );
and \U$8873 ( \10764 , RI2b5e785b3b48_446, \10090 );
and \U$8874 ( \10765 , RI2b5e785b31e8_466, \10092 );
and \U$8875 ( \10766 , RI2b5e785b2888_486, \10094 );
and \U$8876 ( \10767 , RI2b5e785b1898_506, \10096 );
and \U$8877 ( \10768 , RI2b5e785b0f38_526, \10098 );
and \U$8878 ( \10769 , RI2b5e785b05d8_546, \10100 );
and \U$8879 ( \10770 , RI2b5e785afc78_566, \10102 );
and \U$8880 ( \10771 , RI2b5e785af048_586, \10104 );
or \U$8881 ( \10772 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 );
_DC r32db ( \10773_nR32db , \10772 , \10114 );
buf \U$8882 ( \10774 , \10773_nR32db );
and \U$8883 ( \10775 , \10774 , \10217 );
nor \U$8884 ( \10776 , 1'b0 , \10775 );
xnor \U$8885 ( \10777 , \10776 , 1'b0 );
and \U$8886 ( \10778 , \10754 , \10777 );
and \U$8887 ( \10779 , \10709 , \10778 );
and \U$8888 ( \10780 , \10562 , \10778 );
or \U$8889 ( \10781 , \10710 , \10779 , \10780 );
and \U$8891 ( \10782 , \10703 , \10226 );
and \U$8892 ( \10783 , \10637 , \10224 );
nor \U$8893 ( \10784 , \10782 , \10783 );
xnor \U$8894 ( \10785 , \10784 , \10035 );
and \U$8895 ( \10786 , \10751 , \10164 );
and \U$8896 ( \10787 , \10682 , \10162 );
nor \U$8897 ( \10788 , \10786 , \10787 );
xnor \U$8898 ( \10789 , \10788 , \10190 );
xor \U$8899 ( \10790 , \10785 , \10789 );
and \U$8901 ( \10791 , \10730 , \10217 );
nor \U$8902 ( \10792 , 1'b0 , \10791 );
xnor \U$8903 ( \10793 , \10792 , 1'b0 );
xor \U$8904 ( \10794 , \10790 , \10793 );
and \U$8905 ( \10795 , \10553 , \10532 );
and \U$8906 ( \10796 , \10460 , \10530 );
nor \U$8907 ( \10797 , \10795 , \10796 );
xnor \U$8908 ( \10798 , \10797 , \10558 );
and \U$8909 ( \10799 , \10611 , \10590 );
and \U$8910 ( \10800 , \10520 , \10588 );
nor \U$8911 ( \10801 , \10799 , \10800 );
xnor \U$8912 ( \10802 , \10801 , \10616 );
xor \U$8913 ( \10803 , \10798 , \10802 );
and \U$8914 ( \10804 , \10658 , \10291 );
and \U$8915 ( \10805 , \10582 , \10289 );
nor \U$8916 ( \10806 , \10804 , \10805 );
xnor \U$8917 ( \10807 , \10806 , \10296 );
xor \U$8918 ( \10808 , \10803 , \10807 );
and \U$8919 ( \10809 , \10794 , \10808 );
or \U$8921 ( \10810 , 1'b0 , \10809 , 1'b0 );
xor \U$8922 ( \10811 , \10781 , \10810 );
and \U$8923 ( \10812 , \10682 , \10164 );
and \U$8924 ( \10813 , \10703 , \10162 );
nor \U$8925 ( \10814 , \10812 , \10813 );
xnor \U$8926 ( \10815 , \10814 , \10190 );
and \U$8928 ( \10816 , \10751 , \10217 );
nor \U$8929 ( \10817 , 1'b0 , \10816 );
xnor \U$8930 ( \10818 , \10817 , 1'b0 );
xor \U$8931 ( \10819 , \10815 , \10818 );
xor \U$8933 ( \10820 , \10819 , 1'b0 );
and \U$8934 ( \10821 , \10520 , \10590 );
and \U$8935 ( \10822 , \10553 , \10588 );
nor \U$8936 ( \10823 , \10821 , \10822 );
xnor \U$8937 ( \10824 , \10823 , \10616 );
and \U$8938 ( \10825 , \10582 , \10291 );
and \U$8939 ( \10826 , \10611 , \10289 );
nor \U$8940 ( \10827 , \10825 , \10826 );
xnor \U$8941 ( \10828 , \10827 , \10296 );
xor \U$8942 ( \10829 , \10824 , \10828 );
and \U$8943 ( \10830 , \10637 , \10226 );
and \U$8944 ( \10831 , \10658 , \10224 );
nor \U$8945 ( \10832 , \10830 , \10831 );
xnor \U$8946 ( \10833 , \10832 , \10035 );
xor \U$8947 ( \10834 , \10829 , \10833 );
xor \U$8948 ( \10835 , \10820 , \10834 );
and \U$8949 ( \10836 , \10344 , \10436 );
and \U$8950 ( \10837 , \10212 , \10433 );
nor \U$8951 ( \10838 , \10836 , \10837 );
xnor \U$8952 ( \10839 , \10838 , \10430 );
and \U$8953 ( \10840 , \10367 , \10472 );
and \U$8954 ( \10841 , \10323 , \10470 );
nor \U$8955 ( \10842 , \10840 , \10841 );
xnor \U$8956 ( \10843 , \10842 , \10498 );
xor \U$8957 ( \10844 , \10839 , \10843 );
and \U$8958 ( \10845 , \10460 , \10532 );
and \U$8959 ( \10846 , \10493 , \10530 );
nor \U$8960 ( \10847 , \10845 , \10846 );
xnor \U$8961 ( \10848 , \10847 , \10558 );
xor \U$8962 ( \10849 , \10844 , \10848 );
xor \U$8963 ( \10850 , \10835 , \10849 );
xor \U$8964 ( \10851 , \10811 , \10850 );
and \U$8966 ( \10852 , \10493 , \10436 );
and \U$8967 ( \10853 , \10367 , \10433 );
nor \U$8968 ( \10854 , \10852 , \10853 );
xnor \U$8969 ( \10855 , \10854 , \10430 );
and \U$8970 ( \10856 , \10553 , \10472 );
and \U$8971 ( \10857 , \10460 , \10470 );
nor \U$8972 ( \10858 , \10856 , \10857 );
xnor \U$8973 ( \10859 , \10858 , \10498 );
and \U$8974 ( \10860 , \10855 , \10859 );
or \U$8976 ( \10861 , 1'b0 , \10860 , 1'b0 );
and \U$8977 ( \10862 , \10611 , \10532 );
and \U$8978 ( \10863 , \10520 , \10530 );
nor \U$8979 ( \10864 , \10862 , \10863 );
xnor \U$8980 ( \10865 , \10864 , \10558 );
and \U$8981 ( \10866 , \10658 , \10590 );
and \U$8982 ( \10867 , \10582 , \10588 );
nor \U$8983 ( \10868 , \10866 , \10867 );
xnor \U$8984 ( \10869 , \10868 , \10616 );
and \U$8985 ( \10870 , \10865 , \10869 );
and \U$8986 ( \10871 , \10703 , \10291 );
and \U$8987 ( \10872 , \10637 , \10289 );
nor \U$8988 ( \10873 , \10871 , \10872 );
xnor \U$8989 ( \10874 , \10873 , \10296 );
and \U$8990 ( \10875 , \10869 , \10874 );
and \U$8991 ( \10876 , \10865 , \10874 );
or \U$8992 ( \10877 , \10870 , \10875 , \10876 );
and \U$8993 ( \10878 , \10861 , \10877 );
and \U$8994 ( \10879 , \10751 , \10226 );
and \U$8995 ( \10880 , \10682 , \10224 );
nor \U$8996 ( \10881 , \10879 , \10880 );
xnor \U$8997 ( \10882 , \10881 , \10035 );
and \U$8998 ( \10883 , \10774 , \10164 );
and \U$8999 ( \10884 , \10730 , \10162 );
nor \U$9000 ( \10885 , \10883 , \10884 );
xnor \U$9001 ( \10886 , \10885 , \10190 );
and \U$9002 ( \10887 , \10882 , \10886 );
and \U$9003 ( \10888 , RI2b5e785c0550_267, \10069 );
and \U$9004 ( \10889 , RI2b5e785bc590_287, \10071 );
and \U$9005 ( \10890 , RI2b5e785bbc30_307, \10074 );
and \U$9006 ( \10891 , RI2b5e785b9d40_327, \10077 );
and \U$9007 ( \10892 , RI2b5e785b93e0_347, \10079 );
and \U$9008 ( \10893 , RI2b5e785b78b0_367, \10082 );
and \U$9009 ( \10894 , RI2b5e785b6f50_387, \10084 );
and \U$9010 ( \10895 , RI2b5e785b57e0_407, \10086 );
and \U$9011 ( \10896 , RI2b5e785b4e80_427, \10088 );
and \U$9012 ( \10897 , RI2b5e785b3ad0_447, \10090 );
and \U$9013 ( \10898 , RI2b5e785b3170_467, \10092 );
and \U$9014 ( \10899 , RI2b5e785b2810_487, \10094 );
and \U$9015 ( \10900 , RI2b5e785b1820_507, \10096 );
and \U$9016 ( \10901 , RI2b5e785b0ec0_527, \10098 );
and \U$9017 ( \10902 , RI2b5e785b0560_547, \10100 );
and \U$9018 ( \10903 , RI2b5e785afc00_567, \10102 );
and \U$9019 ( \10904 , RI2b5e785aefd0_587, \10104 );
or \U$9020 ( \10905 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 );
_DC r31e3 ( \10906_nR31e3 , \10905 , \10114 );
buf \U$9021 ( \10907 , \10906_nR31e3 );
nand \U$9022 ( \10908 , \10907 , \10217 );
xnor \U$9023 ( \10909 , \10908 , 1'b0 );
and \U$9024 ( \10910 , \10886 , \10909 );
and \U$9025 ( \10911 , \10882 , \10909 );
or \U$9026 ( \10912 , \10887 , \10910 , \10911 );
and \U$9027 ( \10913 , \10877 , \10912 );
and \U$9028 ( \10914 , \10861 , \10912 );
or \U$9029 ( \10915 , \10878 , \10913 , \10914 );
xor \U$9030 ( \10916 , \10754 , \10777 );
xor \U$9031 ( \10917 , \10617 , \10661 );
xor \U$9032 ( \10918 , \10917 , \10706 );
and \U$9033 ( \10919 , \10916 , \10918 );
xor \U$9034 ( \10920 , \10440 , \10499 );
xor \U$9035 ( \10921 , \10920 , \10559 );
and \U$9036 ( \10922 , \10918 , \10921 );
and \U$9037 ( \10923 , \10916 , \10921 );
or \U$9038 ( \10924 , \10919 , \10922 , \10923 );
and \U$9039 ( \10925 , \10915 , \10924 );
and \U$9041 ( \10926 , \10323 , \10436 );
and \U$9042 ( \10927 , \10344 , \10433 );
nor \U$9043 ( \10928 , \10926 , \10927 );
xnor \U$9044 ( \10929 , \10928 , \10430 );
xor \U$9045 ( \10930 , 1'b0 , \10929 );
and \U$9046 ( \10931 , \10493 , \10472 );
and \U$9047 ( \10932 , \10367 , \10470 );
nor \U$9048 ( \10933 , \10931 , \10932 );
xnor \U$9049 ( \10934 , \10933 , \10498 );
xor \U$9050 ( \10935 , \10930 , \10934 );
and \U$9051 ( \10936 , \10924 , \10935 );
and \U$9052 ( \10937 , \10915 , \10935 );
or \U$9053 ( \10938 , \10925 , \10936 , \10937 );
xor \U$9055 ( \10939 , 1'b0 , \10794 );
xor \U$9056 ( \10940 , \10939 , \10808 );
xor \U$9057 ( \10941 , \10562 , \10709 );
xor \U$9058 ( \10942 , \10941 , \10778 );
and \U$9059 ( \10943 , \10940 , \10942 );
xor \U$9060 ( \10944 , \10938 , \10943 );
and \U$9062 ( \10945 , \10929 , \10934 );
or \U$9064 ( \10946 , 1'b0 , \10945 , 1'b0 );
and \U$9065 ( \10947 , \10798 , \10802 );
and \U$9066 ( \10948 , \10802 , \10807 );
and \U$9067 ( \10949 , \10798 , \10807 );
or \U$9068 ( \10950 , \10947 , \10948 , \10949 );
xor \U$9069 ( \10951 , \10946 , \10950 );
and \U$9070 ( \10952 , \10785 , \10789 );
and \U$9071 ( \10953 , \10789 , \10793 );
and \U$9072 ( \10954 , \10785 , \10793 );
or \U$9073 ( \10955 , \10952 , \10953 , \10954 );
xor \U$9074 ( \10956 , \10951 , \10955 );
xor \U$9075 ( \10957 , \10944 , \10956 );
xor \U$9076 ( \10958 , \10851 , \10957 );
and \U$9077 ( \10959 , \10460 , \10436 );
and \U$9078 ( \10960 , \10493 , \10433 );
nor \U$9079 ( \10961 , \10959 , \10960 );
xnor \U$9080 ( \10962 , \10961 , \10430 );
and \U$9081 ( \10963 , \10520 , \10472 );
and \U$9082 ( \10964 , \10553 , \10470 );
nor \U$9083 ( \10965 , \10963 , \10964 );
xnor \U$9084 ( \10966 , \10965 , \10498 );
and \U$9085 ( \10967 , \10962 , \10966 );
and \U$9086 ( \10968 , \10582 , \10532 );
and \U$9087 ( \10969 , \10611 , \10530 );
nor \U$9088 ( \10970 , \10968 , \10969 );
xnor \U$9089 ( \10971 , \10970 , \10558 );
and \U$9090 ( \10972 , \10966 , \10971 );
and \U$9091 ( \10973 , \10962 , \10971 );
or \U$9092 ( \10974 , \10967 , \10972 , \10973 );
and \U$9093 ( \10975 , \10637 , \10590 );
and \U$9094 ( \10976 , \10658 , \10588 );
nor \U$9095 ( \10977 , \10975 , \10976 );
xnor \U$9096 ( \10978 , \10977 , \10616 );
and \U$9097 ( \10979 , \10682 , \10291 );
and \U$9098 ( \10980 , \10703 , \10289 );
nor \U$9099 ( \10981 , \10979 , \10980 );
xnor \U$9100 ( \10982 , \10981 , \10296 );
and \U$9101 ( \10983 , \10978 , \10982 );
and \U$9102 ( \10984 , \10730 , \10226 );
and \U$9103 ( \10985 , \10751 , \10224 );
nor \U$9104 ( \10986 , \10984 , \10985 );
xnor \U$9105 ( \10987 , \10986 , \10035 );
and \U$9106 ( \10988 , \10982 , \10987 );
and \U$9107 ( \10989 , \10978 , \10987 );
or \U$9108 ( \10990 , \10983 , \10988 , \10989 );
and \U$9109 ( \10991 , \10974 , \10990 );
xor \U$9110 ( \10992 , \10882 , \10886 );
xor \U$9111 ( \10993 , \10992 , \10909 );
and \U$9112 ( \10994 , \10990 , \10993 );
and \U$9113 ( \10995 , \10974 , \10993 );
or \U$9114 ( \10996 , \10991 , \10994 , \10995 );
xor \U$9115 ( \10997 , \10865 , \10869 );
xor \U$9116 ( \10998 , \10997 , \10874 );
xor \U$9117 ( \10999 , 1'b0 , \10855 );
xor \U$9118 ( \11000 , \10999 , \10859 );
and \U$9119 ( \11001 , \10998 , \11000 );
and \U$9120 ( \11002 , \10996 , \11001 );
xor \U$9121 ( \11003 , \10916 , \10918 );
xor \U$9122 ( \11004 , \11003 , \10921 );
and \U$9123 ( \11005 , \11001 , \11004 );
and \U$9124 ( \11006 , \10996 , \11004 );
or \U$9125 ( \11007 , \11002 , \11005 , \11006 );
xor \U$9126 ( \11008 , \10940 , \10942 );
and \U$9127 ( \11009 , \11007 , \11008 );
xor \U$9128 ( \11010 , \10915 , \10924 );
xor \U$9129 ( \11011 , \11010 , \10935 );
and \U$9130 ( \11012 , \11008 , \11011 );
and \U$9131 ( \11013 , \11007 , \11011 );
or \U$9132 ( \11014 , \11009 , \11012 , \11013 );
nor \U$9133 ( \11015 , \10958 , \11014 );
and \U$9134 ( \11016 , \10938 , \10943 );
and \U$9135 ( \11017 , \10943 , \10956 );
and \U$9136 ( \11018 , \10938 , \10956 );
or \U$9137 ( \11019 , \11016 , \11017 , \11018 );
and \U$9138 ( \11020 , \10781 , \10810 );
and \U$9139 ( \11021 , \10810 , \10850 );
and \U$9140 ( \11022 , \10781 , \10850 );
or \U$9141 ( \11023 , \11020 , \11021 , \11022 );
and \U$9143 ( \11024 , \10212 , \10436 );
and \U$9144 ( \11025 , \10116 , \10433 );
nor \U$9145 ( \11026 , \11024 , \11025 );
xnor \U$9146 ( \11027 , \11026 , \10430 );
xor \U$9147 ( \11028 , 1'b0 , \11027 );
and \U$9148 ( \11029 , \10323 , \10472 );
and \U$9149 ( \11030 , \10344 , \10470 );
nor \U$9150 ( \11031 , \11029 , \11030 );
xnor \U$9151 ( \11032 , \11031 , \10498 );
xor \U$9152 ( \11033 , \11028 , \11032 );
and \U$9154 ( \11034 , \10658 , \10226 );
and \U$9155 ( \11035 , \10582 , \10224 );
nor \U$9156 ( \11036 , \11034 , \11035 );
xnor \U$9157 ( \11037 , \11036 , \10035 );
and \U$9158 ( \11038 , \10703 , \10164 );
and \U$9159 ( \11039 , \10637 , \10162 );
nor \U$9160 ( \11040 , \11038 , \11039 );
xnor \U$9161 ( \11041 , \11040 , \10190 );
xor \U$9162 ( \11042 , \11037 , \11041 );
and \U$9164 ( \11043 , \10682 , \10217 );
nor \U$9165 ( \11044 , 1'b0 , \11043 );
xnor \U$9166 ( \11045 , \11044 , 1'b0 );
xor \U$9167 ( \11046 , \11042 , \11045 );
xor \U$9168 ( \11047 , 1'b0 , \11046 );
xor \U$9169 ( \11048 , \11033 , \11047 );
and \U$9170 ( \11049 , \10839 , \10843 );
and \U$9171 ( \11050 , \10843 , \10848 );
and \U$9172 ( \11051 , \10839 , \10848 );
or \U$9173 ( \11052 , \11049 , \11050 , \11051 );
and \U$9174 ( \11053 , \10824 , \10828 );
and \U$9175 ( \11054 , \10828 , \10833 );
and \U$9176 ( \11055 , \10824 , \10833 );
or \U$9177 ( \11056 , \11053 , \11054 , \11055 );
xor \U$9178 ( \11057 , \11052 , \11056 );
and \U$9179 ( \11058 , \10815 , \10818 );
or \U$9182 ( \11059 , \11058 , 1'b0 , 1'b0 );
xor \U$9183 ( \11060 , \11057 , \11059 );
xor \U$9184 ( \11061 , \11048 , \11060 );
xor \U$9185 ( \11062 , \11023 , \11061 );
and \U$9186 ( \11063 , \10946 , \10950 );
and \U$9187 ( \11064 , \10950 , \10955 );
and \U$9188 ( \11065 , \10946 , \10955 );
or \U$9189 ( \11066 , \11063 , \11064 , \11065 );
and \U$9190 ( \11067 , \10820 , \10834 );
and \U$9191 ( \11068 , \10834 , \10849 );
and \U$9192 ( \11069 , \10820 , \10849 );
or \U$9193 ( \11070 , \11067 , \11068 , \11069 );
xor \U$9194 ( \11071 , \11066 , \11070 );
and \U$9195 ( \11072 , \10493 , \10532 );
and \U$9196 ( \11073 , \10367 , \10530 );
nor \U$9197 ( \11074 , \11072 , \11073 );
xnor \U$9198 ( \11075 , \11074 , \10558 );
and \U$9199 ( \11076 , \10553 , \10590 );
and \U$9200 ( \11077 , \10460 , \10588 );
nor \U$9201 ( \11078 , \11076 , \11077 );
xnor \U$9202 ( \11079 , \11078 , \10616 );
xor \U$9203 ( \11080 , \11075 , \11079 );
and \U$9204 ( \11081 , \10611 , \10291 );
and \U$9205 ( \11082 , \10520 , \10289 );
nor \U$9206 ( \11083 , \11081 , \11082 );
xnor \U$9207 ( \11084 , \11083 , \10296 );
xor \U$9208 ( \11085 , \11080 , \11084 );
xor \U$9209 ( \11086 , \11071 , \11085 );
xor \U$9210 ( \11087 , \11062 , \11086 );
xor \U$9211 ( \11088 , \11019 , \11087 );
and \U$9212 ( \11089 , \10851 , \10957 );
nor \U$9213 ( \11090 , \11088 , \11089 );
nor \U$9214 ( \11091 , \11015 , \11090 );
and \U$9215 ( \11092 , \11023 , \11061 );
and \U$9216 ( \11093 , \11061 , \11086 );
and \U$9217 ( \11094 , \11023 , \11086 );
or \U$9218 ( \11095 , \11092 , \11093 , \11094 );
and \U$9220 ( \11096 , \11027 , \11032 );
or \U$9222 ( \11097 , 1'b0 , \11096 , 1'b0 );
and \U$9223 ( \11098 , \11075 , \11079 );
and \U$9224 ( \11099 , \11079 , \11084 );
and \U$9225 ( \11100 , \11075 , \11084 );
or \U$9226 ( \11101 , \11098 , \11099 , \11100 );
xor \U$9227 ( \11102 , \11097 , \11101 );
and \U$9228 ( \11103 , \11037 , \11041 );
and \U$9229 ( \11104 , \11041 , \11045 );
and \U$9230 ( \11105 , \11037 , \11045 );
or \U$9231 ( \11106 , \11103 , \11104 , \11105 );
xor \U$9232 ( \11107 , \11102 , \11106 );
and \U$9233 ( \11108 , \11052 , \11056 );
and \U$9234 ( \11109 , \11056 , \11059 );
and \U$9235 ( \11110 , \11052 , \11059 );
or \U$9236 ( \11111 , \11108 , \11109 , \11110 );
xor \U$9238 ( \11112 , \11111 , 1'b0 );
and \U$9239 ( \11113 , \10116 , \10436 );
and \U$9240 ( \11114 , \10185 , \10433 );
nor \U$9241 ( \11115 , \11113 , \11114 );
xnor \U$9242 ( \11116 , \11115 , \10430 );
and \U$9243 ( \11117 , \10344 , \10472 );
and \U$9244 ( \11118 , \10212 , \10470 );
nor \U$9245 ( \11119 , \11117 , \11118 );
xnor \U$9246 ( \11120 , \11119 , \10498 );
xor \U$9247 ( \11121 , \11116 , \11120 );
and \U$9248 ( \11122 , \10367 , \10532 );
and \U$9249 ( \11123 , \10323 , \10530 );
nor \U$9250 ( \11124 , \11122 , \11123 );
xnor \U$9251 ( \11125 , \11124 , \10558 );
xor \U$9252 ( \11126 , \11121 , \11125 );
xor \U$9253 ( \11127 , \11112 , \11126 );
xor \U$9254 ( \11128 , \11107 , \11127 );
xor \U$9255 ( \11129 , \11095 , \11128 );
and \U$9256 ( \11130 , \11066 , \11070 );
and \U$9257 ( \11131 , \11070 , \11085 );
and \U$9258 ( \11132 , \11066 , \11085 );
or \U$9259 ( \11133 , \11130 , \11131 , \11132 );
and \U$9260 ( \11134 , \11033 , \11047 );
and \U$9261 ( \11135 , \11047 , \11060 );
and \U$9262 ( \11136 , \11033 , \11060 );
or \U$9263 ( \11137 , \11134 , \11135 , \11136 );
xor \U$9264 ( \11138 , \11133 , \11137 );
and \U$9266 ( \11139 , \10637 , \10164 );
and \U$9267 ( \11140 , \10658 , \10162 );
nor \U$9268 ( \11141 , \11139 , \11140 );
xnor \U$9269 ( \11142 , \11141 , \10190 );
and \U$9271 ( \11143 , \10703 , \10217 );
nor \U$9272 ( \11144 , 1'b0 , \11143 );
xnor \U$9273 ( \11145 , \11144 , 1'b0 );
xor \U$9274 ( \11146 , \11142 , \11145 );
xor \U$9276 ( \11147 , \11146 , 1'b0 );
xor \U$9277 ( \11148 , 1'b0 , \11147 );
and \U$9278 ( \11149 , \10460 , \10590 );
and \U$9279 ( \11150 , \10493 , \10588 );
nor \U$9280 ( \11151 , \11149 , \11150 );
xnor \U$9281 ( \11152 , \11151 , \10616 );
and \U$9282 ( \11153 , \10520 , \10291 );
and \U$9283 ( \11154 , \10553 , \10289 );
nor \U$9284 ( \11155 , \11153 , \11154 );
xnor \U$9285 ( \11156 , \11155 , \10296 );
xor \U$9286 ( \11157 , \11152 , \11156 );
and \U$9287 ( \11158 , \10582 , \10226 );
and \U$9288 ( \11159 , \10611 , \10224 );
nor \U$9289 ( \11160 , \11158 , \11159 );
xnor \U$9290 ( \11161 , \11160 , \10035 );
xor \U$9291 ( \11162 , \11157 , \11161 );
xor \U$9292 ( \11163 , \11148 , \11162 );
xor \U$9293 ( \11164 , \11138 , \11163 );
xor \U$9294 ( \11165 , \11129 , \11164 );
and \U$9295 ( \11166 , \11019 , \11087 );
nor \U$9296 ( \11167 , \11165 , \11166 );
and \U$9297 ( \11168 , \11133 , \11137 );
and \U$9298 ( \11169 , \11137 , \11163 );
and \U$9299 ( \11170 , \11133 , \11163 );
or \U$9300 ( \11171 , \11168 , \11169 , \11170 );
and \U$9301 ( \11172 , \11107 , \11127 );
xor \U$9302 ( \11173 , \11171 , \11172 );
and \U$9305 ( \11174 , \11111 , \11126 );
or \U$9306 ( \11175 , 1'b0 , 1'b0 , \11174 );
and \U$9308 ( \11176 , \10611 , \10226 );
and \U$9309 ( \11177 , \10520 , \10224 );
nor \U$9310 ( \11178 , \11176 , \11177 );
xnor \U$9311 ( \11179 , \11178 , \10035 );
and \U$9312 ( \11180 , \10658 , \10164 );
and \U$9313 ( \11181 , \10582 , \10162 );
nor \U$9314 ( \11182 , \11180 , \11181 );
xnor \U$9315 ( \11183 , \11182 , \10190 );
xor \U$9316 ( \11184 , \11179 , \11183 );
and \U$9318 ( \11185 , \10637 , \10217 );
nor \U$9319 ( \11186 , 1'b0 , \11185 );
xnor \U$9320 ( \11187 , \11186 , 1'b0 );
xor \U$9321 ( \11188 , \11184 , \11187 );
xor \U$9322 ( \11189 , 1'b0 , \11188 );
and \U$9323 ( \11190 , \10323 , \10532 );
and \U$9324 ( \11191 , \10344 , \10530 );
nor \U$9325 ( \11192 , \11190 , \11191 );
xnor \U$9326 ( \11193 , \11192 , \10558 );
and \U$9327 ( \11194 , \10493 , \10590 );
and \U$9328 ( \11195 , \10367 , \10588 );
nor \U$9329 ( \11196 , \11194 , \11195 );
xnor \U$9330 ( \11197 , \11196 , \10616 );
xor \U$9331 ( \11198 , \11193 , \11197 );
and \U$9332 ( \11199 , \10553 , \10291 );
and \U$9333 ( \11200 , \10460 , \10289 );
nor \U$9334 ( \11201 , \11199 , \11200 );
xnor \U$9335 ( \11202 , \11201 , \10296 );
xor \U$9336 ( \11203 , \11198 , \11202 );
xor \U$9337 ( \11204 , \11189 , \11203 );
and \U$9338 ( \11205 , \11116 , \11120 );
and \U$9339 ( \11206 , \11120 , \11125 );
and \U$9340 ( \11207 , \11116 , \11125 );
or \U$9341 ( \11208 , \11205 , \11206 , \11207 );
and \U$9342 ( \11209 , \11152 , \11156 );
and \U$9343 ( \11210 , \11156 , \11161 );
and \U$9344 ( \11211 , \11152 , \11161 );
or \U$9345 ( \11212 , \11209 , \11210 , \11211 );
xor \U$9346 ( \11213 , \11208 , \11212 );
and \U$9347 ( \11214 , \11142 , \11145 );
or \U$9350 ( \11215 , \11214 , 1'b0 , 1'b0 );
xor \U$9351 ( \11216 , \11213 , \11215 );
xor \U$9352 ( \11217 , \11204 , \11216 );
xor \U$9353 ( \11218 , \11175 , \11217 );
and \U$9354 ( \11219 , \11097 , \11101 );
and \U$9355 ( \11220 , \11101 , \11106 );
and \U$9356 ( \11221 , \11097 , \11106 );
or \U$9357 ( \11222 , \11219 , \11220 , \11221 );
and \U$9359 ( \11223 , \11147 , \11162 );
or \U$9361 ( \11224 , 1'b0 , \11223 , 1'b0 );
xor \U$9362 ( \11225 , \11222 , \11224 );
and \U$9364 ( \11226 , \10185 , \10436 );
not \U$9365 ( \11227 , \11226 );
xnor \U$9366 ( \11228 , \11227 , \10430 );
xor \U$9367 ( \11229 , 1'b0 , \11228 );
and \U$9368 ( \11230 , \10212 , \10472 );
and \U$9369 ( \11231 , \10116 , \10470 );
nor \U$9370 ( \11232 , \11230 , \11231 );
xnor \U$9371 ( \11233 , \11232 , \10498 );
xor \U$9372 ( \11234 , \11229 , \11233 );
xor \U$9373 ( \11235 , \11225 , \11234 );
xor \U$9374 ( \11236 , \11218 , \11235 );
xor \U$9375 ( \11237 , \11173 , \11236 );
and \U$9376 ( \11238 , \11095 , \11128 );
and \U$9377 ( \11239 , \11128 , \11164 );
and \U$9378 ( \11240 , \11095 , \11164 );
or \U$9379 ( \11241 , \11238 , \11239 , \11240 );
nor \U$9380 ( \11242 , \11237 , \11241 );
nor \U$9381 ( \11243 , \11167 , \11242 );
nand \U$9382 ( \11244 , \11091 , \11243 );
and \U$9383 ( \11245 , \11175 , \11217 );
and \U$9384 ( \11246 , \11217 , \11235 );
and \U$9385 ( \11247 , \11175 , \11235 );
or \U$9386 ( \11248 , \11245 , \11246 , \11247 );
and \U$9387 ( \11249 , \11208 , \11212 );
and \U$9388 ( \11250 , \11212 , \11215 );
and \U$9389 ( \11251 , \11208 , \11215 );
or \U$9390 ( \11252 , \11249 , \11250 , \11251 );
and \U$9392 ( \11253 , \11188 , \11203 );
or \U$9394 ( \11254 , 1'b0 , \11253 , 1'b0 );
xor \U$9395 ( \11255 , \11252 , \11254 );
and \U$9396 ( \11256 , \10367 , \10590 );
and \U$9397 ( \11257 , \10323 , \10588 );
nor \U$9398 ( \11258 , \11256 , \11257 );
xnor \U$9399 ( \11259 , \11258 , \10616 );
and \U$9400 ( \11260 , \10460 , \10291 );
and \U$9401 ( \11261 , \10493 , \10289 );
nor \U$9402 ( \11262 , \11260 , \11261 );
xnor \U$9403 ( \11263 , \11262 , \10296 );
xor \U$9404 ( \11264 , \11259 , \11263 );
and \U$9405 ( \11265 , \10520 , \10226 );
and \U$9406 ( \11266 , \10553 , \10224 );
nor \U$9407 ( \11267 , \11265 , \11266 );
xnor \U$9408 ( \11268 , \11267 , \10035 );
xor \U$9409 ( \11269 , \11264 , \11268 );
xor \U$9410 ( \11270 , \11255 , \11269 );
xor \U$9411 ( \11271 , \11248 , \11270 );
and \U$9412 ( \11272 , \11222 , \11224 );
and \U$9413 ( \11273 , \11224 , \11234 );
and \U$9414 ( \11274 , \11222 , \11234 );
or \U$9415 ( \11275 , \11272 , \11273 , \11274 );
and \U$9416 ( \11276 , \11204 , \11216 );
xor \U$9417 ( \11277 , \11275 , \11276 );
not \U$9418 ( \11278 , \10430 );
and \U$9419 ( \11279 , \10116 , \10472 );
and \U$9420 ( \11280 , \10185 , \10470 );
nor \U$9421 ( \11281 , \11279 , \11280 );
xnor \U$9422 ( \11282 , \11281 , \10498 );
xor \U$9423 ( \11283 , \11278 , \11282 );
and \U$9424 ( \11284 , \10344 , \10532 );
and \U$9425 ( \11285 , \10212 , \10530 );
nor \U$9426 ( \11286 , \11284 , \11285 );
xnor \U$9427 ( \11287 , \11286 , \10558 );
xor \U$9428 ( \11288 , \11283 , \11287 );
and \U$9430 ( \11289 , \10582 , \10164 );
and \U$9431 ( \11290 , \10611 , \10162 );
nor \U$9432 ( \11291 , \11289 , \11290 );
xnor \U$9433 ( \11292 , \11291 , \10190 );
and \U$9435 ( \11293 , \10658 , \10217 );
nor \U$9436 ( \11294 , 1'b0 , \11293 );
xnor \U$9437 ( \11295 , \11294 , 1'b0 );
xor \U$9438 ( \11296 , \11292 , \11295 );
xor \U$9440 ( \11297 , \11296 , 1'b0 );
xor \U$9441 ( \11298 , 1'b1 , \11297 );
xor \U$9442 ( \11299 , \11288 , \11298 );
and \U$9444 ( \11300 , \11228 , \11233 );
or \U$9446 ( \11301 , 1'b0 , \11300 , 1'b0 );
and \U$9447 ( \11302 , \11193 , \11197 );
and \U$9448 ( \11303 , \11197 , \11202 );
and \U$9449 ( \11304 , \11193 , \11202 );
or \U$9450 ( \11305 , \11302 , \11303 , \11304 );
xor \U$9451 ( \11306 , \11301 , \11305 );
and \U$9452 ( \11307 , \11179 , \11183 );
and \U$9453 ( \11308 , \11183 , \11187 );
and \U$9454 ( \11309 , \11179 , \11187 );
or \U$9455 ( \11310 , \11307 , \11308 , \11309 );
xor \U$9456 ( \11311 , \11306 , \11310 );
xor \U$9457 ( \11312 , \11299 , \11311 );
xor \U$9458 ( \11313 , \11277 , \11312 );
xor \U$9459 ( \11314 , \11271 , \11313 );
and \U$9460 ( \11315 , \11171 , \11172 );
and \U$9461 ( \11316 , \11172 , \11236 );
and \U$9462 ( \11317 , \11171 , \11236 );
or \U$9463 ( \11318 , \11315 , \11316 , \11317 );
nor \U$9464 ( \11319 , \11314 , \11318 );
and \U$9465 ( \11320 , \11275 , \11276 );
and \U$9466 ( \11321 , \11276 , \11312 );
and \U$9467 ( \11322 , \11275 , \11312 );
or \U$9468 ( \11323 , \11320 , \11321 , \11322 );
and \U$9469 ( \11324 , \11278 , \11282 );
and \U$9470 ( \11325 , \11282 , \11287 );
and \U$9471 ( \11326 , \11278 , \11287 );
or \U$9472 ( \11327 , \11324 , \11325 , \11326 );
and \U$9473 ( \11328 , \11259 , \11263 );
and \U$9474 ( \11329 , \11263 , \11268 );
and \U$9475 ( \11330 , \11259 , \11268 );
or \U$9476 ( \11331 , \11328 , \11329 , \11330 );
xor \U$9477 ( \11332 , \11327 , \11331 );
and \U$9478 ( \11333 , \11292 , \11295 );
or \U$9481 ( \11334 , \11333 , 1'b0 , 1'b0 );
xor \U$9482 ( \11335 , \11332 , \11334 );
and \U$9483 ( \11336 , \11301 , \11305 );
and \U$9484 ( \11337 , \11305 , \11310 );
and \U$9485 ( \11338 , \11301 , \11310 );
or \U$9486 ( \11339 , \11336 , \11337 , \11338 );
and \U$9489 ( \11340 , 1'b1 , \11297 );
or \U$9491 ( \11341 , 1'b0 , \11340 , 1'b0 );
xor \U$9492 ( \11342 , \11339 , \11341 );
and \U$9493 ( \11343 , \10611 , \10164 );
and \U$9494 ( \11344 , \10520 , \10162 );
nor \U$9495 ( \11345 , \11343 , \11344 );
xnor \U$9496 ( \11346 , \11345 , \10190 );
and \U$9498 ( \11347 , \10582 , \10217 );
nor \U$9499 ( \11348 , 1'b0 , \11347 );
xnor \U$9500 ( \11349 , \11348 , 1'b0 );
xor \U$9501 ( \11350 , \11346 , \11349 );
xor \U$9503 ( \11351 , \11350 , 1'b0 );
and \U$9504 ( \11352 , \10323 , \10590 );
and \U$9505 ( \11353 , \10344 , \10588 );
nor \U$9506 ( \11354 , \11352 , \11353 );
xnor \U$9507 ( \11355 , \11354 , \10616 );
and \U$9508 ( \11356 , \10493 , \10291 );
and \U$9509 ( \11357 , \10367 , \10289 );
nor \U$9510 ( \11358 , \11356 , \11357 );
xnor \U$9511 ( \11359 , \11358 , \10296 );
xor \U$9512 ( \11360 , \11355 , \11359 );
and \U$9513 ( \11361 , \10553 , \10226 );
and \U$9514 ( \11362 , \10460 , \10224 );
nor \U$9515 ( \11363 , \11361 , \11362 );
xnor \U$9516 ( \11364 , \11363 , \10035 );
xor \U$9517 ( \11365 , \11360 , \11364 );
xor \U$9518 ( \11366 , \11351 , \11365 );
and \U$9520 ( \11367 , \10185 , \10472 );
not \U$9521 ( \11368 , \11367 );
xnor \U$9522 ( \11369 , \11368 , \10498 );
xor \U$9523 ( \11370 , 1'b0 , \11369 );
and \U$9524 ( \11371 , \10212 , \10532 );
and \U$9525 ( \11372 , \10116 , \10530 );
nor \U$9526 ( \11373 , \11371 , \11372 );
xnor \U$9527 ( \11374 , \11373 , \10558 );
xor \U$9528 ( \11375 , \11370 , \11374 );
xor \U$9529 ( \11376 , \11366 , \11375 );
xor \U$9530 ( \11377 , \11342 , \11376 );
xor \U$9531 ( \11378 , \11335 , \11377 );
xor \U$9532 ( \11379 , \11323 , \11378 );
and \U$9533 ( \11380 , \11252 , \11254 );
and \U$9534 ( \11381 , \11254 , \11269 );
and \U$9535 ( \11382 , \11252 , \11269 );
or \U$9536 ( \11383 , \11380 , \11381 , \11382 );
and \U$9537 ( \11384 , \11288 , \11298 );
and \U$9538 ( \11385 , \11298 , \11311 );
and \U$9539 ( \11386 , \11288 , \11311 );
or \U$9540 ( \11387 , \11384 , \11385 , \11386 );
xor \U$9541 ( \11388 , \11383 , \11387 );
xor \U$9543 ( \11389 , \11388 , 1'b1 );
xor \U$9544 ( \11390 , \11379 , \11389 );
and \U$9545 ( \11391 , \11248 , \11270 );
and \U$9546 ( \11392 , \11270 , \11313 );
and \U$9547 ( \11393 , \11248 , \11313 );
or \U$9548 ( \11394 , \11391 , \11392 , \11393 );
nor \U$9549 ( \11395 , \11390 , \11394 );
nor \U$9550 ( \11396 , \11319 , \11395 );
and \U$9551 ( \11397 , \11383 , \11387 );
and \U$9552 ( \11398 , \11387 , 1'b1 );
and \U$9553 ( \11399 , \11383 , 1'b1 );
or \U$9554 ( \11400 , \11397 , \11398 , \11399 );
and \U$9555 ( \11401 , \11335 , \11377 );
xor \U$9556 ( \11402 , \11400 , \11401 );
and \U$9557 ( \11403 , \11339 , \11341 );
and \U$9558 ( \11404 , \11341 , \11376 );
and \U$9559 ( \11405 , \11339 , \11376 );
or \U$9560 ( \11406 , \11403 , \11404 , \11405 );
and \U$9562 ( \11407 , \10611 , \10217 );
nor \U$9563 ( \11408 , 1'b0 , \11407 );
xnor \U$9564 ( \11409 , \11408 , 1'b0 );
xor \U$9566 ( \11410 , \11409 , 1'b0 );
xor \U$9568 ( \11411 , \11410 , 1'b0 );
and \U$9569 ( \11412 , \10367 , \10291 );
and \U$9570 ( \11413 , \10323 , \10289 );
nor \U$9571 ( \11414 , \11412 , \11413 );
xnor \U$9572 ( \11415 , \11414 , \10296 );
and \U$9573 ( \11416 , \10460 , \10226 );
and \U$9574 ( \11417 , \10493 , \10224 );
nor \U$9575 ( \11418 , \11416 , \11417 );
xnor \U$9576 ( \11419 , \11418 , \10035 );
xor \U$9577 ( \11420 , \11415 , \11419 );
and \U$9578 ( \11421 , \10520 , \10164 );
and \U$9579 ( \11422 , \10553 , \10162 );
nor \U$9580 ( \11423 , \11421 , \11422 );
xnor \U$9581 ( \11424 , \11423 , \10190 );
xor \U$9582 ( \11425 , \11420 , \11424 );
xor \U$9583 ( \11426 , \11411 , \11425 );
not \U$9584 ( \11427 , \10498 );
and \U$9585 ( \11428 , \10116 , \10532 );
and \U$9586 ( \11429 , \10185 , \10530 );
nor \U$9587 ( \11430 , \11428 , \11429 );
xnor \U$9588 ( \11431 , \11430 , \10558 );
xor \U$9589 ( \11432 , \11427 , \11431 );
and \U$9590 ( \11433 , \10344 , \10590 );
and \U$9591 ( \11434 , \10212 , \10588 );
nor \U$9592 ( \11435 , \11433 , \11434 );
xnor \U$9593 ( \11436 , \11435 , \10616 );
xor \U$9594 ( \11437 , \11432 , \11436 );
xor \U$9595 ( \11438 , \11426 , \11437 );
xor \U$9597 ( \11439 , \11438 , 1'b0 );
and \U$9599 ( \11440 , \11369 , \11374 );
or \U$9601 ( \11441 , 1'b0 , \11440 , 1'b0 );
and \U$9602 ( \11442 , \11355 , \11359 );
and \U$9603 ( \11443 , \11359 , \11364 );
and \U$9604 ( \11444 , \11355 , \11364 );
or \U$9605 ( \11445 , \11442 , \11443 , \11444 );
xor \U$9606 ( \11446 , \11441 , \11445 );
and \U$9607 ( \11447 , \11346 , \11349 );
or \U$9610 ( \11448 , \11447 , 1'b0 , 1'b0 );
xor \U$9611 ( \11449 , \11446 , \11448 );
xor \U$9612 ( \11450 , \11439 , \11449 );
xor \U$9613 ( \11451 , \11406 , \11450 );
and \U$9614 ( \11452 , \11327 , \11331 );
and \U$9615 ( \11453 , \11331 , \11334 );
and \U$9616 ( \11454 , \11327 , \11334 );
or \U$9617 ( \11455 , \11452 , \11453 , \11454 );
xor \U$9619 ( \11456 , \11455 , 1'b0 );
and \U$9620 ( \11457 , \11351 , \11365 );
and \U$9621 ( \11458 , \11365 , \11375 );
and \U$9622 ( \11459 , \11351 , \11375 );
or \U$9623 ( \11460 , \11457 , \11458 , \11459 );
xor \U$9624 ( \11461 , \11456 , \11460 );
xor \U$9625 ( \11462 , \11451 , \11461 );
xor \U$9626 ( \11463 , \11402 , \11462 );
and \U$9627 ( \11464 , \11323 , \11378 );
and \U$9628 ( \11465 , \11378 , \11389 );
and \U$9629 ( \11466 , \11323 , \11389 );
or \U$9630 ( \11467 , \11464 , \11465 , \11466 );
nor \U$9631 ( \11468 , \11463 , \11467 );
and \U$9632 ( \11469 , \11406 , \11450 );
and \U$9633 ( \11470 , \11450 , \11461 );
and \U$9634 ( \11471 , \11406 , \11461 );
or \U$9635 ( \11472 , \11469 , \11470 , \11471 );
and \U$9636 ( \11473 , \11441 , \11445 );
and \U$9637 ( \11474 , \11445 , \11448 );
and \U$9638 ( \11475 , \11441 , \11448 );
or \U$9639 ( \11476 , \11473 , \11474 , \11475 );
xor \U$9641 ( \11477 , \11476 , 1'b0 );
and \U$9642 ( \11478 , \11411 , \11425 );
and \U$9643 ( \11479 , \11425 , \11437 );
and \U$9644 ( \11480 , \11411 , \11437 );
or \U$9645 ( \11481 , \11478 , \11479 , \11480 );
xor \U$9646 ( \11482 , \11477 , \11481 );
xor \U$9647 ( \11483 , \11472 , \11482 );
and \U$9650 ( \11484 , \11455 , \11460 );
or \U$9651 ( \11485 , 1'b0 , 1'b0 , \11484 );
and \U$9654 ( \11486 , \11438 , \11449 );
or \U$9655 ( \11487 , 1'b0 , 1'b0 , \11486 );
xor \U$9656 ( \11488 , \11485 , \11487 );
and \U$9657 ( \11489 , \10323 , \10291 );
and \U$9658 ( \11490 , \10344 , \10289 );
nor \U$9659 ( \11491 , \11489 , \11490 );
xnor \U$9660 ( \11492 , \11491 , \10296 );
and \U$9661 ( \11493 , \10493 , \10226 );
and \U$9662 ( \11494 , \10367 , \10224 );
nor \U$9663 ( \11495 , \11493 , \11494 );
xnor \U$9664 ( \11496 , \11495 , \10035 );
xor \U$9665 ( \11497 , \11492 , \11496 );
and \U$9666 ( \11498 , \10553 , \10164 );
and \U$9667 ( \11499 , \10460 , \10162 );
nor \U$9668 ( \11500 , \11498 , \11499 );
xnor \U$9669 ( \11501 , \11500 , \10190 );
xor \U$9670 ( \11502 , \11497 , \11501 );
and \U$9672 ( \11503 , \10185 , \10532 );
not \U$9673 ( \11504 , \11503 );
xnor \U$9674 ( \11505 , \11504 , \10558 );
xor \U$9675 ( \11506 , 1'b0 , \11505 );
and \U$9676 ( \11507 , \10212 , \10590 );
and \U$9677 ( \11508 , \10116 , \10588 );
nor \U$9678 ( \11509 , \11507 , \11508 );
xnor \U$9679 ( \11510 , \11509 , \10616 );
xor \U$9680 ( \11511 , \11506 , \11510 );
xor \U$9681 ( \11512 , \11502 , \11511 );
and \U$9684 ( \11513 , \10520 , \10217 );
nor \U$9685 ( \11514 , 1'b0 , \11513 );
xnor \U$9686 ( \11515 , \11514 , 1'b0 );
xor \U$9688 ( \11516 , \11515 , 1'b0 );
xor \U$9690 ( \11517 , \11516 , 1'b0 );
xnor \U$9691 ( \11518 , 1'b0 , \11517 );
xor \U$9692 ( \11519 , \11512 , \11518 );
and \U$9693 ( \11520 , \11427 , \11431 );
and \U$9694 ( \11521 , \11431 , \11436 );
and \U$9695 ( \11522 , \11427 , \11436 );
or \U$9696 ( \11523 , \11520 , \11521 , \11522 );
and \U$9697 ( \11524 , \11415 , \11419 );
and \U$9698 ( \11525 , \11419 , \11424 );
and \U$9699 ( \11526 , \11415 , \11424 );
or \U$9700 ( \11527 , \11524 , \11525 , \11526 );
xor \U$9701 ( \11528 , \11523 , \11527 );
xor \U$9703 ( \11529 , \11528 , 1'b0 );
xor \U$9704 ( \11530 , \11519 , \11529 );
xor \U$9705 ( \11531 , \11488 , \11530 );
xor \U$9706 ( \11532 , \11483 , \11531 );
and \U$9707 ( \11533 , \11400 , \11401 );
and \U$9708 ( \11534 , \11401 , \11462 );
and \U$9709 ( \11535 , \11400 , \11462 );
or \U$9710 ( \11536 , \11533 , \11534 , \11535 );
nor \U$9711 ( \11537 , \11532 , \11536 );
nor \U$9712 ( \11538 , \11468 , \11537 );
nand \U$9713 ( \11539 , \11396 , \11538 );
nor \U$9714 ( \11540 , \11244 , \11539 );
and \U$9715 ( \11541 , \11485 , \11487 );
and \U$9716 ( \11542 , \11487 , \11530 );
and \U$9717 ( \11543 , \11485 , \11530 );
or \U$9718 ( \11544 , \11541 , \11542 , \11543 );
and \U$9719 ( \11545 , \11523 , \11527 );
or \U$9722 ( \11546 , \11545 , 1'b0 , 1'b0 );
or \U$9723 ( \11547 , 1'b0 , \11517 );
xor \U$9724 ( \11548 , \11546 , \11547 );
and \U$9725 ( \11549 , \11502 , \11511 );
xor \U$9726 ( \11550 , \11548 , \11549 );
xor \U$9727 ( \11551 , \11544 , \11550 );
and \U$9730 ( \11552 , \11476 , \11481 );
or \U$9731 ( \11553 , 1'b0 , 1'b0 , \11552 );
and \U$9732 ( \11554 , \11512 , \11518 );
and \U$9733 ( \11555 , \11518 , \11529 );
and \U$9734 ( \11556 , \11512 , \11529 );
or \U$9735 ( \11557 , \11554 , \11555 , \11556 );
xor \U$9736 ( \11558 , \11553 , \11557 );
and \U$9738 ( \11559 , \10367 , \10226 );
and \U$9739 ( \11560 , \10323 , \10224 );
nor \U$9740 ( \11561 , \11559 , \11560 );
xnor \U$9741 ( \11562 , \11561 , \10035 );
and \U$9742 ( \11563 , \10460 , \10164 );
and \U$9743 ( \11564 , \10493 , \10162 );
nor \U$9744 ( \11565 , \11563 , \11564 );
xnor \U$9745 ( \11566 , \11565 , \10190 );
xor \U$9746 ( \11567 , \11562 , \11566 );
and \U$9748 ( \11568 , \10553 , \10217 );
nor \U$9749 ( \11569 , 1'b0 , \11568 );
xnor \U$9750 ( \11570 , \11569 , 1'b0 );
xor \U$9751 ( \11571 , \11567 , \11570 );
xor \U$9752 ( \11572 , 1'b0 , \11571 );
not \U$9753 ( \11573 , \10558 );
and \U$9754 ( \11574 , \10116 , \10590 );
and \U$9755 ( \11575 , \10185 , \10588 );
nor \U$9756 ( \11576 , \11574 , \11575 );
xnor \U$9757 ( \11577 , \11576 , \10616 );
xor \U$9758 ( \11578 , \11573 , \11577 );
and \U$9759 ( \11579 , \10344 , \10291 );
and \U$9760 ( \11580 , \10212 , \10289 );
nor \U$9761 ( \11581 , \11579 , \11580 );
xnor \U$9762 ( \11582 , \11581 , \10296 );
xor \U$9763 ( \11583 , \11578 , \11582 );
xor \U$9764 ( \11584 , \11572 , \11583 );
xor \U$9766 ( \11585 , \11584 , 1'b0 );
and \U$9768 ( \11586 , \11505 , \11510 );
or \U$9770 ( \11587 , 1'b0 , \11586 , 1'b0 );
and \U$9771 ( \11588 , \11492 , \11496 );
and \U$9772 ( \11589 , \11496 , \11501 );
and \U$9773 ( \11590 , \11492 , \11501 );
or \U$9774 ( \11591 , \11588 , \11589 , \11590 );
xor \U$9775 ( \11592 , \11587 , \11591 );
xor \U$9777 ( \11593 , \11592 , 1'b0 );
xor \U$9778 ( \11594 , \11585 , \11593 );
xor \U$9779 ( \11595 , \11558 , \11594 );
xor \U$9780 ( \11596 , \11551 , \11595 );
and \U$9781 ( \11597 , \11472 , \11482 );
and \U$9782 ( \11598 , \11482 , \11531 );
and \U$9783 ( \11599 , \11472 , \11531 );
or \U$9784 ( \11600 , \11597 , \11598 , \11599 );
nor \U$9785 ( \11601 , \11596 , \11600 );
and \U$9786 ( \11602 , \11553 , \11557 );
and \U$9787 ( \11603 , \11557 , \11594 );
and \U$9788 ( \11604 , \11553 , \11594 );
or \U$9789 ( \11605 , \11602 , \11603 , \11604 );
and \U$9790 ( \11606 , \11587 , \11591 );
or \U$9793 ( \11607 , \11606 , 1'b0 , 1'b0 );
xor \U$9795 ( \11608 , \11607 , 1'b0 );
and \U$9797 ( \11609 , \11571 , \11583 );
or \U$9799 ( \11610 , 1'b0 , \11609 , 1'b0 );
xor \U$9800 ( \11611 , \11608 , \11610 );
xor \U$9801 ( \11612 , \11605 , \11611 );
and \U$9802 ( \11613 , \11546 , \11547 );
and \U$9803 ( \11614 , \11547 , \11549 );
and \U$9804 ( \11615 , \11546 , \11549 );
or \U$9805 ( \11616 , \11613 , \11614 , \11615 );
and \U$9808 ( \11617 , \11584 , \11593 );
or \U$9809 ( \11618 , 1'b0 , 1'b0 , \11617 );
xor \U$9810 ( \11619 , \11616 , \11618 );
and \U$9811 ( \11620 , \10323 , \10226 );
and \U$9812 ( \11621 , \10344 , \10224 );
nor \U$9813 ( \11622 , \11620 , \11621 );
xnor \U$9814 ( \11623 , \11622 , \10035 );
and \U$9815 ( \11624 , \10493 , \10164 );
and \U$9816 ( \11625 , \10367 , \10162 );
nor \U$9817 ( \11626 , \11624 , \11625 );
xnor \U$9818 ( \11627 , \11626 , \10190 );
xor \U$9819 ( \11628 , \11623 , \11627 );
and \U$9821 ( \11629 , \10460 , \10217 );
nor \U$9822 ( \11630 , 1'b0 , \11629 );
xnor \U$9823 ( \11631 , \11630 , 1'b0 );
xor \U$9824 ( \11632 , \11628 , \11631 );
and \U$9826 ( \11633 , \10185 , \10590 );
not \U$9827 ( \11634 , \11633 );
xnor \U$9828 ( \11635 , \11634 , \10616 );
xor \U$9829 ( \11636 , 1'b0 , \11635 );
and \U$9830 ( \11637 , \10212 , \10291 );
and \U$9831 ( \11638 , \10116 , \10289 );
nor \U$9832 ( \11639 , \11637 , \11638 );
xnor \U$9833 ( \11640 , \11639 , \10296 );
xor \U$9834 ( \11641 , \11636 , \11640 );
xor \U$9835 ( \11642 , \11632 , \11641 );
xor \U$9837 ( \11643 , \11642 , 1'b1 );
and \U$9838 ( \11644 , \11573 , \11577 );
and \U$9839 ( \11645 , \11577 , \11582 );
and \U$9840 ( \11646 , \11573 , \11582 );
or \U$9841 ( \11647 , \11644 , \11645 , \11646 );
and \U$9842 ( \11648 , \11562 , \11566 );
and \U$9843 ( \11649 , \11566 , \11570 );
and \U$9844 ( \11650 , \11562 , \11570 );
or \U$9845 ( \11651 , \11648 , \11649 , \11650 );
xor \U$9846 ( \11652 , \11647 , \11651 );
xor \U$9848 ( \11653 , \11652 , 1'b0 );
xor \U$9849 ( \11654 , \11643 , \11653 );
xor \U$9850 ( \11655 , \11619 , \11654 );
xor \U$9851 ( \11656 , \11612 , \11655 );
and \U$9852 ( \11657 , \11544 , \11550 );
and \U$9853 ( \11658 , \11550 , \11595 );
and \U$9854 ( \11659 , \11544 , \11595 );
or \U$9855 ( \11660 , \11657 , \11658 , \11659 );
nor \U$9856 ( \11661 , \11656 , \11660 );
nor \U$9857 ( \11662 , \11601 , \11661 );
and \U$9858 ( \11663 , \11616 , \11618 );
and \U$9859 ( \11664 , \11618 , \11654 );
and \U$9860 ( \11665 , \11616 , \11654 );
or \U$9861 ( \11666 , \11663 , \11664 , \11665 );
and \U$9862 ( \11667 , \11647 , \11651 );
or \U$9865 ( \11668 , \11667 , 1'b0 , 1'b0 );
xor \U$9867 ( \11669 , \11668 , 1'b0 );
and \U$9868 ( \11670 , \11632 , \11641 );
xor \U$9869 ( \11671 , \11669 , \11670 );
xor \U$9870 ( \11672 , \11666 , \11671 );
and \U$9873 ( \11673 , \11607 , \11610 );
or \U$9874 ( \11674 , 1'b0 , 1'b0 , \11673 );
and \U$9875 ( \11675 , \11642 , 1'b1 );
and \U$9876 ( \11676 , 1'b1 , \11653 );
and \U$9877 ( \11677 , \11642 , \11653 );
or \U$9878 ( \11678 , \11675 , \11676 , \11677 );
xor \U$9879 ( \11679 , \11674 , \11678 );
and \U$9881 ( \11680 , \10367 , \10164 );
and \U$9882 ( \11681 , \10323 , \10162 );
nor \U$9883 ( \11682 , \11680 , \11681 );
xnor \U$9884 ( \11683 , \11682 , \10190 );
and \U$9886 ( \11684 , \10493 , \10217 );
nor \U$9887 ( \11685 , 1'b0 , \11684 );
xnor \U$9888 ( \11686 , \11685 , 1'b0 );
xor \U$9889 ( \11687 , \11683 , \11686 );
xor \U$9891 ( \11688 , \11687 , 1'b0 );
xor \U$9892 ( \11689 , 1'b0 , \11688 );
not \U$9893 ( \11690 , \10616 );
and \U$9894 ( \11691 , \10116 , \10291 );
and \U$9895 ( \11692 , \10185 , \10289 );
nor \U$9896 ( \11693 , \11691 , \11692 );
xnor \U$9897 ( \11694 , \11693 , \10296 );
xor \U$9898 ( \11695 , \11690 , \11694 );
and \U$9899 ( \11696 , \10344 , \10226 );
and \U$9900 ( \11697 , \10212 , \10224 );
nor \U$9901 ( \11698 , \11696 , \11697 );
xnor \U$9902 ( \11699 , \11698 , \10035 );
xor \U$9903 ( \11700 , \11695 , \11699 );
xor \U$9904 ( \11701 , \11689 , \11700 );
xor \U$9906 ( \11702 , \11701 , 1'b0 );
and \U$9908 ( \11703 , \11635 , \11640 );
or \U$9910 ( \11704 , 1'b0 , \11703 , 1'b0 );
and \U$9911 ( \11705 , \11623 , \11627 );
and \U$9912 ( \11706 , \11627 , \11631 );
and \U$9913 ( \11707 , \11623 , \11631 );
or \U$9914 ( \11708 , \11705 , \11706 , \11707 );
xor \U$9915 ( \11709 , \11704 , \11708 );
xor \U$9917 ( \11710 , \11709 , 1'b0 );
xor \U$9918 ( \11711 , \11702 , \11710 );
xor \U$9919 ( \11712 , \11679 , \11711 );
xor \U$9920 ( \11713 , \11672 , \11712 );
and \U$9921 ( \11714 , \11605 , \11611 );
and \U$9922 ( \11715 , \11611 , \11655 );
and \U$9923 ( \11716 , \11605 , \11655 );
or \U$9924 ( \11717 , \11714 , \11715 , \11716 );
nor \U$9925 ( \11718 , \11713 , \11717 );
and \U$9926 ( \11719 , \11674 , \11678 );
and \U$9927 ( \11720 , \11678 , \11711 );
and \U$9928 ( \11721 , \11674 , \11711 );
or \U$9929 ( \11722 , \11719 , \11720 , \11721 );
and \U$9930 ( \11723 , \11704 , \11708 );
or \U$9933 ( \11724 , \11723 , 1'b0 , 1'b0 );
xor \U$9935 ( \11725 , \11724 , 1'b0 );
and \U$9937 ( \11726 , \11688 , \11700 );
or \U$9939 ( \11727 , 1'b0 , \11726 , 1'b0 );
xor \U$9940 ( \11728 , \11725 , \11727 );
xor \U$9941 ( \11729 , \11722 , \11728 );
and \U$9944 ( \11730 , \11668 , \11670 );
or \U$9945 ( \11731 , 1'b0 , 1'b0 , \11730 );
and \U$9948 ( \11732 , \11701 , \11710 );
or \U$9949 ( \11733 , 1'b0 , 1'b0 , \11732 );
xor \U$9950 ( \11734 , \11731 , \11733 );
xor \U$9951 ( \11735 , \10347 , \10370 );
xor \U$9953 ( \11736 , \11735 , 1'b0 );
xor \U$9955 ( \11737 , 1'b0 , \10297 );
xor \U$9956 ( \11738 , \11737 , \10301 );
xor \U$9957 ( \11739 , \11736 , \11738 );
xor \U$9959 ( \11740 , \11739 , 1'b1 );
and \U$9960 ( \11741 , \11690 , \11694 );
and \U$9961 ( \11742 , \11694 , \11699 );
and \U$9962 ( \11743 , \11690 , \11699 );
or \U$9963 ( \11744 , \11741 , \11742 , \11743 );
and \U$9964 ( \11745 , \11683 , \11686 );
or \U$9967 ( \11746 , \11745 , 1'b0 , 1'b0 );
xor \U$9968 ( \11747 , \11744 , \11746 );
xor \U$9970 ( \11748 , \11747 , 1'b0 );
xor \U$9971 ( \11749 , \11740 , \11748 );
xor \U$9972 ( \11750 , \11734 , \11749 );
xor \U$9973 ( \11751 , \11729 , \11750 );
and \U$9974 ( \11752 , \11666 , \11671 );
and \U$9975 ( \11753 , \11671 , \11712 );
and \U$9976 ( \11754 , \11666 , \11712 );
or \U$9977 ( \11755 , \11752 , \11753 , \11754 );
nor \U$9978 ( \11756 , \11751 , \11755 );
nor \U$9979 ( \11757 , \11718 , \11756 );
nand \U$9980 ( \11758 , \11662 , \11757 );
and \U$9981 ( \11759 , \11731 , \11733 );
and \U$9982 ( \11760 , \11733 , \11749 );
and \U$9983 ( \11761 , \11731 , \11749 );
or \U$9984 ( \11762 , \11759 , \11760 , \11761 );
and \U$9985 ( \11763 , \11744 , \11746 );
or \U$9988 ( \11764 , \11763 , 1'b0 , 1'b0 );
xor \U$9990 ( \11765 , \11764 , 1'b0 );
and \U$9991 ( \11766 , \11736 , \11738 );
xor \U$9992 ( \11767 , \11765 , \11766 );
xor \U$9993 ( \11768 , \11762 , \11767 );
and \U$9996 ( \11769 , \11724 , \11727 );
or \U$9997 ( \11770 , 1'b0 , 1'b0 , \11769 );
and \U$9998 ( \11771 , \11739 , 1'b1 );
and \U$9999 ( \11772 , 1'b1 , \11748 );
and \U$10000 ( \11773 , \11739 , \11748 );
or \U$10001 ( \11774 , \11771 , \11772 , \11773 );
xor \U$10002 ( \11775 , \11770 , \11774 );
xor \U$10004 ( \11776 , 1'b0 , \10379 );
xor \U$10005 ( \11777 , \11776 , \10390 );
xor \U$10007 ( \11778 , \11777 , 1'b0 );
xor \U$10008 ( \11779 , \10303 , \10372 );
xor \U$10010 ( \11780 , \11779 , 1'b0 );
xor \U$10011 ( \11781 , \11778 , \11780 );
xor \U$10012 ( \11782 , \11775 , \11781 );
xor \U$10013 ( \11783 , \11768 , \11782 );
and \U$10014 ( \11784 , \11722 , \11728 );
and \U$10015 ( \11785 , \11728 , \11750 );
and \U$10016 ( \11786 , \11722 , \11750 );
or \U$10017 ( \11787 , \11784 , \11785 , \11786 );
nor \U$10018 ( \11788 , \11783 , \11787 );
and \U$10019 ( \11789 , \11770 , \11774 );
and \U$10020 ( \11790 , \11774 , \11781 );
and \U$10021 ( \11791 , \11770 , \11781 );
or \U$10022 ( \11792 , \11789 , \11790 , \11791 );
xor \U$10024 ( \11793 , \10374 , 1'b0 );
xor \U$10025 ( \11794 , \11793 , \10392 );
xor \U$10026 ( \11795 , \11792 , \11794 );
and \U$10029 ( \11796 , \11764 , \11766 );
or \U$10030 ( \11797 , 1'b0 , 1'b0 , \11796 );
and \U$10033 ( \11798 , \11777 , \11780 );
or \U$10034 ( \11799 , 1'b0 , 1'b0 , \11798 );
xor \U$10035 ( \11800 , \11797 , \11799 );
xor \U$10036 ( \11801 , \10402 , 1'b1 );
xor \U$10037 ( \11802 , \11801 , \10409 );
xor \U$10038 ( \11803 , \11800 , \11802 );
xor \U$10039 ( \11804 , \11795 , \11803 );
and \U$10040 ( \11805 , \11762 , \11767 );
and \U$10041 ( \11806 , \11767 , \11782 );
and \U$10042 ( \11807 , \11762 , \11782 );
or \U$10043 ( \11808 , \11805 , \11806 , \11807 );
nor \U$10044 ( \11809 , \11804 , \11808 );
nor \U$10045 ( \11810 , \11788 , \11809 );
and \U$10046 ( \11811 , \11797 , \11799 );
and \U$10047 ( \11812 , \11799 , \11802 );
and \U$10048 ( \11813 , \11797 , \11802 );
or \U$10049 ( \11814 , \11811 , \11812 , \11813 );
and \U$10051 ( \11815 , \10399 , \10401 );
xor \U$10052 ( \11816 , 1'b0 , \11815 );
xor \U$10053 ( \11817 , \11814 , \11816 );
xor \U$10054 ( \11818 , \10394 , \10412 );
xor \U$10055 ( \11819 , \11818 , \10415 );
xor \U$10056 ( \11820 , \11817 , \11819 );
and \U$10057 ( \11821 , \11792 , \11794 );
and \U$10058 ( \11822 , \11794 , \11803 );
and \U$10059 ( \11823 , \11792 , \11803 );
or \U$10060 ( \11824 , \11821 , \11822 , \11823 );
nor \U$10061 ( \11825 , \11820 , \11824 );
xor \U$10063 ( \11826 , \10418 , 1'b0 );
xor \U$10064 ( \11827 , \11826 , \10420 );
and \U$10065 ( \11828 , \11814 , \11816 );
and \U$10066 ( \11829 , \11816 , \11819 );
and \U$10067 ( \11830 , \11814 , \11819 );
or \U$10068 ( \11831 , \11828 , \11829 , \11830 );
nor \U$10069 ( \11832 , \11827 , \11831 );
nor \U$10070 ( \11833 , \11825 , \11832 );
nand \U$10071 ( \11834 , \11810 , \11833 );
nor \U$10072 ( \11835 , \11758 , \11834 );
nand \U$10073 ( \11836 , \11540 , \11835 );
and \U$10074 ( \11837 , \10637 , \10436 );
and \U$10075 ( \11838 , \10658 , \10433 );
nor \U$10076 ( \11839 , \11837 , \11838 );
xnor \U$10077 ( \11840 , \11839 , \10430 );
and \U$10078 ( \11841 , \10682 , \10472 );
and \U$10079 ( \11842 , \10703 , \10470 );
nor \U$10080 ( \11843 , \11841 , \11842 );
xnor \U$10081 ( \11844 , \11843 , \10498 );
and \U$10082 ( \11845 , \11840 , \11844 );
and \U$10083 ( \11846 , \10730 , \10532 );
and \U$10084 ( \11847 , \10751 , \10530 );
nor \U$10085 ( \11848 , \11846 , \11847 );
xnor \U$10086 ( \11849 , \11848 , \10558 );
and \U$10087 ( \11850 , \11844 , \11849 );
and \U$10088 ( \11851 , \11840 , \11849 );
or \U$10089 ( \11852 , \11845 , \11850 , \11851 );
and \U$10090 ( \11853 , \10751 , \10532 );
and \U$10091 ( \11854 , \10682 , \10530 );
nor \U$10092 ( \11855 , \11853 , \11854 );
xnor \U$10093 ( \11856 , \11855 , \10558 );
and \U$10094 ( \11857 , \10774 , \10590 );
and \U$10095 ( \11858 , \10730 , \10588 );
nor \U$10096 ( \11859 , \11857 , \11858 );
xnor \U$10097 ( \11860 , \11859 , \10616 );
xor \U$10098 ( \11861 , \11856 , \11860 );
nand \U$10099 ( \11862 , \10907 , \10289 );
xnor \U$10100 ( \11863 , \11862 , \10296 );
xor \U$10101 ( \11864 , \11861 , \11863 );
and \U$10102 ( \11865 , \11852 , \11864 );
and \U$10103 ( \11866 , \10658 , \10436 );
and \U$10104 ( \11867 , \10582 , \10433 );
nor \U$10105 ( \11868 , \11866 , \11867 );
xnor \U$10106 ( \11869 , \11868 , \10430 );
xor \U$10107 ( \11870 , \10296 , \11869 );
and \U$10108 ( \11871 , \10703 , \10472 );
and \U$10109 ( \11872 , \10637 , \10470 );
nor \U$10110 ( \11873 , \11871 , \11872 );
xnor \U$10111 ( \11874 , \11873 , \10498 );
xor \U$10112 ( \11875 , \11870 , \11874 );
and \U$10113 ( \11876 , \11864 , \11875 );
and \U$10114 ( \11877 , \11852 , \11875 );
or \U$10115 ( \11878 , \11865 , \11876 , \11877 );
and \U$10116 ( \11879 , \10907 , \10291 );
and \U$10117 ( \11880 , \10774 , \10289 );
nor \U$10118 ( \11881 , \11879 , \11880 );
xnor \U$10119 ( \11882 , \11881 , \10296 );
and \U$10120 ( \11883 , \10582 , \10436 );
and \U$10121 ( \11884 , \10611 , \10433 );
nor \U$10122 ( \11885 , \11883 , \11884 );
xnor \U$10123 ( \11886 , \11885 , \10430 );
and \U$10124 ( \11887 , \10637 , \10472 );
and \U$10125 ( \11888 , \10658 , \10470 );
nor \U$10126 ( \11889 , \11887 , \11888 );
xnor \U$10127 ( \11890 , \11889 , \10498 );
xor \U$10128 ( \11891 , \11886 , \11890 );
and \U$10129 ( \11892 , \10682 , \10532 );
and \U$10130 ( \11893 , \10703 , \10530 );
nor \U$10131 ( \11894 , \11892 , \11893 );
xnor \U$10132 ( \11895 , \11894 , \10558 );
xor \U$10133 ( \11896 , \11891 , \11895 );
xor \U$10134 ( \11897 , \11882 , \11896 );
xor \U$10135 ( \11898 , \11878 , \11897 );
and \U$10136 ( \11899 , \10296 , \11869 );
and \U$10137 ( \11900 , \11869 , \11874 );
and \U$10138 ( \11901 , \10296 , \11874 );
or \U$10139 ( \11902 , \11899 , \11900 , \11901 );
and \U$10140 ( \11903 , \11856 , \11860 );
and \U$10141 ( \11904 , \11860 , \11863 );
and \U$10142 ( \11905 , \11856 , \11863 );
or \U$10143 ( \11906 , \11903 , \11904 , \11905 );
xor \U$10144 ( \11907 , \11902 , \11906 );
and \U$10145 ( \11908 , \10730 , \10590 );
and \U$10146 ( \11909 , \10751 , \10588 );
nor \U$10147 ( \11910 , \11908 , \11909 );
xnor \U$10148 ( \11911 , \11910 , \10616 );
xor \U$10149 ( \11912 , \11907 , \11911 );
xor \U$10150 ( \11913 , \11898 , \11912 );
and \U$10151 ( \11914 , \10703 , \10436 );
and \U$10152 ( \11915 , \10637 , \10433 );
nor \U$10153 ( \11916 , \11914 , \11915 );
xnor \U$10154 ( \11917 , \11916 , \10430 );
and \U$10155 ( \11918 , \10616 , \11917 );
and \U$10156 ( \11919 , \10751 , \10472 );
and \U$10157 ( \11920 , \10682 , \10470 );
nor \U$10158 ( \11921 , \11919 , \11920 );
xnor \U$10159 ( \11922 , \11921 , \10498 );
and \U$10160 ( \11923 , \11917 , \11922 );
and \U$10161 ( \11924 , \10616 , \11922 );
or \U$10162 ( \11925 , \11918 , \11923 , \11924 );
and \U$10163 ( \11926 , \10774 , \10532 );
and \U$10164 ( \11927 , \10730 , \10530 );
nor \U$10165 ( \11928 , \11926 , \11927 );
xnor \U$10166 ( \11929 , \11928 , \10558 );
nand \U$10167 ( \11930 , \10907 , \10588 );
xnor \U$10168 ( \11931 , \11930 , \10616 );
and \U$10169 ( \11932 , \11929 , \11931 );
and \U$10170 ( \11933 , \11925 , \11932 );
and \U$10171 ( \11934 , \10907 , \10590 );
and \U$10172 ( \11935 , \10774 , \10588 );
nor \U$10173 ( \11936 , \11934 , \11935 );
xnor \U$10174 ( \11937 , \11936 , \10616 );
and \U$10175 ( \11938 , \11932 , \11937 );
and \U$10176 ( \11939 , \11925 , \11937 );
or \U$10177 ( \11940 , \11933 , \11938 , \11939 );
xor \U$10178 ( \11941 , \11852 , \11864 );
xor \U$10179 ( \11942 , \11941 , \11875 );
and \U$10180 ( \11943 , \11940 , \11942 );
nor \U$10181 ( \11944 , \11913 , \11943 );
and \U$10182 ( \11945 , \11886 , \11890 );
and \U$10183 ( \11946 , \11890 , \11895 );
and \U$10184 ( \11947 , \11886 , \11895 );
or \U$10185 ( \11948 , \11945 , \11946 , \11947 );
nand \U$10186 ( \11949 , \10907 , \10224 );
xnor \U$10187 ( \11950 , \11949 , \10035 );
xor \U$10188 ( \11951 , \11948 , \11950 );
and \U$10189 ( \11952 , \10703 , \10532 );
and \U$10190 ( \11953 , \10637 , \10530 );
nor \U$10191 ( \11954 , \11952 , \11953 );
xnor \U$10192 ( \11955 , \11954 , \10558 );
and \U$10193 ( \11956 , \10751 , \10590 );
and \U$10194 ( \11957 , \10682 , \10588 );
nor \U$10195 ( \11958 , \11956 , \11957 );
xnor \U$10196 ( \11959 , \11958 , \10616 );
xor \U$10197 ( \11960 , \11955 , \11959 );
and \U$10198 ( \11961 , \10774 , \10291 );
and \U$10199 ( \11962 , \10730 , \10289 );
nor \U$10200 ( \11963 , \11961 , \11962 );
xnor \U$10201 ( \11964 , \11963 , \10296 );
xor \U$10202 ( \11965 , \11960 , \11964 );
xor \U$10203 ( \11966 , \11951 , \11965 );
and \U$10204 ( \11967 , \11902 , \11906 );
and \U$10205 ( \11968 , \11906 , \11911 );
and \U$10206 ( \11969 , \11902 , \11911 );
or \U$10207 ( \11970 , \11967 , \11968 , \11969 );
and \U$10208 ( \11971 , \11882 , \11896 );
xor \U$10209 ( \11972 , \11970 , \11971 );
and \U$10210 ( \11973 , \10611 , \10436 );
and \U$10211 ( \11974 , \10520 , \10433 );
nor \U$10212 ( \11975 , \11973 , \11974 );
xnor \U$10213 ( \11976 , \11975 , \10430 );
xor \U$10214 ( \11977 , \10035 , \11976 );
and \U$10215 ( \11978 , \10658 , \10472 );
and \U$10216 ( \11979 , \10582 , \10470 );
nor \U$10217 ( \11980 , \11978 , \11979 );
xnor \U$10218 ( \11981 , \11980 , \10498 );
xor \U$10219 ( \11982 , \11977 , \11981 );
xor \U$10220 ( \11983 , \11972 , \11982 );
xor \U$10221 ( \11984 , \11966 , \11983 );
and \U$10222 ( \11985 , \11878 , \11897 );
and \U$10223 ( \11986 , \11897 , \11912 );
and \U$10224 ( \11987 , \11878 , \11912 );
or \U$10225 ( \11988 , \11985 , \11986 , \11987 );
nor \U$10226 ( \11989 , \11984 , \11988 );
nor \U$10227 ( \11990 , \11944 , \11989 );
and \U$10228 ( \11991 , \11970 , \11971 );
and \U$10229 ( \11992 , \11971 , \11982 );
and \U$10230 ( \11993 , \11970 , \11982 );
or \U$10231 ( \11994 , \11991 , \11992 , \11993 );
and \U$10232 ( \11995 , \11948 , \11950 );
and \U$10233 ( \11996 , \11950 , \11965 );
and \U$10234 ( \11997 , \11948 , \11965 );
or \U$10235 ( \11998 , \11995 , \11996 , \11997 );
and \U$10236 ( \11999 , \10520 , \10436 );
and \U$10237 ( \12000 , \10553 , \10433 );
nor \U$10238 ( \12001 , \11999 , \12000 );
xnor \U$10239 ( \12002 , \12001 , \10430 );
and \U$10240 ( \12003 , \10582 , \10472 );
and \U$10241 ( \12004 , \10611 , \10470 );
nor \U$10242 ( \12005 , \12003 , \12004 );
xnor \U$10243 ( \12006 , \12005 , \10498 );
xor \U$10244 ( \12007 , \12002 , \12006 );
and \U$10245 ( \12008 , \10637 , \10532 );
and \U$10246 ( \12009 , \10658 , \10530 );
nor \U$10247 ( \12010 , \12008 , \12009 );
xnor \U$10248 ( \12011 , \12010 , \10558 );
xor \U$10249 ( \12012 , \12007 , \12011 );
xor \U$10250 ( \12013 , \11998 , \12012 );
and \U$10251 ( \12014 , \10035 , \11976 );
and \U$10252 ( \12015 , \11976 , \11981 );
and \U$10253 ( \12016 , \10035 , \11981 );
or \U$10254 ( \12017 , \12014 , \12015 , \12016 );
and \U$10255 ( \12018 , \11955 , \11959 );
and \U$10256 ( \12019 , \11959 , \11964 );
and \U$10257 ( \12020 , \11955 , \11964 );
or \U$10258 ( \12021 , \12018 , \12019 , \12020 );
xor \U$10259 ( \12022 , \12017 , \12021 );
and \U$10260 ( \12023 , \10682 , \10590 );
and \U$10261 ( \12024 , \10703 , \10588 );
nor \U$10262 ( \12025 , \12023 , \12024 );
xnor \U$10263 ( \12026 , \12025 , \10616 );
and \U$10264 ( \12027 , \10730 , \10291 );
and \U$10265 ( \12028 , \10751 , \10289 );
nor \U$10266 ( \12029 , \12027 , \12028 );
xnor \U$10267 ( \12030 , \12029 , \10296 );
xor \U$10268 ( \12031 , \12026 , \12030 );
and \U$10269 ( \12032 , \10907 , \10226 );
and \U$10270 ( \12033 , \10774 , \10224 );
nor \U$10271 ( \12034 , \12032 , \12033 );
xnor \U$10272 ( \12035 , \12034 , \10035 );
xor \U$10273 ( \12036 , \12031 , \12035 );
xor \U$10274 ( \12037 , \12022 , \12036 );
xor \U$10275 ( \12038 , \12013 , \12037 );
xor \U$10276 ( \12039 , \11994 , \12038 );
and \U$10277 ( \12040 , \11966 , \11983 );
nor \U$10278 ( \12041 , \12039 , \12040 );
and \U$10279 ( \12042 , \11998 , \12012 );
and \U$10280 ( \12043 , \12012 , \12037 );
and \U$10281 ( \12044 , \11998 , \12037 );
or \U$10282 ( \12045 , \12042 , \12043 , \12044 );
and \U$10283 ( \12046 , \12017 , \12021 );
and \U$10284 ( \12047 , \12021 , \12036 );
and \U$10285 ( \12048 , \12017 , \12036 );
or \U$10286 ( \12049 , \12046 , \12047 , \12048 );
nand \U$10287 ( \12050 , \10907 , \10162 );
xnor \U$10288 ( \12051 , \12050 , \10190 );
and \U$10289 ( \12052 , \10658 , \10532 );
and \U$10290 ( \12053 , \10582 , \10530 );
nor \U$10291 ( \12054 , \12052 , \12053 );
xnor \U$10292 ( \12055 , \12054 , \10558 );
and \U$10293 ( \12056 , \10703 , \10590 );
and \U$10294 ( \12057 , \10637 , \10588 );
nor \U$10295 ( \12058 , \12056 , \12057 );
xnor \U$10296 ( \12059 , \12058 , \10616 );
xor \U$10297 ( \12060 , \12055 , \12059 );
and \U$10298 ( \12061 , \10751 , \10291 );
and \U$10299 ( \12062 , \10682 , \10289 );
nor \U$10300 ( \12063 , \12061 , \12062 );
xnor \U$10301 ( \12064 , \12063 , \10296 );
xor \U$10302 ( \12065 , \12060 , \12064 );
xor \U$10303 ( \12066 , \12051 , \12065 );
and \U$10304 ( \12067 , \10553 , \10436 );
and \U$10305 ( \12068 , \10460 , \10433 );
nor \U$10306 ( \12069 , \12067 , \12068 );
xnor \U$10307 ( \12070 , \12069 , \10430 );
xor \U$10308 ( \12071 , \10190 , \12070 );
and \U$10309 ( \12072 , \10611 , \10472 );
and \U$10310 ( \12073 , \10520 , \10470 );
nor \U$10311 ( \12074 , \12072 , \12073 );
xnor \U$10312 ( \12075 , \12074 , \10498 );
xor \U$10313 ( \12076 , \12071 , \12075 );
xor \U$10314 ( \12077 , \12066 , \12076 );
xor \U$10315 ( \12078 , \12049 , \12077 );
and \U$10316 ( \12079 , \12002 , \12006 );
and \U$10317 ( \12080 , \12006 , \12011 );
and \U$10318 ( \12081 , \12002 , \12011 );
or \U$10319 ( \12082 , \12079 , \12080 , \12081 );
and \U$10320 ( \12083 , \12026 , \12030 );
and \U$10321 ( \12084 , \12030 , \12035 );
and \U$10322 ( \12085 , \12026 , \12035 );
or \U$10323 ( \12086 , \12083 , \12084 , \12085 );
xor \U$10324 ( \12087 , \12082 , \12086 );
and \U$10325 ( \12088 , \10774 , \10226 );
and \U$10326 ( \12089 , \10730 , \10224 );
nor \U$10327 ( \12090 , \12088 , \12089 );
xnor \U$10328 ( \12091 , \12090 , \10035 );
xor \U$10329 ( \12092 , \12087 , \12091 );
xor \U$10330 ( \12093 , \12078 , \12092 );
xor \U$10331 ( \12094 , \12045 , \12093 );
and \U$10332 ( \12095 , \11994 , \12038 );
nor \U$10333 ( \12096 , \12094 , \12095 );
nor \U$10334 ( \12097 , \12041 , \12096 );
nand \U$10335 ( \12098 , \11990 , \12097 );
and \U$10336 ( \12099 , \12049 , \12077 );
and \U$10337 ( \12100 , \12077 , \12092 );
and \U$10338 ( \12101 , \12049 , \12092 );
or \U$10339 ( \12102 , \12099 , \12100 , \12101 );
xor \U$10340 ( \12103 , \10962 , \10966 );
xor \U$10341 ( \12104 , \12103 , \10971 );
and \U$10342 ( \12105 , \10190 , \12070 );
and \U$10343 ( \12106 , \12070 , \12075 );
and \U$10344 ( \12107 , \10190 , \12075 );
or \U$10345 ( \12108 , \12105 , \12106 , \12107 );
and \U$10346 ( \12109 , \12055 , \12059 );
and \U$10347 ( \12110 , \12059 , \12064 );
and \U$10348 ( \12111 , \12055 , \12064 );
or \U$10349 ( \12112 , \12109 , \12110 , \12111 );
xor \U$10350 ( \12113 , \12108 , \12112 );
and \U$10351 ( \12114 , \10907 , \10164 );
and \U$10352 ( \12115 , \10774 , \10162 );
nor \U$10353 ( \12116 , \12114 , \12115 );
xnor \U$10354 ( \12117 , \12116 , \10190 );
xor \U$10355 ( \12118 , \12113 , \12117 );
xor \U$10356 ( \12119 , \12104 , \12118 );
xor \U$10357 ( \12120 , \12102 , \12119 );
and \U$10358 ( \12121 , \12082 , \12086 );
and \U$10359 ( \12122 , \12086 , \12091 );
and \U$10360 ( \12123 , \12082 , \12091 );
or \U$10361 ( \12124 , \12121 , \12122 , \12123 );
and \U$10362 ( \12125 , \12051 , \12065 );
and \U$10363 ( \12126 , \12065 , \12076 );
and \U$10364 ( \12127 , \12051 , \12076 );
or \U$10365 ( \12128 , \12125 , \12126 , \12127 );
xor \U$10366 ( \12129 , \12124 , \12128 );
xor \U$10367 ( \12130 , \10978 , \10982 );
xor \U$10368 ( \12131 , \12130 , \10987 );
xor \U$10369 ( \12132 , \12129 , \12131 );
xor \U$10370 ( \12133 , \12120 , \12132 );
and \U$10371 ( \12134 , \12045 , \12093 );
nor \U$10372 ( \12135 , \12133 , \12134 );
and \U$10373 ( \12136 , \12124 , \12128 );
and \U$10374 ( \12137 , \12128 , \12131 );
and \U$10375 ( \12138 , \12124 , \12131 );
or \U$10376 ( \12139 , \12136 , \12137 , \12138 );
and \U$10377 ( \12140 , \12104 , \12118 );
xor \U$10378 ( \12141 , \12139 , \12140 );
and \U$10379 ( \12142 , \12108 , \12112 );
and \U$10380 ( \12143 , \12112 , \12117 );
and \U$10381 ( \12144 , \12108 , \12117 );
or \U$10382 ( \12145 , \12142 , \12143 , \12144 );
xor \U$10383 ( \12146 , \10998 , \11000 );
xor \U$10384 ( \12147 , \12145 , \12146 );
xor \U$10385 ( \12148 , \10974 , \10990 );
xor \U$10386 ( \12149 , \12148 , \10993 );
xor \U$10387 ( \12150 , \12147 , \12149 );
xor \U$10388 ( \12151 , \12141 , \12150 );
and \U$10389 ( \12152 , \12102 , \12119 );
and \U$10390 ( \12153 , \12119 , \12132 );
and \U$10391 ( \12154 , \12102 , \12132 );
or \U$10392 ( \12155 , \12152 , \12153 , \12154 );
nor \U$10393 ( \12156 , \12151 , \12155 );
nor \U$10394 ( \12157 , \12135 , \12156 );
and \U$10395 ( \12158 , \12145 , \12146 );
and \U$10396 ( \12159 , \12146 , \12149 );
and \U$10397 ( \12160 , \12145 , \12149 );
or \U$10398 ( \12161 , \12158 , \12159 , \12160 );
xor \U$10399 ( \12162 , \10861 , \10877 );
xor \U$10400 ( \12163 , \12162 , \10912 );
xor \U$10401 ( \12164 , \12161 , \12163 );
xor \U$10402 ( \12165 , \10996 , \11001 );
xor \U$10403 ( \12166 , \12165 , \11004 );
xor \U$10404 ( \12167 , \12164 , \12166 );
and \U$10405 ( \12168 , \12139 , \12140 );
and \U$10406 ( \12169 , \12140 , \12150 );
and \U$10407 ( \12170 , \12139 , \12150 );
or \U$10408 ( \12171 , \12168 , \12169 , \12170 );
nor \U$10409 ( \12172 , \12167 , \12171 );
xor \U$10410 ( \12173 , \11007 , \11008 );
xor \U$10411 ( \12174 , \12173 , \11011 );
and \U$10412 ( \12175 , \12161 , \12163 );
and \U$10413 ( \12176 , \12163 , \12166 );
and \U$10414 ( \12177 , \12161 , \12166 );
or \U$10415 ( \12178 , \12175 , \12176 , \12177 );
nor \U$10416 ( \12179 , \12174 , \12178 );
nor \U$10417 ( \12180 , \12172 , \12179 );
nand \U$10418 ( \12181 , \12157 , \12180 );
nor \U$10419 ( \12182 , \12098 , \12181 );
and \U$10420 ( \12183 , \10751 , \10436 );
and \U$10421 ( \12184 , \10682 , \10433 );
nor \U$10422 ( \12185 , \12183 , \12184 );
xnor \U$10423 ( \12186 , \12185 , \10430 );
and \U$10424 ( \12187 , \10558 , \12186 );
and \U$10425 ( \12188 , \10774 , \10472 );
and \U$10426 ( \12189 , \10730 , \10470 );
nor \U$10427 ( \12190 , \12188 , \12189 );
xnor \U$10428 ( \12191 , \12190 , \10498 );
and \U$10429 ( \12192 , \12186 , \12191 );
and \U$10430 ( \12193 , \10558 , \12191 );
or \U$10431 ( \12194 , \12187 , \12192 , \12193 );
and \U$10432 ( \12195 , \10682 , \10436 );
and \U$10433 ( \12196 , \10703 , \10433 );
nor \U$10434 ( \12197 , \12195 , \12196 );
xnor \U$10435 ( \12198 , \12197 , \10430 );
and \U$10436 ( \12199 , \10730 , \10472 );
and \U$10437 ( \12200 , \10751 , \10470 );
nor \U$10438 ( \12201 , \12199 , \12200 );
xnor \U$10439 ( \12202 , \12201 , \10498 );
xor \U$10440 ( \12203 , \12198 , \12202 );
and \U$10441 ( \12204 , \10907 , \10532 );
and \U$10442 ( \12205 , \10774 , \10530 );
nor \U$10443 ( \12206 , \12204 , \12205 );
xnor \U$10444 ( \12207 , \12206 , \10558 );
xor \U$10445 ( \12208 , \12203 , \12207 );
xor \U$10446 ( \12209 , \12194 , \12208 );
nand \U$10447 ( \12210 , \10907 , \10530 );
xnor \U$10448 ( \12211 , \12210 , \10558 );
xor \U$10449 ( \12212 , \10558 , \12186 );
xor \U$10450 ( \12213 , \12212 , \12191 );
and \U$10451 ( \12214 , \12211 , \12213 );
nor \U$10452 ( \12215 , \12209 , \12214 );
and \U$10453 ( \12216 , \12198 , \12202 );
and \U$10454 ( \12217 , \12202 , \12207 );
and \U$10455 ( \12218 , \12198 , \12207 );
or \U$10456 ( \12219 , \12216 , \12217 , \12218 );
xor \U$10457 ( \12220 , \11929 , \11931 );
xor \U$10458 ( \12221 , \12219 , \12220 );
xor \U$10459 ( \12222 , \10616 , \11917 );
xor \U$10460 ( \12223 , \12222 , \11922 );
xor \U$10461 ( \12224 , \12221 , \12223 );
and \U$10462 ( \12225 , \12194 , \12208 );
nor \U$10463 ( \12226 , \12224 , \12225 );
nor \U$10464 ( \12227 , \12215 , \12226 );
xor \U$10465 ( \12228 , \11840 , \11844 );
xor \U$10466 ( \12229 , \12228 , \11849 );
xor \U$10467 ( \12230 , \11925 , \11932 );
xor \U$10468 ( \12231 , \12230 , \11937 );
xor \U$10469 ( \12232 , \12229 , \12231 );
and \U$10470 ( \12233 , \12219 , \12220 );
and \U$10471 ( \12234 , \12220 , \12223 );
and \U$10472 ( \12235 , \12219 , \12223 );
or \U$10473 ( \12236 , \12233 , \12234 , \12235 );
nor \U$10474 ( \12237 , \12232 , \12236 );
xor \U$10475 ( \12238 , \11940 , \11942 );
and \U$10476 ( \12239 , \12229 , \12231 );
nor \U$10477 ( \12240 , \12238 , \12239 );
nor \U$10478 ( \12241 , \12237 , \12240 );
nand \U$10479 ( \12242 , \12227 , \12241 );
and \U$10480 ( \12243 , \10730 , \10436 );
and \U$10481 ( \12244 , \10751 , \10433 );
nor \U$10482 ( \12245 , \12243 , \12244 );
xnor \U$10483 ( \12246 , \12245 , \10430 );
and \U$10484 ( \12247 , \10907 , \10472 );
and \U$10485 ( \12248 , \10774 , \10470 );
nor \U$10486 ( \12249 , \12247 , \12248 );
xnor \U$10487 ( \12250 , \12249 , \10498 );
xor \U$10488 ( \12251 , \12246 , \12250 );
and \U$10489 ( \12252 , \10774 , \10436 );
and \U$10490 ( \12253 , \10730 , \10433 );
nor \U$10491 ( \12254 , \12252 , \12253 );
xnor \U$10492 ( \12255 , \12254 , \10430 );
and \U$10493 ( \12256 , \12255 , \10498 );
nor \U$10494 ( \12257 , \12251 , \12256 );
xor \U$10495 ( \12258 , \12211 , \12213 );
and \U$10496 ( \12259 , \12246 , \12250 );
nor \U$10497 ( \12260 , \12258 , \12259 );
nor \U$10498 ( \12261 , \12257 , \12260 );
xor \U$10499 ( \12262 , \12255 , \10498 );
nand \U$10500 ( \12263 , \10907 , \10470 );
xnor \U$10501 ( \12264 , \12263 , \10498 );
nor \U$10502 ( \12265 , \12262 , \12264 );
and \U$10503 ( \12266 , \10907 , \10436 );
and \U$10504 ( \12267 , \10774 , \10433 );
nor \U$10505 ( \12268 , \12266 , \12267 );
xnor \U$10506 ( \12269 , \12268 , \10430 );
nand \U$10507 ( \12270 , \10907 , \10433 );
xnor \U$10508 ( \12271 , \12270 , \10430 );
and \U$10509 ( \12272 , \12271 , \10430 );
nand \U$10510 ( \12273 , \12269 , \12272 );
or \U$10511 ( \12274 , \12265 , \12273 );
nand \U$10512 ( \12275 , \12262 , \12264 );
nand \U$10513 ( \12276 , \12274 , \12275 );
and \U$10514 ( \12277 , \12261 , \12276 );
nand \U$10515 ( \12278 , \12251 , \12256 );
or \U$10516 ( \12279 , \12260 , \12278 );
nand \U$10517 ( \12280 , \12258 , \12259 );
nand \U$10518 ( \12281 , \12279 , \12280 );
nor \U$10519 ( \12282 , \12277 , \12281 );
or \U$10520 ( \12283 , \12242 , \12282 );
nand \U$10521 ( \12284 , \12209 , \12214 );
or \U$10522 ( \12285 , \12226 , \12284 );
nand \U$10523 ( \12286 , \12224 , \12225 );
nand \U$10524 ( \12287 , \12285 , \12286 );
and \U$10525 ( \12288 , \12241 , \12287 );
nand \U$10526 ( \12289 , \12232 , \12236 );
or \U$10527 ( \12290 , \12240 , \12289 );
nand \U$10528 ( \12291 , \12238 , \12239 );
nand \U$10529 ( \12292 , \12290 , \12291 );
nor \U$10530 ( \12293 , \12288 , \12292 );
nand \U$10531 ( \12294 , \12283 , \12293 );
and \U$10532 ( \12295 , \12182 , \12294 );
nand \U$10533 ( \12296 , \11913 , \11943 );
or \U$10534 ( \12297 , \11989 , \12296 );
nand \U$10535 ( \12298 , \11984 , \11988 );
nand \U$10536 ( \12299 , \12297 , \12298 );
and \U$10537 ( \12300 , \12097 , \12299 );
nand \U$10538 ( \12301 , \12039 , \12040 );
or \U$10539 ( \12302 , \12096 , \12301 );
nand \U$10540 ( \12303 , \12094 , \12095 );
nand \U$10541 ( \12304 , \12302 , \12303 );
nor \U$10542 ( \12305 , \12300 , \12304 );
or \U$10543 ( \12306 , \12181 , \12305 );
nand \U$10544 ( \12307 , \12133 , \12134 );
or \U$10545 ( \12308 , \12156 , \12307 );
nand \U$10546 ( \12309 , \12151 , \12155 );
nand \U$10547 ( \12310 , \12308 , \12309 );
and \U$10548 ( \12311 , \12180 , \12310 );
nand \U$10549 ( \12312 , \12167 , \12171 );
or \U$10550 ( \12313 , \12179 , \12312 );
nand \U$10551 ( \12314 , \12174 , \12178 );
nand \U$10552 ( \12315 , \12313 , \12314 );
nor \U$10553 ( \12316 , \12311 , \12315 );
nand \U$10554 ( \12317 , \12306 , \12316 );
nor \U$10555 ( \12318 , \12295 , \12317 );
or \U$10556 ( \12319 , \11836 , \12318 );
nand \U$10557 ( \12320 , \10958 , \11014 );
or \U$10558 ( \12321 , \11090 , \12320 );
nand \U$10559 ( \12322 , \11088 , \11089 );
nand \U$10560 ( \12323 , \12321 , \12322 );
and \U$10561 ( \12324 , \11243 , \12323 );
nand \U$10562 ( \12325 , \11165 , \11166 );
or \U$10563 ( \12326 , \11242 , \12325 );
nand \U$10564 ( \12327 , \11237 , \11241 );
nand \U$10565 ( \12328 , \12326 , \12327 );
nor \U$10566 ( \12329 , \12324 , \12328 );
or \U$10567 ( \12330 , \11539 , \12329 );
nand \U$10568 ( \12331 , \11314 , \11318 );
or \U$10569 ( \12332 , \11395 , \12331 );
nand \U$10570 ( \12333 , \11390 , \11394 );
nand \U$10571 ( \12334 , \12332 , \12333 );
and \U$10572 ( \12335 , \11538 , \12334 );
nand \U$10573 ( \12336 , \11463 , \11467 );
or \U$10574 ( \12337 , \11537 , \12336 );
nand \U$10575 ( \12338 , \11532 , \11536 );
nand \U$10576 ( \12339 , \12337 , \12338 );
nor \U$10577 ( \12340 , \12335 , \12339 );
nand \U$10578 ( \12341 , \12330 , \12340 );
and \U$10579 ( \12342 , \11835 , \12341 );
nand \U$10580 ( \12343 , \11596 , \11600 );
or \U$10581 ( \12344 , \11661 , \12343 );
nand \U$10582 ( \12345 , \11656 , \11660 );
nand \U$10583 ( \12346 , \12344 , \12345 );
and \U$10584 ( \12347 , \11757 , \12346 );
nand \U$10585 ( \12348 , \11713 , \11717 );
or \U$10586 ( \12349 , \11756 , \12348 );
nand \U$10587 ( \12350 , \11751 , \11755 );
nand \U$10588 ( \12351 , \12349 , \12350 );
nor \U$10589 ( \12352 , \12347 , \12351 );
or \U$10590 ( \12353 , \11834 , \12352 );
nand \U$10591 ( \12354 , \11783 , \11787 );
or \U$10592 ( \12355 , \11809 , \12354 );
nand \U$10593 ( \12356 , \11804 , \11808 );
nand \U$10594 ( \12357 , \12355 , \12356 );
and \U$10595 ( \12358 , \11833 , \12357 );
nand \U$10596 ( \12359 , \11820 , \11824 );
or \U$10597 ( \12360 , \11832 , \12359 );
nand \U$10598 ( \12361 , \11827 , \11831 );
nand \U$10599 ( \12362 , \12360 , \12361 );
nor \U$10600 ( \12363 , \12358 , \12362 );
nand \U$10601 ( \12364 , \12353 , \12363 );
nor \U$10602 ( \12365 , \12342 , \12364 );
nand \U$10603 ( \12366 , \12319 , \12365 );
not \U$10604 ( \12367 , \12366 );
xor \U$10605 ( \12368 , \10426 , \12367 );
buf \U$10606 ( \12369 , \12368 );
buf \U$10611 ( \12370 , RI2b5e785db058_15);
buf \U$10612 ( \12371 , RI2b5e785dafe0_16);
buf \U$10613 ( \12372 , RI2b5e785daf68_17);
buf \U$10614 ( \12373 , RI2b5e785daef0_18);
buf \U$10615 ( \12374 , RI2b5e785dae78_19);
buf \U$10616 ( \12375 , RI2b5e785dae00_20);
buf \U$10617 ( \12376 , RI2b5e785dad88_21);
buf \U$10618 ( \12377 , RI2b5e785dad10_22);
buf \U$10619 ( \12378 , RI2b5e785dac98_23);
buf \U$10620 ( \12379 , RI2b5e785dac20_24);
buf \U$10621 ( \12380 , RI2b5e785daba8_25);
and \U$10622 ( \12381 , \12379 , \12380 );
and \U$10623 ( \12382 , \12378 , \12381 );
and \U$10624 ( \12383 , \12377 , \12382 );
and \U$10625 ( \12384 , \12376 , \12383 );
and \U$10626 ( \12385 , \12375 , \12384 );
and \U$10627 ( \12386 , \12374 , \12385 );
and \U$10628 ( \12387 , \12373 , \12386 );
and \U$10629 ( \12388 , \12372 , \12387 );
and \U$10630 ( \12389 , \12371 , \12388 );
xor \U$10631 ( \12390 , \12370 , \12389 );
buf \U$10632 ( \12391 , \12390 );
buf \U$10633 ( \12392 , \12391 );
buf \U$10634 ( \12393 , RI2b5e785ae3a0_613);
buf \U$10635 ( \12394 , RI2b5e785ae580_609);
buf \U$10636 ( \12395 , RI2b5e785ae5f8_608);
buf \U$10637 ( \12396 , RI2b5e785ae670_607);
buf \U$10638 ( \12397 , RI2b5e785ae6e8_606);
buf \U$10639 ( \12398 , RI2b5e785ae760_605);
buf \U$10640 ( \12399 , RI2b5e785ae7d8_604);
buf \U$10641 ( \12400 , RI2b5e785ae850_603);
buf \U$10642 ( \12401 , RI2b5e785ae8c8_602);
buf \U$10643 ( \12402 , RI2b5e785ae940_601);
buf \U$10644 ( \12403 , RI2b5e785ae3a0_613);
buf \U$10645 ( \12404 , RI2b5e785ae418_612);
buf \U$10646 ( \12405 , RI2b5e785ae490_611);
buf \U$10647 ( \12406 , RI2b5e785ae508_610);
and \U$10648 ( \12407 , \12403 , \12404 , \12405 , \12406 );
nor \U$10649 ( \12408 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12407 );
buf \U$10650 ( \12409 , \12408 );
buf \U$10651 ( \12410 , \12409 );
xor \U$10652 ( \12411 , \12393 , \12410 );
buf \U$10653 ( \12412 , \12411 );
buf \U$10654 ( \12413 , RI2b5e785ae418_612);
and \U$10655 ( \12414 , \12393 , \12410 );
xor \U$10656 ( \12415 , \12413 , \12414 );
buf \U$10657 ( \12416 , \12415 );
buf \U$10658 ( \12417 , RI2b5e785ae490_611);
and \U$10659 ( \12418 , \12413 , \12414 );
xor \U$10660 ( \12419 , \12417 , \12418 );
buf \U$10661 ( \12420 , \12419 );
buf \U$10662 ( \12421 , RI2b5e785ae508_610);
and \U$10663 ( \12422 , \12417 , \12418 );
xor \U$10664 ( \12423 , \12421 , \12422 );
buf \U$10665 ( \12424 , \12423 );
buf \U$10666 ( \12425 , RI2b5e785ae580_609);
and \U$10667 ( \12426 , \12421 , \12422 );
xor \U$10668 ( \12427 , \12425 , \12426 );
buf \U$10669 ( \12428 , \12427 );
not \U$10670 ( \12429 , \12428 );
nor \U$10671 ( \12430 , \12412 , \12416 , \12420 , \12424 , \12429 );
and \U$10672 ( \12431 , RI2b5e785daa40_28, \12430 );
and \U$10673 ( \12432 , \12412 , \12416 , \12420 , \12424 , \12429 );
and \U$10674 ( \12433 , RI2b5e78549540_41, \12432 );
not \U$10675 ( \12434 , \12412 );
and \U$10676 ( \12435 , \12434 , \12416 , \12420 , \12424 , \12429 );
and \U$10677 ( \12436 , RI2b5e785388a8_54, \12435 );
not \U$10678 ( \12437 , \12416 );
and \U$10679 ( \12438 , \12412 , \12437 , \12420 , \12424 , \12429 );
and \U$10680 ( \12439 , RI2b5e784a6330_67, \12438 );
and \U$10681 ( \12440 , \12434 , \12437 , \12420 , \12424 , \12429 );
and \U$10682 ( \12441 , RI2b5e78495698_80, \12440 );
not \U$10683 ( \12442 , \12420 );
and \U$10684 ( \12443 , \12412 , \12416 , \12442 , \12424 , \12429 );
and \U$10685 ( \12444 , RI2b5e78495080_93, \12443 );
and \U$10686 ( \12445 , \12434 , \12416 , \12442 , \12424 , \12429 );
and \U$10687 ( \12446 , RI2b5e78403b80_106, \12445 );
and \U$10688 ( \12447 , \12412 , \12437 , \12442 , \12424 , \12429 );
and \U$10689 ( \12448 , RI2b5e775b1e60_119, \12447 );
and \U$10690 ( \12449 , \12434 , \12437 , \12442 , \12424 , \12429 );
and \U$10691 ( \12450 , RI2b5e7750bdf8_132, \12449 );
nor \U$10692 ( \12451 , \12434 , \12437 , \12442 , \12424 , \12428 );
and \U$10693 ( \12452 , RI2b5e774ff5d0_145, \12451 );
nor \U$10694 ( \12453 , \12412 , \12437 , \12442 , \12424 , \12428 );
and \U$10695 ( \12454 , RI2b5e774f65e8_158, \12453 );
nor \U$10696 ( \12455 , \12434 , \12416 , \12442 , \12424 , \12428 );
and \U$10697 ( \12456 , RI2b5e774eabd0_171, \12455 );
nor \U$10698 ( \12457 , \12412 , \12416 , \12442 , \12424 , \12428 );
and \U$10699 ( \12458 , RI2b5e774de3a8_184, \12457 );
nor \U$10700 ( \12459 , \12434 , \12437 , \12420 , \12424 , \12428 );
and \U$10701 ( \12460 , RI2b5e774d53c0_197, \12459 );
nor \U$10702 ( \12461 , \12412 , \12437 , \12420 , \12424 , \12428 );
and \U$10703 ( \12462 , RI2b5e785f4300_210, \12461 );
nor \U$10704 ( \12463 , \12434 , \12416 , \12420 , \12424 , \12428 );
and \U$10705 ( \12464 , RI2b5e785f3ce8_223, \12463 );
nor \U$10706 ( \12465 , \12412 , \12416 , \12420 , \12424 , \12428 );
and \U$10707 ( \12466 , RI2b5e785eb0c0_236, \12465 );
or \U$10708 ( \12467 , \12431 , \12433 , \12436 , \12439 , \12441 , \12444 , \12446 , \12448 , \12450 , \12452 , \12454 , \12456 , \12458 , \12460 , \12462 , \12464 , \12466 );
buf \U$10709 ( \12468 , \12428 );
buf \U$10710 ( \12469 , \12412 );
buf \U$10711 ( \12470 , \12416 );
buf \U$10712 ( \12471 , \12420 );
buf \U$10713 ( \12472 , \12424 );
or \U$10714 ( \12473 , \12469 , \12470 , \12471 , \12472 );
and \U$10715 ( \12474 , \12468 , \12473 );
buf \U$10716 ( \12475 , \12474 );
_DC r39aa ( \12476_nR39aa , \12467 , \12475 );
buf \U$10717 ( \12477 , \12476_nR39aa );
not \U$10718 ( \12478 , \12477 );
xor \U$10719 ( \12479 , \12392 , \12478 );
xor \U$10720 ( \12480 , \12371 , \12388 );
buf \U$10721 ( \12481 , \12480 );
buf \U$10722 ( \12482 , \12481 );
and \U$10723 ( \12483 , RI2b5e785da9c8_29, \12430 );
and \U$10724 ( \12484 , RI2b5e785494c8_42, \12432 );
and \U$10725 ( \12485 , RI2b5e78538830_55, \12435 );
and \U$10726 ( \12486 , RI2b5e784a62b8_68, \12438 );
and \U$10727 ( \12487 , RI2b5e78495620_81, \12440 );
and \U$10728 ( \12488 , RI2b5e78495008_94, \12443 );
and \U$10729 ( \12489 , RI2b5e78403b08_107, \12445 );
and \U$10730 ( \12490 , RI2b5e775b1de8_120, \12447 );
and \U$10731 ( \12491 , RI2b5e7750bd80_133, \12449 );
and \U$10732 ( \12492 , RI2b5e774ff558_146, \12451 );
and \U$10733 ( \12493 , RI2b5e774f6570_159, \12453 );
and \U$10734 ( \12494 , RI2b5e774eab58_172, \12455 );
and \U$10735 ( \12495 , RI2b5e774de330_185, \12457 );
and \U$10736 ( \12496 , RI2b5e774d5348_198, \12459 );
and \U$10737 ( \12497 , RI2b5e785f4288_211, \12461 );
and \U$10738 ( \12498 , RI2b5e785f3658_224, \12463 );
and \U$10739 ( \12499 , RI2b5e785eb048_237, \12465 );
or \U$10740 ( \12500 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 );
_DC r3986 ( \12501_nR3986 , \12500 , \12475 );
buf \U$10741 ( \12502 , \12501_nR3986 );
not \U$10742 ( \12503 , \12502 );
and \U$10743 ( \12504 , \12482 , \12503 );
xor \U$10744 ( \12505 , \12372 , \12387 );
buf \U$10745 ( \12506 , \12505 );
buf \U$10746 ( \12507 , \12506 );
and \U$10747 ( \12508 , RI2b5e785da950_30, \12430 );
and \U$10748 ( \12509 , RI2b5e78549450_43, \12432 );
and \U$10749 ( \12510 , RI2b5e785387b8_56, \12435 );
and \U$10750 ( \12511 , RI2b5e784a6240_69, \12438 );
and \U$10751 ( \12512 , RI2b5e784955a8_82, \12440 );
and \U$10752 ( \12513 , RI2b5e78494f90_95, \12443 );
and \U$10753 ( \12514 , RI2b5e78403a90_108, \12445 );
and \U$10754 ( \12515 , RI2b5e775b1d70_121, \12447 );
and \U$10755 ( \12516 , RI2b5e7750bd08_134, \12449 );
and \U$10756 ( \12517 , RI2b5e774ff4e0_147, \12451 );
and \U$10757 ( \12518 , RI2b5e774f64f8_160, \12453 );
and \U$10758 ( \12519 , RI2b5e774eaae0_173, \12455 );
and \U$10759 ( \12520 , RI2b5e774de2b8_186, \12457 );
and \U$10760 ( \12521 , RI2b5e774d52d0_199, \12459 );
and \U$10761 ( \12522 , RI2b5e785f4210_212, \12461 );
and \U$10762 ( \12523 , RI2b5e785eb5e8_225, \12463 );
and \U$10763 ( \12524 , RI2b5e785e6c50_238, \12465 );
or \U$10764 ( \12525 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 );
_DC r37f3 ( \12526_nR37f3 , \12525 , \12475 );
buf \U$10765 ( \12527 , \12526_nR37f3 );
not \U$10766 ( \12528 , \12527 );
and \U$10767 ( \12529 , \12507 , \12528 );
xor \U$10768 ( \12530 , \12373 , \12386 );
buf \U$10769 ( \12531 , \12530 );
buf \U$10770 ( \12532 , \12531 );
and \U$10771 ( \12533 , RI2b5e785da8d8_31, \12430 );
and \U$10772 ( \12534 , RI2b5e785493d8_44, \12432 );
and \U$10773 ( \12535 , RI2b5e78538740_57, \12435 );
and \U$10774 ( \12536 , RI2b5e784a61c8_70, \12438 );
and \U$10775 ( \12537 , RI2b5e78495530_83, \12440 );
and \U$10776 ( \12538 , RI2b5e78494f18_96, \12443 );
and \U$10777 ( \12539 , RI2b5e78403a18_109, \12445 );
and \U$10778 ( \12540 , RI2b5e775b1cf8_122, \12447 );
and \U$10779 ( \12541 , RI2b5e7750bc90_135, \12449 );
and \U$10780 ( \12542 , RI2b5e774ff468_148, \12451 );
and \U$10781 ( \12543 , RI2b5e774f6480_161, \12453 );
and \U$10782 ( \12544 , RI2b5e774eaa68_174, \12455 );
and \U$10783 ( \12545 , RI2b5e774de240_187, \12457 );
and \U$10784 ( \12546 , RI2b5e774d5258_200, \12459 );
and \U$10785 ( \12547 , RI2b5e785f4198_213, \12461 );
and \U$10786 ( \12548 , RI2b5e785eb570_226, \12463 );
and \U$10787 ( \12549 , RI2b5e785e6bd8_239, \12465 );
or \U$10788 ( \12550 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 );
_DC r37cf ( \12551_nR37cf , \12550 , \12475 );
buf \U$10789 ( \12552 , \12551_nR37cf );
not \U$10790 ( \12553 , \12552 );
and \U$10791 ( \12554 , \12532 , \12553 );
xor \U$10792 ( \12555 , \12374 , \12385 );
buf \U$10793 ( \12556 , \12555 );
buf \U$10794 ( \12557 , \12556 );
and \U$10795 ( \12558 , RI2b5e785da860_32, \12430 );
and \U$10796 ( \12559 , RI2b5e78549360_45, \12432 );
and \U$10797 ( \12560 , RI2b5e785386c8_58, \12435 );
and \U$10798 ( \12561 , RI2b5e784a6150_71, \12438 );
and \U$10799 ( \12562 , RI2b5e784954b8_84, \12440 );
and \U$10800 ( \12563 , RI2b5e78494ea0_97, \12443 );
and \U$10801 ( \12564 , RI2b5e784039a0_110, \12445 );
and \U$10802 ( \12565 , RI2b5e775b1c80_123, \12447 );
and \U$10803 ( \12566 , RI2b5e7750bc18_136, \12449 );
and \U$10804 ( \12567 , RI2b5e774ff3f0_149, \12451 );
and \U$10805 ( \12568 , RI2b5e774f6408_162, \12453 );
and \U$10806 ( \12569 , RI2b5e774ea9f0_175, \12455 );
and \U$10807 ( \12570 , RI2b5e774de1c8_188, \12457 );
and \U$10808 ( \12571 , RI2b5e774d51e0_201, \12459 );
and \U$10809 ( \12572 , RI2b5e785f4120_214, \12461 );
and \U$10810 ( \12573 , RI2b5e785eb4f8_227, \12463 );
and \U$10811 ( \12574 , RI2b5e785e64d0_240, \12465 );
or \U$10812 ( \12575 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 );
_DC r3650 ( \12576_nR3650 , \12575 , \12475 );
buf \U$10813 ( \12577 , \12576_nR3650 );
not \U$10814 ( \12578 , \12577 );
and \U$10815 ( \12579 , \12557 , \12578 );
xor \U$10816 ( \12580 , \12375 , \12384 );
buf \U$10817 ( \12581 , \12580 );
buf \U$10818 ( \12582 , \12581 );
and \U$10819 ( \12583 , RI2b5e78549900_33, \12430 );
and \U$10820 ( \12584 , RI2b5e78538c68_46, \12432 );
and \U$10821 ( \12585 , RI2b5e78538650_59, \12435 );
and \U$10822 ( \12586 , RI2b5e784a60d8_72, \12438 );
and \U$10823 ( \12587 , RI2b5e78495440_85, \12440 );
and \U$10824 ( \12588 , RI2b5e78494e28_98, \12443 );
and \U$10825 ( \12589 , RI2b5e78403928_111, \12445 );
and \U$10826 ( \12590 , RI2b5e775b1c08_124, \12447 );
and \U$10827 ( \12591 , RI2b5e7750bba0_137, \12449 );
and \U$10828 ( \12592 , RI2b5e774ff378_150, \12451 );
and \U$10829 ( \12593 , RI2b5e774f6390_163, \12453 );
and \U$10830 ( \12594 , RI2b5e774ea978_176, \12455 );
and \U$10831 ( \12595 , RI2b5e774de150_189, \12457 );
and \U$10832 ( \12596 , RI2b5e774d5168_202, \12459 );
and \U$10833 ( \12597 , RI2b5e785f40a8_215, \12461 );
and \U$10834 ( \12598 , RI2b5e785eb480_228, \12463 );
and \U$10835 ( \12599 , RI2b5e785da608_241, \12465 );
or \U$10836 ( \12600 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 );
_DC r362c ( \12601_nR362c , \12600 , \12475 );
buf \U$10837 ( \12602 , \12601_nR362c );
not \U$10838 ( \12603 , \12602 );
and \U$10839 ( \12604 , \12582 , \12603 );
xor \U$10840 ( \12605 , \12376 , \12383 );
buf \U$10841 ( \12606 , \12605 );
buf \U$10842 ( \12607 , \12606 );
and \U$10843 ( \12608 , RI2b5e78549888_34, \12430 );
and \U$10844 ( \12609 , RI2b5e78538bf0_47, \12432 );
and \U$10845 ( \12610 , RI2b5e785385d8_60, \12435 );
and \U$10846 ( \12611 , RI2b5e784a6060_73, \12438 );
and \U$10847 ( \12612 , RI2b5e784953c8_86, \12440 );
and \U$10848 ( \12613 , RI2b5e78403ec8_99, \12443 );
and \U$10849 ( \12614 , RI2b5e775b21a8_112, \12445 );
and \U$10850 ( \12615 , RI2b5e775b1b90_125, \12447 );
and \U$10851 ( \12616 , RI2b5e7750bb28_138, \12449 );
and \U$10852 ( \12617 , RI2b5e774ff300_151, \12451 );
and \U$10853 ( \12618 , RI2b5e774f6318_164, \12453 );
and \U$10854 ( \12619 , RI2b5e774ea900_177, \12455 );
and \U$10855 ( \12620 , RI2b5e774de0d8_190, \12457 );
and \U$10856 ( \12621 , RI2b5e774d50f0_203, \12459 );
and \U$10857 ( \12622 , RI2b5e785f4030_216, \12461 );
and \U$10858 ( \12623 , RI2b5e785eb408_229, \12463 );
and \U$10859 ( \12624 , RI2b5e785da590_242, \12465 );
or \U$10860 ( \12625 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 );
_DC r34e1 ( \12626_nR34e1 , \12625 , \12475 );
buf \U$10861 ( \12627 , \12626_nR34e1 );
not \U$10862 ( \12628 , \12627 );
and \U$10863 ( \12629 , \12607 , \12628 );
xor \U$10864 ( \12630 , \12377 , \12382 );
buf \U$10865 ( \12631 , \12630 );
buf \U$10866 ( \12632 , \12631 );
and \U$10867 ( \12633 , RI2b5e78549810_35, \12430 );
and \U$10868 ( \12634 , RI2b5e78538b78_48, \12432 );
and \U$10869 ( \12635 , RI2b5e78538560_61, \12435 );
and \U$10870 ( \12636 , RI2b5e784a5fe8_74, \12438 );
and \U$10871 ( \12637 , RI2b5e78495350_87, \12440 );
and \U$10872 ( \12638 , RI2b5e78403e50_100, \12443 );
and \U$10873 ( \12639 , RI2b5e775b2130_113, \12445 );
and \U$10874 ( \12640 , RI2b5e775b1b18_126, \12447 );
and \U$10875 ( \12641 , RI2b5e7750bab0_139, \12449 );
and \U$10876 ( \12642 , RI2b5e774ff288_152, \12451 );
and \U$10877 ( \12643 , RI2b5e774f62a0_165, \12453 );
and \U$10878 ( \12644 , RI2b5e774ea888_178, \12455 );
and \U$10879 ( \12645 , RI2b5e774de060_191, \12457 );
and \U$10880 ( \12646 , RI2b5e774d5078_204, \12459 );
and \U$10881 ( \12647 , RI2b5e785f3fb8_217, \12461 );
and \U$10882 ( \12648 , RI2b5e785eb390_230, \12463 );
and \U$10883 ( \12649 , RI2b5e785da518_243, \12465 );
or \U$10884 ( \12650 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 );
_DC r34bd ( \12651_nR34bd , \12650 , \12475 );
buf \U$10885 ( \12652 , \12651_nR34bd );
not \U$10886 ( \12653 , \12652 );
and \U$10887 ( \12654 , \12632 , \12653 );
xor \U$10888 ( \12655 , \12378 , \12381 );
buf \U$10889 ( \12656 , \12655 );
buf \U$10890 ( \12657 , \12656 );
and \U$10891 ( \12658 , RI2b5e78549798_36, \12430 );
and \U$10892 ( \12659 , RI2b5e78538b00_49, \12432 );
and \U$10893 ( \12660 , RI2b5e785384e8_62, \12435 );
and \U$10894 ( \12661 , RI2b5e784a5f70_75, \12438 );
and \U$10895 ( \12662 , RI2b5e784952d8_88, \12440 );
and \U$10896 ( \12663 , RI2b5e78403dd8_101, \12443 );
and \U$10897 ( \12664 , RI2b5e775b20b8_114, \12445 );
and \U$10898 ( \12665 , RI2b5e775b1aa0_127, \12447 );
and \U$10899 ( \12666 , RI2b5e7750ba38_140, \12449 );
and \U$10900 ( \12667 , RI2b5e774ff210_153, \12451 );
and \U$10901 ( \12668 , RI2b5e774f6228_166, \12453 );
and \U$10902 ( \12669 , RI2b5e774ea810_179, \12455 );
and \U$10903 ( \12670 , RI2b5e774ddfe8_192, \12457 );
and \U$10904 ( \12671 , RI2b5e774d5000_205, \12459 );
and \U$10905 ( \12672 , RI2b5e785f3f40_218, \12461 );
and \U$10906 ( \12673 , RI2b5e785eb318_231, \12463 );
and \U$10907 ( \12674 , RI2b5e785da4a0_244, \12465 );
or \U$10908 ( \12675 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 );
_DC r33a2 ( \12676_nR33a2 , \12675 , \12475 );
buf \U$10909 ( \12677 , \12676_nR33a2 );
not \U$10910 ( \12678 , \12677 );
and \U$10911 ( \12679 , \12657 , \12678 );
xor \U$10912 ( \12680 , \12379 , \12380 );
buf \U$10913 ( \12681 , \12680 );
buf \U$10914 ( \12682 , \12681 );
and \U$10915 ( \12683 , RI2b5e78549720_37, \12430 );
and \U$10916 ( \12684 , RI2b5e78538a88_50, \12432 );
and \U$10917 ( \12685 , RI2b5e78538470_63, \12435 );
and \U$10918 ( \12686 , RI2b5e784a5ef8_76, \12438 );
and \U$10919 ( \12687 , RI2b5e78495260_89, \12440 );
and \U$10920 ( \12688 , RI2b5e78403d60_102, \12443 );
and \U$10921 ( \12689 , RI2b5e775b2040_115, \12445 );
and \U$10922 ( \12690 , RI2b5e775b1a28_128, \12447 );
and \U$10923 ( \12691 , RI2b5e7750b9c0_141, \12449 );
and \U$10924 ( \12692 , RI2b5e774ff198_154, \12451 );
and \U$10925 ( \12693 , RI2b5e774f61b0_167, \12453 );
and \U$10926 ( \12694 , RI2b5e774ea798_180, \12455 );
and \U$10927 ( \12695 , RI2b5e774ddf70_193, \12457 );
and \U$10928 ( \12696 , RI2b5e774d4f88_206, \12459 );
and \U$10929 ( \12697 , RI2b5e785f3ec8_219, \12461 );
and \U$10930 ( \12698 , RI2b5e785eb2a0_232, \12463 );
and \U$10931 ( \12699 , RI2b5e785da428_245, \12465 );
or \U$10932 ( \12700 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 );
_DC r33bb ( \12701_nR33bb , \12700 , \12475 );
buf \U$10933 ( \12702 , \12701_nR33bb );
not \U$10934 ( \12703 , \12702 );
and \U$10935 ( \12704 , \12682 , \12703 );
not \U$10936 ( \12705 , \12380 );
buf \U$10937 ( \12706 , \12705 );
buf \U$10938 ( \12707 , \12706 );
and \U$10939 ( \12708 , RI2b5e785496a8_38, \12430 );
and \U$10940 ( \12709 , RI2b5e78538a10_51, \12432 );
and \U$10941 ( \12710 , RI2b5e785383f8_64, \12435 );
and \U$10942 ( \12711 , RI2b5e784a5e80_77, \12438 );
and \U$10943 ( \12712 , RI2b5e784951e8_90, \12440 );
and \U$10944 ( \12713 , RI2b5e78403ce8_103, \12443 );
and \U$10945 ( \12714 , RI2b5e775b1fc8_116, \12445 );
and \U$10946 ( \12715 , RI2b5e775b19b0_129, \12447 );
and \U$10947 ( \12716 , RI2b5e7750b948_142, \12449 );
and \U$10948 ( \12717 , RI2b5e774ff120_155, \12451 );
and \U$10949 ( \12718 , RI2b5e774f6138_168, \12453 );
and \U$10950 ( \12719 , RI2b5e774ea720_181, \12455 );
and \U$10951 ( \12720 , RI2b5e774ddef8_194, \12457 );
and \U$10952 ( \12721 , RI2b5e774d4f10_207, \12459 );
and \U$10953 ( \12722 , RI2b5e785f3e50_220, \12461 );
and \U$10954 ( \12723 , RI2b5e785eb228_233, \12463 );
and \U$10955 ( \12724 , RI2b5e785da3b0_246, \12465 );
or \U$10956 ( \12725 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 );
_DC r32b8 ( \12726_nR32b8 , \12725 , \12475 );
buf \U$10957 ( \12727 , \12726_nR32b8 );
not \U$10958 ( \12728 , \12727 );
and \U$10959 ( \12729 , \12707 , \12728 );
buf \U$10960 ( \12730 , RI2b5e785dab30_26);
buf \U$10963 ( \12731 , \12730 );
and \U$10964 ( \12732 , RI2b5e78549630_39, \12430 );
and \U$10965 ( \12733 , RI2b5e78538998_52, \12432 );
and \U$10966 ( \12734 , RI2b5e78538380_65, \12435 );
and \U$10967 ( \12735 , RI2b5e784a5e08_78, \12438 );
and \U$10968 ( \12736 , RI2b5e78495170_91, \12440 );
and \U$10969 ( \12737 , RI2b5e78403c70_104, \12443 );
and \U$10970 ( \12738 , RI2b5e775b1f50_117, \12445 );
and \U$10971 ( \12739 , RI2b5e775b1938_130, \12447 );
and \U$10972 ( \12740 , RI2b5e7750b8d0_143, \12449 );
and \U$10973 ( \12741 , RI2b5e774ff0a8_156, \12451 );
and \U$10974 ( \12742 , RI2b5e774f60c0_169, \12453 );
and \U$10975 ( \12743 , RI2b5e774ea6a8_182, \12455 );
and \U$10976 ( \12744 , RI2b5e774dde80_195, \12457 );
and \U$10977 ( \12745 , RI2b5e774d4e98_208, \12459 );
and \U$10978 ( \12746 , RI2b5e785f3dd8_221, \12461 );
and \U$10979 ( \12747 , RI2b5e785eb1b0_234, \12463 );
and \U$10980 ( \12748 , RI2b5e785da338_247, \12465 );
or \U$10981 ( \12749 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 );
_DC r329c ( \12750_nR329c , \12749 , \12475 );
buf \U$10982 ( \12751 , \12750_nR329c );
not \U$10983 ( \12752 , \12751 );
or \U$10984 ( \12753 , \12731 , \12752 );
and \U$10985 ( \12754 , \12728 , \12753 );
and \U$10986 ( \12755 , \12707 , \12753 );
or \U$10987 ( \12756 , \12729 , \12754 , \12755 );
and \U$10988 ( \12757 , \12703 , \12756 );
and \U$10989 ( \12758 , \12682 , \12756 );
or \U$10990 ( \12759 , \12704 , \12757 , \12758 );
and \U$10991 ( \12760 , \12678 , \12759 );
and \U$10992 ( \12761 , \12657 , \12759 );
or \U$10993 ( \12762 , \12679 , \12760 , \12761 );
and \U$10994 ( \12763 , \12653 , \12762 );
and \U$10995 ( \12764 , \12632 , \12762 );
or \U$10996 ( \12765 , \12654 , \12763 , \12764 );
and \U$10997 ( \12766 , \12628 , \12765 );
and \U$10998 ( \12767 , \12607 , \12765 );
or \U$10999 ( \12768 , \12629 , \12766 , \12767 );
and \U$11000 ( \12769 , \12603 , \12768 );
and \U$11001 ( \12770 , \12582 , \12768 );
or \U$11002 ( \12771 , \12604 , \12769 , \12770 );
and \U$11003 ( \12772 , \12578 , \12771 );
and \U$11004 ( \12773 , \12557 , \12771 );
or \U$11005 ( \12774 , \12579 , \12772 , \12773 );
and \U$11006 ( \12775 , \12553 , \12774 );
and \U$11007 ( \12776 , \12532 , \12774 );
or \U$11008 ( \12777 , \12554 , \12775 , \12776 );
and \U$11009 ( \12778 , \12528 , \12777 );
and \U$11010 ( \12779 , \12507 , \12777 );
or \U$11011 ( \12780 , \12529 , \12778 , \12779 );
and \U$11012 ( \12781 , \12503 , \12780 );
and \U$11013 ( \12782 , \12482 , \12780 );
or \U$11014 ( \12783 , \12504 , \12781 , \12782 );
xor \U$11015 ( \12784 , \12479 , \12783 );
buf \U$11016 ( \12785 , \12784 );
buf \U$11017 ( \12786 , \12785 );
xor \U$11018 ( \12787 , \12482 , \12503 );
xor \U$11019 ( \12788 , \12787 , \12780 );
buf \U$11020 ( \12789 , \12788 );
buf \U$11021 ( \12790 , \12789 );
xor \U$11022 ( \12791 , \12507 , \12528 );
xor \U$11023 ( \12792 , \12791 , \12777 );
buf \U$11024 ( \12793 , \12792 );
buf \U$11025 ( \12794 , \12793 );
and \U$11026 ( \12795 , \12790 , \12794 );
not \U$11027 ( \12796 , \12795 );
and \U$11028 ( \12797 , \12786 , \12796 );
not \U$11029 ( \12798 , \12797 );
buf \U$11030 ( \12799 , \12412 );
buf \U$11031 ( \12800 , RI2b5e785ae5f8_608);
and \U$11032 ( \12801 , \12425 , \12426 );
xor \U$11033 ( \12802 , \12800 , \12801 );
buf \U$11034 ( \12803 , \12802 );
buf \U$11035 ( \12804 , \12803 );
buf \U$11036 ( \12805 , RI2b5e785ae670_607);
and \U$11037 ( \12806 , \12800 , \12801 );
xor \U$11038 ( \12807 , \12805 , \12806 );
buf \U$11039 ( \12808 , \12807 );
buf \U$11040 ( \12809 , \12808 );
buf \U$11041 ( \12810 , RI2b5e785ae6e8_606);
and \U$11042 ( \12811 , \12805 , \12806 );
xor \U$11043 ( \12812 , \12810 , \12811 );
buf \U$11044 ( \12813 , \12812 );
buf \U$11045 ( \12814 , \12813 );
buf \U$11046 ( \12815 , RI2b5e785ae760_605);
and \U$11047 ( \12816 , \12810 , \12811 );
xor \U$11048 ( \12817 , \12815 , \12816 );
buf \U$11049 ( \12818 , \12817 );
buf \U$11050 ( \12819 , \12818 );
buf \U$11051 ( \12820 , RI2b5e785ae7d8_604);
and \U$11052 ( \12821 , \12815 , \12816 );
xor \U$11053 ( \12822 , \12820 , \12821 );
buf \U$11054 ( \12823 , \12822 );
buf \U$11055 ( \12824 , \12823 );
buf \U$11056 ( \12825 , RI2b5e785ae850_603);
and \U$11057 ( \12826 , \12820 , \12821 );
xor \U$11058 ( \12827 , \12825 , \12826 );
buf \U$11059 ( \12828 , \12827 );
buf \U$11060 ( \12829 , \12828 );
buf \U$11061 ( \12830 , RI2b5e785ae8c8_602);
and \U$11062 ( \12831 , \12825 , \12826 );
xor \U$11063 ( \12832 , \12830 , \12831 );
buf \U$11064 ( \12833 , \12832 );
buf \U$11065 ( \12834 , \12833 );
buf \U$11066 ( \12835 , RI2b5e785ae940_601);
and \U$11067 ( \12836 , \12830 , \12831 );
xor \U$11068 ( \12837 , \12835 , \12836 );
buf \U$11069 ( \12838 , \12837 );
buf \U$11070 ( \12839 , \12838 );
buf \U$11071 ( \12840 , \12428 );
nor \U$11072 ( \12841 , \12804 , \12809 , \12814 , \12819 , \12824 , \12829 , \12834 , \12839 , \12840 );
buf \U$11073 ( \12842 , \12841 );
buf \U$11074 ( \12843 , \12842 );
xor \U$11075 ( \12844 , \12799 , \12843 );
buf \U$11076 ( \12845 , \12844 );
buf \U$11077 ( \12846 , \12416 );
and \U$11078 ( \12847 , \12799 , \12843 );
xor \U$11079 ( \12848 , \12846 , \12847 );
buf \U$11080 ( \12849 , \12848 );
buf \U$11081 ( \12850 , \12420 );
and \U$11082 ( \12851 , \12846 , \12847 );
xor \U$11083 ( \12852 , \12850 , \12851 );
buf \U$11084 ( \12853 , \12852 );
buf \U$11085 ( \12854 , \12424 );
and \U$11086 ( \12855 , \12850 , \12851 );
xor \U$11087 ( \12856 , \12854 , \12855 );
buf \U$11088 ( \12857 , \12856 );
buf \U$11089 ( \12858 , \12428 );
and \U$11090 ( \12859 , \12854 , \12855 );
xor \U$11091 ( \12860 , \12858 , \12859 );
buf \U$11092 ( \12861 , \12860 );
not \U$11093 ( \12862 , \12861 );
nor \U$11094 ( \12863 , \12845 , \12849 , \12853 , \12857 , \12862 );
and \U$11095 ( \12864 , RI2b5e785da248_249, \12863 );
and \U$11096 ( \12865 , \12845 , \12849 , \12853 , \12857 , \12862 );
and \U$11097 ( \12866 , RI2b5e785be750_269, \12865 );
not \U$11098 ( \12867 , \12845 );
and \U$11099 ( \12868 , \12867 , \12849 , \12853 , \12857 , \12862 );
and \U$11100 ( \12869 , RI2b5e785bc4a0_289, \12868 );
not \U$11101 ( \12870 , \12849 );
and \U$11102 ( \12871 , \12845 , \12870 , \12853 , \12857 , \12862 );
and \U$11103 ( \12872 , RI2b5e785bbb40_309, \12871 );
and \U$11104 ( \12873 , \12867 , \12870 , \12853 , \12857 , \12862 );
and \U$11105 ( \12874 , RI2b5e785b9c50_329, \12873 );
not \U$11106 ( \12875 , \12853 );
and \U$11107 ( \12876 , \12845 , \12849 , \12875 , \12857 , \12862 );
and \U$11108 ( \12877 , RI2b5e785b8120_349, \12876 );
and \U$11109 ( \12878 , \12867 , \12849 , \12875 , \12857 , \12862 );
and \U$11110 ( \12879 , RI2b5e785b77c0_369, \12878 );
and \U$11111 ( \12880 , \12845 , \12870 , \12875 , \12857 , \12862 );
and \U$11112 ( \12881 , RI2b5e785b6e60_389, \12880 );
and \U$11113 ( \12882 , \12867 , \12870 , \12875 , \12857 , \12862 );
and \U$11114 ( \12883 , RI2b5e785b56f0_409, \12882 );
nor \U$11115 ( \12884 , \12867 , \12870 , \12875 , \12857 , \12861 );
and \U$11116 ( \12885 , RI2b5e785b4d90_429, \12884 );
nor \U$11117 ( \12886 , \12845 , \12870 , \12875 , \12857 , \12861 );
and \U$11118 ( \12887 , RI2b5e785b39e0_449, \12886 );
nor \U$11119 ( \12888 , \12867 , \12849 , \12875 , \12857 , \12861 );
and \U$11120 ( \12889 , RI2b5e785b3080_469, \12888 );
nor \U$11121 ( \12890 , \12845 , \12849 , \12875 , \12857 , \12861 );
and \U$11122 ( \12891 , RI2b5e785b2720_489, \12890 );
nor \U$11123 ( \12892 , \12867 , \12870 , \12853 , \12857 , \12861 );
and \U$11124 ( \12893 , RI2b5e785b1730_509, \12892 );
nor \U$11125 ( \12894 , \12845 , \12870 , \12853 , \12857 , \12861 );
and \U$11126 ( \12895 , RI2b5e785b0dd0_529, \12894 );
nor \U$11127 ( \12896 , \12867 , \12849 , \12853 , \12857 , \12861 );
and \U$11128 ( \12897 , RI2b5e785b0470_549, \12896 );
nor \U$11129 ( \12898 , \12845 , \12849 , \12853 , \12857 , \12861 );
and \U$11130 ( \12899 , RI2b5e785af840_569, \12898 );
or \U$11131 ( \12900 , \12864 , \12866 , \12869 , \12872 , \12874 , \12877 , \12879 , \12881 , \12883 , \12885 , \12887 , \12889 , \12891 , \12893 , \12895 , \12897 , \12899 );
buf \U$11132 ( \12901 , \12861 );
buf \U$11133 ( \12902 , \12845 );
buf \U$11134 ( \12903 , \12849 );
buf \U$11135 ( \12904 , \12853 );
buf \U$11136 ( \12905 , \12857 );
or \U$11137 ( \12906 , \12902 , \12903 , \12904 , \12905 );
and \U$11138 ( \12907 , \12901 , \12906 );
buf \U$11139 ( \12908 , \12907 );
_DC r4084 ( \12909_nR4084 , \12900 , \12908 );
buf \U$11140 ( \12910 , \12909_nR4084 );
buf \U$11141 ( \12911 , RI2b5e785db0d0_14);
and \U$11142 ( \12912 , \12370 , \12389 );
and \U$11143 ( \12913 , \12911 , \12912 );
buf \U$11144 ( \12914 , \12913 );
buf \U$11145 ( \12915 , \12914 );
xor \U$11146 ( \12916 , \12911 , \12912 );
buf \U$11147 ( \12917 , \12916 );
buf \U$11148 ( \12918 , \12917 );
and \U$11149 ( \12919 , RI2b5e785daab8_27, \12430 );
and \U$11150 ( \12920 , RI2b5e785495b8_40, \12432 );
and \U$11151 ( \12921 , RI2b5e78538920_53, \12435 );
and \U$11152 ( \12922 , RI2b5e784a63a8_66, \12438 );
and \U$11153 ( \12923 , RI2b5e78495710_79, \12440 );
and \U$11154 ( \12924 , RI2b5e784950f8_92, \12443 );
and \U$11155 ( \12925 , RI2b5e78403bf8_105, \12445 );
and \U$11156 ( \12926 , RI2b5e775b1ed8_118, \12447 );
and \U$11157 ( \12927 , RI2b5e775b18c0_131, \12449 );
and \U$11158 ( \12928 , RI2b5e7750b858_144, \12451 );
and \U$11159 ( \12929 , RI2b5e774ff030_157, \12453 );
and \U$11160 ( \12930 , RI2b5e774f6048_170, \12455 );
and \U$11161 ( \12931 , RI2b5e774ea630_183, \12457 );
and \U$11162 ( \12932 , RI2b5e774dde08_196, \12459 );
and \U$11163 ( \12933 , RI2b5e774d4e20_209, \12461 );
and \U$11164 ( \12934 , RI2b5e785f3d60_222, \12463 );
and \U$11165 ( \12935 , RI2b5e785eb138_235, \12465 );
or \U$11166 ( \12936 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 );
_DC r3b65 ( \12937_nR3b65 , \12936 , \12475 );
buf \U$11167 ( \12938 , \12937_nR3b65 );
not \U$11168 ( \12939 , \12938 );
and \U$11169 ( \12940 , \12918 , \12939 );
and \U$11170 ( \12941 , \12392 , \12478 );
and \U$11171 ( \12942 , \12478 , \12783 );
and \U$11172 ( \12943 , \12392 , \12783 );
or \U$11173 ( \12944 , \12941 , \12942 , \12943 );
and \U$11174 ( \12945 , \12939 , \12944 );
and \U$11175 ( \12946 , \12918 , \12944 );
or \U$11176 ( \12947 , \12940 , \12945 , \12946 );
xnor \U$11177 ( \12948 , \12915 , \12947 );
buf \U$11178 ( \12949 , \12948 );
buf \U$11179 ( \12950 , \12949 );
xor \U$11180 ( \12951 , \12918 , \12939 );
xor \U$11181 ( \12952 , \12951 , \12944 );
buf \U$11182 ( \12953 , \12952 );
buf \U$11183 ( \12954 , \12953 );
xor \U$11184 ( \12955 , \12950 , \12954 );
xor \U$11185 ( \12956 , \12954 , \12786 );
not \U$11186 ( \12957 , \12956 );
and \U$11187 ( \12958 , \12955 , \12957 );
and \U$11188 ( \12959 , \12910 , \12958 );
and \U$11189 ( \12960 , RI2b5e785da2c0_248, \12863 );
and \U$11190 ( \12961 , RI2b5e785be7c8_268, \12865 );
and \U$11191 ( \12962 , RI2b5e785bc518_288, \12868 );
and \U$11192 ( \12963 , RI2b5e785bbbb8_308, \12871 );
and \U$11193 ( \12964 , RI2b5e785b9cc8_328, \12873 );
and \U$11194 ( \12965 , RI2b5e785b9368_348, \12876 );
and \U$11195 ( \12966 , RI2b5e785b7838_368, \12878 );
and \U$11196 ( \12967 , RI2b5e785b6ed8_388, \12880 );
and \U$11197 ( \12968 , RI2b5e785b5768_408, \12882 );
and \U$11198 ( \12969 , RI2b5e785b4e08_428, \12884 );
and \U$11199 ( \12970 , RI2b5e785b3a58_448, \12886 );
and \U$11200 ( \12971 , RI2b5e785b30f8_468, \12888 );
and \U$11201 ( \12972 , RI2b5e785b2798_488, \12890 );
and \U$11202 ( \12973 , RI2b5e785b17a8_508, \12892 );
and \U$11203 ( \12974 , RI2b5e785b0e48_528, \12894 );
and \U$11204 ( \12975 , RI2b5e785b04e8_548, \12896 );
and \U$11205 ( \12976 , RI2b5e785afb88_568, \12898 );
or \U$11206 ( \12977 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 );
_DC r4179 ( \12978_nR4179 , \12977 , \12908 );
buf \U$11207 ( \12979 , \12978_nR4179 );
and \U$11208 ( \12980 , \12979 , \12956 );
nor \U$11209 ( \12981 , \12959 , \12980 );
and \U$11210 ( \12982 , \12954 , \12786 );
not \U$11211 ( \12983 , \12982 );
and \U$11212 ( \12984 , \12950 , \12983 );
xnor \U$11213 ( \12985 , \12981 , \12984 );
xor \U$11214 ( \12986 , \12798 , \12985 );
and \U$11216 ( \12987 , RI2b5e785da1d0_250, \12863 );
and \U$11217 ( \12988 , RI2b5e785be6d8_270, \12865 );
and \U$11218 ( \12989 , RI2b5e785bc428_290, \12868 );
and \U$11219 ( \12990 , RI2b5e785bbac8_310, \12871 );
and \U$11220 ( \12991 , RI2b5e785b9bd8_330, \12873 );
and \U$11221 ( \12992 , RI2b5e785b80a8_350, \12876 );
and \U$11222 ( \12993 , RI2b5e785b7748_370, \12878 );
and \U$11223 ( \12994 , RI2b5e785b6de8_390, \12880 );
and \U$11224 ( \12995 , RI2b5e785b5678_410, \12882 );
and \U$11225 ( \12996 , RI2b5e785b4d18_430, \12884 );
and \U$11226 ( \12997 , RI2b5e785b3968_450, \12886 );
and \U$11227 ( \12998 , RI2b5e785b3008_470, \12888 );
and \U$11228 ( \12999 , RI2b5e785b26a8_490, \12890 );
and \U$11229 ( \13000 , RI2b5e785b16b8_510, \12892 );
and \U$11230 ( \13001 , RI2b5e785b0d58_530, \12894 );
and \U$11231 ( \13002 , RI2b5e785b03f8_550, \12896 );
and \U$11232 ( \13003 , RI2b5e785af7c8_570, \12898 );
or \U$11233 ( \13004 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 );
_DC r3fbb ( \13005_nR3fbb , \13004 , \12908 );
buf \U$11234 ( \13006 , \13005_nR3fbb );
or \U$11235 ( \13007 , \12915 , \12947 );
not \U$11236 ( \13008 , \13007 );
buf \U$11237 ( \13009 , \13008 );
buf \U$11238 ( \13010 , \13009 );
xor \U$11239 ( \13011 , \13010 , \12950 );
and \U$11240 ( \13012 , \13006 , \13011 );
nor \U$11241 ( \13013 , 1'b0 , \13012 );
xnor \U$11243 ( \13014 , \13013 , 1'b0 );
xor \U$11244 ( \13015 , \12986 , \13014 );
xor \U$11245 ( \13016 , 1'b0 , \13015 );
xor \U$11247 ( \13017 , \12786 , \12790 );
xor \U$11248 ( \13018 , \12790 , \12794 );
not \U$11249 ( \13019 , \13018 );
and \U$11250 ( \13020 , \13017 , \13019 );
and \U$11251 ( \13021 , \12979 , \13020 );
not \U$11252 ( \13022 , \13021 );
xnor \U$11253 ( \13023 , \13022 , \12797 );
and \U$11254 ( \13024 , \13006 , \12958 );
and \U$11255 ( \13025 , \12910 , \12956 );
nor \U$11256 ( \13026 , \13024 , \13025 );
xnor \U$11257 ( \13027 , \13026 , \12984 );
and \U$11258 ( \13028 , \13023 , \13027 );
or \U$11260 ( \13029 , 1'b0 , \13028 , 1'b0 );
xor \U$11262 ( \13030 , \13029 , 1'b0 );
xor \U$11264 ( \13031 , \13030 , 1'b0 );
and \U$11265 ( \13032 , \13016 , \13031 );
or \U$11266 ( \13033 , 1'b0 , 1'b0 , \13032 );
and \U$11269 ( \13034 , \12979 , \12958 );
not \U$11270 ( \13035 , \13034 );
xnor \U$11271 ( \13036 , \13035 , \12984 );
xor \U$11272 ( \13037 , 1'b0 , \13036 );
and \U$11274 ( \13038 , \12910 , \13011 );
nor \U$11275 ( \13039 , 1'b0 , \13038 );
xnor \U$11276 ( \13040 , \13039 , 1'b0 );
xor \U$11277 ( \13041 , \13037 , \13040 );
xor \U$11278 ( \13042 , 1'b0 , \13041 );
xor \U$11280 ( \13043 , \13042 , 1'b1 );
and \U$11281 ( \13044 , \12798 , \12985 );
and \U$11282 ( \13045 , \12985 , \13014 );
and \U$11283 ( \13046 , \12798 , \13014 );
or \U$11284 ( \13047 , \13044 , \13045 , \13046 );
xor \U$11286 ( \13048 , \13047 , 1'b0 );
xor \U$11288 ( \13049 , \13048 , 1'b0 );
xor \U$11289 ( \13050 , \13043 , \13049 );
and \U$11290 ( \13051 , \13033 , \13050 );
or \U$11292 ( \13052 , 1'b0 , \13051 , 1'b0 );
xor \U$11294 ( \13053 , \13052 , 1'b0 );
and \U$11296 ( \13054 , \13042 , 1'b1 );
and \U$11297 ( \13055 , 1'b1 , \13049 );
and \U$11298 ( \13056 , \13042 , \13049 );
or \U$11299 ( \13057 , \13054 , \13055 , \13056 );
xor \U$11300 ( \13058 , 1'b0 , \13057 );
not \U$11302 ( \13059 , \12984 );
and \U$11304 ( \13060 , \12979 , \13011 );
nor \U$11305 ( \13061 , 1'b0 , \13060 );
xnor \U$11306 ( \13062 , \13061 , 1'b0 );
xor \U$11307 ( \13063 , \13059 , \13062 );
xor \U$11309 ( \13064 , \13063 , 1'b0 );
xor \U$11310 ( \13065 , 1'b0 , \13064 );
xor \U$11312 ( \13066 , \13065 , 1'b0 );
and \U$11314 ( \13067 , \13036 , \13040 );
or \U$11316 ( \13068 , 1'b0 , \13067 , 1'b0 );
xor \U$11318 ( \13069 , \13068 , 1'b0 );
xor \U$11320 ( \13070 , \13069 , 1'b0 );
xor \U$11321 ( \13071 , \13066 , \13070 );
xor \U$11322 ( \13072 , \13058 , \13071 );
xor \U$11323 ( \13073 , \13053 , \13072 );
xor \U$11329 ( \13074 , \12532 , \12553 );
xor \U$11330 ( \13075 , \13074 , \12774 );
buf \U$11331 ( \13076 , \13075 );
buf \U$11332 ( \13077 , \13076 );
xor \U$11333 ( \13078 , \12794 , \13077 );
xor \U$11334 ( \13079 , \12557 , \12578 );
xor \U$11335 ( \13080 , \13079 , \12771 );
buf \U$11336 ( \13081 , \13080 );
buf \U$11337 ( \13082 , \13081 );
xor \U$11338 ( \13083 , \13077 , \13082 );
not \U$11339 ( \13084 , \13083 );
and \U$11340 ( \13085 , \13078 , \13084 );
and \U$11341 ( \13086 , \12979 , \13085 );
not \U$11342 ( \13087 , \13086 );
and \U$11343 ( \13088 , \13077 , \13082 );
not \U$11344 ( \13089 , \13088 );
and \U$11345 ( \13090 , \12794 , \13089 );
xnor \U$11346 ( \13091 , \13087 , \13090 );
and \U$11347 ( \13092 , \13006 , \13020 );
and \U$11348 ( \13093 , \12910 , \13018 );
nor \U$11349 ( \13094 , \13092 , \13093 );
xnor \U$11350 ( \13095 , \13094 , \12797 );
and \U$11351 ( \13096 , \13091 , \13095 );
or \U$11353 ( \13097 , 1'b0 , \13096 , 1'b0 );
and \U$11354 ( \13098 , RI2b5e785da0e0_252, \12863 );
and \U$11355 ( \13099 , RI2b5e785be5e8_272, \12865 );
and \U$11356 ( \13100 , RI2b5e785bc338_292, \12868 );
and \U$11357 ( \13101 , RI2b5e785bb9d8_312, \12871 );
and \U$11358 ( \13102 , RI2b5e785b9ae8_332, \12873 );
and \U$11359 ( \13103 , RI2b5e785b7fb8_352, \12876 );
and \U$11360 ( \13104 , RI2b5e785b7658_372, \12878 );
and \U$11361 ( \13105 , RI2b5e785b5ee8_392, \12880 );
and \U$11362 ( \13106 , RI2b5e785b5588_412, \12882 );
and \U$11363 ( \13107 , RI2b5e785b4c28_432, \12884 );
and \U$11364 ( \13108 , RI2b5e785b3878_452, \12886 );
and \U$11365 ( \13109 , RI2b5e785b2f18_472, \12888 );
and \U$11366 ( \13110 , RI2b5e785b25b8_492, \12890 );
and \U$11367 ( \13111 , RI2b5e785b15c8_512, \12892 );
and \U$11368 ( \13112 , RI2b5e785b0c68_532, \12894 );
and \U$11369 ( \13113 , RI2b5e785b0308_552, \12896 );
and \U$11370 ( \13114 , RI2b5e785af6d8_572, \12898 );
or \U$11371 ( \13115 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 );
_DC r3e1c ( \13116_nR3e1c , \13115 , \12908 );
buf \U$11372 ( \13117 , \13116_nR3e1c );
and \U$11373 ( \13118 , \13117 , \12958 );
and \U$11374 ( \13119 , RI2b5e785da158_251, \12863 );
and \U$11375 ( \13120 , RI2b5e785be660_271, \12865 );
and \U$11376 ( \13121 , RI2b5e785bc3b0_291, \12868 );
and \U$11377 ( \13122 , RI2b5e785bba50_311, \12871 );
and \U$11378 ( \13123 , RI2b5e785b9b60_331, \12873 );
and \U$11379 ( \13124 , RI2b5e785b8030_351, \12876 );
and \U$11380 ( \13125 , RI2b5e785b76d0_371, \12878 );
and \U$11381 ( \13126 , RI2b5e785b6d70_391, \12880 );
and \U$11382 ( \13127 , RI2b5e785b5600_411, \12882 );
and \U$11383 ( \13128 , RI2b5e785b4ca0_431, \12884 );
and \U$11384 ( \13129 , RI2b5e785b38f0_451, \12886 );
and \U$11385 ( \13130 , RI2b5e785b2f90_471, \12888 );
and \U$11386 ( \13131 , RI2b5e785b2630_491, \12890 );
and \U$11387 ( \13132 , RI2b5e785b1640_511, \12892 );
and \U$11388 ( \13133 , RI2b5e785b0ce0_531, \12894 );
and \U$11389 ( \13134 , RI2b5e785b0380_551, \12896 );
and \U$11390 ( \13135 , RI2b5e785af750_571, \12898 );
or \U$11391 ( \13136 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 );
_DC r3efa ( \13137_nR3efa , \13136 , \12908 );
buf \U$11392 ( \13138 , \13137_nR3efa );
and \U$11393 ( \13139 , \13138 , \12956 );
nor \U$11394 ( \13140 , \13118 , \13139 );
xnor \U$11395 ( \13141 , \13140 , \12984 );
and \U$11397 ( \13142 , RI2b5e785da068_253, \12863 );
and \U$11398 ( \13143 , RI2b5e785be570_273, \12865 );
and \U$11399 ( \13144 , RI2b5e785bc2c0_293, \12868 );
and \U$11400 ( \13145 , RI2b5e785bb960_313, \12871 );
and \U$11401 ( \13146 , RI2b5e785b9a70_333, \12873 );
and \U$11402 ( \13147 , RI2b5e785b7f40_353, \12876 );
and \U$11403 ( \13148 , RI2b5e785b75e0_373, \12878 );
and \U$11404 ( \13149 , RI2b5e785b5e70_393, \12880 );
and \U$11405 ( \13150 , RI2b5e785b5510_413, \12882 );
and \U$11406 ( \13151 , RI2b5e785b4bb0_433, \12884 );
and \U$11407 ( \13152 , RI2b5e785b3800_453, \12886 );
and \U$11408 ( \13153 , RI2b5e785b2ea0_473, \12888 );
and \U$11409 ( \13154 , RI2b5e785b2540_493, \12890 );
and \U$11410 ( \13155 , RI2b5e785b1550_513, \12892 );
and \U$11411 ( \13156 , RI2b5e785b0bf0_533, \12894 );
and \U$11412 ( \13157 , RI2b5e785b0290_553, \12896 );
and \U$11413 ( \13158 , RI2b5e785af660_573, \12898 );
or \U$11414 ( \13159 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 );
_DC r3d33 ( \13160_nR3d33 , \13159 , \12908 );
buf \U$11415 ( \13161 , \13160_nR3d33 );
and \U$11416 ( \13162 , \13161 , \13011 );
nor \U$11417 ( \13163 , 1'b0 , \13162 );
xnor \U$11418 ( \13164 , \13163 , 1'b0 );
and \U$11419 ( \13165 , \13141 , \13164 );
or \U$11422 ( \13166 , \13165 , 1'b0 , 1'b0 );
and \U$11423 ( \13167 , \13097 , \13166 );
or \U$11426 ( \13168 , \13167 , 1'b0 , 1'b0 );
and \U$11429 ( \13169 , \13117 , \13011 );
nor \U$11430 ( \13170 , 1'b0 , \13169 );
xnor \U$11431 ( \13171 , \13170 , 1'b0 );
xor \U$11433 ( \13172 , \13171 , 1'b0 );
xor \U$11435 ( \13173 , \13172 , 1'b0 );
not \U$11436 ( \13174 , \13090 );
and \U$11437 ( \13175 , \12910 , \13020 );
and \U$11438 ( \13176 , \12979 , \13018 );
nor \U$11439 ( \13177 , \13175 , \13176 );
xnor \U$11440 ( \13178 , \13177 , \12797 );
xor \U$11441 ( \13179 , \13174 , \13178 );
and \U$11442 ( \13180 , \13138 , \12958 );
and \U$11443 ( \13181 , \13006 , \12956 );
nor \U$11444 ( \13182 , \13180 , \13181 );
xnor \U$11445 ( \13183 , \13182 , \12984 );
xor \U$11446 ( \13184 , \13179 , \13183 );
and \U$11447 ( \13185 , \13173 , \13184 );
or \U$11449 ( \13186 , 1'b0 , \13185 , 1'b0 );
and \U$11450 ( \13187 , \13168 , \13186 );
or \U$11451 ( \13188 , 1'b0 , 1'b0 , \13187 );
and \U$11453 ( \13189 , \13138 , \13011 );
nor \U$11454 ( \13190 , 1'b0 , \13189 );
xnor \U$11455 ( \13191 , \13190 , 1'b0 );
xor \U$11457 ( \13192 , \13191 , 1'b0 );
xor \U$11459 ( \13193 , \13192 , 1'b0 );
xor \U$11461 ( \13194 , 1'b0 , \13023 );
xor \U$11462 ( \13195 , \13194 , \13027 );
xor \U$11463 ( \13196 , \13193 , \13195 );
and \U$11465 ( \13197 , \13196 , 1'b1 );
and \U$11466 ( \13198 , \13174 , \13178 );
and \U$11467 ( \13199 , \13178 , \13183 );
and \U$11468 ( \13200 , \13174 , \13183 );
or \U$11469 ( \13201 , \13198 , \13199 , \13200 );
xor \U$11471 ( \13202 , \13201 , 1'b0 );
xor \U$11473 ( \13203 , \13202 , 1'b0 );
and \U$11474 ( \13204 , 1'b1 , \13203 );
and \U$11475 ( \13205 , \13196 , \13203 );
or \U$11476 ( \13206 , \13197 , \13204 , \13205 );
and \U$11477 ( \13207 , \13188 , \13206 );
xor \U$11479 ( \13208 , \13016 , 1'b0 );
xor \U$11480 ( \13209 , \13208 , \13031 );
and \U$11481 ( \13210 , \13206 , \13209 );
and \U$11482 ( \13211 , \13188 , \13209 );
or \U$11483 ( \13212 , \13207 , \13210 , \13211 );
xor \U$11485 ( \13213 , 1'b0 , \13033 );
xor \U$11486 ( \13214 , \13213 , \13050 );
and \U$11487 ( \13215 , \13212 , \13214 );
or \U$11488 ( \13216 , 1'b0 , 1'b0 , \13215 );
nand \U$11489 ( \13217 , \13073 , \13216 );
nor \U$11490 ( \13218 , \13073 , \13216 );
not \U$11491 ( \13219 , \13218 );
nand \U$11492 ( \13220 , \13217 , \13219 );
xor \U$11493 ( \13221 , \12707 , \12728 );
xor \U$11494 ( \13222 , \13221 , \12753 );
buf \U$11495 ( \13223 , \13222 );
buf \U$11496 ( \13224 , \13223 );
xor \U$11497 ( \13225 , \12731 , \12751 );
buf \U$11498 ( \13226 , \13225 );
buf \U$11499 ( \13227 , \13226 );
xor \U$11500 ( \13228 , \13224 , \13227 );
not \U$11501 ( \13229 , \13227 );
and \U$11502 ( \13230 , \13228 , \13229 );
and \U$11503 ( \13231 , \13161 , \13230 );
and \U$11504 ( \13232 , \13117 , \13227 );
nor \U$11505 ( \13233 , \13231 , \13232 );
xnor \U$11506 ( \13234 , \13233 , \13224 );
and \U$11507 ( \13235 , RI2b5e785c2bc0_255, \12863 );
and \U$11508 ( \13236 , RI2b5e785be480_275, \12865 );
and \U$11509 ( \13237 , RI2b5e785bc1d0_295, \12868 );
and \U$11510 ( \13238 , RI2b5e785ba2e0_315, \12871 );
and \U$11511 ( \13239 , RI2b5e785b9980_335, \12873 );
and \U$11512 ( \13240 , RI2b5e785b7e50_355, \12876 );
and \U$11513 ( \13241 , RI2b5e785b74f0_375, \12878 );
and \U$11514 ( \13242 , RI2b5e785b5d80_395, \12880 );
and \U$11515 ( \13243 , RI2b5e785b5420_415, \12882 );
and \U$11516 ( \13244 , RI2b5e785b4ac0_435, \12884 );
and \U$11517 ( \13245 , RI2b5e785b3710_455, \12886 );
and \U$11518 ( \13246 , RI2b5e785b2db0_475, \12888 );
and \U$11519 ( \13247 , RI2b5e785b2450_495, \12890 );
and \U$11520 ( \13248 , RI2b5e785b1460_515, \12892 );
and \U$11521 ( \13249 , RI2b5e785b0b00_535, \12894 );
and \U$11522 ( \13250 , RI2b5e785b01a0_555, \12896 );
and \U$11523 ( \13251 , RI2b5e785af570_575, \12898 );
or \U$11524 ( \13252 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 );
_DC r3ba2 ( \13253_nR3ba2 , \13252 , \12908 );
buf \U$11525 ( \13254 , \13253_nR3ba2 );
xor \U$11526 ( \13255 , \12657 , \12678 );
xor \U$11527 ( \13256 , \13255 , \12759 );
buf \U$11528 ( \13257 , \13256 );
buf \U$11529 ( \13258 , \13257 );
xor \U$11530 ( \13259 , \12682 , \12703 );
xor \U$11531 ( \13260 , \13259 , \12756 );
buf \U$11532 ( \13261 , \13260 );
buf \U$11533 ( \13262 , \13261 );
xor \U$11534 ( \13263 , \13258 , \13262 );
xor \U$11535 ( \13264 , \13262 , \13224 );
not \U$11536 ( \13265 , \13264 );
and \U$11537 ( \13266 , \13263 , \13265 );
and \U$11538 ( \13267 , \13254 , \13266 );
and \U$11539 ( \13268 , RI2b5e785c2c38_254, \12863 );
and \U$11540 ( \13269 , RI2b5e785be4f8_274, \12865 );
and \U$11541 ( \13270 , RI2b5e785bc248_294, \12868 );
and \U$11542 ( \13271 , RI2b5e785ba358_314, \12871 );
and \U$11543 ( \13272 , RI2b5e785b99f8_334, \12873 );
and \U$11544 ( \13273 , RI2b5e785b7ec8_354, \12876 );
and \U$11545 ( \13274 , RI2b5e785b7568_374, \12878 );
and \U$11546 ( \13275 , RI2b5e785b5df8_394, \12880 );
and \U$11547 ( \13276 , RI2b5e785b5498_414, \12882 );
and \U$11548 ( \13277 , RI2b5e785b4b38_434, \12884 );
and \U$11549 ( \13278 , RI2b5e785b3788_454, \12886 );
and \U$11550 ( \13279 , RI2b5e785b2e28_474, \12888 );
and \U$11551 ( \13280 , RI2b5e785b24c8_494, \12890 );
and \U$11552 ( \13281 , RI2b5e785b14d8_514, \12892 );
and \U$11553 ( \13282 , RI2b5e785b0b78_534, \12894 );
and \U$11554 ( \13283 , RI2b5e785b0218_554, \12896 );
and \U$11555 ( \13284 , RI2b5e785af5e8_574, \12898 );
or \U$11556 ( \13285 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 );
_DC r3c4f ( \13286_nR3c4f , \13285 , \12908 );
buf \U$11557 ( \13287 , \13286_nR3c4f );
and \U$11558 ( \13288 , \13287 , \13264 );
nor \U$11559 ( \13289 , \13267 , \13288 );
and \U$11560 ( \13290 , \13262 , \13224 );
not \U$11561 ( \13291 , \13290 );
and \U$11562 ( \13292 , \13258 , \13291 );
xnor \U$11563 ( \13293 , \13289 , \13292 );
and \U$11564 ( \13294 , \13234 , \13293 );
and \U$11565 ( \13295 , RI2b5e785c0a00_257, \12863 );
and \U$11566 ( \13296 , RI2b5e785be390_277, \12865 );
and \U$11567 ( \13297 , RI2b5e785bc0e0_297, \12868 );
and \U$11568 ( \13298 , RI2b5e785ba1f0_317, \12871 );
and \U$11569 ( \13299 , RI2b5e785b9890_337, \12873 );
and \U$11570 ( \13300 , RI2b5e785b7d60_357, \12876 );
and \U$11571 ( \13301 , RI2b5e785b7400_377, \12878 );
and \U$11572 ( \13302 , RI2b5e785b5c90_397, \12880 );
and \U$11573 ( \13303 , RI2b5e785b5330_417, \12882 );
and \U$11574 ( \13304 , RI2b5e785b49d0_437, \12884 );
and \U$11575 ( \13305 , RI2b5e785b3620_457, \12886 );
and \U$11576 ( \13306 , RI2b5e785b2cc0_477, \12888 );
and \U$11577 ( \13307 , RI2b5e785b2360_497, \12890 );
and \U$11578 ( \13308 , RI2b5e785b1370_517, \12892 );
and \U$11579 ( \13309 , RI2b5e785b0a10_537, \12894 );
and \U$11580 ( \13310 , RI2b5e785b00b0_557, \12896 );
and \U$11581 ( \13311 , RI2b5e785af480_577, \12898 );
or \U$11582 ( \13312 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 );
_DC r39e2 ( \13313_nR39e2 , \13312 , \12908 );
buf \U$11583 ( \13314 , \13313_nR39e2 );
xor \U$11584 ( \13315 , \12607 , \12628 );
xor \U$11585 ( \13316 , \13315 , \12765 );
buf \U$11586 ( \13317 , \13316 );
buf \U$11587 ( \13318 , \13317 );
xor \U$11588 ( \13319 , \12632 , \12653 );
xor \U$11589 ( \13320 , \13319 , \12762 );
buf \U$11590 ( \13321 , \13320 );
buf \U$11591 ( \13322 , \13321 );
xor \U$11592 ( \13323 , \13318 , \13322 );
xor \U$11593 ( \13324 , \13322 , \13258 );
not \U$11594 ( \13325 , \13324 );
and \U$11595 ( \13326 , \13323 , \13325 );
and \U$11596 ( \13327 , \13314 , \13326 );
and \U$11597 ( \13328 , RI2b5e785c2b48_256, \12863 );
and \U$11598 ( \13329 , RI2b5e785be408_276, \12865 );
and \U$11599 ( \13330 , RI2b5e785bc158_296, \12868 );
and \U$11600 ( \13331 , RI2b5e785ba268_316, \12871 );
and \U$11601 ( \13332 , RI2b5e785b9908_336, \12873 );
and \U$11602 ( \13333 , RI2b5e785b7dd8_356, \12876 );
and \U$11603 ( \13334 , RI2b5e785b7478_376, \12878 );
and \U$11604 ( \13335 , RI2b5e785b5d08_396, \12880 );
and \U$11605 ( \13336 , RI2b5e785b53a8_416, \12882 );
and \U$11606 ( \13337 , RI2b5e785b4a48_436, \12884 );
and \U$11607 ( \13338 , RI2b5e785b3698_456, \12886 );
and \U$11608 ( \13339 , RI2b5e785b2d38_476, \12888 );
and \U$11609 ( \13340 , RI2b5e785b23d8_496, \12890 );
and \U$11610 ( \13341 , RI2b5e785b13e8_516, \12892 );
and \U$11611 ( \13342 , RI2b5e785b0a88_536, \12894 );
and \U$11612 ( \13343 , RI2b5e785b0128_556, \12896 );
and \U$11613 ( \13344 , RI2b5e785af4f8_576, \12898 );
or \U$11614 ( \13345 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 );
_DC r3a7a ( \13346_nR3a7a , \13345 , \12908 );
buf \U$11615 ( \13347 , \13346_nR3a7a );
and \U$11616 ( \13348 , \13347 , \13324 );
nor \U$11617 ( \13349 , \13327 , \13348 );
and \U$11618 ( \13350 , \13322 , \13258 );
not \U$11619 ( \13351 , \13350 );
and \U$11620 ( \13352 , \13318 , \13351 );
xnor \U$11621 ( \13353 , \13349 , \13352 );
and \U$11622 ( \13354 , \13293 , \13353 );
and \U$11623 ( \13355 , \13234 , \13353 );
or \U$11624 ( \13356 , \13294 , \13354 , \13355 );
and \U$11625 ( \13357 , RI2b5e785c0910_259, \12863 );
and \U$11626 ( \13358 , RI2b5e785be2a0_279, \12865 );
and \U$11627 ( \13359 , RI2b5e785bbff0_299, \12868 );
and \U$11628 ( \13360 , RI2b5e785ba100_319, \12871 );
and \U$11629 ( \13361 , RI2b5e785b97a0_339, \12873 );
and \U$11630 ( \13362 , RI2b5e785b7c70_359, \12876 );
and \U$11631 ( \13363 , RI2b5e785b7310_379, \12878 );
and \U$11632 ( \13364 , RI2b5e785b5ba0_399, \12880 );
and \U$11633 ( \13365 , RI2b5e785b5240_419, \12882 );
and \U$11634 ( \13366 , RI2b5e785b48e0_439, \12884 );
and \U$11635 ( \13367 , RI2b5e785b3530_459, \12886 );
and \U$11636 ( \13368 , RI2b5e785b2bd0_479, \12888 );
and \U$11637 ( \13369 , RI2b5e785b2270_499, \12890 );
and \U$11638 ( \13370 , RI2b5e785b1280_519, \12892 );
and \U$11639 ( \13371 , RI2b5e785b0920_539, \12894 );
and \U$11640 ( \13372 , RI2b5e785affc0_559, \12896 );
and \U$11641 ( \13373 , RI2b5e785af390_579, \12898 );
or \U$11642 ( \13374 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 );
_DC r3817 ( \13375_nR3817 , \13374 , \12908 );
buf \U$11643 ( \13376 , \13375_nR3817 );
xor \U$11644 ( \13377 , \12582 , \12603 );
xor \U$11645 ( \13378 , \13377 , \12768 );
buf \U$11646 ( \13379 , \13378 );
buf \U$11647 ( \13380 , \13379 );
xor \U$11648 ( \13381 , \13082 , \13380 );
xor \U$11649 ( \13382 , \13380 , \13318 );
not \U$11650 ( \13383 , \13382 );
and \U$11651 ( \13384 , \13381 , \13383 );
and \U$11652 ( \13385 , \13376 , \13384 );
and \U$11653 ( \13386 , RI2b5e785c0988_258, \12863 );
and \U$11654 ( \13387 , RI2b5e785be318_278, \12865 );
and \U$11655 ( \13388 , RI2b5e785bc068_298, \12868 );
and \U$11656 ( \13389 , RI2b5e785ba178_318, \12871 );
and \U$11657 ( \13390 , RI2b5e785b9818_338, \12873 );
and \U$11658 ( \13391 , RI2b5e785b7ce8_358, \12876 );
and \U$11659 ( \13392 , RI2b5e785b7388_378, \12878 );
and \U$11660 ( \13393 , RI2b5e785b5c18_398, \12880 );
and \U$11661 ( \13394 , RI2b5e785b52b8_418, \12882 );
and \U$11662 ( \13395 , RI2b5e785b4958_438, \12884 );
and \U$11663 ( \13396 , RI2b5e785b35a8_458, \12886 );
and \U$11664 ( \13397 , RI2b5e785b2c48_478, \12888 );
and \U$11665 ( \13398 , RI2b5e785b22e8_498, \12890 );
and \U$11666 ( \13399 , RI2b5e785b12f8_518, \12892 );
and \U$11667 ( \13400 , RI2b5e785b0998_538, \12894 );
and \U$11668 ( \13401 , RI2b5e785b0038_558, \12896 );
and \U$11669 ( \13402 , RI2b5e785af408_578, \12898 );
or \U$11670 ( \13403 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 );
_DC r38a1 ( \13404_nR38a1 , \13403 , \12908 );
buf \U$11671 ( \13405 , \13404_nR38a1 );
and \U$11672 ( \13406 , \13405 , \13382 );
nor \U$11673 ( \13407 , \13385 , \13406 );
and \U$11674 ( \13408 , \13380 , \13318 );
not \U$11675 ( \13409 , \13408 );
and \U$11676 ( \13410 , \13082 , \13409 );
xnor \U$11677 ( \13411 , \13407 , \13410 );
and \U$11678 ( \13412 , RI2b5e785c0820_261, \12863 );
and \U$11679 ( \13413 , RI2b5e785be1b0_281, \12865 );
and \U$11680 ( \13414 , RI2b5e785bbf00_301, \12868 );
and \U$11681 ( \13415 , RI2b5e785ba010_321, \12871 );
and \U$11682 ( \13416 , RI2b5e785b96b0_341, \12873 );
and \U$11683 ( \13417 , RI2b5e785b7b80_361, \12876 );
and \U$11684 ( \13418 , RI2b5e785b7220_381, \12878 );
and \U$11685 ( \13419 , RI2b5e785b5ab0_401, \12880 );
and \U$11686 ( \13420 , RI2b5e785b5150_421, \12882 );
and \U$11687 ( \13421 , RI2b5e785b47f0_441, \12884 );
and \U$11688 ( \13422 , RI2b5e785b3440_461, \12886 );
and \U$11689 ( \13423 , RI2b5e785b2ae0_481, \12888 );
and \U$11690 ( \13424 , RI2b5e785b2180_501, \12890 );
and \U$11691 ( \13425 , RI2b5e785b1190_521, \12892 );
and \U$11692 ( \13426 , RI2b5e785b0830_541, \12894 );
and \U$11693 ( \13427 , RI2b5e785afed0_561, \12896 );
and \U$11694 ( \13428 , RI2b5e785af2a0_581, \12898 );
or \U$11695 ( \13429 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 );
_DC r3674 ( \13430_nR3674 , \13429 , \12908 );
buf \U$11696 ( \13431 , \13430_nR3674 );
and \U$11697 ( \13432 , \13431 , \13085 );
and \U$11698 ( \13433 , RI2b5e785c0898_260, \12863 );
and \U$11699 ( \13434 , RI2b5e785be228_280, \12865 );
and \U$11700 ( \13435 , RI2b5e785bbf78_300, \12868 );
and \U$11701 ( \13436 , RI2b5e785ba088_320, \12871 );
and \U$11702 ( \13437 , RI2b5e785b9728_340, \12873 );
and \U$11703 ( \13438 , RI2b5e785b7bf8_360, \12876 );
and \U$11704 ( \13439 , RI2b5e785b7298_380, \12878 );
and \U$11705 ( \13440 , RI2b5e785b5b28_400, \12880 );
and \U$11706 ( \13441 , RI2b5e785b51c8_420, \12882 );
and \U$11707 ( \13442 , RI2b5e785b4868_440, \12884 );
and \U$11708 ( \13443 , RI2b5e785b34b8_460, \12886 );
and \U$11709 ( \13444 , RI2b5e785b2b58_480, \12888 );
and \U$11710 ( \13445 , RI2b5e785b21f8_500, \12890 );
and \U$11711 ( \13446 , RI2b5e785b1208_520, \12892 );
and \U$11712 ( \13447 , RI2b5e785b08a8_540, \12894 );
and \U$11713 ( \13448 , RI2b5e785aff48_560, \12896 );
and \U$11714 ( \13449 , RI2b5e785af318_580, \12898 );
or \U$11715 ( \13450 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 );
_DC r36e8 ( \13451_nR36e8 , \13450 , \12908 );
buf \U$11716 ( \13452 , \13451_nR36e8 );
and \U$11717 ( \13453 , \13452 , \13083 );
nor \U$11718 ( \13454 , \13432 , \13453 );
xnor \U$11719 ( \13455 , \13454 , \13090 );
and \U$11720 ( \13456 , \13411 , \13455 );
and \U$11721 ( \13457 , RI2b5e785c0730_263, \12863 );
and \U$11722 ( \13458 , RI2b5e785be0c0_283, \12865 );
and \U$11723 ( \13459 , RI2b5e785bbe10_303, \12868 );
and \U$11724 ( \13460 , RI2b5e785b9f20_323, \12871 );
and \U$11725 ( \13461 , RI2b5e785b95c0_343, \12873 );
and \U$11726 ( \13462 , RI2b5e785b7a90_363, \12876 );
and \U$11727 ( \13463 , RI2b5e785b7130_383, \12878 );
and \U$11728 ( \13464 , RI2b5e785b59c0_403, \12880 );
and \U$11729 ( \13465 , RI2b5e785b5060_423, \12882 );
and \U$11730 ( \13466 , RI2b5e785b3cb0_443, \12884 );
and \U$11731 ( \13467 , RI2b5e785b3350_463, \12886 );
and \U$11732 ( \13468 , RI2b5e785b29f0_483, \12888 );
and \U$11733 ( \13469 , RI2b5e785b1a00_503, \12890 );
and \U$11734 ( \13470 , RI2b5e785b10a0_523, \12892 );
and \U$11735 ( \13471 , RI2b5e785b0740_543, \12894 );
and \U$11736 ( \13472 , RI2b5e785afde0_563, \12896 );
and \U$11737 ( \13473 , RI2b5e785af1b0_583, \12898 );
or \U$11738 ( \13474 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 );
_DC r3503 ( \13475_nR3503 , \13474 , \12908 );
buf \U$11739 ( \13476 , \13475_nR3503 );
and \U$11740 ( \13477 , \13476 , \13020 );
and \U$11741 ( \13478 , RI2b5e785c07a8_262, \12863 );
and \U$11742 ( \13479 , RI2b5e785be138_282, \12865 );
and \U$11743 ( \13480 , RI2b5e785bbe88_302, \12868 );
and \U$11744 ( \13481 , RI2b5e785b9f98_322, \12871 );
and \U$11745 ( \13482 , RI2b5e785b9638_342, \12873 );
and \U$11746 ( \13483 , RI2b5e785b7b08_362, \12876 );
and \U$11747 ( \13484 , RI2b5e785b71a8_382, \12878 );
and \U$11748 ( \13485 , RI2b5e785b5a38_402, \12880 );
and \U$11749 ( \13486 , RI2b5e785b50d8_422, \12882 );
and \U$11750 ( \13487 , RI2b5e785b4778_442, \12884 );
and \U$11751 ( \13488 , RI2b5e785b33c8_462, \12886 );
and \U$11752 ( \13489 , RI2b5e785b2a68_482, \12888 );
and \U$11753 ( \13490 , RI2b5e785b1a78_502, \12890 );
and \U$11754 ( \13491 , RI2b5e785b1118_522, \12892 );
and \U$11755 ( \13492 , RI2b5e785b07b8_542, \12894 );
and \U$11756 ( \13493 , RI2b5e785afe58_562, \12896 );
and \U$11757 ( \13494 , RI2b5e785af228_582, \12898 );
or \U$11758 ( \13495 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 );
_DC r356a ( \13496_nR356a , \13495 , \12908 );
buf \U$11759 ( \13497 , \13496_nR356a );
and \U$11760 ( \13498 , \13497 , \13018 );
nor \U$11761 ( \13499 , \13477 , \13498 );
xnor \U$11762 ( \13500 , \13499 , \12797 );
and \U$11763 ( \13501 , \13455 , \13500 );
and \U$11764 ( \13502 , \13411 , \13500 );
or \U$11765 ( \13503 , \13456 , \13501 , \13502 );
and \U$11766 ( \13504 , \13356 , \13503 );
and \U$11767 ( \13505 , RI2b5e785c0640_265, \12863 );
and \U$11768 ( \13506 , RI2b5e785bdfd0_285, \12865 );
and \U$11769 ( \13507 , RI2b5e785bbd20_305, \12868 );
and \U$11770 ( \13508 , RI2b5e785b9e30_325, \12871 );
and \U$11771 ( \13509 , RI2b5e785b94d0_345, \12873 );
and \U$11772 ( \13510 , RI2b5e785b79a0_365, \12876 );
and \U$11773 ( \13511 , RI2b5e785b7040_385, \12878 );
and \U$11774 ( \13512 , RI2b5e785b58d0_405, \12880 );
and \U$11775 ( \13513 , RI2b5e785b4f70_425, \12882 );
and \U$11776 ( \13514 , RI2b5e785b3bc0_445, \12884 );
and \U$11777 ( \13515 , RI2b5e785b3260_465, \12886 );
and \U$11778 ( \13516 , RI2b5e785b2900_485, \12888 );
and \U$11779 ( \13517 , RI2b5e785b1910_505, \12890 );
and \U$11780 ( \13518 , RI2b5e785b0fb0_525, \12892 );
and \U$11781 ( \13519 , RI2b5e785b0650_545, \12894 );
and \U$11782 ( \13520 , RI2b5e785afcf0_565, \12896 );
and \U$11783 ( \13521 , RI2b5e785af0c0_585, \12898 );
or \U$11784 ( \13522 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 );
_DC r3385 ( \13523_nR3385 , \13522 , \12908 );
buf \U$11785 ( \13524 , \13523_nR3385 );
and \U$11786 ( \13525 , \13524 , \12958 );
and \U$11787 ( \13526 , RI2b5e785c06b8_264, \12863 );
and \U$11788 ( \13527 , RI2b5e785be048_284, \12865 );
and \U$11789 ( \13528 , RI2b5e785bbd98_304, \12868 );
and \U$11790 ( \13529 , RI2b5e785b9ea8_324, \12871 );
and \U$11791 ( \13530 , RI2b5e785b9548_344, \12873 );
and \U$11792 ( \13531 , RI2b5e785b7a18_364, \12876 );
and \U$11793 ( \13532 , RI2b5e785b70b8_384, \12878 );
and \U$11794 ( \13533 , RI2b5e785b5948_404, \12880 );
and \U$11795 ( \13534 , RI2b5e785b4fe8_424, \12882 );
and \U$11796 ( \13535 , RI2b5e785b3c38_444, \12884 );
and \U$11797 ( \13536 , RI2b5e785b32d8_464, \12886 );
and \U$11798 ( \13537 , RI2b5e785b2978_484, \12888 );
and \U$11799 ( \13538 , RI2b5e785b1988_504, \12890 );
and \U$11800 ( \13539 , RI2b5e785b1028_524, \12892 );
and \U$11801 ( \13540 , RI2b5e785b06c8_544, \12894 );
and \U$11802 ( \13541 , RI2b5e785afd68_564, \12896 );
and \U$11803 ( \13542 , RI2b5e785af138_584, \12898 );
or \U$11804 ( \13543 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 );
_DC r3418 ( \13544_nR3418 , \13543 , \12908 );
buf \U$11805 ( \13545 , \13544_nR3418 );
and \U$11806 ( \13546 , \13545 , \12956 );
nor \U$11807 ( \13547 , \13525 , \13546 );
xnor \U$11808 ( \13548 , \13547 , \12984 );
and \U$11810 ( \13549 , RI2b5e785c05c8_266, \12863 );
and \U$11811 ( \13550 , RI2b5e785bdf58_286, \12865 );
and \U$11812 ( \13551 , RI2b5e785bbca8_306, \12868 );
and \U$11813 ( \13552 , RI2b5e785b9db8_326, \12871 );
and \U$11814 ( \13553 , RI2b5e785b9458_346, \12873 );
and \U$11815 ( \13554 , RI2b5e785b7928_366, \12876 );
and \U$11816 ( \13555 , RI2b5e785b6fc8_386, \12878 );
and \U$11817 ( \13556 , RI2b5e785b5858_406, \12880 );
and \U$11818 ( \13557 , RI2b5e785b4ef8_426, \12882 );
and \U$11819 ( \13558 , RI2b5e785b3b48_446, \12884 );
and \U$11820 ( \13559 , RI2b5e785b31e8_466, \12886 );
and \U$11821 ( \13560 , RI2b5e785b2888_486, \12888 );
and \U$11822 ( \13561 , RI2b5e785b1898_506, \12890 );
and \U$11823 ( \13562 , RI2b5e785b0f38_526, \12892 );
and \U$11824 ( \13563 , RI2b5e785b05d8_546, \12894 );
and \U$11825 ( \13564 , RI2b5e785afc78_566, \12896 );
and \U$11826 ( \13565 , RI2b5e785af048_586, \12898 );
or \U$11827 ( \13566 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 );
_DC r32fd ( \13567_nR32fd , \13566 , \12908 );
buf \U$11828 ( \13568 , \13567_nR32fd );
and \U$11829 ( \13569 , \13568 , \13011 );
nor \U$11830 ( \13570 , 1'b0 , \13569 );
xnor \U$11831 ( \13571 , \13570 , 1'b0 );
and \U$11832 ( \13572 , \13548 , \13571 );
and \U$11833 ( \13573 , \13503 , \13572 );
and \U$11834 ( \13574 , \13356 , \13572 );
or \U$11835 ( \13575 , \13504 , \13573 , \13574 );
and \U$11837 ( \13576 , \13497 , \13020 );
and \U$11838 ( \13577 , \13431 , \13018 );
nor \U$11839 ( \13578 , \13576 , \13577 );
xnor \U$11840 ( \13579 , \13578 , \12797 );
and \U$11841 ( \13580 , \13545 , \12958 );
and \U$11842 ( \13581 , \13476 , \12956 );
nor \U$11843 ( \13582 , \13580 , \13581 );
xnor \U$11844 ( \13583 , \13582 , \12984 );
xor \U$11845 ( \13584 , \13579 , \13583 );
and \U$11847 ( \13585 , \13524 , \13011 );
nor \U$11848 ( \13586 , 1'b0 , \13585 );
xnor \U$11849 ( \13587 , \13586 , 1'b0 );
xor \U$11850 ( \13588 , \13584 , \13587 );
and \U$11851 ( \13589 , \13347 , \13326 );
and \U$11852 ( \13590 , \13254 , \13324 );
nor \U$11853 ( \13591 , \13589 , \13590 );
xnor \U$11854 ( \13592 , \13591 , \13352 );
and \U$11855 ( \13593 , \13405 , \13384 );
and \U$11856 ( \13594 , \13314 , \13382 );
nor \U$11857 ( \13595 , \13593 , \13594 );
xnor \U$11858 ( \13596 , \13595 , \13410 );
xor \U$11859 ( \13597 , \13592 , \13596 );
and \U$11860 ( \13598 , \13452 , \13085 );
and \U$11861 ( \13599 , \13376 , \13083 );
nor \U$11862 ( \13600 , \13598 , \13599 );
xnor \U$11863 ( \13601 , \13600 , \13090 );
xor \U$11864 ( \13602 , \13597 , \13601 );
and \U$11865 ( \13603 , \13588 , \13602 );
or \U$11867 ( \13604 , 1'b0 , \13603 , 1'b0 );
xor \U$11868 ( \13605 , \13575 , \13604 );
and \U$11869 ( \13606 , \13476 , \12958 );
and \U$11870 ( \13607 , \13497 , \12956 );
nor \U$11871 ( \13608 , \13606 , \13607 );
xnor \U$11872 ( \13609 , \13608 , \12984 );
and \U$11874 ( \13610 , \13545 , \13011 );
nor \U$11875 ( \13611 , 1'b0 , \13610 );
xnor \U$11876 ( \13612 , \13611 , 1'b0 );
xor \U$11877 ( \13613 , \13609 , \13612 );
xor \U$11879 ( \13614 , \13613 , 1'b0 );
and \U$11880 ( \13615 , \13314 , \13384 );
and \U$11881 ( \13616 , \13347 , \13382 );
nor \U$11882 ( \13617 , \13615 , \13616 );
xnor \U$11883 ( \13618 , \13617 , \13410 );
and \U$11884 ( \13619 , \13376 , \13085 );
and \U$11885 ( \13620 , \13405 , \13083 );
nor \U$11886 ( \13621 , \13619 , \13620 );
xnor \U$11887 ( \13622 , \13621 , \13090 );
xor \U$11888 ( \13623 , \13618 , \13622 );
and \U$11889 ( \13624 , \13431 , \13020 );
and \U$11890 ( \13625 , \13452 , \13018 );
nor \U$11891 ( \13626 , \13624 , \13625 );
xnor \U$11892 ( \13627 , \13626 , \12797 );
xor \U$11893 ( \13628 , \13623 , \13627 );
xor \U$11894 ( \13629 , \13614 , \13628 );
and \U$11895 ( \13630 , \13138 , \13230 );
and \U$11896 ( \13631 , \13006 , \13227 );
nor \U$11897 ( \13632 , \13630 , \13631 );
xnor \U$11898 ( \13633 , \13632 , \13224 );
and \U$11899 ( \13634 , \13161 , \13266 );
and \U$11900 ( \13635 , \13117 , \13264 );
nor \U$11901 ( \13636 , \13634 , \13635 );
xnor \U$11902 ( \13637 , \13636 , \13292 );
xor \U$11903 ( \13638 , \13633 , \13637 );
and \U$11904 ( \13639 , \13254 , \13326 );
and \U$11905 ( \13640 , \13287 , \13324 );
nor \U$11906 ( \13641 , \13639 , \13640 );
xnor \U$11907 ( \13642 , \13641 , \13352 );
xor \U$11908 ( \13643 , \13638 , \13642 );
xor \U$11909 ( \13644 , \13629 , \13643 );
xor \U$11910 ( \13645 , \13605 , \13644 );
and \U$11912 ( \13646 , \13287 , \13230 );
and \U$11913 ( \13647 , \13161 , \13227 );
nor \U$11914 ( \13648 , \13646 , \13647 );
xnor \U$11915 ( \13649 , \13648 , \13224 );
and \U$11916 ( \13650 , \13347 , \13266 );
and \U$11917 ( \13651 , \13254 , \13264 );
nor \U$11918 ( \13652 , \13650 , \13651 );
xnor \U$11919 ( \13653 , \13652 , \13292 );
and \U$11920 ( \13654 , \13649 , \13653 );
or \U$11922 ( \13655 , 1'b0 , \13654 , 1'b0 );
and \U$11923 ( \13656 , \13405 , \13326 );
and \U$11924 ( \13657 , \13314 , \13324 );
nor \U$11925 ( \13658 , \13656 , \13657 );
xnor \U$11926 ( \13659 , \13658 , \13352 );
and \U$11927 ( \13660 , \13452 , \13384 );
and \U$11928 ( \13661 , \13376 , \13382 );
nor \U$11929 ( \13662 , \13660 , \13661 );
xnor \U$11930 ( \13663 , \13662 , \13410 );
and \U$11931 ( \13664 , \13659 , \13663 );
and \U$11932 ( \13665 , \13497 , \13085 );
and \U$11933 ( \13666 , \13431 , \13083 );
nor \U$11934 ( \13667 , \13665 , \13666 );
xnor \U$11935 ( \13668 , \13667 , \13090 );
and \U$11936 ( \13669 , \13663 , \13668 );
and \U$11937 ( \13670 , \13659 , \13668 );
or \U$11938 ( \13671 , \13664 , \13669 , \13670 );
and \U$11939 ( \13672 , \13655 , \13671 );
and \U$11940 ( \13673 , \13545 , \13020 );
and \U$11941 ( \13674 , \13476 , \13018 );
nor \U$11942 ( \13675 , \13673 , \13674 );
xnor \U$11943 ( \13676 , \13675 , \12797 );
and \U$11944 ( \13677 , \13568 , \12958 );
and \U$11945 ( \13678 , \13524 , \12956 );
nor \U$11946 ( \13679 , \13677 , \13678 );
xnor \U$11947 ( \13680 , \13679 , \12984 );
and \U$11948 ( \13681 , \13676 , \13680 );
and \U$11949 ( \13682 , RI2b5e785c0550_267, \12863 );
and \U$11950 ( \13683 , RI2b5e785bc590_287, \12865 );
and \U$11951 ( \13684 , RI2b5e785bbc30_307, \12868 );
and \U$11952 ( \13685 , RI2b5e785b9d40_327, \12871 );
and \U$11953 ( \13686 , RI2b5e785b93e0_347, \12873 );
and \U$11954 ( \13687 , RI2b5e785b78b0_367, \12876 );
and \U$11955 ( \13688 , RI2b5e785b6f50_387, \12878 );
and \U$11956 ( \13689 , RI2b5e785b57e0_407, \12880 );
and \U$11957 ( \13690 , RI2b5e785b4e80_427, \12882 );
and \U$11958 ( \13691 , RI2b5e785b3ad0_447, \12884 );
and \U$11959 ( \13692 , RI2b5e785b3170_467, \12886 );
and \U$11960 ( \13693 , RI2b5e785b2810_487, \12888 );
and \U$11961 ( \13694 , RI2b5e785b1820_507, \12890 );
and \U$11962 ( \13695 , RI2b5e785b0ec0_527, \12892 );
and \U$11963 ( \13696 , RI2b5e785b0560_547, \12894 );
and \U$11964 ( \13697 , RI2b5e785afc00_567, \12896 );
and \U$11965 ( \13698 , RI2b5e785aefd0_587, \12898 );
or \U$11966 ( \13699 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 );
_DC r326b ( \13700_nR326b , \13699 , \12908 );
buf \U$11967 ( \13701 , \13700_nR326b );
nand \U$11968 ( \13702 , \13701 , \13011 );
xnor \U$11969 ( \13703 , \13702 , 1'b0 );
and \U$11970 ( \13704 , \13680 , \13703 );
and \U$11971 ( \13705 , \13676 , \13703 );
or \U$11972 ( \13706 , \13681 , \13704 , \13705 );
and \U$11973 ( \13707 , \13671 , \13706 );
and \U$11974 ( \13708 , \13655 , \13706 );
or \U$11975 ( \13709 , \13672 , \13707 , \13708 );
xor \U$11976 ( \13710 , \13548 , \13571 );
xor \U$11977 ( \13711 , \13411 , \13455 );
xor \U$11978 ( \13712 , \13711 , \13500 );
and \U$11979 ( \13713 , \13710 , \13712 );
xor \U$11980 ( \13714 , \13234 , \13293 );
xor \U$11981 ( \13715 , \13714 , \13353 );
and \U$11982 ( \13716 , \13712 , \13715 );
and \U$11983 ( \13717 , \13710 , \13715 );
or \U$11984 ( \13718 , \13713 , \13716 , \13717 );
and \U$11985 ( \13719 , \13709 , \13718 );
and \U$11987 ( \13720 , \13117 , \13230 );
and \U$11988 ( \13721 , \13138 , \13227 );
nor \U$11989 ( \13722 , \13720 , \13721 );
xnor \U$11990 ( \13723 , \13722 , \13224 );
xor \U$11991 ( \13724 , 1'b0 , \13723 );
and \U$11992 ( \13725 , \13287 , \13266 );
and \U$11993 ( \13726 , \13161 , \13264 );
nor \U$11994 ( \13727 , \13725 , \13726 );
xnor \U$11995 ( \13728 , \13727 , \13292 );
xor \U$11996 ( \13729 , \13724 , \13728 );
and \U$11997 ( \13730 , \13718 , \13729 );
and \U$11998 ( \13731 , \13709 , \13729 );
or \U$11999 ( \13732 , \13719 , \13730 , \13731 );
xor \U$12001 ( \13733 , 1'b0 , \13588 );
xor \U$12002 ( \13734 , \13733 , \13602 );
xor \U$12003 ( \13735 , \13356 , \13503 );
xor \U$12004 ( \13736 , \13735 , \13572 );
and \U$12005 ( \13737 , \13734 , \13736 );
xor \U$12006 ( \13738 , \13732 , \13737 );
and \U$12008 ( \13739 , \13723 , \13728 );
or \U$12010 ( \13740 , 1'b0 , \13739 , 1'b0 );
and \U$12011 ( \13741 , \13592 , \13596 );
and \U$12012 ( \13742 , \13596 , \13601 );
and \U$12013 ( \13743 , \13592 , \13601 );
or \U$12014 ( \13744 , \13741 , \13742 , \13743 );
xor \U$12015 ( \13745 , \13740 , \13744 );
and \U$12016 ( \13746 , \13579 , \13583 );
and \U$12017 ( \13747 , \13583 , \13587 );
and \U$12018 ( \13748 , \13579 , \13587 );
or \U$12019 ( \13749 , \13746 , \13747 , \13748 );
xor \U$12020 ( \13750 , \13745 , \13749 );
xor \U$12021 ( \13751 , \13738 , \13750 );
xor \U$12022 ( \13752 , \13645 , \13751 );
and \U$12023 ( \13753 , \13254 , \13230 );
and \U$12024 ( \13754 , \13287 , \13227 );
nor \U$12025 ( \13755 , \13753 , \13754 );
xnor \U$12026 ( \13756 , \13755 , \13224 );
and \U$12027 ( \13757 , \13314 , \13266 );
and \U$12028 ( \13758 , \13347 , \13264 );
nor \U$12029 ( \13759 , \13757 , \13758 );
xnor \U$12030 ( \13760 , \13759 , \13292 );
and \U$12031 ( \13761 , \13756 , \13760 );
and \U$12032 ( \13762 , \13376 , \13326 );
and \U$12033 ( \13763 , \13405 , \13324 );
nor \U$12034 ( \13764 , \13762 , \13763 );
xnor \U$12035 ( \13765 , \13764 , \13352 );
and \U$12036 ( \13766 , \13760 , \13765 );
and \U$12037 ( \13767 , \13756 , \13765 );
or \U$12038 ( \13768 , \13761 , \13766 , \13767 );
and \U$12039 ( \13769 , \13431 , \13384 );
and \U$12040 ( \13770 , \13452 , \13382 );
nor \U$12041 ( \13771 , \13769 , \13770 );
xnor \U$12042 ( \13772 , \13771 , \13410 );
and \U$12043 ( \13773 , \13476 , \13085 );
and \U$12044 ( \13774 , \13497 , \13083 );
nor \U$12045 ( \13775 , \13773 , \13774 );
xnor \U$12046 ( \13776 , \13775 , \13090 );
and \U$12047 ( \13777 , \13772 , \13776 );
and \U$12048 ( \13778 , \13524 , \13020 );
and \U$12049 ( \13779 , \13545 , \13018 );
nor \U$12050 ( \13780 , \13778 , \13779 );
xnor \U$12051 ( \13781 , \13780 , \12797 );
and \U$12052 ( \13782 , \13776 , \13781 );
and \U$12053 ( \13783 , \13772 , \13781 );
or \U$12054 ( \13784 , \13777 , \13782 , \13783 );
and \U$12055 ( \13785 , \13768 , \13784 );
xor \U$12056 ( \13786 , \13676 , \13680 );
xor \U$12057 ( \13787 , \13786 , \13703 );
and \U$12058 ( \13788 , \13784 , \13787 );
and \U$12059 ( \13789 , \13768 , \13787 );
or \U$12060 ( \13790 , \13785 , \13788 , \13789 );
xor \U$12061 ( \13791 , \13659 , \13663 );
xor \U$12062 ( \13792 , \13791 , \13668 );
xor \U$12063 ( \13793 , 1'b0 , \13649 );
xor \U$12064 ( \13794 , \13793 , \13653 );
and \U$12065 ( \13795 , \13792 , \13794 );
and \U$12066 ( \13796 , \13790 , \13795 );
xor \U$12067 ( \13797 , \13710 , \13712 );
xor \U$12068 ( \13798 , \13797 , \13715 );
and \U$12069 ( \13799 , \13795 , \13798 );
and \U$12070 ( \13800 , \13790 , \13798 );
or \U$12071 ( \13801 , \13796 , \13799 , \13800 );
xor \U$12072 ( \13802 , \13734 , \13736 );
and \U$12073 ( \13803 , \13801 , \13802 );
xor \U$12074 ( \13804 , \13709 , \13718 );
xor \U$12075 ( \13805 , \13804 , \13729 );
and \U$12076 ( \13806 , \13802 , \13805 );
and \U$12077 ( \13807 , \13801 , \13805 );
or \U$12078 ( \13808 , \13803 , \13806 , \13807 );
nor \U$12079 ( \13809 , \13752 , \13808 );
and \U$12080 ( \13810 , \13732 , \13737 );
and \U$12081 ( \13811 , \13737 , \13750 );
and \U$12082 ( \13812 , \13732 , \13750 );
or \U$12083 ( \13813 , \13810 , \13811 , \13812 );
and \U$12084 ( \13814 , \13575 , \13604 );
and \U$12085 ( \13815 , \13604 , \13644 );
and \U$12086 ( \13816 , \13575 , \13644 );
or \U$12087 ( \13817 , \13814 , \13815 , \13816 );
and \U$12089 ( \13818 , \13006 , \13230 );
and \U$12090 ( \13819 , \12910 , \13227 );
nor \U$12091 ( \13820 , \13818 , \13819 );
xnor \U$12092 ( \13821 , \13820 , \13224 );
xor \U$12093 ( \13822 , 1'b0 , \13821 );
and \U$12094 ( \13823 , \13117 , \13266 );
and \U$12095 ( \13824 , \13138 , \13264 );
nor \U$12096 ( \13825 , \13823 , \13824 );
xnor \U$12097 ( \13826 , \13825 , \13292 );
xor \U$12098 ( \13827 , \13822 , \13826 );
and \U$12100 ( \13828 , \13452 , \13020 );
and \U$12101 ( \13829 , \13376 , \13018 );
nor \U$12102 ( \13830 , \13828 , \13829 );
xnor \U$12103 ( \13831 , \13830 , \12797 );
and \U$12104 ( \13832 , \13497 , \12958 );
and \U$12105 ( \13833 , \13431 , \12956 );
nor \U$12106 ( \13834 , \13832 , \13833 );
xnor \U$12107 ( \13835 , \13834 , \12984 );
xor \U$12108 ( \13836 , \13831 , \13835 );
and \U$12110 ( \13837 , \13476 , \13011 );
nor \U$12111 ( \13838 , 1'b0 , \13837 );
xnor \U$12112 ( \13839 , \13838 , 1'b0 );
xor \U$12113 ( \13840 , \13836 , \13839 );
xor \U$12114 ( \13841 , 1'b0 , \13840 );
xor \U$12115 ( \13842 , \13827 , \13841 );
and \U$12116 ( \13843 , \13633 , \13637 );
and \U$12117 ( \13844 , \13637 , \13642 );
and \U$12118 ( \13845 , \13633 , \13642 );
or \U$12119 ( \13846 , \13843 , \13844 , \13845 );
and \U$12120 ( \13847 , \13618 , \13622 );
and \U$12121 ( \13848 , \13622 , \13627 );
and \U$12122 ( \13849 , \13618 , \13627 );
or \U$12123 ( \13850 , \13847 , \13848 , \13849 );
xor \U$12124 ( \13851 , \13846 , \13850 );
and \U$12125 ( \13852 , \13609 , \13612 );
or \U$12128 ( \13853 , \13852 , 1'b0 , 1'b0 );
xor \U$12129 ( \13854 , \13851 , \13853 );
xor \U$12130 ( \13855 , \13842 , \13854 );
xor \U$12131 ( \13856 , \13817 , \13855 );
and \U$12132 ( \13857 , \13740 , \13744 );
and \U$12133 ( \13858 , \13744 , \13749 );
and \U$12134 ( \13859 , \13740 , \13749 );
or \U$12135 ( \13860 , \13857 , \13858 , \13859 );
and \U$12136 ( \13861 , \13614 , \13628 );
and \U$12137 ( \13862 , \13628 , \13643 );
and \U$12138 ( \13863 , \13614 , \13643 );
or \U$12139 ( \13864 , \13861 , \13862 , \13863 );
xor \U$12140 ( \13865 , \13860 , \13864 );
and \U$12141 ( \13866 , \13287 , \13326 );
and \U$12142 ( \13867 , \13161 , \13324 );
nor \U$12143 ( \13868 , \13866 , \13867 );
xnor \U$12144 ( \13869 , \13868 , \13352 );
and \U$12145 ( \13870 , \13347 , \13384 );
and \U$12146 ( \13871 , \13254 , \13382 );
nor \U$12147 ( \13872 , \13870 , \13871 );
xnor \U$12148 ( \13873 , \13872 , \13410 );
xor \U$12149 ( \13874 , \13869 , \13873 );
and \U$12150 ( \13875 , \13405 , \13085 );
and \U$12151 ( \13876 , \13314 , \13083 );
nor \U$12152 ( \13877 , \13875 , \13876 );
xnor \U$12153 ( \13878 , \13877 , \13090 );
xor \U$12154 ( \13879 , \13874 , \13878 );
xor \U$12155 ( \13880 , \13865 , \13879 );
xor \U$12156 ( \13881 , \13856 , \13880 );
xor \U$12157 ( \13882 , \13813 , \13881 );
and \U$12158 ( \13883 , \13645 , \13751 );
nor \U$12159 ( \13884 , \13882 , \13883 );
nor \U$12160 ( \13885 , \13809 , \13884 );
and \U$12161 ( \13886 , \13817 , \13855 );
and \U$12162 ( \13887 , \13855 , \13880 );
and \U$12163 ( \13888 , \13817 , \13880 );
or \U$12164 ( \13889 , \13886 , \13887 , \13888 );
and \U$12166 ( \13890 , \13821 , \13826 );
or \U$12168 ( \13891 , 1'b0 , \13890 , 1'b0 );
and \U$12169 ( \13892 , \13869 , \13873 );
and \U$12170 ( \13893 , \13873 , \13878 );
and \U$12171 ( \13894 , \13869 , \13878 );
or \U$12172 ( \13895 , \13892 , \13893 , \13894 );
xor \U$12173 ( \13896 , \13891 , \13895 );
and \U$12174 ( \13897 , \13831 , \13835 );
and \U$12175 ( \13898 , \13835 , \13839 );
and \U$12176 ( \13899 , \13831 , \13839 );
or \U$12177 ( \13900 , \13897 , \13898 , \13899 );
xor \U$12178 ( \13901 , \13896 , \13900 );
and \U$12179 ( \13902 , \13846 , \13850 );
and \U$12180 ( \13903 , \13850 , \13853 );
and \U$12181 ( \13904 , \13846 , \13853 );
or \U$12182 ( \13905 , \13902 , \13903 , \13904 );
xor \U$12184 ( \13906 , \13905 , 1'b0 );
and \U$12185 ( \13907 , \12910 , \13230 );
and \U$12186 ( \13908 , \12979 , \13227 );
nor \U$12187 ( \13909 , \13907 , \13908 );
xnor \U$12188 ( \13910 , \13909 , \13224 );
and \U$12189 ( \13911 , \13138 , \13266 );
and \U$12190 ( \13912 , \13006 , \13264 );
nor \U$12191 ( \13913 , \13911 , \13912 );
xnor \U$12192 ( \13914 , \13913 , \13292 );
xor \U$12193 ( \13915 , \13910 , \13914 );
and \U$12194 ( \13916 , \13161 , \13326 );
and \U$12195 ( \13917 , \13117 , \13324 );
nor \U$12196 ( \13918 , \13916 , \13917 );
xnor \U$12197 ( \13919 , \13918 , \13352 );
xor \U$12198 ( \13920 , \13915 , \13919 );
xor \U$12199 ( \13921 , \13906 , \13920 );
xor \U$12200 ( \13922 , \13901 , \13921 );
xor \U$12201 ( \13923 , \13889 , \13922 );
and \U$12202 ( \13924 , \13860 , \13864 );
and \U$12203 ( \13925 , \13864 , \13879 );
and \U$12204 ( \13926 , \13860 , \13879 );
or \U$12205 ( \13927 , \13924 , \13925 , \13926 );
and \U$12206 ( \13928 , \13827 , \13841 );
and \U$12207 ( \13929 , \13841 , \13854 );
and \U$12208 ( \13930 , \13827 , \13854 );
or \U$12209 ( \13931 , \13928 , \13929 , \13930 );
xor \U$12210 ( \13932 , \13927 , \13931 );
and \U$12212 ( \13933 , \13431 , \12958 );
and \U$12213 ( \13934 , \13452 , \12956 );
nor \U$12214 ( \13935 , \13933 , \13934 );
xnor \U$12215 ( \13936 , \13935 , \12984 );
and \U$12217 ( \13937 , \13497 , \13011 );
nor \U$12218 ( \13938 , 1'b0 , \13937 );
xnor \U$12219 ( \13939 , \13938 , 1'b0 );
xor \U$12220 ( \13940 , \13936 , \13939 );
xor \U$12222 ( \13941 , \13940 , 1'b0 );
xor \U$12223 ( \13942 , 1'b0 , \13941 );
and \U$12224 ( \13943 , \13254 , \13384 );
and \U$12225 ( \13944 , \13287 , \13382 );
nor \U$12226 ( \13945 , \13943 , \13944 );
xnor \U$12227 ( \13946 , \13945 , \13410 );
and \U$12228 ( \13947 , \13314 , \13085 );
and \U$12229 ( \13948 , \13347 , \13083 );
nor \U$12230 ( \13949 , \13947 , \13948 );
xnor \U$12231 ( \13950 , \13949 , \13090 );
xor \U$12232 ( \13951 , \13946 , \13950 );
and \U$12233 ( \13952 , \13376 , \13020 );
and \U$12234 ( \13953 , \13405 , \13018 );
nor \U$12235 ( \13954 , \13952 , \13953 );
xnor \U$12236 ( \13955 , \13954 , \12797 );
xor \U$12237 ( \13956 , \13951 , \13955 );
xor \U$12238 ( \13957 , \13942 , \13956 );
xor \U$12239 ( \13958 , \13932 , \13957 );
xor \U$12240 ( \13959 , \13923 , \13958 );
and \U$12241 ( \13960 , \13813 , \13881 );
nor \U$12242 ( \13961 , \13959 , \13960 );
and \U$12243 ( \13962 , \13927 , \13931 );
and \U$12244 ( \13963 , \13931 , \13957 );
and \U$12245 ( \13964 , \13927 , \13957 );
or \U$12246 ( \13965 , \13962 , \13963 , \13964 );
and \U$12247 ( \13966 , \13901 , \13921 );
xor \U$12248 ( \13967 , \13965 , \13966 );
and \U$12251 ( \13968 , \13905 , \13920 );
or \U$12252 ( \13969 , 1'b0 , 1'b0 , \13968 );
and \U$12254 ( \13970 , \13405 , \13020 );
and \U$12255 ( \13971 , \13314 , \13018 );
nor \U$12256 ( \13972 , \13970 , \13971 );
xnor \U$12257 ( \13973 , \13972 , \12797 );
and \U$12258 ( \13974 , \13452 , \12958 );
and \U$12259 ( \13975 , \13376 , \12956 );
nor \U$12260 ( \13976 , \13974 , \13975 );
xnor \U$12261 ( \13977 , \13976 , \12984 );
xor \U$12262 ( \13978 , \13973 , \13977 );
and \U$12264 ( \13979 , \13431 , \13011 );
nor \U$12265 ( \13980 , 1'b0 , \13979 );
xnor \U$12266 ( \13981 , \13980 , 1'b0 );
xor \U$12267 ( \13982 , \13978 , \13981 );
xor \U$12268 ( \13983 , 1'b0 , \13982 );
and \U$12269 ( \13984 , \13117 , \13326 );
and \U$12270 ( \13985 , \13138 , \13324 );
nor \U$12271 ( \13986 , \13984 , \13985 );
xnor \U$12272 ( \13987 , \13986 , \13352 );
and \U$12273 ( \13988 , \13287 , \13384 );
and \U$12274 ( \13989 , \13161 , \13382 );
nor \U$12275 ( \13990 , \13988 , \13989 );
xnor \U$12276 ( \13991 , \13990 , \13410 );
xor \U$12277 ( \13992 , \13987 , \13991 );
and \U$12278 ( \13993 , \13347 , \13085 );
and \U$12279 ( \13994 , \13254 , \13083 );
nor \U$12280 ( \13995 , \13993 , \13994 );
xnor \U$12281 ( \13996 , \13995 , \13090 );
xor \U$12282 ( \13997 , \13992 , \13996 );
xor \U$12283 ( \13998 , \13983 , \13997 );
and \U$12284 ( \13999 , \13910 , \13914 );
and \U$12285 ( \14000 , \13914 , \13919 );
and \U$12286 ( \14001 , \13910 , \13919 );
or \U$12287 ( \14002 , \13999 , \14000 , \14001 );
and \U$12288 ( \14003 , \13946 , \13950 );
and \U$12289 ( \14004 , \13950 , \13955 );
and \U$12290 ( \14005 , \13946 , \13955 );
or \U$12291 ( \14006 , \14003 , \14004 , \14005 );
xor \U$12292 ( \14007 , \14002 , \14006 );
and \U$12293 ( \14008 , \13936 , \13939 );
or \U$12296 ( \14009 , \14008 , 1'b0 , 1'b0 );
xor \U$12297 ( \14010 , \14007 , \14009 );
xor \U$12298 ( \14011 , \13998 , \14010 );
xor \U$12299 ( \14012 , \13969 , \14011 );
and \U$12300 ( \14013 , \13891 , \13895 );
and \U$12301 ( \14014 , \13895 , \13900 );
and \U$12302 ( \14015 , \13891 , \13900 );
or \U$12303 ( \14016 , \14013 , \14014 , \14015 );
and \U$12305 ( \14017 , \13941 , \13956 );
or \U$12307 ( \14018 , 1'b0 , \14017 , 1'b0 );
xor \U$12308 ( \14019 , \14016 , \14018 );
and \U$12310 ( \14020 , \12979 , \13230 );
not \U$12311 ( \14021 , \14020 );
xnor \U$12312 ( \14022 , \14021 , \13224 );
xor \U$12313 ( \14023 , 1'b0 , \14022 );
and \U$12314 ( \14024 , \13006 , \13266 );
and \U$12315 ( \14025 , \12910 , \13264 );
nor \U$12316 ( \14026 , \14024 , \14025 );
xnor \U$12317 ( \14027 , \14026 , \13292 );
xor \U$12318 ( \14028 , \14023 , \14027 );
xor \U$12319 ( \14029 , \14019 , \14028 );
xor \U$12320 ( \14030 , \14012 , \14029 );
xor \U$12321 ( \14031 , \13967 , \14030 );
and \U$12322 ( \14032 , \13889 , \13922 );
and \U$12323 ( \14033 , \13922 , \13958 );
and \U$12324 ( \14034 , \13889 , \13958 );
or \U$12325 ( \14035 , \14032 , \14033 , \14034 );
nor \U$12326 ( \14036 , \14031 , \14035 );
nor \U$12327 ( \14037 , \13961 , \14036 );
nand \U$12328 ( \14038 , \13885 , \14037 );
and \U$12329 ( \14039 , \13969 , \14011 );
and \U$12330 ( \14040 , \14011 , \14029 );
and \U$12331 ( \14041 , \13969 , \14029 );
or \U$12332 ( \14042 , \14039 , \14040 , \14041 );
and \U$12333 ( \14043 , \14002 , \14006 );
and \U$12334 ( \14044 , \14006 , \14009 );
and \U$12335 ( \14045 , \14002 , \14009 );
or \U$12336 ( \14046 , \14043 , \14044 , \14045 );
and \U$12338 ( \14047 , \13982 , \13997 );
or \U$12340 ( \14048 , 1'b0 , \14047 , 1'b0 );
xor \U$12341 ( \14049 , \14046 , \14048 );
and \U$12342 ( \14050 , \13161 , \13384 );
and \U$12343 ( \14051 , \13117 , \13382 );
nor \U$12344 ( \14052 , \14050 , \14051 );
xnor \U$12345 ( \14053 , \14052 , \13410 );
and \U$12346 ( \14054 , \13254 , \13085 );
and \U$12347 ( \14055 , \13287 , \13083 );
nor \U$12348 ( \14056 , \14054 , \14055 );
xnor \U$12349 ( \14057 , \14056 , \13090 );
xor \U$12350 ( \14058 , \14053 , \14057 );
and \U$12351 ( \14059 , \13314 , \13020 );
and \U$12352 ( \14060 , \13347 , \13018 );
nor \U$12353 ( \14061 , \14059 , \14060 );
xnor \U$12354 ( \14062 , \14061 , \12797 );
xor \U$12355 ( \14063 , \14058 , \14062 );
xor \U$12356 ( \14064 , \14049 , \14063 );
xor \U$12357 ( \14065 , \14042 , \14064 );
and \U$12358 ( \14066 , \14016 , \14018 );
and \U$12359 ( \14067 , \14018 , \14028 );
and \U$12360 ( \14068 , \14016 , \14028 );
or \U$12361 ( \14069 , \14066 , \14067 , \14068 );
and \U$12362 ( \14070 , \13998 , \14010 );
xor \U$12363 ( \14071 , \14069 , \14070 );
not \U$12364 ( \14072 , \13224 );
and \U$12365 ( \14073 , \12910 , \13266 );
and \U$12366 ( \14074 , \12979 , \13264 );
nor \U$12367 ( \14075 , \14073 , \14074 );
xnor \U$12368 ( \14076 , \14075 , \13292 );
xor \U$12369 ( \14077 , \14072 , \14076 );
and \U$12370 ( \14078 , \13138 , \13326 );
and \U$12371 ( \14079 , \13006 , \13324 );
nor \U$12372 ( \14080 , \14078 , \14079 );
xnor \U$12373 ( \14081 , \14080 , \13352 );
xor \U$12374 ( \14082 , \14077 , \14081 );
and \U$12376 ( \14083 , \13376 , \12958 );
and \U$12377 ( \14084 , \13405 , \12956 );
nor \U$12378 ( \14085 , \14083 , \14084 );
xnor \U$12379 ( \14086 , \14085 , \12984 );
and \U$12381 ( \14087 , \13452 , \13011 );
nor \U$12382 ( \14088 , 1'b0 , \14087 );
xnor \U$12383 ( \14089 , \14088 , 1'b0 );
xor \U$12384 ( \14090 , \14086 , \14089 );
xor \U$12386 ( \14091 , \14090 , 1'b0 );
xor \U$12387 ( \14092 , 1'b1 , \14091 );
xor \U$12388 ( \14093 , \14082 , \14092 );
and \U$12390 ( \14094 , \14022 , \14027 );
or \U$12392 ( \14095 , 1'b0 , \14094 , 1'b0 );
and \U$12393 ( \14096 , \13987 , \13991 );
and \U$12394 ( \14097 , \13991 , \13996 );
and \U$12395 ( \14098 , \13987 , \13996 );
or \U$12396 ( \14099 , \14096 , \14097 , \14098 );
xor \U$12397 ( \14100 , \14095 , \14099 );
and \U$12398 ( \14101 , \13973 , \13977 );
and \U$12399 ( \14102 , \13977 , \13981 );
and \U$12400 ( \14103 , \13973 , \13981 );
or \U$12401 ( \14104 , \14101 , \14102 , \14103 );
xor \U$12402 ( \14105 , \14100 , \14104 );
xor \U$12403 ( \14106 , \14093 , \14105 );
xor \U$12404 ( \14107 , \14071 , \14106 );
xor \U$12405 ( \14108 , \14065 , \14107 );
and \U$12406 ( \14109 , \13965 , \13966 );
and \U$12407 ( \14110 , \13966 , \14030 );
and \U$12408 ( \14111 , \13965 , \14030 );
or \U$12409 ( \14112 , \14109 , \14110 , \14111 );
nor \U$12410 ( \14113 , \14108 , \14112 );
and \U$12411 ( \14114 , \14069 , \14070 );
and \U$12412 ( \14115 , \14070 , \14106 );
and \U$12413 ( \14116 , \14069 , \14106 );
or \U$12414 ( \14117 , \14114 , \14115 , \14116 );
and \U$12415 ( \14118 , \14072 , \14076 );
and \U$12416 ( \14119 , \14076 , \14081 );
and \U$12417 ( \14120 , \14072 , \14081 );
or \U$12418 ( \14121 , \14118 , \14119 , \14120 );
and \U$12419 ( \14122 , \14053 , \14057 );
and \U$12420 ( \14123 , \14057 , \14062 );
and \U$12421 ( \14124 , \14053 , \14062 );
or \U$12422 ( \14125 , \14122 , \14123 , \14124 );
xor \U$12423 ( \14126 , \14121 , \14125 );
and \U$12424 ( \14127 , \14086 , \14089 );
or \U$12427 ( \14128 , \14127 , 1'b0 , 1'b0 );
xor \U$12428 ( \14129 , \14126 , \14128 );
and \U$12429 ( \14130 , \14095 , \14099 );
and \U$12430 ( \14131 , \14099 , \14104 );
and \U$12431 ( \14132 , \14095 , \14104 );
or \U$12432 ( \14133 , \14130 , \14131 , \14132 );
and \U$12435 ( \14134 , 1'b1 , \14091 );
or \U$12437 ( \14135 , 1'b0 , \14134 , 1'b0 );
xor \U$12438 ( \14136 , \14133 , \14135 );
and \U$12439 ( \14137 , \13405 , \12958 );
and \U$12440 ( \14138 , \13314 , \12956 );
nor \U$12441 ( \14139 , \14137 , \14138 );
xnor \U$12442 ( \14140 , \14139 , \12984 );
and \U$12444 ( \14141 , \13376 , \13011 );
nor \U$12445 ( \14142 , 1'b0 , \14141 );
xnor \U$12446 ( \14143 , \14142 , 1'b0 );
xor \U$12447 ( \14144 , \14140 , \14143 );
xor \U$12449 ( \14145 , \14144 , 1'b0 );
and \U$12450 ( \14146 , \13117 , \13384 );
and \U$12451 ( \14147 , \13138 , \13382 );
nor \U$12452 ( \14148 , \14146 , \14147 );
xnor \U$12453 ( \14149 , \14148 , \13410 );
and \U$12454 ( \14150 , \13287 , \13085 );
and \U$12455 ( \14151 , \13161 , \13083 );
nor \U$12456 ( \14152 , \14150 , \14151 );
xnor \U$12457 ( \14153 , \14152 , \13090 );
xor \U$12458 ( \14154 , \14149 , \14153 );
and \U$12459 ( \14155 , \13347 , \13020 );
and \U$12460 ( \14156 , \13254 , \13018 );
nor \U$12461 ( \14157 , \14155 , \14156 );
xnor \U$12462 ( \14158 , \14157 , \12797 );
xor \U$12463 ( \14159 , \14154 , \14158 );
xor \U$12464 ( \14160 , \14145 , \14159 );
and \U$12466 ( \14161 , \12979 , \13266 );
not \U$12467 ( \14162 , \14161 );
xnor \U$12468 ( \14163 , \14162 , \13292 );
xor \U$12469 ( \14164 , 1'b0 , \14163 );
and \U$12470 ( \14165 , \13006 , \13326 );
and \U$12471 ( \14166 , \12910 , \13324 );
nor \U$12472 ( \14167 , \14165 , \14166 );
xnor \U$12473 ( \14168 , \14167 , \13352 );
xor \U$12474 ( \14169 , \14164 , \14168 );
xor \U$12475 ( \14170 , \14160 , \14169 );
xor \U$12476 ( \14171 , \14136 , \14170 );
xor \U$12477 ( \14172 , \14129 , \14171 );
xor \U$12478 ( \14173 , \14117 , \14172 );
and \U$12479 ( \14174 , \14046 , \14048 );
and \U$12480 ( \14175 , \14048 , \14063 );
and \U$12481 ( \14176 , \14046 , \14063 );
or \U$12482 ( \14177 , \14174 , \14175 , \14176 );
and \U$12483 ( \14178 , \14082 , \14092 );
and \U$12484 ( \14179 , \14092 , \14105 );
and \U$12485 ( \14180 , \14082 , \14105 );
or \U$12486 ( \14181 , \14178 , \14179 , \14180 );
xor \U$12487 ( \14182 , \14177 , \14181 );
xor \U$12489 ( \14183 , \14182 , 1'b1 );
xor \U$12490 ( \14184 , \14173 , \14183 );
and \U$12491 ( \14185 , \14042 , \14064 );
and \U$12492 ( \14186 , \14064 , \14107 );
and \U$12493 ( \14187 , \14042 , \14107 );
or \U$12494 ( \14188 , \14185 , \14186 , \14187 );
nor \U$12495 ( \14189 , \14184 , \14188 );
nor \U$12496 ( \14190 , \14113 , \14189 );
and \U$12497 ( \14191 , \14177 , \14181 );
and \U$12498 ( \14192 , \14181 , 1'b1 );
and \U$12499 ( \14193 , \14177 , 1'b1 );
or \U$12500 ( \14194 , \14191 , \14192 , \14193 );
and \U$12501 ( \14195 , \14129 , \14171 );
xor \U$12502 ( \14196 , \14194 , \14195 );
and \U$12503 ( \14197 , \14133 , \14135 );
and \U$12504 ( \14198 , \14135 , \14170 );
and \U$12505 ( \14199 , \14133 , \14170 );
or \U$12506 ( \14200 , \14197 , \14198 , \14199 );
and \U$12508 ( \14201 , \13405 , \13011 );
nor \U$12509 ( \14202 , 1'b0 , \14201 );
xnor \U$12510 ( \14203 , \14202 , 1'b0 );
xor \U$12512 ( \14204 , \14203 , 1'b0 );
xor \U$12514 ( \14205 , \14204 , 1'b0 );
and \U$12515 ( \14206 , \13161 , \13085 );
and \U$12516 ( \14207 , \13117 , \13083 );
nor \U$12517 ( \14208 , \14206 , \14207 );
xnor \U$12518 ( \14209 , \14208 , \13090 );
and \U$12519 ( \14210 , \13254 , \13020 );
and \U$12520 ( \14211 , \13287 , \13018 );
nor \U$12521 ( \14212 , \14210 , \14211 );
xnor \U$12522 ( \14213 , \14212 , \12797 );
xor \U$12523 ( \14214 , \14209 , \14213 );
and \U$12524 ( \14215 , \13314 , \12958 );
and \U$12525 ( \14216 , \13347 , \12956 );
nor \U$12526 ( \14217 , \14215 , \14216 );
xnor \U$12527 ( \14218 , \14217 , \12984 );
xor \U$12528 ( \14219 , \14214 , \14218 );
xor \U$12529 ( \14220 , \14205 , \14219 );
not \U$12530 ( \14221 , \13292 );
and \U$12531 ( \14222 , \12910 , \13326 );
and \U$12532 ( \14223 , \12979 , \13324 );
nor \U$12533 ( \14224 , \14222 , \14223 );
xnor \U$12534 ( \14225 , \14224 , \13352 );
xor \U$12535 ( \14226 , \14221 , \14225 );
and \U$12536 ( \14227 , \13138 , \13384 );
and \U$12537 ( \14228 , \13006 , \13382 );
nor \U$12538 ( \14229 , \14227 , \14228 );
xnor \U$12539 ( \14230 , \14229 , \13410 );
xor \U$12540 ( \14231 , \14226 , \14230 );
xor \U$12541 ( \14232 , \14220 , \14231 );
xor \U$12543 ( \14233 , \14232 , 1'b0 );
and \U$12545 ( \14234 , \14163 , \14168 );
or \U$12547 ( \14235 , 1'b0 , \14234 , 1'b0 );
and \U$12548 ( \14236 , \14149 , \14153 );
and \U$12549 ( \14237 , \14153 , \14158 );
and \U$12550 ( \14238 , \14149 , \14158 );
or \U$12551 ( \14239 , \14236 , \14237 , \14238 );
xor \U$12552 ( \14240 , \14235 , \14239 );
and \U$12553 ( \14241 , \14140 , \14143 );
or \U$12556 ( \14242 , \14241 , 1'b0 , 1'b0 );
xor \U$12557 ( \14243 , \14240 , \14242 );
xor \U$12558 ( \14244 , \14233 , \14243 );
xor \U$12559 ( \14245 , \14200 , \14244 );
and \U$12560 ( \14246 , \14121 , \14125 );
and \U$12561 ( \14247 , \14125 , \14128 );
and \U$12562 ( \14248 , \14121 , \14128 );
or \U$12563 ( \14249 , \14246 , \14247 , \14248 );
xor \U$12565 ( \14250 , \14249 , 1'b0 );
and \U$12566 ( \14251 , \14145 , \14159 );
and \U$12567 ( \14252 , \14159 , \14169 );
and \U$12568 ( \14253 , \14145 , \14169 );
or \U$12569 ( \14254 , \14251 , \14252 , \14253 );
xor \U$12570 ( \14255 , \14250 , \14254 );
xor \U$12571 ( \14256 , \14245 , \14255 );
xor \U$12572 ( \14257 , \14196 , \14256 );
and \U$12573 ( \14258 , \14117 , \14172 );
and \U$12574 ( \14259 , \14172 , \14183 );
and \U$12575 ( \14260 , \14117 , \14183 );
or \U$12576 ( \14261 , \14258 , \14259 , \14260 );
nor \U$12577 ( \14262 , \14257 , \14261 );
and \U$12578 ( \14263 , \14200 , \14244 );
and \U$12579 ( \14264 , \14244 , \14255 );
and \U$12580 ( \14265 , \14200 , \14255 );
or \U$12581 ( \14266 , \14263 , \14264 , \14265 );
and \U$12582 ( \14267 , \14235 , \14239 );
and \U$12583 ( \14268 , \14239 , \14242 );
and \U$12584 ( \14269 , \14235 , \14242 );
or \U$12585 ( \14270 , \14267 , \14268 , \14269 );
xor \U$12587 ( \14271 , \14270 , 1'b0 );
and \U$12588 ( \14272 , \14205 , \14219 );
and \U$12589 ( \14273 , \14219 , \14231 );
and \U$12590 ( \14274 , \14205 , \14231 );
or \U$12591 ( \14275 , \14272 , \14273 , \14274 );
xor \U$12592 ( \14276 , \14271 , \14275 );
xor \U$12593 ( \14277 , \14266 , \14276 );
and \U$12596 ( \14278 , \14249 , \14254 );
or \U$12597 ( \14279 , 1'b0 , 1'b0 , \14278 );
and \U$12600 ( \14280 , \14232 , \14243 );
or \U$12601 ( \14281 , 1'b0 , 1'b0 , \14280 );
xor \U$12602 ( \14282 , \14279 , \14281 );
and \U$12603 ( \14283 , \13117 , \13085 );
and \U$12604 ( \14284 , \13138 , \13083 );
nor \U$12605 ( \14285 , \14283 , \14284 );
xnor \U$12606 ( \14286 , \14285 , \13090 );
and \U$12607 ( \14287 , \13287 , \13020 );
and \U$12608 ( \14288 , \13161 , \13018 );
nor \U$12609 ( \14289 , \14287 , \14288 );
xnor \U$12610 ( \14290 , \14289 , \12797 );
xor \U$12611 ( \14291 , \14286 , \14290 );
and \U$12612 ( \14292 , \13347 , \12958 );
and \U$12613 ( \14293 , \13254 , \12956 );
nor \U$12614 ( \14294 , \14292 , \14293 );
xnor \U$12615 ( \14295 , \14294 , \12984 );
xor \U$12616 ( \14296 , \14291 , \14295 );
and \U$12618 ( \14297 , \12979 , \13326 );
not \U$12619 ( \14298 , \14297 );
xnor \U$12620 ( \14299 , \14298 , \13352 );
xor \U$12621 ( \14300 , 1'b0 , \14299 );
and \U$12622 ( \14301 , \13006 , \13384 );
and \U$12623 ( \14302 , \12910 , \13382 );
nor \U$12624 ( \14303 , \14301 , \14302 );
xnor \U$12625 ( \14304 , \14303 , \13410 );
xor \U$12626 ( \14305 , \14300 , \14304 );
xor \U$12627 ( \14306 , \14296 , \14305 );
and \U$12630 ( \14307 , \13314 , \13011 );
nor \U$12631 ( \14308 , 1'b0 , \14307 );
xnor \U$12632 ( \14309 , \14308 , 1'b0 );
xor \U$12634 ( \14310 , \14309 , 1'b0 );
xor \U$12636 ( \14311 , \14310 , 1'b0 );
xnor \U$12637 ( \14312 , 1'b0 , \14311 );
xor \U$12638 ( \14313 , \14306 , \14312 );
and \U$12639 ( \14314 , \14221 , \14225 );
and \U$12640 ( \14315 , \14225 , \14230 );
and \U$12641 ( \14316 , \14221 , \14230 );
or \U$12642 ( \14317 , \14314 , \14315 , \14316 );
and \U$12643 ( \14318 , \14209 , \14213 );
and \U$12644 ( \14319 , \14213 , \14218 );
and \U$12645 ( \14320 , \14209 , \14218 );
or \U$12646 ( \14321 , \14318 , \14319 , \14320 );
xor \U$12647 ( \14322 , \14317 , \14321 );
xor \U$12649 ( \14323 , \14322 , 1'b0 );
xor \U$12650 ( \14324 , \14313 , \14323 );
xor \U$12651 ( \14325 , \14282 , \14324 );
xor \U$12652 ( \14326 , \14277 , \14325 );
and \U$12653 ( \14327 , \14194 , \14195 );
and \U$12654 ( \14328 , \14195 , \14256 );
and \U$12655 ( \14329 , \14194 , \14256 );
or \U$12656 ( \14330 , \14327 , \14328 , \14329 );
nor \U$12657 ( \14331 , \14326 , \14330 );
nor \U$12658 ( \14332 , \14262 , \14331 );
nand \U$12659 ( \14333 , \14190 , \14332 );
nor \U$12660 ( \14334 , \14038 , \14333 );
and \U$12661 ( \14335 , \14279 , \14281 );
and \U$12662 ( \14336 , \14281 , \14324 );
and \U$12663 ( \14337 , \14279 , \14324 );
or \U$12664 ( \14338 , \14335 , \14336 , \14337 );
and \U$12665 ( \14339 , \14317 , \14321 );
or \U$12668 ( \14340 , \14339 , 1'b0 , 1'b0 );
or \U$12669 ( \14341 , 1'b0 , \14311 );
xor \U$12670 ( \14342 , \14340 , \14341 );
and \U$12671 ( \14343 , \14296 , \14305 );
xor \U$12672 ( \14344 , \14342 , \14343 );
xor \U$12673 ( \14345 , \14338 , \14344 );
and \U$12676 ( \14346 , \14270 , \14275 );
or \U$12677 ( \14347 , 1'b0 , 1'b0 , \14346 );
and \U$12678 ( \14348 , \14306 , \14312 );
and \U$12679 ( \14349 , \14312 , \14323 );
and \U$12680 ( \14350 , \14306 , \14323 );
or \U$12681 ( \14351 , \14348 , \14349 , \14350 );
xor \U$12682 ( \14352 , \14347 , \14351 );
and \U$12684 ( \14353 , \13161 , \13020 );
and \U$12685 ( \14354 , \13117 , \13018 );
nor \U$12686 ( \14355 , \14353 , \14354 );
xnor \U$12687 ( \14356 , \14355 , \12797 );
and \U$12688 ( \14357 , \13254 , \12958 );
and \U$12689 ( \14358 , \13287 , \12956 );
nor \U$12690 ( \14359 , \14357 , \14358 );
xnor \U$12691 ( \14360 , \14359 , \12984 );
xor \U$12692 ( \14361 , \14356 , \14360 );
and \U$12694 ( \14362 , \13347 , \13011 );
nor \U$12695 ( \14363 , 1'b0 , \14362 );
xnor \U$12696 ( \14364 , \14363 , 1'b0 );
xor \U$12697 ( \14365 , \14361 , \14364 );
xor \U$12698 ( \14366 , 1'b0 , \14365 );
not \U$12699 ( \14367 , \13352 );
and \U$12700 ( \14368 , \12910 , \13384 );
and \U$12701 ( \14369 , \12979 , \13382 );
nor \U$12702 ( \14370 , \14368 , \14369 );
xnor \U$12703 ( \14371 , \14370 , \13410 );
xor \U$12704 ( \14372 , \14367 , \14371 );
and \U$12705 ( \14373 , \13138 , \13085 );
and \U$12706 ( \14374 , \13006 , \13083 );
nor \U$12707 ( \14375 , \14373 , \14374 );
xnor \U$12708 ( \14376 , \14375 , \13090 );
xor \U$12709 ( \14377 , \14372 , \14376 );
xor \U$12710 ( \14378 , \14366 , \14377 );
xor \U$12712 ( \14379 , \14378 , 1'b0 );
and \U$12714 ( \14380 , \14299 , \14304 );
or \U$12716 ( \14381 , 1'b0 , \14380 , 1'b0 );
and \U$12717 ( \14382 , \14286 , \14290 );
and \U$12718 ( \14383 , \14290 , \14295 );
and \U$12719 ( \14384 , \14286 , \14295 );
or \U$12720 ( \14385 , \14382 , \14383 , \14384 );
xor \U$12721 ( \14386 , \14381 , \14385 );
xor \U$12723 ( \14387 , \14386 , 1'b0 );
xor \U$12724 ( \14388 , \14379 , \14387 );
xor \U$12725 ( \14389 , \14352 , \14388 );
xor \U$12726 ( \14390 , \14345 , \14389 );
and \U$12727 ( \14391 , \14266 , \14276 );
and \U$12728 ( \14392 , \14276 , \14325 );
and \U$12729 ( \14393 , \14266 , \14325 );
or \U$12730 ( \14394 , \14391 , \14392 , \14393 );
nor \U$12731 ( \14395 , \14390 , \14394 );
and \U$12732 ( \14396 , \14347 , \14351 );
and \U$12733 ( \14397 , \14351 , \14388 );
and \U$12734 ( \14398 , \14347 , \14388 );
or \U$12735 ( \14399 , \14396 , \14397 , \14398 );
and \U$12736 ( \14400 , \14381 , \14385 );
or \U$12739 ( \14401 , \14400 , 1'b0 , 1'b0 );
xor \U$12741 ( \14402 , \14401 , 1'b0 );
and \U$12743 ( \14403 , \14365 , \14377 );
or \U$12745 ( \14404 , 1'b0 , \14403 , 1'b0 );
xor \U$12746 ( \14405 , \14402 , \14404 );
xor \U$12747 ( \14406 , \14399 , \14405 );
and \U$12748 ( \14407 , \14340 , \14341 );
and \U$12749 ( \14408 , \14341 , \14343 );
and \U$12750 ( \14409 , \14340 , \14343 );
or \U$12751 ( \14410 , \14407 , \14408 , \14409 );
and \U$12754 ( \14411 , \14378 , \14387 );
or \U$12755 ( \14412 , 1'b0 , 1'b0 , \14411 );
xor \U$12756 ( \14413 , \14410 , \14412 );
and \U$12757 ( \14414 , \13117 , \13020 );
and \U$12758 ( \14415 , \13138 , \13018 );
nor \U$12759 ( \14416 , \14414 , \14415 );
xnor \U$12760 ( \14417 , \14416 , \12797 );
and \U$12761 ( \14418 , \13287 , \12958 );
and \U$12762 ( \14419 , \13161 , \12956 );
nor \U$12763 ( \14420 , \14418 , \14419 );
xnor \U$12764 ( \14421 , \14420 , \12984 );
xor \U$12765 ( \14422 , \14417 , \14421 );
and \U$12767 ( \14423 , \13254 , \13011 );
nor \U$12768 ( \14424 , 1'b0 , \14423 );
xnor \U$12769 ( \14425 , \14424 , 1'b0 );
xor \U$12770 ( \14426 , \14422 , \14425 );
and \U$12772 ( \14427 , \12979 , \13384 );
not \U$12773 ( \14428 , \14427 );
xnor \U$12774 ( \14429 , \14428 , \13410 );
xor \U$12775 ( \14430 , 1'b0 , \14429 );
and \U$12776 ( \14431 , \13006 , \13085 );
and \U$12777 ( \14432 , \12910 , \13083 );
nor \U$12778 ( \14433 , \14431 , \14432 );
xnor \U$12779 ( \14434 , \14433 , \13090 );
xor \U$12780 ( \14435 , \14430 , \14434 );
xor \U$12781 ( \14436 , \14426 , \14435 );
xor \U$12783 ( \14437 , \14436 , 1'b1 );
and \U$12784 ( \14438 , \14367 , \14371 );
and \U$12785 ( \14439 , \14371 , \14376 );
and \U$12786 ( \14440 , \14367 , \14376 );
or \U$12787 ( \14441 , \14438 , \14439 , \14440 );
and \U$12788 ( \14442 , \14356 , \14360 );
and \U$12789 ( \14443 , \14360 , \14364 );
and \U$12790 ( \14444 , \14356 , \14364 );
or \U$12791 ( \14445 , \14442 , \14443 , \14444 );
xor \U$12792 ( \14446 , \14441 , \14445 );
xor \U$12794 ( \14447 , \14446 , 1'b0 );
xor \U$12795 ( \14448 , \14437 , \14447 );
xor \U$12796 ( \14449 , \14413 , \14448 );
xor \U$12797 ( \14450 , \14406 , \14449 );
and \U$12798 ( \14451 , \14338 , \14344 );
and \U$12799 ( \14452 , \14344 , \14389 );
and \U$12800 ( \14453 , \14338 , \14389 );
or \U$12801 ( \14454 , \14451 , \14452 , \14453 );
nor \U$12802 ( \14455 , \14450 , \14454 );
nor \U$12803 ( \14456 , \14395 , \14455 );
and \U$12804 ( \14457 , \14410 , \14412 );
and \U$12805 ( \14458 , \14412 , \14448 );
and \U$12806 ( \14459 , \14410 , \14448 );
or \U$12807 ( \14460 , \14457 , \14458 , \14459 );
and \U$12808 ( \14461 , \14441 , \14445 );
or \U$12811 ( \14462 , \14461 , 1'b0 , 1'b0 );
xor \U$12813 ( \14463 , \14462 , 1'b0 );
and \U$12814 ( \14464 , \14426 , \14435 );
xor \U$12815 ( \14465 , \14463 , \14464 );
xor \U$12816 ( \14466 , \14460 , \14465 );
and \U$12819 ( \14467 , \14401 , \14404 );
or \U$12820 ( \14468 , 1'b0 , 1'b0 , \14467 );
and \U$12821 ( \14469 , \14436 , 1'b1 );
and \U$12822 ( \14470 , 1'b1 , \14447 );
and \U$12823 ( \14471 , \14436 , \14447 );
or \U$12824 ( \14472 , \14469 , \14470 , \14471 );
xor \U$12825 ( \14473 , \14468 , \14472 );
and \U$12827 ( \14474 , \13161 , \12958 );
and \U$12828 ( \14475 , \13117 , \12956 );
nor \U$12829 ( \14476 , \14474 , \14475 );
xnor \U$12830 ( \14477 , \14476 , \12984 );
and \U$12832 ( \14478 , \13287 , \13011 );
nor \U$12833 ( \14479 , 1'b0 , \14478 );
xnor \U$12834 ( \14480 , \14479 , 1'b0 );
xor \U$12835 ( \14481 , \14477 , \14480 );
xor \U$12837 ( \14482 , \14481 , 1'b0 );
xor \U$12838 ( \14483 , 1'b0 , \14482 );
not \U$12839 ( \14484 , \13410 );
and \U$12840 ( \14485 , \12910 , \13085 );
and \U$12841 ( \14486 , \12979 , \13083 );
nor \U$12842 ( \14487 , \14485 , \14486 );
xnor \U$12843 ( \14488 , \14487 , \13090 );
xor \U$12844 ( \14489 , \14484 , \14488 );
and \U$12845 ( \14490 , \13138 , \13020 );
and \U$12846 ( \14491 , \13006 , \13018 );
nor \U$12847 ( \14492 , \14490 , \14491 );
xnor \U$12848 ( \14493 , \14492 , \12797 );
xor \U$12849 ( \14494 , \14489 , \14493 );
xor \U$12850 ( \14495 , \14483 , \14494 );
xor \U$12852 ( \14496 , \14495 , 1'b0 );
and \U$12854 ( \14497 , \14429 , \14434 );
or \U$12856 ( \14498 , 1'b0 , \14497 , 1'b0 );
and \U$12857 ( \14499 , \14417 , \14421 );
and \U$12858 ( \14500 , \14421 , \14425 );
and \U$12859 ( \14501 , \14417 , \14425 );
or \U$12860 ( \14502 , \14499 , \14500 , \14501 );
xor \U$12861 ( \14503 , \14498 , \14502 );
xor \U$12863 ( \14504 , \14503 , 1'b0 );
xor \U$12864 ( \14505 , \14496 , \14504 );
xor \U$12865 ( \14506 , \14473 , \14505 );
xor \U$12866 ( \14507 , \14466 , \14506 );
and \U$12867 ( \14508 , \14399 , \14405 );
and \U$12868 ( \14509 , \14405 , \14449 );
and \U$12869 ( \14510 , \14399 , \14449 );
or \U$12870 ( \14511 , \14508 , \14509 , \14510 );
nor \U$12871 ( \14512 , \14507 , \14511 );
and \U$12872 ( \14513 , \14468 , \14472 );
and \U$12873 ( \14514 , \14472 , \14505 );
and \U$12874 ( \14515 , \14468 , \14505 );
or \U$12875 ( \14516 , \14513 , \14514 , \14515 );
and \U$12876 ( \14517 , \14498 , \14502 );
or \U$12879 ( \14518 , \14517 , 1'b0 , 1'b0 );
xor \U$12881 ( \14519 , \14518 , 1'b0 );
and \U$12883 ( \14520 , \14482 , \14494 );
or \U$12885 ( \14521 , 1'b0 , \14520 , 1'b0 );
xor \U$12886 ( \14522 , \14519 , \14521 );
xor \U$12887 ( \14523 , \14516 , \14522 );
and \U$12890 ( \14524 , \14462 , \14464 );
or \U$12891 ( \14525 , 1'b0 , 1'b0 , \14524 );
and \U$12894 ( \14526 , \14495 , \14504 );
or \U$12895 ( \14527 , 1'b0 , 1'b0 , \14526 );
xor \U$12896 ( \14528 , \14525 , \14527 );
xor \U$12897 ( \14529 , \13141 , \13164 );
xor \U$12899 ( \14530 , \14529 , 1'b0 );
xor \U$12901 ( \14531 , 1'b0 , \13091 );
xor \U$12902 ( \14532 , \14531 , \13095 );
xor \U$12903 ( \14533 , \14530 , \14532 );
xor \U$12905 ( \14534 , \14533 , 1'b1 );
and \U$12906 ( \14535 , \14484 , \14488 );
and \U$12907 ( \14536 , \14488 , \14493 );
and \U$12908 ( \14537 , \14484 , \14493 );
or \U$12909 ( \14538 , \14535 , \14536 , \14537 );
and \U$12910 ( \14539 , \14477 , \14480 );
or \U$12913 ( \14540 , \14539 , 1'b0 , 1'b0 );
xor \U$12914 ( \14541 , \14538 , \14540 );
xor \U$12916 ( \14542 , \14541 , 1'b0 );
xor \U$12917 ( \14543 , \14534 , \14542 );
xor \U$12918 ( \14544 , \14528 , \14543 );
xor \U$12919 ( \14545 , \14523 , \14544 );
and \U$12920 ( \14546 , \14460 , \14465 );
and \U$12921 ( \14547 , \14465 , \14506 );
and \U$12922 ( \14548 , \14460 , \14506 );
or \U$12923 ( \14549 , \14546 , \14547 , \14548 );
nor \U$12924 ( \14550 , \14545 , \14549 );
nor \U$12925 ( \14551 , \14512 , \14550 );
nand \U$12926 ( \14552 , \14456 , \14551 );
and \U$12927 ( \14553 , \14525 , \14527 );
and \U$12928 ( \14554 , \14527 , \14543 );
and \U$12929 ( \14555 , \14525 , \14543 );
or \U$12930 ( \14556 , \14553 , \14554 , \14555 );
and \U$12931 ( \14557 , \14538 , \14540 );
or \U$12934 ( \14558 , \14557 , 1'b0 , 1'b0 );
xor \U$12936 ( \14559 , \14558 , 1'b0 );
and \U$12937 ( \14560 , \14530 , \14532 );
xor \U$12938 ( \14561 , \14559 , \14560 );
xor \U$12939 ( \14562 , \14556 , \14561 );
and \U$12942 ( \14563 , \14518 , \14521 );
or \U$12943 ( \14564 , 1'b0 , 1'b0 , \14563 );
and \U$12944 ( \14565 , \14533 , 1'b1 );
and \U$12945 ( \14566 , 1'b1 , \14542 );
and \U$12946 ( \14567 , \14533 , \14542 );
or \U$12947 ( \14568 , \14565 , \14566 , \14567 );
xor \U$12948 ( \14569 , \14564 , \14568 );
xor \U$12950 ( \14570 , 1'b0 , \13173 );
xor \U$12951 ( \14571 , \14570 , \13184 );
xor \U$12953 ( \14572 , \14571 , 1'b0 );
xor \U$12954 ( \14573 , \13097 , \13166 );
xor \U$12956 ( \14574 , \14573 , 1'b0 );
xor \U$12957 ( \14575 , \14572 , \14574 );
xor \U$12958 ( \14576 , \14569 , \14575 );
xor \U$12959 ( \14577 , \14562 , \14576 );
and \U$12960 ( \14578 , \14516 , \14522 );
and \U$12961 ( \14579 , \14522 , \14544 );
and \U$12962 ( \14580 , \14516 , \14544 );
or \U$12963 ( \14581 , \14578 , \14579 , \14580 );
nor \U$12964 ( \14582 , \14577 , \14581 );
and \U$12965 ( \14583 , \14564 , \14568 );
and \U$12966 ( \14584 , \14568 , \14575 );
and \U$12967 ( \14585 , \14564 , \14575 );
or \U$12968 ( \14586 , \14583 , \14584 , \14585 );
xor \U$12970 ( \14587 , \13168 , 1'b0 );
xor \U$12971 ( \14588 , \14587 , \13186 );
xor \U$12972 ( \14589 , \14586 , \14588 );
and \U$12975 ( \14590 , \14558 , \14560 );
or \U$12976 ( \14591 , 1'b0 , 1'b0 , \14590 );
and \U$12979 ( \14592 , \14571 , \14574 );
or \U$12980 ( \14593 , 1'b0 , 1'b0 , \14592 );
xor \U$12981 ( \14594 , \14591 , \14593 );
xor \U$12982 ( \14595 , \13196 , 1'b1 );
xor \U$12983 ( \14596 , \14595 , \13203 );
xor \U$12984 ( \14597 , \14594 , \14596 );
xor \U$12985 ( \14598 , \14589 , \14597 );
and \U$12986 ( \14599 , \14556 , \14561 );
and \U$12987 ( \14600 , \14561 , \14576 );
and \U$12988 ( \14601 , \14556 , \14576 );
or \U$12989 ( \14602 , \14599 , \14600 , \14601 );
nor \U$12990 ( \14603 , \14598 , \14602 );
nor \U$12991 ( \14604 , \14582 , \14603 );
and \U$12992 ( \14605 , \14591 , \14593 );
and \U$12993 ( \14606 , \14593 , \14596 );
and \U$12994 ( \14607 , \14591 , \14596 );
or \U$12995 ( \14608 , \14605 , \14606 , \14607 );
and \U$12997 ( \14609 , \13193 , \13195 );
xor \U$12998 ( \14610 , 1'b0 , \14609 );
xor \U$12999 ( \14611 , \14608 , \14610 );
xor \U$13000 ( \14612 , \13188 , \13206 );
xor \U$13001 ( \14613 , \14612 , \13209 );
xor \U$13002 ( \14614 , \14611 , \14613 );
and \U$13003 ( \14615 , \14586 , \14588 );
and \U$13004 ( \14616 , \14588 , \14597 );
and \U$13005 ( \14617 , \14586 , \14597 );
or \U$13006 ( \14618 , \14615 , \14616 , \14617 );
nor \U$13007 ( \14619 , \14614 , \14618 );
xor \U$13009 ( \14620 , \13212 , 1'b0 );
xor \U$13010 ( \14621 , \14620 , \13214 );
and \U$13011 ( \14622 , \14608 , \14610 );
and \U$13012 ( \14623 , \14610 , \14613 );
and \U$13013 ( \14624 , \14608 , \14613 );
or \U$13014 ( \14625 , \14622 , \14623 , \14624 );
nor \U$13015 ( \14626 , \14621 , \14625 );
nor \U$13016 ( \14627 , \14619 , \14626 );
nand \U$13017 ( \14628 , \14604 , \14627 );
nor \U$13018 ( \14629 , \14552 , \14628 );
nand \U$13019 ( \14630 , \14334 , \14629 );
and \U$13020 ( \14631 , \13431 , \13230 );
and \U$13021 ( \14632 , \13452 , \13227 );
nor \U$13022 ( \14633 , \14631 , \14632 );
xnor \U$13023 ( \14634 , \14633 , \13224 );
and \U$13024 ( \14635 , \13476 , \13266 );
and \U$13025 ( \14636 , \13497 , \13264 );
nor \U$13026 ( \14637 , \14635 , \14636 );
xnor \U$13027 ( \14638 , \14637 , \13292 );
and \U$13028 ( \14639 , \14634 , \14638 );
and \U$13029 ( \14640 , \13524 , \13326 );
and \U$13030 ( \14641 , \13545 , \13324 );
nor \U$13031 ( \14642 , \14640 , \14641 );
xnor \U$13032 ( \14643 , \14642 , \13352 );
and \U$13033 ( \14644 , \14638 , \14643 );
and \U$13034 ( \14645 , \14634 , \14643 );
or \U$13035 ( \14646 , \14639 , \14644 , \14645 );
and \U$13036 ( \14647 , \13545 , \13326 );
and \U$13037 ( \14648 , \13476 , \13324 );
nor \U$13038 ( \14649 , \14647 , \14648 );
xnor \U$13039 ( \14650 , \14649 , \13352 );
and \U$13040 ( \14651 , \13568 , \13384 );
and \U$13041 ( \14652 , \13524 , \13382 );
nor \U$13042 ( \14653 , \14651 , \14652 );
xnor \U$13043 ( \14654 , \14653 , \13410 );
xor \U$13044 ( \14655 , \14650 , \14654 );
nand \U$13045 ( \14656 , \13701 , \13083 );
xnor \U$13046 ( \14657 , \14656 , \13090 );
xor \U$13047 ( \14658 , \14655 , \14657 );
and \U$13048 ( \14659 , \14646 , \14658 );
and \U$13049 ( \14660 , \13452 , \13230 );
and \U$13050 ( \14661 , \13376 , \13227 );
nor \U$13051 ( \14662 , \14660 , \14661 );
xnor \U$13052 ( \14663 , \14662 , \13224 );
xor \U$13053 ( \14664 , \13090 , \14663 );
and \U$13054 ( \14665 , \13497 , \13266 );
and \U$13055 ( \14666 , \13431 , \13264 );
nor \U$13056 ( \14667 , \14665 , \14666 );
xnor \U$13057 ( \14668 , \14667 , \13292 );
xor \U$13058 ( \14669 , \14664 , \14668 );
and \U$13059 ( \14670 , \14658 , \14669 );
and \U$13060 ( \14671 , \14646 , \14669 );
or \U$13061 ( \14672 , \14659 , \14670 , \14671 );
and \U$13062 ( \14673 , \13701 , \13085 );
and \U$13063 ( \14674 , \13568 , \13083 );
nor \U$13064 ( \14675 , \14673 , \14674 );
xnor \U$13065 ( \14676 , \14675 , \13090 );
and \U$13066 ( \14677 , \13376 , \13230 );
and \U$13067 ( \14678 , \13405 , \13227 );
nor \U$13068 ( \14679 , \14677 , \14678 );
xnor \U$13069 ( \14680 , \14679 , \13224 );
and \U$13070 ( \14681 , \13431 , \13266 );
and \U$13071 ( \14682 , \13452 , \13264 );
nor \U$13072 ( \14683 , \14681 , \14682 );
xnor \U$13073 ( \14684 , \14683 , \13292 );
xor \U$13074 ( \14685 , \14680 , \14684 );
and \U$13075 ( \14686 , \13476 , \13326 );
and \U$13076 ( \14687 , \13497 , \13324 );
nor \U$13077 ( \14688 , \14686 , \14687 );
xnor \U$13078 ( \14689 , \14688 , \13352 );
xor \U$13079 ( \14690 , \14685 , \14689 );
xor \U$13080 ( \14691 , \14676 , \14690 );
xor \U$13081 ( \14692 , \14672 , \14691 );
and \U$13082 ( \14693 , \13090 , \14663 );
and \U$13083 ( \14694 , \14663 , \14668 );
and \U$13084 ( \14695 , \13090 , \14668 );
or \U$13085 ( \14696 , \14693 , \14694 , \14695 );
and \U$13086 ( \14697 , \14650 , \14654 );
and \U$13087 ( \14698 , \14654 , \14657 );
and \U$13088 ( \14699 , \14650 , \14657 );
or \U$13089 ( \14700 , \14697 , \14698 , \14699 );
xor \U$13090 ( \14701 , \14696 , \14700 );
and \U$13091 ( \14702 , \13524 , \13384 );
and \U$13092 ( \14703 , \13545 , \13382 );
nor \U$13093 ( \14704 , \14702 , \14703 );
xnor \U$13094 ( \14705 , \14704 , \13410 );
xor \U$13095 ( \14706 , \14701 , \14705 );
xor \U$13096 ( \14707 , \14692 , \14706 );
and \U$13097 ( \14708 , \13497 , \13230 );
and \U$13098 ( \14709 , \13431 , \13227 );
nor \U$13099 ( \14710 , \14708 , \14709 );
xnor \U$13100 ( \14711 , \14710 , \13224 );
and \U$13101 ( \14712 , \13410 , \14711 );
and \U$13102 ( \14713 , \13545 , \13266 );
and \U$13103 ( \14714 , \13476 , \13264 );
nor \U$13104 ( \14715 , \14713 , \14714 );
xnor \U$13105 ( \14716 , \14715 , \13292 );
and \U$13106 ( \14717 , \14711 , \14716 );
and \U$13107 ( \14718 , \13410 , \14716 );
or \U$13108 ( \14719 , \14712 , \14717 , \14718 );
and \U$13109 ( \14720 , \13568 , \13326 );
and \U$13110 ( \14721 , \13524 , \13324 );
nor \U$13111 ( \14722 , \14720 , \14721 );
xnor \U$13112 ( \14723 , \14722 , \13352 );
nand \U$13113 ( \14724 , \13701 , \13382 );
xnor \U$13114 ( \14725 , \14724 , \13410 );
and \U$13115 ( \14726 , \14723 , \14725 );
and \U$13116 ( \14727 , \14719 , \14726 );
and \U$13117 ( \14728 , \13701 , \13384 );
and \U$13118 ( \14729 , \13568 , \13382 );
nor \U$13119 ( \14730 , \14728 , \14729 );
xnor \U$13120 ( \14731 , \14730 , \13410 );
and \U$13121 ( \14732 , \14726 , \14731 );
and \U$13122 ( \14733 , \14719 , \14731 );
or \U$13123 ( \14734 , \14727 , \14732 , \14733 );
xor \U$13124 ( \14735 , \14646 , \14658 );
xor \U$13125 ( \14736 , \14735 , \14669 );
and \U$13126 ( \14737 , \14734 , \14736 );
nor \U$13127 ( \14738 , \14707 , \14737 );
and \U$13128 ( \14739 , \14680 , \14684 );
and \U$13129 ( \14740 , \14684 , \14689 );
and \U$13130 ( \14741 , \14680 , \14689 );
or \U$13131 ( \14742 , \14739 , \14740 , \14741 );
nand \U$13132 ( \14743 , \13701 , \13018 );
xnor \U$13133 ( \14744 , \14743 , \12797 );
xor \U$13134 ( \14745 , \14742 , \14744 );
and \U$13135 ( \14746 , \13497 , \13326 );
and \U$13136 ( \14747 , \13431 , \13324 );
nor \U$13137 ( \14748 , \14746 , \14747 );
xnor \U$13138 ( \14749 , \14748 , \13352 );
and \U$13139 ( \14750 , \13545 , \13384 );
and \U$13140 ( \14751 , \13476 , \13382 );
nor \U$13141 ( \14752 , \14750 , \14751 );
xnor \U$13142 ( \14753 , \14752 , \13410 );
xor \U$13143 ( \14754 , \14749 , \14753 );
and \U$13144 ( \14755 , \13568 , \13085 );
and \U$13145 ( \14756 , \13524 , \13083 );
nor \U$13146 ( \14757 , \14755 , \14756 );
xnor \U$13147 ( \14758 , \14757 , \13090 );
xor \U$13148 ( \14759 , \14754 , \14758 );
xor \U$13149 ( \14760 , \14745 , \14759 );
and \U$13150 ( \14761 , \14696 , \14700 );
and \U$13151 ( \14762 , \14700 , \14705 );
and \U$13152 ( \14763 , \14696 , \14705 );
or \U$13153 ( \14764 , \14761 , \14762 , \14763 );
and \U$13154 ( \14765 , \14676 , \14690 );
xor \U$13155 ( \14766 , \14764 , \14765 );
and \U$13156 ( \14767 , \13405 , \13230 );
and \U$13157 ( \14768 , \13314 , \13227 );
nor \U$13158 ( \14769 , \14767 , \14768 );
xnor \U$13159 ( \14770 , \14769 , \13224 );
xor \U$13160 ( \14771 , \12797 , \14770 );
and \U$13161 ( \14772 , \13452 , \13266 );
and \U$13162 ( \14773 , \13376 , \13264 );
nor \U$13163 ( \14774 , \14772 , \14773 );
xnor \U$13164 ( \14775 , \14774 , \13292 );
xor \U$13165 ( \14776 , \14771 , \14775 );
xor \U$13166 ( \14777 , \14766 , \14776 );
xor \U$13167 ( \14778 , \14760 , \14777 );
and \U$13168 ( \14779 , \14672 , \14691 );
and \U$13169 ( \14780 , \14691 , \14706 );
and \U$13170 ( \14781 , \14672 , \14706 );
or \U$13171 ( \14782 , \14779 , \14780 , \14781 );
nor \U$13172 ( \14783 , \14778 , \14782 );
nor \U$13173 ( \14784 , \14738 , \14783 );
and \U$13174 ( \14785 , \14764 , \14765 );
and \U$13175 ( \14786 , \14765 , \14776 );
and \U$13176 ( \14787 , \14764 , \14776 );
or \U$13177 ( \14788 , \14785 , \14786 , \14787 );
and \U$13178 ( \14789 , \14742 , \14744 );
and \U$13179 ( \14790 , \14744 , \14759 );
and \U$13180 ( \14791 , \14742 , \14759 );
or \U$13181 ( \14792 , \14789 , \14790 , \14791 );
and \U$13182 ( \14793 , \13314 , \13230 );
and \U$13183 ( \14794 , \13347 , \13227 );
nor \U$13184 ( \14795 , \14793 , \14794 );
xnor \U$13185 ( \14796 , \14795 , \13224 );
and \U$13186 ( \14797 , \13376 , \13266 );
and \U$13187 ( \14798 , \13405 , \13264 );
nor \U$13188 ( \14799 , \14797 , \14798 );
xnor \U$13189 ( \14800 , \14799 , \13292 );
xor \U$13190 ( \14801 , \14796 , \14800 );
and \U$13191 ( \14802 , \13431 , \13326 );
and \U$13192 ( \14803 , \13452 , \13324 );
nor \U$13193 ( \14804 , \14802 , \14803 );
xnor \U$13194 ( \14805 , \14804 , \13352 );
xor \U$13195 ( \14806 , \14801 , \14805 );
xor \U$13196 ( \14807 , \14792 , \14806 );
and \U$13197 ( \14808 , \12797 , \14770 );
and \U$13198 ( \14809 , \14770 , \14775 );
and \U$13199 ( \14810 , \12797 , \14775 );
or \U$13200 ( \14811 , \14808 , \14809 , \14810 );
and \U$13201 ( \14812 , \14749 , \14753 );
and \U$13202 ( \14813 , \14753 , \14758 );
and \U$13203 ( \14814 , \14749 , \14758 );
or \U$13204 ( \14815 , \14812 , \14813 , \14814 );
xor \U$13205 ( \14816 , \14811 , \14815 );
and \U$13206 ( \14817 , \13476 , \13384 );
and \U$13207 ( \14818 , \13497 , \13382 );
nor \U$13208 ( \14819 , \14817 , \14818 );
xnor \U$13209 ( \14820 , \14819 , \13410 );
and \U$13210 ( \14821 , \13524 , \13085 );
and \U$13211 ( \14822 , \13545 , \13083 );
nor \U$13212 ( \14823 , \14821 , \14822 );
xnor \U$13213 ( \14824 , \14823 , \13090 );
xor \U$13214 ( \14825 , \14820 , \14824 );
and \U$13215 ( \14826 , \13701 , \13020 );
and \U$13216 ( \14827 , \13568 , \13018 );
nor \U$13217 ( \14828 , \14826 , \14827 );
xnor \U$13218 ( \14829 , \14828 , \12797 );
xor \U$13219 ( \14830 , \14825 , \14829 );
xor \U$13220 ( \14831 , \14816 , \14830 );
xor \U$13221 ( \14832 , \14807 , \14831 );
xor \U$13222 ( \14833 , \14788 , \14832 );
and \U$13223 ( \14834 , \14760 , \14777 );
nor \U$13224 ( \14835 , \14833 , \14834 );
and \U$13225 ( \14836 , \14792 , \14806 );
and \U$13226 ( \14837 , \14806 , \14831 );
and \U$13227 ( \14838 , \14792 , \14831 );
or \U$13228 ( \14839 , \14836 , \14837 , \14838 );
and \U$13229 ( \14840 , \14811 , \14815 );
and \U$13230 ( \14841 , \14815 , \14830 );
and \U$13231 ( \14842 , \14811 , \14830 );
or \U$13232 ( \14843 , \14840 , \14841 , \14842 );
nand \U$13233 ( \14844 , \13701 , \12956 );
xnor \U$13234 ( \14845 , \14844 , \12984 );
and \U$13235 ( \14846 , \13452 , \13326 );
and \U$13236 ( \14847 , \13376 , \13324 );
nor \U$13237 ( \14848 , \14846 , \14847 );
xnor \U$13238 ( \14849 , \14848 , \13352 );
and \U$13239 ( \14850 , \13497 , \13384 );
and \U$13240 ( \14851 , \13431 , \13382 );
nor \U$13241 ( \14852 , \14850 , \14851 );
xnor \U$13242 ( \14853 , \14852 , \13410 );
xor \U$13243 ( \14854 , \14849 , \14853 );
and \U$13244 ( \14855 , \13545 , \13085 );
and \U$13245 ( \14856 , \13476 , \13083 );
nor \U$13246 ( \14857 , \14855 , \14856 );
xnor \U$13247 ( \14858 , \14857 , \13090 );
xor \U$13248 ( \14859 , \14854 , \14858 );
xor \U$13249 ( \14860 , \14845 , \14859 );
and \U$13250 ( \14861 , \13347 , \13230 );
and \U$13251 ( \14862 , \13254 , \13227 );
nor \U$13252 ( \14863 , \14861 , \14862 );
xnor \U$13253 ( \14864 , \14863 , \13224 );
xor \U$13254 ( \14865 , \12984 , \14864 );
and \U$13255 ( \14866 , \13405 , \13266 );
and \U$13256 ( \14867 , \13314 , \13264 );
nor \U$13257 ( \14868 , \14866 , \14867 );
xnor \U$13258 ( \14869 , \14868 , \13292 );
xor \U$13259 ( \14870 , \14865 , \14869 );
xor \U$13260 ( \14871 , \14860 , \14870 );
xor \U$13261 ( \14872 , \14843 , \14871 );
and \U$13262 ( \14873 , \14796 , \14800 );
and \U$13263 ( \14874 , \14800 , \14805 );
and \U$13264 ( \14875 , \14796 , \14805 );
or \U$13265 ( \14876 , \14873 , \14874 , \14875 );
and \U$13266 ( \14877 , \14820 , \14824 );
and \U$13267 ( \14878 , \14824 , \14829 );
and \U$13268 ( \14879 , \14820 , \14829 );
or \U$13269 ( \14880 , \14877 , \14878 , \14879 );
xor \U$13270 ( \14881 , \14876 , \14880 );
and \U$13271 ( \14882 , \13568 , \13020 );
and \U$13272 ( \14883 , \13524 , \13018 );
nor \U$13273 ( \14884 , \14882 , \14883 );
xnor \U$13274 ( \14885 , \14884 , \12797 );
xor \U$13275 ( \14886 , \14881 , \14885 );
xor \U$13276 ( \14887 , \14872 , \14886 );
xor \U$13277 ( \14888 , \14839 , \14887 );
and \U$13278 ( \14889 , \14788 , \14832 );
nor \U$13279 ( \14890 , \14888 , \14889 );
nor \U$13280 ( \14891 , \14835 , \14890 );
nand \U$13281 ( \14892 , \14784 , \14891 );
and \U$13282 ( \14893 , \14843 , \14871 );
and \U$13283 ( \14894 , \14871 , \14886 );
and \U$13284 ( \14895 , \14843 , \14886 );
or \U$13285 ( \14896 , \14893 , \14894 , \14895 );
xor \U$13286 ( \14897 , \13756 , \13760 );
xor \U$13287 ( \14898 , \14897 , \13765 );
and \U$13288 ( \14899 , \12984 , \14864 );
and \U$13289 ( \14900 , \14864 , \14869 );
and \U$13290 ( \14901 , \12984 , \14869 );
or \U$13291 ( \14902 , \14899 , \14900 , \14901 );
and \U$13292 ( \14903 , \14849 , \14853 );
and \U$13293 ( \14904 , \14853 , \14858 );
and \U$13294 ( \14905 , \14849 , \14858 );
or \U$13295 ( \14906 , \14903 , \14904 , \14905 );
xor \U$13296 ( \14907 , \14902 , \14906 );
and \U$13297 ( \14908 , \13701 , \12958 );
and \U$13298 ( \14909 , \13568 , \12956 );
nor \U$13299 ( \14910 , \14908 , \14909 );
xnor \U$13300 ( \14911 , \14910 , \12984 );
xor \U$13301 ( \14912 , \14907 , \14911 );
xor \U$13302 ( \14913 , \14898 , \14912 );
xor \U$13303 ( \14914 , \14896 , \14913 );
and \U$13304 ( \14915 , \14876 , \14880 );
and \U$13305 ( \14916 , \14880 , \14885 );
and \U$13306 ( \14917 , \14876 , \14885 );
or \U$13307 ( \14918 , \14915 , \14916 , \14917 );
and \U$13308 ( \14919 , \14845 , \14859 );
and \U$13309 ( \14920 , \14859 , \14870 );
and \U$13310 ( \14921 , \14845 , \14870 );
or \U$13311 ( \14922 , \14919 , \14920 , \14921 );
xor \U$13312 ( \14923 , \14918 , \14922 );
xor \U$13313 ( \14924 , \13772 , \13776 );
xor \U$13314 ( \14925 , \14924 , \13781 );
xor \U$13315 ( \14926 , \14923 , \14925 );
xor \U$13316 ( \14927 , \14914 , \14926 );
and \U$13317 ( \14928 , \14839 , \14887 );
nor \U$13318 ( \14929 , \14927 , \14928 );
and \U$13319 ( \14930 , \14918 , \14922 );
and \U$13320 ( \14931 , \14922 , \14925 );
and \U$13321 ( \14932 , \14918 , \14925 );
or \U$13322 ( \14933 , \14930 , \14931 , \14932 );
and \U$13323 ( \14934 , \14898 , \14912 );
xor \U$13324 ( \14935 , \14933 , \14934 );
and \U$13325 ( \14936 , \14902 , \14906 );
and \U$13326 ( \14937 , \14906 , \14911 );
and \U$13327 ( \14938 , \14902 , \14911 );
or \U$13328 ( \14939 , \14936 , \14937 , \14938 );
xor \U$13329 ( \14940 , \13792 , \13794 );
xor \U$13330 ( \14941 , \14939 , \14940 );
xor \U$13331 ( \14942 , \13768 , \13784 );
xor \U$13332 ( \14943 , \14942 , \13787 );
xor \U$13333 ( \14944 , \14941 , \14943 );
xor \U$13334 ( \14945 , \14935 , \14944 );
and \U$13335 ( \14946 , \14896 , \14913 );
and \U$13336 ( \14947 , \14913 , \14926 );
and \U$13337 ( \14948 , \14896 , \14926 );
or \U$13338 ( \14949 , \14946 , \14947 , \14948 );
nor \U$13339 ( \14950 , \14945 , \14949 );
nor \U$13340 ( \14951 , \14929 , \14950 );
and \U$13341 ( \14952 , \14939 , \14940 );
and \U$13342 ( \14953 , \14940 , \14943 );
and \U$13343 ( \14954 , \14939 , \14943 );
or \U$13344 ( \14955 , \14952 , \14953 , \14954 );
xor \U$13345 ( \14956 , \13655 , \13671 );
xor \U$13346 ( \14957 , \14956 , \13706 );
xor \U$13347 ( \14958 , \14955 , \14957 );
xor \U$13348 ( \14959 , \13790 , \13795 );
xor \U$13349 ( \14960 , \14959 , \13798 );
xor \U$13350 ( \14961 , \14958 , \14960 );
and \U$13351 ( \14962 , \14933 , \14934 );
and \U$13352 ( \14963 , \14934 , \14944 );
and \U$13353 ( \14964 , \14933 , \14944 );
or \U$13354 ( \14965 , \14962 , \14963 , \14964 );
nor \U$13355 ( \14966 , \14961 , \14965 );
xor \U$13356 ( \14967 , \13801 , \13802 );
xor \U$13357 ( \14968 , \14967 , \13805 );
and \U$13358 ( \14969 , \14955 , \14957 );
and \U$13359 ( \14970 , \14957 , \14960 );
and \U$13360 ( \14971 , \14955 , \14960 );
or \U$13361 ( \14972 , \14969 , \14970 , \14971 );
nor \U$13362 ( \14973 , \14968 , \14972 );
nor \U$13363 ( \14974 , \14966 , \14973 );
nand \U$13364 ( \14975 , \14951 , \14974 );
nor \U$13365 ( \14976 , \14892 , \14975 );
and \U$13366 ( \14977 , \13545 , \13230 );
and \U$13367 ( \14978 , \13476 , \13227 );
nor \U$13368 ( \14979 , \14977 , \14978 );
xnor \U$13369 ( \14980 , \14979 , \13224 );
and \U$13370 ( \14981 , \13352 , \14980 );
and \U$13371 ( \14982 , \13568 , \13266 );
and \U$13372 ( \14983 , \13524 , \13264 );
nor \U$13373 ( \14984 , \14982 , \14983 );
xnor \U$13374 ( \14985 , \14984 , \13292 );
and \U$13375 ( \14986 , \14980 , \14985 );
and \U$13376 ( \14987 , \13352 , \14985 );
or \U$13377 ( \14988 , \14981 , \14986 , \14987 );
and \U$13378 ( \14989 , \13476 , \13230 );
and \U$13379 ( \14990 , \13497 , \13227 );
nor \U$13380 ( \14991 , \14989 , \14990 );
xnor \U$13381 ( \14992 , \14991 , \13224 );
and \U$13382 ( \14993 , \13524 , \13266 );
and \U$13383 ( \14994 , \13545 , \13264 );
nor \U$13384 ( \14995 , \14993 , \14994 );
xnor \U$13385 ( \14996 , \14995 , \13292 );
xor \U$13386 ( \14997 , \14992 , \14996 );
and \U$13387 ( \14998 , \13701 , \13326 );
and \U$13388 ( \14999 , \13568 , \13324 );
nor \U$13389 ( \15000 , \14998 , \14999 );
xnor \U$13390 ( \15001 , \15000 , \13352 );
xor \U$13391 ( \15002 , \14997 , \15001 );
xor \U$13392 ( \15003 , \14988 , \15002 );
nand \U$13393 ( \15004 , \13701 , \13324 );
xnor \U$13394 ( \15005 , \15004 , \13352 );
xor \U$13395 ( \15006 , \13352 , \14980 );
xor \U$13396 ( \15007 , \15006 , \14985 );
and \U$13397 ( \15008 , \15005 , \15007 );
nor \U$13398 ( \15009 , \15003 , \15008 );
and \U$13399 ( \15010 , \14992 , \14996 );
and \U$13400 ( \15011 , \14996 , \15001 );
and \U$13401 ( \15012 , \14992 , \15001 );
or \U$13402 ( \15013 , \15010 , \15011 , \15012 );
xor \U$13403 ( \15014 , \14723 , \14725 );
xor \U$13404 ( \15015 , \15013 , \15014 );
xor \U$13405 ( \15016 , \13410 , \14711 );
xor \U$13406 ( \15017 , \15016 , \14716 );
xor \U$13407 ( \15018 , \15015 , \15017 );
and \U$13408 ( \15019 , \14988 , \15002 );
nor \U$13409 ( \15020 , \15018 , \15019 );
nor \U$13410 ( \15021 , \15009 , \15020 );
xor \U$13411 ( \15022 , \14634 , \14638 );
xor \U$13412 ( \15023 , \15022 , \14643 );
xor \U$13413 ( \15024 , \14719 , \14726 );
xor \U$13414 ( \15025 , \15024 , \14731 );
xor \U$13415 ( \15026 , \15023 , \15025 );
and \U$13416 ( \15027 , \15013 , \15014 );
and \U$13417 ( \15028 , \15014 , \15017 );
and \U$13418 ( \15029 , \15013 , \15017 );
or \U$13419 ( \15030 , \15027 , \15028 , \15029 );
nor \U$13420 ( \15031 , \15026 , \15030 );
xor \U$13421 ( \15032 , \14734 , \14736 );
and \U$13422 ( \15033 , \15023 , \15025 );
nor \U$13423 ( \15034 , \15032 , \15033 );
nor \U$13424 ( \15035 , \15031 , \15034 );
nand \U$13425 ( \15036 , \15021 , \15035 );
and \U$13426 ( \15037 , \13524 , \13230 );
and \U$13427 ( \15038 , \13545 , \13227 );
nor \U$13428 ( \15039 , \15037 , \15038 );
xnor \U$13429 ( \15040 , \15039 , \13224 );
and \U$13430 ( \15041 , \13701 , \13266 );
and \U$13431 ( \15042 , \13568 , \13264 );
nor \U$13432 ( \15043 , \15041 , \15042 );
xnor \U$13433 ( \15044 , \15043 , \13292 );
xor \U$13434 ( \15045 , \15040 , \15044 );
and \U$13435 ( \15046 , \13568 , \13230 );
and \U$13436 ( \15047 , \13524 , \13227 );
nor \U$13437 ( \15048 , \15046 , \15047 );
xnor \U$13438 ( \15049 , \15048 , \13224 );
and \U$13439 ( \15050 , \15049 , \13292 );
nor \U$13440 ( \15051 , \15045 , \15050 );
xor \U$13441 ( \15052 , \15005 , \15007 );
and \U$13442 ( \15053 , \15040 , \15044 );
nor \U$13443 ( \15054 , \15052 , \15053 );
nor \U$13444 ( \15055 , \15051 , \15054 );
xor \U$13445 ( \15056 , \15049 , \13292 );
nand \U$13446 ( \15057 , \13701 , \13264 );
xnor \U$13447 ( \15058 , \15057 , \13292 );
nor \U$13448 ( \15059 , \15056 , \15058 );
and \U$13449 ( \15060 , \13701 , \13230 );
and \U$13450 ( \15061 , \13568 , \13227 );
nor \U$13451 ( \15062 , \15060 , \15061 );
xnor \U$13452 ( \15063 , \15062 , \13224 );
nand \U$13453 ( \15064 , \13701 , \13227 );
xnor \U$13454 ( \15065 , \15064 , \13224 );
and \U$13455 ( \15066 , \15065 , \13224 );
nand \U$13456 ( \15067 , \15063 , \15066 );
or \U$13457 ( \15068 , \15059 , \15067 );
nand \U$13458 ( \15069 , \15056 , \15058 );
nand \U$13459 ( \15070 , \15068 , \15069 );
and \U$13460 ( \15071 , \15055 , \15070 );
nand \U$13461 ( \15072 , \15045 , \15050 );
or \U$13462 ( \15073 , \15054 , \15072 );
nand \U$13463 ( \15074 , \15052 , \15053 );
nand \U$13464 ( \15075 , \15073 , \15074 );
nor \U$13465 ( \15076 , \15071 , \15075 );
or \U$13466 ( \15077 , \15036 , \15076 );
nand \U$13467 ( \15078 , \15003 , \15008 );
or \U$13468 ( \15079 , \15020 , \15078 );
nand \U$13469 ( \15080 , \15018 , \15019 );
nand \U$13470 ( \15081 , \15079 , \15080 );
and \U$13471 ( \15082 , \15035 , \15081 );
nand \U$13472 ( \15083 , \15026 , \15030 );
or \U$13473 ( \15084 , \15034 , \15083 );
nand \U$13474 ( \15085 , \15032 , \15033 );
nand \U$13475 ( \15086 , \15084 , \15085 );
nor \U$13476 ( \15087 , \15082 , \15086 );
nand \U$13477 ( \15088 , \15077 , \15087 );
and \U$13478 ( \15089 , \14976 , \15088 );
nand \U$13479 ( \15090 , \14707 , \14737 );
or \U$13480 ( \15091 , \14783 , \15090 );
nand \U$13481 ( \15092 , \14778 , \14782 );
nand \U$13482 ( \15093 , \15091 , \15092 );
and \U$13483 ( \15094 , \14891 , \15093 );
nand \U$13484 ( \15095 , \14833 , \14834 );
or \U$13485 ( \15096 , \14890 , \15095 );
nand \U$13486 ( \15097 , \14888 , \14889 );
nand \U$13487 ( \15098 , \15096 , \15097 );
nor \U$13488 ( \15099 , \15094 , \15098 );
or \U$13489 ( \15100 , \14975 , \15099 );
nand \U$13490 ( \15101 , \14927 , \14928 );
or \U$13491 ( \15102 , \14950 , \15101 );
nand \U$13492 ( \15103 , \14945 , \14949 );
nand \U$13493 ( \15104 , \15102 , \15103 );
and \U$13494 ( \15105 , \14974 , \15104 );
nand \U$13495 ( \15106 , \14961 , \14965 );
or \U$13496 ( \15107 , \14973 , \15106 );
nand \U$13497 ( \15108 , \14968 , \14972 );
nand \U$13498 ( \15109 , \15107 , \15108 );
nor \U$13499 ( \15110 , \15105 , \15109 );
nand \U$13500 ( \15111 , \15100 , \15110 );
nor \U$13501 ( \15112 , \15089 , \15111 );
or \U$13502 ( \15113 , \14630 , \15112 );
nand \U$13503 ( \15114 , \13752 , \13808 );
or \U$13504 ( \15115 , \13884 , \15114 );
nand \U$13505 ( \15116 , \13882 , \13883 );
nand \U$13506 ( \15117 , \15115 , \15116 );
and \U$13507 ( \15118 , \14037 , \15117 );
nand \U$13508 ( \15119 , \13959 , \13960 );
or \U$13509 ( \15120 , \14036 , \15119 );
nand \U$13510 ( \15121 , \14031 , \14035 );
nand \U$13511 ( \15122 , \15120 , \15121 );
nor \U$13512 ( \15123 , \15118 , \15122 );
or \U$13513 ( \15124 , \14333 , \15123 );
nand \U$13514 ( \15125 , \14108 , \14112 );
or \U$13515 ( \15126 , \14189 , \15125 );
nand \U$13516 ( \15127 , \14184 , \14188 );
nand \U$13517 ( \15128 , \15126 , \15127 );
and \U$13518 ( \15129 , \14332 , \15128 );
nand \U$13519 ( \15130 , \14257 , \14261 );
or \U$13520 ( \15131 , \14331 , \15130 );
nand \U$13521 ( \15132 , \14326 , \14330 );
nand \U$13522 ( \15133 , \15131 , \15132 );
nor \U$13523 ( \15134 , \15129 , \15133 );
nand \U$13524 ( \15135 , \15124 , \15134 );
and \U$13525 ( \15136 , \14629 , \15135 );
nand \U$13526 ( \15137 , \14390 , \14394 );
or \U$13527 ( \15138 , \14455 , \15137 );
nand \U$13528 ( \15139 , \14450 , \14454 );
nand \U$13529 ( \15140 , \15138 , \15139 );
and \U$13530 ( \15141 , \14551 , \15140 );
nand \U$13531 ( \15142 , \14507 , \14511 );
or \U$13532 ( \15143 , \14550 , \15142 );
nand \U$13533 ( \15144 , \14545 , \14549 );
nand \U$13534 ( \15145 , \15143 , \15144 );
nor \U$13535 ( \15146 , \15141 , \15145 );
or \U$13536 ( \15147 , \14628 , \15146 );
nand \U$13537 ( \15148 , \14577 , \14581 );
or \U$13538 ( \15149 , \14603 , \15148 );
nand \U$13539 ( \15150 , \14598 , \14602 );
nand \U$13540 ( \15151 , \15149 , \15150 );
and \U$13541 ( \15152 , \14627 , \15151 );
nand \U$13542 ( \15153 , \14614 , \14618 );
or \U$13543 ( \15154 , \14626 , \15153 );
nand \U$13544 ( \15155 , \14621 , \14625 );
nand \U$13545 ( \15156 , \15154 , \15155 );
nor \U$13546 ( \15157 , \15152 , \15156 );
nand \U$13547 ( \15158 , \15147 , \15157 );
nor \U$13548 ( \15159 , \15136 , \15158 );
nand \U$13549 ( \15160 , \15113 , \15159 );
not \U$13550 ( \15161 , \15160 );
xor \U$13551 ( \15162 , \13220 , \15161 );
buf \U$13552 ( \15163 , \15162 );
buf \U$13553 ( \15164 , RI2b5e785db0d0_14);
buf \U$13554 ( \15165 , RI2b5e785db058_15);
buf \U$13555 ( \15166 , RI2b5e785dafe0_16);
buf \U$13556 ( \15167 , RI2b5e785daf68_17);
buf \U$13557 ( \15168 , RI2b5e785daef0_18);
buf \U$13558 ( \15169 , RI2b5e785dae78_19);
buf \U$13559 ( \15170 , RI2b5e785dae00_20);
buf \U$13560 ( \15171 , RI2b5e785dad88_21);
buf \U$13561 ( \15172 , RI2b5e785dad10_22);
buf \U$13562 ( \15173 , RI2b5e785dac98_23);
buf \U$13563 ( \15174 , RI2b5e785dac20_24);
buf \U$13564 ( \15175 , RI2b5e785daba8_25);
not \U$13565 ( \15176 , RI2b5e785ae328_614);
buf \U$13566 ( \15177 , \15176 );
and \U$13567 ( \15178 , \15175 , \15177 );
and \U$13568 ( \15179 , \15174 , \15178 );
and \U$13569 ( \15180 , \15173 , \15179 );
and \U$13570 ( \15181 , \15172 , \15180 );
and \U$13571 ( \15182 , \15171 , \15181 );
and \U$13572 ( \15183 , \15170 , \15182 );
and \U$13573 ( \15184 , \15169 , \15183 );
and \U$13574 ( \15185 , \15168 , \15184 );
and \U$13575 ( \15186 , \15167 , \15185 );
and \U$13576 ( \15187 , \15166 , \15186 );
and \U$13577 ( \15188 , \15165 , \15187 );
xor \U$13578 ( \15189 , \15164 , \15188 );
buf \U$13579 ( \15190 , \15189 );
buf \U$13580 ( \15191 , \15190 );
not \U$13581 ( \15192 , \15191 );
nor \U$13582 ( \15193 , \12412 , \12416 , \12420 , \12424 , \12429 );
and \U$13583 ( \15194 , RI2b5e785daab8_27, \15193 );
and \U$13584 ( \15195 , \12412 , \12416 , \12420 , \12424 , \12429 );
and \U$13585 ( \15196 , RI2b5e785495b8_40, \15195 );
and \U$13586 ( \15197 , \12434 , \12416 , \12420 , \12424 , \12429 );
and \U$13587 ( \15198 , RI2b5e78538920_53, \15197 );
and \U$13588 ( \15199 , \12412 , \12437 , \12420 , \12424 , \12429 );
and \U$13589 ( \15200 , RI2b5e784a63a8_66, \15199 );
and \U$13590 ( \15201 , \12434 , \12437 , \12420 , \12424 , \12429 );
and \U$13591 ( \15202 , RI2b5e78495710_79, \15201 );
and \U$13592 ( \15203 , \12412 , \12416 , \12442 , \12424 , \12429 );
and \U$13593 ( \15204 , RI2b5e784950f8_92, \15203 );
and \U$13594 ( \15205 , \12434 , \12416 , \12442 , \12424 , \12429 );
and \U$13595 ( \15206 , RI2b5e78403bf8_105, \15205 );
and \U$13596 ( \15207 , \12412 , \12437 , \12442 , \12424 , \12429 );
and \U$13597 ( \15208 , RI2b5e775b1ed8_118, \15207 );
and \U$13598 ( \15209 , \12434 , \12437 , \12442 , \12424 , \12429 );
and \U$13599 ( \15210 , RI2b5e775b18c0_131, \15209 );
nor \U$13600 ( \15211 , \12434 , \12437 , \12442 , \12424 , \12428 );
and \U$13601 ( \15212 , RI2b5e7750b858_144, \15211 );
nor \U$13602 ( \15213 , \12412 , \12437 , \12442 , \12424 , \12428 );
and \U$13603 ( \15214 , RI2b5e774ff030_157, \15213 );
nor \U$13604 ( \15215 , \12434 , \12416 , \12442 , \12424 , \12428 );
and \U$13605 ( \15216 , RI2b5e774f6048_170, \15215 );
nor \U$13606 ( \15217 , \12412 , \12416 , \12442 , \12424 , \12428 );
and \U$13607 ( \15218 , RI2b5e774ea630_183, \15217 );
nor \U$13608 ( \15219 , \12434 , \12437 , \12420 , \12424 , \12428 );
and \U$13609 ( \15220 , RI2b5e774dde08_196, \15219 );
nor \U$13610 ( \15221 , \12412 , \12437 , \12420 , \12424 , \12428 );
and \U$13611 ( \15222 , RI2b5e774d4e20_209, \15221 );
nor \U$13612 ( \15223 , \12434 , \12416 , \12420 , \12424 , \12428 );
and \U$13613 ( \15224 , RI2b5e785f3d60_222, \15223 );
nor \U$13614 ( \15225 , \12412 , \12416 , \12420 , \12424 , \12428 );
and \U$13615 ( \15226 , RI2b5e785eb138_235, \15225 );
or \U$13616 ( \15227 , \15194 , \15196 , \15198 , \15200 , \15202 , \15204 , \15206 , \15208 , \15210 , \15212 , \15214 , \15216 , \15218 , \15220 , \15222 , \15224 , \15226 );
buf \U$13617 ( \15228 , \12428 );
buf \U$13618 ( \15229 , \12412 );
buf \U$13619 ( \15230 , \12416 );
buf \U$13620 ( \15231 , \12420 );
buf \U$13621 ( \15232 , \12424 );
or \U$13622 ( \15233 , \15229 , \15230 , \15231 , \15232 );
and \U$13623 ( \15234 , \15228 , \15233 );
buf \U$13624 ( \15235 , \15234 );
_DC r143b ( \15236_nR143b , \15227 , \15235 );
buf \U$13625 ( \15237 , \15236_nR143b );
and \U$13626 ( \15238 , \15192 , \15237 );
xor \U$13627 ( \15239 , \15165 , \15187 );
buf \U$13628 ( \15240 , \15239 );
buf \U$13629 ( \15241 , \15240 );
not \U$13630 ( \15242 , \15241 );
and \U$13631 ( \15243 , RI2b5e785daa40_28, \15193 );
and \U$13632 ( \15244 , RI2b5e78549540_41, \15195 );
and \U$13633 ( \15245 , RI2b5e785388a8_54, \15197 );
and \U$13634 ( \15246 , RI2b5e784a6330_67, \15199 );
and \U$13635 ( \15247 , RI2b5e78495698_80, \15201 );
and \U$13636 ( \15248 , RI2b5e78495080_93, \15203 );
and \U$13637 ( \15249 , RI2b5e78403b80_106, \15205 );
and \U$13638 ( \15250 , RI2b5e775b1e60_119, \15207 );
and \U$13639 ( \15251 , RI2b5e7750bdf8_132, \15209 );
and \U$13640 ( \15252 , RI2b5e774ff5d0_145, \15211 );
and \U$13641 ( \15253 , RI2b5e774f65e8_158, \15213 );
and \U$13642 ( \15254 , RI2b5e774eabd0_171, \15215 );
and \U$13643 ( \15255 , RI2b5e774de3a8_184, \15217 );
and \U$13644 ( \15256 , RI2b5e774d53c0_197, \15219 );
and \U$13645 ( \15257 , RI2b5e785f4300_210, \15221 );
and \U$13646 ( \15258 , RI2b5e785f3ce8_223, \15223 );
and \U$13647 ( \15259 , RI2b5e785eb0c0_236, \15225 );
or \U$13648 ( \15260 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 );
_DC r1454 ( \15261_nR1454 , \15260 , \15235 );
buf \U$13649 ( \15262 , \15261_nR1454 );
and \U$13650 ( \15263 , \15242 , \15262 );
xor \U$13651 ( \15264 , \15166 , \15186 );
buf \U$13652 ( \15265 , \15264 );
buf \U$13653 ( \15266 , \15265 );
not \U$13654 ( \15267 , \15266 );
and \U$13655 ( \15268 , RI2b5e785da9c8_29, \15193 );
and \U$13656 ( \15269 , RI2b5e785494c8_42, \15195 );
and \U$13657 ( \15270 , RI2b5e78538830_55, \15197 );
and \U$13658 ( \15271 , RI2b5e784a62b8_68, \15199 );
and \U$13659 ( \15272 , RI2b5e78495620_81, \15201 );
and \U$13660 ( \15273 , RI2b5e78495008_94, \15203 );
and \U$13661 ( \15274 , RI2b5e78403b08_107, \15205 );
and \U$13662 ( \15275 , RI2b5e775b1de8_120, \15207 );
and \U$13663 ( \15276 , RI2b5e7750bd80_133, \15209 );
and \U$13664 ( \15277 , RI2b5e774ff558_146, \15211 );
and \U$13665 ( \15278 , RI2b5e774f6570_159, \15213 );
and \U$13666 ( \15279 , RI2b5e774eab58_172, \15215 );
and \U$13667 ( \15280 , RI2b5e774de330_185, \15217 );
and \U$13668 ( \15281 , RI2b5e774d5348_198, \15219 );
and \U$13669 ( \15282 , RI2b5e785f4288_211, \15221 );
and \U$13670 ( \15283 , RI2b5e785f3658_224, \15223 );
and \U$13671 ( \15284 , RI2b5e785eb048_237, \15225 );
or \U$13672 ( \15285 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 );
_DC r146d ( \15286_nR146d , \15285 , \15235 );
buf \U$13673 ( \15287 , \15286_nR146d );
and \U$13674 ( \15288 , \15267 , \15287 );
xor \U$13675 ( \15289 , \15167 , \15185 );
buf \U$13676 ( \15290 , \15289 );
buf \U$13677 ( \15291 , \15290 );
not \U$13678 ( \15292 , \15291 );
and \U$13679 ( \15293 , RI2b5e785da950_30, \15193 );
and \U$13680 ( \15294 , RI2b5e78549450_43, \15195 );
and \U$13681 ( \15295 , RI2b5e785387b8_56, \15197 );
and \U$13682 ( \15296 , RI2b5e784a6240_69, \15199 );
and \U$13683 ( \15297 , RI2b5e784955a8_82, \15201 );
and \U$13684 ( \15298 , RI2b5e78494f90_95, \15203 );
and \U$13685 ( \15299 , RI2b5e78403a90_108, \15205 );
and \U$13686 ( \15300 , RI2b5e775b1d70_121, \15207 );
and \U$13687 ( \15301 , RI2b5e7750bd08_134, \15209 );
and \U$13688 ( \15302 , RI2b5e774ff4e0_147, \15211 );
and \U$13689 ( \15303 , RI2b5e774f64f8_160, \15213 );
and \U$13690 ( \15304 , RI2b5e774eaae0_173, \15215 );
and \U$13691 ( \15305 , RI2b5e774de2b8_186, \15217 );
and \U$13692 ( \15306 , RI2b5e774d52d0_199, \15219 );
and \U$13693 ( \15307 , RI2b5e785f4210_212, \15221 );
and \U$13694 ( \15308 , RI2b5e785eb5e8_225, \15223 );
and \U$13695 ( \15309 , RI2b5e785e6c50_238, \15225 );
or \U$13696 ( \15310 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 );
_DC r1486 ( \15311_nR1486 , \15310 , \15235 );
buf \U$13697 ( \15312 , \15311_nR1486 );
and \U$13698 ( \15313 , \15292 , \15312 );
xor \U$13699 ( \15314 , \15168 , \15184 );
buf \U$13700 ( \15315 , \15314 );
buf \U$13701 ( \15316 , \15315 );
not \U$13702 ( \15317 , \15316 );
and \U$13703 ( \15318 , RI2b5e785da8d8_31, \15193 );
and \U$13704 ( \15319 , RI2b5e785493d8_44, \15195 );
and \U$13705 ( \15320 , RI2b5e78538740_57, \15197 );
and \U$13706 ( \15321 , RI2b5e784a61c8_70, \15199 );
and \U$13707 ( \15322 , RI2b5e78495530_83, \15201 );
and \U$13708 ( \15323 , RI2b5e78494f18_96, \15203 );
and \U$13709 ( \15324 , RI2b5e78403a18_109, \15205 );
and \U$13710 ( \15325 , RI2b5e775b1cf8_122, \15207 );
and \U$13711 ( \15326 , RI2b5e7750bc90_135, \15209 );
and \U$13712 ( \15327 , RI2b5e774ff468_148, \15211 );
and \U$13713 ( \15328 , RI2b5e774f6480_161, \15213 );
and \U$13714 ( \15329 , RI2b5e774eaa68_174, \15215 );
and \U$13715 ( \15330 , RI2b5e774de240_187, \15217 );
and \U$13716 ( \15331 , RI2b5e774d5258_200, \15219 );
and \U$13717 ( \15332 , RI2b5e785f4198_213, \15221 );
and \U$13718 ( \15333 , RI2b5e785eb570_226, \15223 );
and \U$13719 ( \15334 , RI2b5e785e6bd8_239, \15225 );
or \U$13720 ( \15335 , \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 );
_DC r149f ( \15336_nR149f , \15335 , \15235 );
buf \U$13721 ( \15337 , \15336_nR149f );
and \U$13722 ( \15338 , \15317 , \15337 );
xor \U$13723 ( \15339 , \15169 , \15183 );
buf \U$13724 ( \15340 , \15339 );
buf \U$13725 ( \15341 , \15340 );
not \U$13726 ( \15342 , \15341 );
and \U$13727 ( \15343 , RI2b5e785da860_32, \15193 );
and \U$13728 ( \15344 , RI2b5e78549360_45, \15195 );
and \U$13729 ( \15345 , RI2b5e785386c8_58, \15197 );
and \U$13730 ( \15346 , RI2b5e784a6150_71, \15199 );
and \U$13731 ( \15347 , RI2b5e784954b8_84, \15201 );
and \U$13732 ( \15348 , RI2b5e78494ea0_97, \15203 );
and \U$13733 ( \15349 , RI2b5e784039a0_110, \15205 );
and \U$13734 ( \15350 , RI2b5e775b1c80_123, \15207 );
and \U$13735 ( \15351 , RI2b5e7750bc18_136, \15209 );
and \U$13736 ( \15352 , RI2b5e774ff3f0_149, \15211 );
and \U$13737 ( \15353 , RI2b5e774f6408_162, \15213 );
and \U$13738 ( \15354 , RI2b5e774ea9f0_175, \15215 );
and \U$13739 ( \15355 , RI2b5e774de1c8_188, \15217 );
and \U$13740 ( \15356 , RI2b5e774d51e0_201, \15219 );
and \U$13741 ( \15357 , RI2b5e785f4120_214, \15221 );
and \U$13742 ( \15358 , RI2b5e785eb4f8_227, \15223 );
and \U$13743 ( \15359 , RI2b5e785e64d0_240, \15225 );
or \U$13744 ( \15360 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 );
_DC r14b8 ( \15361_nR14b8 , \15360 , \15235 );
buf \U$13745 ( \15362 , \15361_nR14b8 );
and \U$13746 ( \15363 , \15342 , \15362 );
xor \U$13747 ( \15364 , \15170 , \15182 );
buf \U$13748 ( \15365 , \15364 );
buf \U$13749 ( \15366 , \15365 );
not \U$13750 ( \15367 , \15366 );
and \U$13751 ( \15368 , RI2b5e78549900_33, \15193 );
and \U$13752 ( \15369 , RI2b5e78538c68_46, \15195 );
and \U$13753 ( \15370 , RI2b5e78538650_59, \15197 );
and \U$13754 ( \15371 , RI2b5e784a60d8_72, \15199 );
and \U$13755 ( \15372 , RI2b5e78495440_85, \15201 );
and \U$13756 ( \15373 , RI2b5e78494e28_98, \15203 );
and \U$13757 ( \15374 , RI2b5e78403928_111, \15205 );
and \U$13758 ( \15375 , RI2b5e775b1c08_124, \15207 );
and \U$13759 ( \15376 , RI2b5e7750bba0_137, \15209 );
and \U$13760 ( \15377 , RI2b5e774ff378_150, \15211 );
and \U$13761 ( \15378 , RI2b5e774f6390_163, \15213 );
and \U$13762 ( \15379 , RI2b5e774ea978_176, \15215 );
and \U$13763 ( \15380 , RI2b5e774de150_189, \15217 );
and \U$13764 ( \15381 , RI2b5e774d5168_202, \15219 );
and \U$13765 ( \15382 , RI2b5e785f40a8_215, \15221 );
and \U$13766 ( \15383 , RI2b5e785eb480_228, \15223 );
and \U$13767 ( \15384 , RI2b5e785da608_241, \15225 );
or \U$13768 ( \15385 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 );
_DC r14d1 ( \15386_nR14d1 , \15385 , \15235 );
buf \U$13769 ( \15387 , \15386_nR14d1 );
and \U$13770 ( \15388 , \15367 , \15387 );
xor \U$13771 ( \15389 , \15171 , \15181 );
buf \U$13772 ( \15390 , \15389 );
buf \U$13773 ( \15391 , \15390 );
not \U$13774 ( \15392 , \15391 );
and \U$13775 ( \15393 , RI2b5e78549888_34, \15193 );
and \U$13776 ( \15394 , RI2b5e78538bf0_47, \15195 );
and \U$13777 ( \15395 , RI2b5e785385d8_60, \15197 );
and \U$13778 ( \15396 , RI2b5e784a6060_73, \15199 );
and \U$13779 ( \15397 , RI2b5e784953c8_86, \15201 );
and \U$13780 ( \15398 , RI2b5e78403ec8_99, \15203 );
and \U$13781 ( \15399 , RI2b5e775b21a8_112, \15205 );
and \U$13782 ( \15400 , RI2b5e775b1b90_125, \15207 );
and \U$13783 ( \15401 , RI2b5e7750bb28_138, \15209 );
and \U$13784 ( \15402 , RI2b5e774ff300_151, \15211 );
and \U$13785 ( \15403 , RI2b5e774f6318_164, \15213 );
and \U$13786 ( \15404 , RI2b5e774ea900_177, \15215 );
and \U$13787 ( \15405 , RI2b5e774de0d8_190, \15217 );
and \U$13788 ( \15406 , RI2b5e774d50f0_203, \15219 );
and \U$13789 ( \15407 , RI2b5e785f4030_216, \15221 );
and \U$13790 ( \15408 , RI2b5e785eb408_229, \15223 );
and \U$13791 ( \15409 , RI2b5e785da590_242, \15225 );
or \U$13792 ( \15410 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 );
_DC r14ea ( \15411_nR14ea , \15410 , \15235 );
buf \U$13793 ( \15412 , \15411_nR14ea );
and \U$13794 ( \15413 , \15392 , \15412 );
xor \U$13795 ( \15414 , \15172 , \15180 );
buf \U$13796 ( \15415 , \15414 );
buf \U$13797 ( \15416 , \15415 );
not \U$13798 ( \15417 , \15416 );
and \U$13799 ( \15418 , RI2b5e78549810_35, \15193 );
and \U$13800 ( \15419 , RI2b5e78538b78_48, \15195 );
and \U$13801 ( \15420 , RI2b5e78538560_61, \15197 );
and \U$13802 ( \15421 , RI2b5e784a5fe8_74, \15199 );
and \U$13803 ( \15422 , RI2b5e78495350_87, \15201 );
and \U$13804 ( \15423 , RI2b5e78403e50_100, \15203 );
and \U$13805 ( \15424 , RI2b5e775b2130_113, \15205 );
and \U$13806 ( \15425 , RI2b5e775b1b18_126, \15207 );
and \U$13807 ( \15426 , RI2b5e7750bab0_139, \15209 );
and \U$13808 ( \15427 , RI2b5e774ff288_152, \15211 );
and \U$13809 ( \15428 , RI2b5e774f62a0_165, \15213 );
and \U$13810 ( \15429 , RI2b5e774ea888_178, \15215 );
and \U$13811 ( \15430 , RI2b5e774de060_191, \15217 );
and \U$13812 ( \15431 , RI2b5e774d5078_204, \15219 );
and \U$13813 ( \15432 , RI2b5e785f3fb8_217, \15221 );
and \U$13814 ( \15433 , RI2b5e785eb390_230, \15223 );
and \U$13815 ( \15434 , RI2b5e785da518_243, \15225 );
or \U$13816 ( \15435 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 );
_DC r1503 ( \15436_nR1503 , \15435 , \15235 );
buf \U$13817 ( \15437 , \15436_nR1503 );
and \U$13818 ( \15438 , \15417 , \15437 );
xor \U$13819 ( \15439 , \15173 , \15179 );
buf \U$13820 ( \15440 , \15439 );
buf \U$13821 ( \15441 , \15440 );
not \U$13822 ( \15442 , \15441 );
and \U$13823 ( \15443 , RI2b5e78549798_36, \15193 );
and \U$13824 ( \15444 , RI2b5e78538b00_49, \15195 );
and \U$13825 ( \15445 , RI2b5e785384e8_62, \15197 );
and \U$13826 ( \15446 , RI2b5e784a5f70_75, \15199 );
and \U$13827 ( \15447 , RI2b5e784952d8_88, \15201 );
and \U$13828 ( \15448 , RI2b5e78403dd8_101, \15203 );
and \U$13829 ( \15449 , RI2b5e775b20b8_114, \15205 );
and \U$13830 ( \15450 , RI2b5e775b1aa0_127, \15207 );
and \U$13831 ( \15451 , RI2b5e7750ba38_140, \15209 );
and \U$13832 ( \15452 , RI2b5e774ff210_153, \15211 );
and \U$13833 ( \15453 , RI2b5e774f6228_166, \15213 );
and \U$13834 ( \15454 , RI2b5e774ea810_179, \15215 );
and \U$13835 ( \15455 , RI2b5e774ddfe8_192, \15217 );
and \U$13836 ( \15456 , RI2b5e774d5000_205, \15219 );
and \U$13837 ( \15457 , RI2b5e785f3f40_218, \15221 );
and \U$13838 ( \15458 , RI2b5e785eb318_231, \15223 );
and \U$13839 ( \15459 , RI2b5e785da4a0_244, \15225 );
or \U$13840 ( \15460 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 );
_DC r151c ( \15461_nR151c , \15460 , \15235 );
buf \U$13841 ( \15462 , \15461_nR151c );
and \U$13842 ( \15463 , \15442 , \15462 );
xor \U$13843 ( \15464 , \15174 , \15178 );
buf \U$13844 ( \15465 , \15464 );
buf \U$13845 ( \15466 , \15465 );
not \U$13846 ( \15467 , \15466 );
and \U$13847 ( \15468 , RI2b5e78549720_37, \15193 );
and \U$13848 ( \15469 , RI2b5e78538a88_50, \15195 );
and \U$13849 ( \15470 , RI2b5e78538470_63, \15197 );
and \U$13850 ( \15471 , RI2b5e784a5ef8_76, \15199 );
and \U$13851 ( \15472 , RI2b5e78495260_89, \15201 );
and \U$13852 ( \15473 , RI2b5e78403d60_102, \15203 );
and \U$13853 ( \15474 , RI2b5e775b2040_115, \15205 );
and \U$13854 ( \15475 , RI2b5e775b1a28_128, \15207 );
and \U$13855 ( \15476 , RI2b5e7750b9c0_141, \15209 );
and \U$13856 ( \15477 , RI2b5e774ff198_154, \15211 );
and \U$13857 ( \15478 , RI2b5e774f61b0_167, \15213 );
and \U$13858 ( \15479 , RI2b5e774ea798_180, \15215 );
and \U$13859 ( \15480 , RI2b5e774ddf70_193, \15217 );
and \U$13860 ( \15481 , RI2b5e774d4f88_206, \15219 );
and \U$13861 ( \15482 , RI2b5e785f3ec8_219, \15221 );
and \U$13862 ( \15483 , RI2b5e785eb2a0_232, \15223 );
and \U$13863 ( \15484 , RI2b5e785da428_245, \15225 );
or \U$13864 ( \15485 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 );
_DC r1535 ( \15486_nR1535 , \15485 , \15235 );
buf \U$13865 ( \15487 , \15486_nR1535 );
and \U$13866 ( \15488 , \15467 , \15487 );
xor \U$13867 ( \15489 , \15175 , \15177 );
buf \U$13868 ( \15490 , \15489 );
buf \U$13869 ( \15491 , \15490 );
not \U$13870 ( \15492 , \15491 );
and \U$13871 ( \15493 , RI2b5e785496a8_38, \15193 );
and \U$13872 ( \15494 , RI2b5e78538a10_51, \15195 );
and \U$13873 ( \15495 , RI2b5e785383f8_64, \15197 );
and \U$13874 ( \15496 , RI2b5e784a5e80_77, \15199 );
and \U$13875 ( \15497 , RI2b5e784951e8_90, \15201 );
and \U$13876 ( \15498 , RI2b5e78403ce8_103, \15203 );
and \U$13877 ( \15499 , RI2b5e775b1fc8_116, \15205 );
and \U$13878 ( \15500 , RI2b5e775b19b0_129, \15207 );
and \U$13879 ( \15501 , RI2b5e7750b948_142, \15209 );
and \U$13880 ( \15502 , RI2b5e774ff120_155, \15211 );
and \U$13881 ( \15503 , RI2b5e774f6138_168, \15213 );
and \U$13882 ( \15504 , RI2b5e774ea720_181, \15215 );
and \U$13883 ( \15505 , RI2b5e774ddef8_194, \15217 );
and \U$13884 ( \15506 , RI2b5e774d4f10_207, \15219 );
and \U$13885 ( \15507 , RI2b5e785f3e50_220, \15221 );
and \U$13886 ( \15508 , RI2b5e785eb228_233, \15223 );
and \U$13887 ( \15509 , RI2b5e785da3b0_246, \15225 );
or \U$13888 ( \15510 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 );
_DC r154e ( \15511_nR154e , \15510 , \15235 );
buf \U$13889 ( \15512 , \15511_nR154e );
and \U$13890 ( \15513 , \15492 , \15512 );
buf \U$13891 ( \15514 , RI2b5e785dab30_26);
buf \U$13894 ( \15515 , \15514 );
not \U$13895 ( \15516 , \15515 );
and \U$13896 ( \15517 , RI2b5e78549630_39, \15193 );
and \U$13897 ( \15518 , RI2b5e78538998_52, \15195 );
and \U$13898 ( \15519 , RI2b5e78538380_65, \15197 );
and \U$13899 ( \15520 , RI2b5e784a5e08_78, \15199 );
and \U$13900 ( \15521 , RI2b5e78495170_91, \15201 );
and \U$13901 ( \15522 , RI2b5e78403c70_104, \15203 );
and \U$13902 ( \15523 , RI2b5e775b1f50_117, \15205 );
and \U$13903 ( \15524 , RI2b5e775b1938_130, \15207 );
and \U$13904 ( \15525 , RI2b5e7750b8d0_143, \15209 );
and \U$13905 ( \15526 , RI2b5e774ff0a8_156, \15211 );
and \U$13906 ( \15527 , RI2b5e774f60c0_169, \15213 );
and \U$13907 ( \15528 , RI2b5e774ea6a8_182, \15215 );
and \U$13908 ( \15529 , RI2b5e774dde80_195, \15217 );
and \U$13909 ( \15530 , RI2b5e774d4e98_208, \15219 );
and \U$13910 ( \15531 , RI2b5e785f3dd8_221, \15221 );
and \U$13911 ( \15532 , RI2b5e785eb1b0_234, \15223 );
and \U$13912 ( \15533 , RI2b5e785da338_247, \15225 );
or \U$13913 ( \15534 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 );
_DC r1568 ( \15535_nR1568 , \15534 , \15235 );
buf \U$13914 ( \15536 , \15535_nR1568 );
and \U$13915 ( \15537 , \15516 , \15536 );
xnor \U$13916 ( \15538 , \15491 , \15512 );
and \U$13917 ( \15539 , \15537 , \15538 );
or \U$13918 ( \15540 , \15513 , \15539 );
xnor \U$13919 ( \15541 , \15466 , \15487 );
and \U$13920 ( \15542 , \15540 , \15541 );
or \U$13921 ( \15543 , \15488 , \15542 );
xnor \U$13922 ( \15544 , \15441 , \15462 );
and \U$13923 ( \15545 , \15543 , \15544 );
or \U$13924 ( \15546 , \15463 , \15545 );
xnor \U$13925 ( \15547 , \15416 , \15437 );
and \U$13926 ( \15548 , \15546 , \15547 );
or \U$13927 ( \15549 , \15438 , \15548 );
xnor \U$13928 ( \15550 , \15391 , \15412 );
and \U$13929 ( \15551 , \15549 , \15550 );
or \U$13930 ( \15552 , \15413 , \15551 );
xnor \U$13931 ( \15553 , \15366 , \15387 );
and \U$13932 ( \15554 , \15552 , \15553 );
or \U$13933 ( \15555 , \15388 , \15554 );
xnor \U$13934 ( \15556 , \15341 , \15362 );
and \U$13935 ( \15557 , \15555 , \15556 );
or \U$13936 ( \15558 , \15363 , \15557 );
xnor \U$13937 ( \15559 , \15316 , \15337 );
and \U$13938 ( \15560 , \15558 , \15559 );
or \U$13939 ( \15561 , \15338 , \15560 );
xnor \U$13940 ( \15562 , \15291 , \15312 );
and \U$13941 ( \15563 , \15561 , \15562 );
or \U$13942 ( \15564 , \15313 , \15563 );
xnor \U$13943 ( \15565 , \15266 , \15287 );
and \U$13944 ( \15566 , \15564 , \15565 );
or \U$13945 ( \15567 , \15288 , \15566 );
xnor \U$13946 ( \15568 , \15241 , \15262 );
and \U$13947 ( \15569 , \15567 , \15568 );
or \U$13948 ( \15570 , \15263 , \15569 );
xnor \U$13949 ( \15571 , \15191 , \15237 );
and \U$13950 ( \15572 , \15570 , \15571 );
or \U$13951 ( \15573 , \15238 , \15572 );
not \U$13952 ( \15574 , \15573 );
buf \U$13953 ( \15575 , \15574 );
buf \U$13954 ( \15576 , RI2b5e785ae580_609);
buf \U$13955 ( \15577 , RI2b5e785ae5f8_608);
buf \U$13956 ( \15578 , RI2b5e785ae670_607);
buf \U$13957 ( \15579 , RI2b5e785ae6e8_606);
buf \U$13958 ( \15580 , RI2b5e785ae760_605);
buf \U$13959 ( \15581 , RI2b5e785ae7d8_604);
buf \U$13960 ( \15582 , RI2b5e785ae850_603);
buf \U$13961 ( \15583 , RI2b5e785ae8c8_602);
buf \U$13962 ( \15584 , RI2b5e785ae940_601);
buf \U$13963 ( \15585 , RI2b5e785ae3a0_613);
buf \U$13964 ( \15586 , RI2b5e785ae418_612);
buf \U$13965 ( \15587 , RI2b5e785ae490_611);
buf \U$13966 ( \15588 , RI2b5e785ae508_610);
and \U$13967 ( \15589 , \15585 , \15586 , \15587 , \15588 );
nor \U$13968 ( \15590 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15589 );
buf \U$13969 ( \15591 , \15590 );
and \U$13970 ( \15592 , \15575 , \15591 );
nor \U$13971 ( \15593 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$13972 ( \15594 , RI2b5e785daab8_27, \15593 );
and \U$13973 ( \15595 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$13974 ( \15596 , RI2b5e785495b8_40, \15595 );
and \U$13975 ( \15597 , \9672 , RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$13976 ( \15598 , RI2b5e78538920_53, \15597 );
and \U$13977 ( \15599 , RI2b5e785ae3a0_613, \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$13978 ( \15600 , RI2b5e784a63a8_66, \15599 );
and \U$13979 ( \15601 , \9672 , \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, \9667 );
and \U$13980 ( \15602 , RI2b5e78495710_79, \15601 );
and \U$13981 ( \15603 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, \9667 );
and \U$13982 ( \15604 , RI2b5e784950f8_92, \15603 );
and \U$13983 ( \15605 , \9672 , RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, \9667 );
and \U$13984 ( \15606 , RI2b5e78403bf8_105, \15605 );
and \U$13985 ( \15607 , RI2b5e785ae3a0_613, \9675 , \9680 , RI2b5e785ae508_610, \9667 );
and \U$13986 ( \15608 , RI2b5e775b1ed8_118, \15607 );
and \U$13987 ( \15609 , \9672 , \9675 , \9680 , RI2b5e785ae508_610, \9667 );
and \U$13988 ( \15610 , RI2b5e775b18c0_131, \15609 );
nor \U$13989 ( \15611 , \9672 , \9675 , \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$13990 ( \15612 , RI2b5e7750b858_144, \15611 );
nor \U$13991 ( \15613 , RI2b5e785ae3a0_613, \9675 , \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$13992 ( \15614 , RI2b5e774ff030_157, \15613 );
nor \U$13993 ( \15615 , \9672 , RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$13994 ( \15616 , RI2b5e774f6048_170, \15615 );
nor \U$13995 ( \15617 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, \9680 , RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$13996 ( \15618 , RI2b5e774ea630_183, \15617 );
nor \U$13997 ( \15619 , \9672 , \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$13998 ( \15620 , RI2b5e774dde08_196, \15619 );
nor \U$13999 ( \15621 , RI2b5e785ae3a0_613, \9675 , RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$14000 ( \15622 , RI2b5e774d4e20_209, \15621 );
nor \U$14001 ( \15623 , \9672 , RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$14002 ( \15624 , RI2b5e785f3d60_222, \15623 );
nor \U$14003 ( \15625 , RI2b5e785ae3a0_613, RI2b5e785ae418_612, RI2b5e785ae490_611, RI2b5e785ae508_610, RI2b5e785ae580_609);
and \U$14004 ( \15626 , RI2b5e785eb138_235, \15625 );
or \U$14005 ( \15627 , \15594 , \15596 , \15598 , \15600 , \15602 , \15604 , \15606 , \15608 , \15610 , \15612 , \15614 , \15616 , \15618 , \15620 , \15622 , \15624 , \15626 );
buf \U$14006 ( \15628 , RI2b5e785ae580_609);
buf \U$14007 ( \15629 , RI2b5e785ae3a0_613);
buf \U$14008 ( \15630 , RI2b5e785ae418_612);
buf \U$14009 ( \15631 , RI2b5e785ae490_611);
buf \U$14010 ( \15632 , RI2b5e785ae508_610);
or \U$14011 ( \15633 , \15629 , \15630 , \15631 , \15632 );
and \U$14012 ( \15634 , \15628 , \15633 );
buf \U$14013 ( \15635 , \15634 );
_DC r15d1 ( \15636_nR15d1 , \15627 , \15635 );
buf \U$14014 ( \15637 , \15636_nR15d1 );
not \U$14015 ( \15638 , \15637 );
nor \U$14016 ( \15639 , \12412 , \12416 , \12420 , \12424 , \12429 );
and \U$14017 ( \15640 , RI2b5e785daab8_27, \15639 );
and \U$14018 ( \15641 , \12412 , \12416 , \12420 , \12424 , \12429 );
and \U$14019 ( \15642 , RI2b5e785495b8_40, \15641 );
and \U$14020 ( \15643 , \12434 , \12416 , \12420 , \12424 , \12429 );
and \U$14021 ( \15644 , RI2b5e78538920_53, \15643 );
and \U$14022 ( \15645 , \12412 , \12437 , \12420 , \12424 , \12429 );
and \U$14023 ( \15646 , RI2b5e784a63a8_66, \15645 );
and \U$14024 ( \15647 , \12434 , \12437 , \12420 , \12424 , \12429 );
and \U$14025 ( \15648 , RI2b5e78495710_79, \15647 );
and \U$14026 ( \15649 , \12412 , \12416 , \12442 , \12424 , \12429 );
and \U$14027 ( \15650 , RI2b5e784950f8_92, \15649 );
and \U$14028 ( \15651 , \12434 , \12416 , \12442 , \12424 , \12429 );
and \U$14029 ( \15652 , RI2b5e78403bf8_105, \15651 );
and \U$14030 ( \15653 , \12412 , \12437 , \12442 , \12424 , \12429 );
and \U$14031 ( \15654 , RI2b5e775b1ed8_118, \15653 );
and \U$14032 ( \15655 , \12434 , \12437 , \12442 , \12424 , \12429 );
and \U$14033 ( \15656 , RI2b5e775b18c0_131, \15655 );
nor \U$14034 ( \15657 , \12434 , \12437 , \12442 , \12424 , \12428 );
and \U$14035 ( \15658 , RI2b5e7750b858_144, \15657 );
nor \U$14036 ( \15659 , \12412 , \12437 , \12442 , \12424 , \12428 );
and \U$14037 ( \15660 , RI2b5e774ff030_157, \15659 );
nor \U$14038 ( \15661 , \12434 , \12416 , \12442 , \12424 , \12428 );
and \U$14039 ( \15662 , RI2b5e774f6048_170, \15661 );
nor \U$14040 ( \15663 , \12412 , \12416 , \12442 , \12424 , \12428 );
and \U$14041 ( \15664 , RI2b5e774ea630_183, \15663 );
nor \U$14042 ( \15665 , \12434 , \12437 , \12420 , \12424 , \12428 );
and \U$14043 ( \15666 , RI2b5e774dde08_196, \15665 );
nor \U$14044 ( \15667 , \12412 , \12437 , \12420 , \12424 , \12428 );
and \U$14045 ( \15668 , RI2b5e774d4e20_209, \15667 );
nor \U$14046 ( \15669 , \12434 , \12416 , \12420 , \12424 , \12428 );
and \U$14047 ( \15670 , RI2b5e785f3d60_222, \15669 );
nor \U$14048 ( \15671 , \12412 , \12416 , \12420 , \12424 , \12428 );
and \U$14049 ( \15672 , RI2b5e785eb138_235, \15671 );
or \U$14050 ( \15673 , \15640 , \15642 , \15644 , \15646 , \15648 , \15650 , \15652 , \15654 , \15656 , \15658 , \15660 , \15662 , \15664 , \15666 , \15668 , \15670 , \15672 );
buf \U$14051 ( \15674 , \12428 );
buf \U$14052 ( \15675 , \12412 );
buf \U$14053 ( \15676 , \12416 );
buf \U$14054 ( \15677 , \12420 );
buf \U$14055 ( \15678 , \12424 );
or \U$14056 ( \15679 , \15675 , \15676 , \15677 , \15678 );
and \U$14057 ( \15680 , \15674 , \15679 );
buf \U$14058 ( \15681 , \15680 );
_DC r15ff ( \15682_nR15ff , \15673 , \15681 );
buf \U$14059 ( \15683 , \15682_nR15ff );
and \U$14060 ( \15684 , \15638 , \15683 );
and \U$14061 ( \15685 , RI2b5e785daa40_28, \15593 );
and \U$14062 ( \15686 , RI2b5e78549540_41, \15595 );
and \U$14063 ( \15687 , RI2b5e785388a8_54, \15597 );
and \U$14064 ( \15688 , RI2b5e784a6330_67, \15599 );
and \U$14065 ( \15689 , RI2b5e78495698_80, \15601 );
and \U$14066 ( \15690 , RI2b5e78495080_93, \15603 );
and \U$14067 ( \15691 , RI2b5e78403b80_106, \15605 );
and \U$14068 ( \15692 , RI2b5e775b1e60_119, \15607 );
and \U$14069 ( \15693 , RI2b5e7750bdf8_132, \15609 );
and \U$14070 ( \15694 , RI2b5e774ff5d0_145, \15611 );
and \U$14071 ( \15695 , RI2b5e774f65e8_158, \15613 );
and \U$14072 ( \15696 , RI2b5e774eabd0_171, \15615 );
and \U$14073 ( \15697 , RI2b5e774de3a8_184, \15617 );
and \U$14074 ( \15698 , RI2b5e774d53c0_197, \15619 );
and \U$14075 ( \15699 , RI2b5e785f4300_210, \15621 );
and \U$14076 ( \15700 , RI2b5e785f3ce8_223, \15623 );
and \U$14077 ( \15701 , RI2b5e785eb0c0_236, \15625 );
or \U$14078 ( \15702 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 );
_DC r1614 ( \15703_nR1614 , \15702 , \15635 );
buf \U$14079 ( \15704 , \15703_nR1614 );
not \U$14080 ( \15705 , \15704 );
and \U$14081 ( \15706 , RI2b5e785daa40_28, \15639 );
and \U$14082 ( \15707 , RI2b5e78549540_41, \15641 );
and \U$14083 ( \15708 , RI2b5e785388a8_54, \15643 );
and \U$14084 ( \15709 , RI2b5e784a6330_67, \15645 );
and \U$14085 ( \15710 , RI2b5e78495698_80, \15647 );
and \U$14086 ( \15711 , RI2b5e78495080_93, \15649 );
and \U$14087 ( \15712 , RI2b5e78403b80_106, \15651 );
and \U$14088 ( \15713 , RI2b5e775b1e60_119, \15653 );
and \U$14089 ( \15714 , RI2b5e7750bdf8_132, \15655 );
and \U$14090 ( \15715 , RI2b5e774ff5d0_145, \15657 );
and \U$14091 ( \15716 , RI2b5e774f65e8_158, \15659 );
and \U$14092 ( \15717 , RI2b5e774eabd0_171, \15661 );
and \U$14093 ( \15718 , RI2b5e774de3a8_184, \15663 );
and \U$14094 ( \15719 , RI2b5e774d53c0_197, \15665 );
and \U$14095 ( \15720 , RI2b5e785f4300_210, \15667 );
and \U$14096 ( \15721 , RI2b5e785f3ce8_223, \15669 );
and \U$14097 ( \15722 , RI2b5e785eb0c0_236, \15671 );
or \U$14098 ( \15723 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 );
_DC r1629 ( \15724_nR1629 , \15723 , \15681 );
buf \U$14099 ( \15725 , \15724_nR1629 );
and \U$14100 ( \15726 , \15705 , \15725 );
and \U$14101 ( \15727 , RI2b5e785da9c8_29, \15593 );
and \U$14102 ( \15728 , RI2b5e785494c8_42, \15595 );
and \U$14103 ( \15729 , RI2b5e78538830_55, \15597 );
and \U$14104 ( \15730 , RI2b5e784a62b8_68, \15599 );
and \U$14105 ( \15731 , RI2b5e78495620_81, \15601 );
and \U$14106 ( \15732 , RI2b5e78495008_94, \15603 );
and \U$14107 ( \15733 , RI2b5e78403b08_107, \15605 );
and \U$14108 ( \15734 , RI2b5e775b1de8_120, \15607 );
and \U$14109 ( \15735 , RI2b5e7750bd80_133, \15609 );
and \U$14110 ( \15736 , RI2b5e774ff558_146, \15611 );
and \U$14111 ( \15737 , RI2b5e774f6570_159, \15613 );
and \U$14112 ( \15738 , RI2b5e774eab58_172, \15615 );
and \U$14113 ( \15739 , RI2b5e774de330_185, \15617 );
and \U$14114 ( \15740 , RI2b5e774d5348_198, \15619 );
and \U$14115 ( \15741 , RI2b5e785f4288_211, \15621 );
and \U$14116 ( \15742 , RI2b5e785f3658_224, \15623 );
and \U$14117 ( \15743 , RI2b5e785eb048_237, \15625 );
or \U$14118 ( \15744 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 );
_DC r163e ( \15745_nR163e , \15744 , \15635 );
buf \U$14119 ( \15746 , \15745_nR163e );
not \U$14120 ( \15747 , \15746 );
and \U$14121 ( \15748 , RI2b5e785da9c8_29, \15639 );
and \U$14122 ( \15749 , RI2b5e785494c8_42, \15641 );
and \U$14123 ( \15750 , RI2b5e78538830_55, \15643 );
and \U$14124 ( \15751 , RI2b5e784a62b8_68, \15645 );
and \U$14125 ( \15752 , RI2b5e78495620_81, \15647 );
and \U$14126 ( \15753 , RI2b5e78495008_94, \15649 );
and \U$14127 ( \15754 , RI2b5e78403b08_107, \15651 );
and \U$14128 ( \15755 , RI2b5e775b1de8_120, \15653 );
and \U$14129 ( \15756 , RI2b5e7750bd80_133, \15655 );
and \U$14130 ( \15757 , RI2b5e774ff558_146, \15657 );
and \U$14131 ( \15758 , RI2b5e774f6570_159, \15659 );
and \U$14132 ( \15759 , RI2b5e774eab58_172, \15661 );
and \U$14133 ( \15760 , RI2b5e774de330_185, \15663 );
and \U$14134 ( \15761 , RI2b5e774d5348_198, \15665 );
and \U$14135 ( \15762 , RI2b5e785f4288_211, \15667 );
and \U$14136 ( \15763 , RI2b5e785f3658_224, \15669 );
and \U$14137 ( \15764 , RI2b5e785eb048_237, \15671 );
or \U$14138 ( \15765 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 );
_DC r1653 ( \15766_nR1653 , \15765 , \15681 );
buf \U$14139 ( \15767 , \15766_nR1653 );
and \U$14140 ( \15768 , \15747 , \15767 );
and \U$14141 ( \15769 , RI2b5e785da950_30, \15593 );
and \U$14142 ( \15770 , RI2b5e78549450_43, \15595 );
and \U$14143 ( \15771 , RI2b5e785387b8_56, \15597 );
and \U$14144 ( \15772 , RI2b5e784a6240_69, \15599 );
and \U$14145 ( \15773 , RI2b5e784955a8_82, \15601 );
and \U$14146 ( \15774 , RI2b5e78494f90_95, \15603 );
and \U$14147 ( \15775 , RI2b5e78403a90_108, \15605 );
and \U$14148 ( \15776 , RI2b5e775b1d70_121, \15607 );
and \U$14149 ( \15777 , RI2b5e7750bd08_134, \15609 );
and \U$14150 ( \15778 , RI2b5e774ff4e0_147, \15611 );
and \U$14151 ( \15779 , RI2b5e774f64f8_160, \15613 );
and \U$14152 ( \15780 , RI2b5e774eaae0_173, \15615 );
and \U$14153 ( \15781 , RI2b5e774de2b8_186, \15617 );
and \U$14154 ( \15782 , RI2b5e774d52d0_199, \15619 );
and \U$14155 ( \15783 , RI2b5e785f4210_212, \15621 );
and \U$14156 ( \15784 , RI2b5e785eb5e8_225, \15623 );
and \U$14157 ( \15785 , RI2b5e785e6c50_238, \15625 );
or \U$14158 ( \15786 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 );
_DC r1668 ( \15787_nR1668 , \15786 , \15635 );
buf \U$14159 ( \15788 , \15787_nR1668 );
not \U$14160 ( \15789 , \15788 );
and \U$14161 ( \15790 , RI2b5e785da950_30, \15639 );
and \U$14162 ( \15791 , RI2b5e78549450_43, \15641 );
and \U$14163 ( \15792 , RI2b5e785387b8_56, \15643 );
and \U$14164 ( \15793 , RI2b5e784a6240_69, \15645 );
and \U$14165 ( \15794 , RI2b5e784955a8_82, \15647 );
and \U$14166 ( \15795 , RI2b5e78494f90_95, \15649 );
and \U$14167 ( \15796 , RI2b5e78403a90_108, \15651 );
and \U$14168 ( \15797 , RI2b5e775b1d70_121, \15653 );
and \U$14169 ( \15798 , RI2b5e7750bd08_134, \15655 );
and \U$14170 ( \15799 , RI2b5e774ff4e0_147, \15657 );
and \U$14171 ( \15800 , RI2b5e774f64f8_160, \15659 );
and \U$14172 ( \15801 , RI2b5e774eaae0_173, \15661 );
and \U$14173 ( \15802 , RI2b5e774de2b8_186, \15663 );
and \U$14174 ( \15803 , RI2b5e774d52d0_199, \15665 );
and \U$14175 ( \15804 , RI2b5e785f4210_212, \15667 );
and \U$14176 ( \15805 , RI2b5e785eb5e8_225, \15669 );
and \U$14177 ( \15806 , RI2b5e785e6c50_238, \15671 );
or \U$14178 ( \15807 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 );
_DC r167d ( \15808_nR167d , \15807 , \15681 );
buf \U$14179 ( \15809 , \15808_nR167d );
and \U$14180 ( \15810 , \15789 , \15809 );
and \U$14181 ( \15811 , RI2b5e785da8d8_31, \15593 );
and \U$14182 ( \15812 , RI2b5e785493d8_44, \15595 );
and \U$14183 ( \15813 , RI2b5e78538740_57, \15597 );
and \U$14184 ( \15814 , RI2b5e784a61c8_70, \15599 );
and \U$14185 ( \15815 , RI2b5e78495530_83, \15601 );
and \U$14186 ( \15816 , RI2b5e78494f18_96, \15603 );
and \U$14187 ( \15817 , RI2b5e78403a18_109, \15605 );
and \U$14188 ( \15818 , RI2b5e775b1cf8_122, \15607 );
and \U$14189 ( \15819 , RI2b5e7750bc90_135, \15609 );
and \U$14190 ( \15820 , RI2b5e774ff468_148, \15611 );
and \U$14191 ( \15821 , RI2b5e774f6480_161, \15613 );
and \U$14192 ( \15822 , RI2b5e774eaa68_174, \15615 );
and \U$14193 ( \15823 , RI2b5e774de240_187, \15617 );
and \U$14194 ( \15824 , RI2b5e774d5258_200, \15619 );
and \U$14195 ( \15825 , RI2b5e785f4198_213, \15621 );
and \U$14196 ( \15826 , RI2b5e785eb570_226, \15623 );
and \U$14197 ( \15827 , RI2b5e785e6bd8_239, \15625 );
or \U$14198 ( \15828 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 );
_DC r1692 ( \15829_nR1692 , \15828 , \15635 );
buf \U$14199 ( \15830 , \15829_nR1692 );
not \U$14200 ( \15831 , \15830 );
and \U$14201 ( \15832 , RI2b5e785da8d8_31, \15639 );
and \U$14202 ( \15833 , RI2b5e785493d8_44, \15641 );
and \U$14203 ( \15834 , RI2b5e78538740_57, \15643 );
and \U$14204 ( \15835 , RI2b5e784a61c8_70, \15645 );
and \U$14205 ( \15836 , RI2b5e78495530_83, \15647 );
and \U$14206 ( \15837 , RI2b5e78494f18_96, \15649 );
and \U$14207 ( \15838 , RI2b5e78403a18_109, \15651 );
and \U$14208 ( \15839 , RI2b5e775b1cf8_122, \15653 );
and \U$14209 ( \15840 , RI2b5e7750bc90_135, \15655 );
and \U$14210 ( \15841 , RI2b5e774ff468_148, \15657 );
and \U$14211 ( \15842 , RI2b5e774f6480_161, \15659 );
and \U$14212 ( \15843 , RI2b5e774eaa68_174, \15661 );
and \U$14213 ( \15844 , RI2b5e774de240_187, \15663 );
and \U$14214 ( \15845 , RI2b5e774d5258_200, \15665 );
and \U$14215 ( \15846 , RI2b5e785f4198_213, \15667 );
and \U$14216 ( \15847 , RI2b5e785eb570_226, \15669 );
and \U$14217 ( \15848 , RI2b5e785e6bd8_239, \15671 );
or \U$14218 ( \15849 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 );
_DC r16a7 ( \15850_nR16a7 , \15849 , \15681 );
buf \U$14219 ( \15851 , \15850_nR16a7 );
and \U$14220 ( \15852 , \15831 , \15851 );
and \U$14221 ( \15853 , RI2b5e785da860_32, \15593 );
and \U$14222 ( \15854 , RI2b5e78549360_45, \15595 );
and \U$14223 ( \15855 , RI2b5e785386c8_58, \15597 );
and \U$14224 ( \15856 , RI2b5e784a6150_71, \15599 );
and \U$14225 ( \15857 , RI2b5e784954b8_84, \15601 );
and \U$14226 ( \15858 , RI2b5e78494ea0_97, \15603 );
and \U$14227 ( \15859 , RI2b5e784039a0_110, \15605 );
and \U$14228 ( \15860 , RI2b5e775b1c80_123, \15607 );
and \U$14229 ( \15861 , RI2b5e7750bc18_136, \15609 );
and \U$14230 ( \15862 , RI2b5e774ff3f0_149, \15611 );
and \U$14231 ( \15863 , RI2b5e774f6408_162, \15613 );
and \U$14232 ( \15864 , RI2b5e774ea9f0_175, \15615 );
and \U$14233 ( \15865 , RI2b5e774de1c8_188, \15617 );
and \U$14234 ( \15866 , RI2b5e774d51e0_201, \15619 );
and \U$14235 ( \15867 , RI2b5e785f4120_214, \15621 );
and \U$14236 ( \15868 , RI2b5e785eb4f8_227, \15623 );
and \U$14237 ( \15869 , RI2b5e785e64d0_240, \15625 );
or \U$14238 ( \15870 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 );
_DC r16bc ( \15871_nR16bc , \15870 , \15635 );
buf \U$14239 ( \15872 , \15871_nR16bc );
not \U$14240 ( \15873 , \15872 );
and \U$14241 ( \15874 , RI2b5e785da860_32, \15639 );
and \U$14242 ( \15875 , RI2b5e78549360_45, \15641 );
and \U$14243 ( \15876 , RI2b5e785386c8_58, \15643 );
and \U$14244 ( \15877 , RI2b5e784a6150_71, \15645 );
and \U$14245 ( \15878 , RI2b5e784954b8_84, \15647 );
and \U$14246 ( \15879 , RI2b5e78494ea0_97, \15649 );
and \U$14247 ( \15880 , RI2b5e784039a0_110, \15651 );
and \U$14248 ( \15881 , RI2b5e775b1c80_123, \15653 );
and \U$14249 ( \15882 , RI2b5e7750bc18_136, \15655 );
and \U$14250 ( \15883 , RI2b5e774ff3f0_149, \15657 );
and \U$14251 ( \15884 , RI2b5e774f6408_162, \15659 );
and \U$14252 ( \15885 , RI2b5e774ea9f0_175, \15661 );
and \U$14253 ( \15886 , RI2b5e774de1c8_188, \15663 );
and \U$14254 ( \15887 , RI2b5e774d51e0_201, \15665 );
and \U$14255 ( \15888 , RI2b5e785f4120_214, \15667 );
and \U$14256 ( \15889 , RI2b5e785eb4f8_227, \15669 );
and \U$14257 ( \15890 , RI2b5e785e64d0_240, \15671 );
or \U$14258 ( \15891 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 );
_DC r16d1 ( \15892_nR16d1 , \15891 , \15681 );
buf \U$14259 ( \15893 , \15892_nR16d1 );
and \U$14260 ( \15894 , \15873 , \15893 );
and \U$14261 ( \15895 , RI2b5e78549900_33, \15593 );
and \U$14262 ( \15896 , RI2b5e78538c68_46, \15595 );
and \U$14263 ( \15897 , RI2b5e78538650_59, \15597 );
and \U$14264 ( \15898 , RI2b5e784a60d8_72, \15599 );
and \U$14265 ( \15899 , RI2b5e78495440_85, \15601 );
and \U$14266 ( \15900 , RI2b5e78494e28_98, \15603 );
and \U$14267 ( \15901 , RI2b5e78403928_111, \15605 );
and \U$14268 ( \15902 , RI2b5e775b1c08_124, \15607 );
and \U$14269 ( \15903 , RI2b5e7750bba0_137, \15609 );
and \U$14270 ( \15904 , RI2b5e774ff378_150, \15611 );
and \U$14271 ( \15905 , RI2b5e774f6390_163, \15613 );
and \U$14272 ( \15906 , RI2b5e774ea978_176, \15615 );
and \U$14273 ( \15907 , RI2b5e774de150_189, \15617 );
and \U$14274 ( \15908 , RI2b5e774d5168_202, \15619 );
and \U$14275 ( \15909 , RI2b5e785f40a8_215, \15621 );
and \U$14276 ( \15910 , RI2b5e785eb480_228, \15623 );
and \U$14277 ( \15911 , RI2b5e785da608_241, \15625 );
or \U$14278 ( \15912 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 );
_DC r16e6 ( \15913_nR16e6 , \15912 , \15635 );
buf \U$14279 ( \15914 , \15913_nR16e6 );
not \U$14280 ( \15915 , \15914 );
and \U$14281 ( \15916 , RI2b5e78549900_33, \15639 );
and \U$14282 ( \15917 , RI2b5e78538c68_46, \15641 );
and \U$14283 ( \15918 , RI2b5e78538650_59, \15643 );
and \U$14284 ( \15919 , RI2b5e784a60d8_72, \15645 );
and \U$14285 ( \15920 , RI2b5e78495440_85, \15647 );
and \U$14286 ( \15921 , RI2b5e78494e28_98, \15649 );
and \U$14287 ( \15922 , RI2b5e78403928_111, \15651 );
and \U$14288 ( \15923 , RI2b5e775b1c08_124, \15653 );
and \U$14289 ( \15924 , RI2b5e7750bba0_137, \15655 );
and \U$14290 ( \15925 , RI2b5e774ff378_150, \15657 );
and \U$14291 ( \15926 , RI2b5e774f6390_163, \15659 );
and \U$14292 ( \15927 , RI2b5e774ea978_176, \15661 );
and \U$14293 ( \15928 , RI2b5e774de150_189, \15663 );
and \U$14294 ( \15929 , RI2b5e774d5168_202, \15665 );
and \U$14295 ( \15930 , RI2b5e785f40a8_215, \15667 );
and \U$14296 ( \15931 , RI2b5e785eb480_228, \15669 );
and \U$14297 ( \15932 , RI2b5e785da608_241, \15671 );
or \U$14298 ( \15933 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 );
_DC r16fb ( \15934_nR16fb , \15933 , \15681 );
buf \U$14299 ( \15935 , \15934_nR16fb );
and \U$14300 ( \15936 , \15915 , \15935 );
and \U$14301 ( \15937 , RI2b5e78549888_34, \15593 );
and \U$14302 ( \15938 , RI2b5e78538bf0_47, \15595 );
and \U$14303 ( \15939 , RI2b5e785385d8_60, \15597 );
and \U$14304 ( \15940 , RI2b5e784a6060_73, \15599 );
and \U$14305 ( \15941 , RI2b5e784953c8_86, \15601 );
and \U$14306 ( \15942 , RI2b5e78403ec8_99, \15603 );
and \U$14307 ( \15943 , RI2b5e775b21a8_112, \15605 );
and \U$14308 ( \15944 , RI2b5e775b1b90_125, \15607 );
and \U$14309 ( \15945 , RI2b5e7750bb28_138, \15609 );
and \U$14310 ( \15946 , RI2b5e774ff300_151, \15611 );
and \U$14311 ( \15947 , RI2b5e774f6318_164, \15613 );
and \U$14312 ( \15948 , RI2b5e774ea900_177, \15615 );
and \U$14313 ( \15949 , RI2b5e774de0d8_190, \15617 );
and \U$14314 ( \15950 , RI2b5e774d50f0_203, \15619 );
and \U$14315 ( \15951 , RI2b5e785f4030_216, \15621 );
and \U$14316 ( \15952 , RI2b5e785eb408_229, \15623 );
and \U$14317 ( \15953 , RI2b5e785da590_242, \15625 );
or \U$14318 ( \15954 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 );
_DC r1710 ( \15955_nR1710 , \15954 , \15635 );
buf \U$14319 ( \15956 , \15955_nR1710 );
not \U$14320 ( \15957 , \15956 );
and \U$14321 ( \15958 , RI2b5e78549888_34, \15639 );
and \U$14322 ( \15959 , RI2b5e78538bf0_47, \15641 );
and \U$14323 ( \15960 , RI2b5e785385d8_60, \15643 );
and \U$14324 ( \15961 , RI2b5e784a6060_73, \15645 );
and \U$14325 ( \15962 , RI2b5e784953c8_86, \15647 );
and \U$14326 ( \15963 , RI2b5e78403ec8_99, \15649 );
and \U$14327 ( \15964 , RI2b5e775b21a8_112, \15651 );
and \U$14328 ( \15965 , RI2b5e775b1b90_125, \15653 );
and \U$14329 ( \15966 , RI2b5e7750bb28_138, \15655 );
and \U$14330 ( \15967 , RI2b5e774ff300_151, \15657 );
and \U$14331 ( \15968 , RI2b5e774f6318_164, \15659 );
and \U$14332 ( \15969 , RI2b5e774ea900_177, \15661 );
and \U$14333 ( \15970 , RI2b5e774de0d8_190, \15663 );
and \U$14334 ( \15971 , RI2b5e774d50f0_203, \15665 );
and \U$14335 ( \15972 , RI2b5e785f4030_216, \15667 );
and \U$14336 ( \15973 , RI2b5e785eb408_229, \15669 );
and \U$14337 ( \15974 , RI2b5e785da590_242, \15671 );
or \U$14338 ( \15975 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 );
_DC r1725 ( \15976_nR1725 , \15975 , \15681 );
buf \U$14339 ( \15977 , \15976_nR1725 );
and \U$14340 ( \15978 , \15957 , \15977 );
and \U$14341 ( \15979 , RI2b5e78549810_35, \15593 );
and \U$14342 ( \15980 , RI2b5e78538b78_48, \15595 );
and \U$14343 ( \15981 , RI2b5e78538560_61, \15597 );
and \U$14344 ( \15982 , RI2b5e784a5fe8_74, \15599 );
and \U$14345 ( \15983 , RI2b5e78495350_87, \15601 );
and \U$14346 ( \15984 , RI2b5e78403e50_100, \15603 );
and \U$14347 ( \15985 , RI2b5e775b2130_113, \15605 );
and \U$14348 ( \15986 , RI2b5e775b1b18_126, \15607 );
and \U$14349 ( \15987 , RI2b5e7750bab0_139, \15609 );
and \U$14350 ( \15988 , RI2b5e774ff288_152, \15611 );
and \U$14351 ( \15989 , RI2b5e774f62a0_165, \15613 );
and \U$14352 ( \15990 , RI2b5e774ea888_178, \15615 );
and \U$14353 ( \15991 , RI2b5e774de060_191, \15617 );
and \U$14354 ( \15992 , RI2b5e774d5078_204, \15619 );
and \U$14355 ( \15993 , RI2b5e785f3fb8_217, \15621 );
and \U$14356 ( \15994 , RI2b5e785eb390_230, \15623 );
and \U$14357 ( \15995 , RI2b5e785da518_243, \15625 );
or \U$14358 ( \15996 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 );
_DC r173a ( \15997_nR173a , \15996 , \15635 );
buf \U$14359 ( \15998 , \15997_nR173a );
not \U$14360 ( \15999 , \15998 );
and \U$14361 ( \16000 , RI2b5e78549810_35, \15639 );
and \U$14362 ( \16001 , RI2b5e78538b78_48, \15641 );
and \U$14363 ( \16002 , RI2b5e78538560_61, \15643 );
and \U$14364 ( \16003 , RI2b5e784a5fe8_74, \15645 );
and \U$14365 ( \16004 , RI2b5e78495350_87, \15647 );
and \U$14366 ( \16005 , RI2b5e78403e50_100, \15649 );
and \U$14367 ( \16006 , RI2b5e775b2130_113, \15651 );
and \U$14368 ( \16007 , RI2b5e775b1b18_126, \15653 );
and \U$14369 ( \16008 , RI2b5e7750bab0_139, \15655 );
and \U$14370 ( \16009 , RI2b5e774ff288_152, \15657 );
and \U$14371 ( \16010 , RI2b5e774f62a0_165, \15659 );
and \U$14372 ( \16011 , RI2b5e774ea888_178, \15661 );
and \U$14373 ( \16012 , RI2b5e774de060_191, \15663 );
and \U$14374 ( \16013 , RI2b5e774d5078_204, \15665 );
and \U$14375 ( \16014 , RI2b5e785f3fb8_217, \15667 );
and \U$14376 ( \16015 , RI2b5e785eb390_230, \15669 );
and \U$14377 ( \16016 , RI2b5e785da518_243, \15671 );
or \U$14378 ( \16017 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 );
_DC r174f ( \16018_nR174f , \16017 , \15681 );
buf \U$14379 ( \16019 , \16018_nR174f );
and \U$14380 ( \16020 , \15999 , \16019 );
and \U$14381 ( \16021 , RI2b5e78549798_36, \15593 );
and \U$14382 ( \16022 , RI2b5e78538b00_49, \15595 );
and \U$14383 ( \16023 , RI2b5e785384e8_62, \15597 );
and \U$14384 ( \16024 , RI2b5e784a5f70_75, \15599 );
and \U$14385 ( \16025 , RI2b5e784952d8_88, \15601 );
and \U$14386 ( \16026 , RI2b5e78403dd8_101, \15603 );
and \U$14387 ( \16027 , RI2b5e775b20b8_114, \15605 );
and \U$14388 ( \16028 , RI2b5e775b1aa0_127, \15607 );
and \U$14389 ( \16029 , RI2b5e7750ba38_140, \15609 );
and \U$14390 ( \16030 , RI2b5e774ff210_153, \15611 );
and \U$14391 ( \16031 , RI2b5e774f6228_166, \15613 );
and \U$14392 ( \16032 , RI2b5e774ea810_179, \15615 );
and \U$14393 ( \16033 , RI2b5e774ddfe8_192, \15617 );
and \U$14394 ( \16034 , RI2b5e774d5000_205, \15619 );
and \U$14395 ( \16035 , RI2b5e785f3f40_218, \15621 );
and \U$14396 ( \16036 , RI2b5e785eb318_231, \15623 );
and \U$14397 ( \16037 , RI2b5e785da4a0_244, \15625 );
or \U$14398 ( \16038 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 );
_DC r1764 ( \16039_nR1764 , \16038 , \15635 );
buf \U$14399 ( \16040 , \16039_nR1764 );
not \U$14400 ( \16041 , \16040 );
and \U$14401 ( \16042 , RI2b5e78549798_36, \15639 );
and \U$14402 ( \16043 , RI2b5e78538b00_49, \15641 );
and \U$14403 ( \16044 , RI2b5e785384e8_62, \15643 );
and \U$14404 ( \16045 , RI2b5e784a5f70_75, \15645 );
and \U$14405 ( \16046 , RI2b5e784952d8_88, \15647 );
and \U$14406 ( \16047 , RI2b5e78403dd8_101, \15649 );
and \U$14407 ( \16048 , RI2b5e775b20b8_114, \15651 );
and \U$14408 ( \16049 , RI2b5e775b1aa0_127, \15653 );
and \U$14409 ( \16050 , RI2b5e7750ba38_140, \15655 );
and \U$14410 ( \16051 , RI2b5e774ff210_153, \15657 );
and \U$14411 ( \16052 , RI2b5e774f6228_166, \15659 );
and \U$14412 ( \16053 , RI2b5e774ea810_179, \15661 );
and \U$14413 ( \16054 , RI2b5e774ddfe8_192, \15663 );
and \U$14414 ( \16055 , RI2b5e774d5000_205, \15665 );
and \U$14415 ( \16056 , RI2b5e785f3f40_218, \15667 );
and \U$14416 ( \16057 , RI2b5e785eb318_231, \15669 );
and \U$14417 ( \16058 , RI2b5e785da4a0_244, \15671 );
or \U$14418 ( \16059 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 );
_DC r1779 ( \16060_nR1779 , \16059 , \15681 );
buf \U$14419 ( \16061 , \16060_nR1779 );
and \U$14420 ( \16062 , \16041 , \16061 );
and \U$14421 ( \16063 , RI2b5e78549720_37, \15593 );
and \U$14422 ( \16064 , RI2b5e78538a88_50, \15595 );
and \U$14423 ( \16065 , RI2b5e78538470_63, \15597 );
and \U$14424 ( \16066 , RI2b5e784a5ef8_76, \15599 );
and \U$14425 ( \16067 , RI2b5e78495260_89, \15601 );
and \U$14426 ( \16068 , RI2b5e78403d60_102, \15603 );
and \U$14427 ( \16069 , RI2b5e775b2040_115, \15605 );
and \U$14428 ( \16070 , RI2b5e775b1a28_128, \15607 );
and \U$14429 ( \16071 , RI2b5e7750b9c0_141, \15609 );
and \U$14430 ( \16072 , RI2b5e774ff198_154, \15611 );
and \U$14431 ( \16073 , RI2b5e774f61b0_167, \15613 );
and \U$14432 ( \16074 , RI2b5e774ea798_180, \15615 );
and \U$14433 ( \16075 , RI2b5e774ddf70_193, \15617 );
and \U$14434 ( \16076 , RI2b5e774d4f88_206, \15619 );
and \U$14435 ( \16077 , RI2b5e785f3ec8_219, \15621 );
and \U$14436 ( \16078 , RI2b5e785eb2a0_232, \15623 );
and \U$14437 ( \16079 , RI2b5e785da428_245, \15625 );
or \U$14438 ( \16080 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 );
_DC r178e ( \16081_nR178e , \16080 , \15635 );
buf \U$14439 ( \16082 , \16081_nR178e );
not \U$14440 ( \16083 , \16082 );
and \U$14441 ( \16084 , RI2b5e78549720_37, \15639 );
and \U$14442 ( \16085 , RI2b5e78538a88_50, \15641 );
and \U$14443 ( \16086 , RI2b5e78538470_63, \15643 );
and \U$14444 ( \16087 , RI2b5e784a5ef8_76, \15645 );
and \U$14445 ( \16088 , RI2b5e78495260_89, \15647 );
and \U$14446 ( \16089 , RI2b5e78403d60_102, \15649 );
and \U$14447 ( \16090 , RI2b5e775b2040_115, \15651 );
and \U$14448 ( \16091 , RI2b5e775b1a28_128, \15653 );
and \U$14449 ( \16092 , RI2b5e7750b9c0_141, \15655 );
and \U$14450 ( \16093 , RI2b5e774ff198_154, \15657 );
and \U$14451 ( \16094 , RI2b5e774f61b0_167, \15659 );
and \U$14452 ( \16095 , RI2b5e774ea798_180, \15661 );
and \U$14453 ( \16096 , RI2b5e774ddf70_193, \15663 );
and \U$14454 ( \16097 , RI2b5e774d4f88_206, \15665 );
and \U$14455 ( \16098 , RI2b5e785f3ec8_219, \15667 );
and \U$14456 ( \16099 , RI2b5e785eb2a0_232, \15669 );
and \U$14457 ( \16100 , RI2b5e785da428_245, \15671 );
or \U$14458 ( \16101 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 );
_DC r17a3 ( \16102_nR17a3 , \16101 , \15681 );
buf \U$14459 ( \16103 , \16102_nR17a3 );
and \U$14460 ( \16104 , \16083 , \16103 );
and \U$14461 ( \16105 , RI2b5e785496a8_38, \15593 );
and \U$14462 ( \16106 , RI2b5e78538a10_51, \15595 );
and \U$14463 ( \16107 , RI2b5e785383f8_64, \15597 );
and \U$14464 ( \16108 , RI2b5e784a5e80_77, \15599 );
and \U$14465 ( \16109 , RI2b5e784951e8_90, \15601 );
and \U$14466 ( \16110 , RI2b5e78403ce8_103, \15603 );
and \U$14467 ( \16111 , RI2b5e775b1fc8_116, \15605 );
and \U$14468 ( \16112 , RI2b5e775b19b0_129, \15607 );
and \U$14469 ( \16113 , RI2b5e7750b948_142, \15609 );
and \U$14470 ( \16114 , RI2b5e774ff120_155, \15611 );
and \U$14471 ( \16115 , RI2b5e774f6138_168, \15613 );
and \U$14472 ( \16116 , RI2b5e774ea720_181, \15615 );
and \U$14473 ( \16117 , RI2b5e774ddef8_194, \15617 );
and \U$14474 ( \16118 , RI2b5e774d4f10_207, \15619 );
and \U$14475 ( \16119 , RI2b5e785f3e50_220, \15621 );
and \U$14476 ( \16120 , RI2b5e785eb228_233, \15623 );
and \U$14477 ( \16121 , RI2b5e785da3b0_246, \15625 );
or \U$14478 ( \16122 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 );
_DC r17b8 ( \16123_nR17b8 , \16122 , \15635 );
buf \U$14479 ( \16124 , \16123_nR17b8 );
not \U$14480 ( \16125 , \16124 );
and \U$14481 ( \16126 , RI2b5e785496a8_38, \15639 );
and \U$14482 ( \16127 , RI2b5e78538a10_51, \15641 );
and \U$14483 ( \16128 , RI2b5e785383f8_64, \15643 );
and \U$14484 ( \16129 , RI2b5e784a5e80_77, \15645 );
and \U$14485 ( \16130 , RI2b5e784951e8_90, \15647 );
and \U$14486 ( \16131 , RI2b5e78403ce8_103, \15649 );
and \U$14487 ( \16132 , RI2b5e775b1fc8_116, \15651 );
and \U$14488 ( \16133 , RI2b5e775b19b0_129, \15653 );
and \U$14489 ( \16134 , RI2b5e7750b948_142, \15655 );
and \U$14490 ( \16135 , RI2b5e774ff120_155, \15657 );
and \U$14491 ( \16136 , RI2b5e774f6138_168, \15659 );
and \U$14492 ( \16137 , RI2b5e774ea720_181, \15661 );
and \U$14493 ( \16138 , RI2b5e774ddef8_194, \15663 );
and \U$14494 ( \16139 , RI2b5e774d4f10_207, \15665 );
and \U$14495 ( \16140 , RI2b5e785f3e50_220, \15667 );
and \U$14496 ( \16141 , RI2b5e785eb228_233, \15669 );
and \U$14497 ( \16142 , RI2b5e785da3b0_246, \15671 );
or \U$14498 ( \16143 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 );
_DC r17cd ( \16144_nR17cd , \16143 , \15681 );
buf \U$14499 ( \16145 , \16144_nR17cd );
and \U$14500 ( \16146 , \16125 , \16145 );
and \U$14501 ( \16147 , RI2b5e78549630_39, \15593 );
and \U$14502 ( \16148 , RI2b5e78538998_52, \15595 );
and \U$14503 ( \16149 , RI2b5e78538380_65, \15597 );
and \U$14504 ( \16150 , RI2b5e784a5e08_78, \15599 );
and \U$14505 ( \16151 , RI2b5e78495170_91, \15601 );
and \U$14506 ( \16152 , RI2b5e78403c70_104, \15603 );
and \U$14507 ( \16153 , RI2b5e775b1f50_117, \15605 );
and \U$14508 ( \16154 , RI2b5e775b1938_130, \15607 );
and \U$14509 ( \16155 , RI2b5e7750b8d0_143, \15609 );
and \U$14510 ( \16156 , RI2b5e774ff0a8_156, \15611 );
and \U$14511 ( \16157 , RI2b5e774f60c0_169, \15613 );
and \U$14512 ( \16158 , RI2b5e774ea6a8_182, \15615 );
and \U$14513 ( \16159 , RI2b5e774dde80_195, \15617 );
and \U$14514 ( \16160 , RI2b5e774d4e98_208, \15619 );
and \U$14515 ( \16161 , RI2b5e785f3dd8_221, \15621 );
and \U$14516 ( \16162 , RI2b5e785eb1b0_234, \15623 );
and \U$14517 ( \16163 , RI2b5e785da338_247, \15625 );
or \U$14518 ( \16164 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 );
_DC r17e2 ( \16165_nR17e2 , \16164 , \15635 );
buf \U$14519 ( \16166 , \16165_nR17e2 );
not \U$14520 ( \16167 , \16166 );
and \U$14521 ( \16168 , RI2b5e78549630_39, \15639 );
and \U$14522 ( \16169 , RI2b5e78538998_52, \15641 );
and \U$14523 ( \16170 , RI2b5e78538380_65, \15643 );
and \U$14524 ( \16171 , RI2b5e784a5e08_78, \15645 );
and \U$14525 ( \16172 , RI2b5e78495170_91, \15647 );
and \U$14526 ( \16173 , RI2b5e78403c70_104, \15649 );
and \U$14527 ( \16174 , RI2b5e775b1f50_117, \15651 );
and \U$14528 ( \16175 , RI2b5e775b1938_130, \15653 );
and \U$14529 ( \16176 , RI2b5e7750b8d0_143, \15655 );
and \U$14530 ( \16177 , RI2b5e774ff0a8_156, \15657 );
and \U$14531 ( \16178 , RI2b5e774f60c0_169, \15659 );
and \U$14532 ( \16179 , RI2b5e774ea6a8_182, \15661 );
and \U$14533 ( \16180 , RI2b5e774dde80_195, \15663 );
and \U$14534 ( \16181 , RI2b5e774d4e98_208, \15665 );
and \U$14535 ( \16182 , RI2b5e785f3dd8_221, \15667 );
and \U$14536 ( \16183 , RI2b5e785eb1b0_234, \15669 );
and \U$14537 ( \16184 , RI2b5e785da338_247, \15671 );
or \U$14538 ( \16185 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 );
_DC r17f7 ( \16186_nR17f7 , \16185 , \15681 );
buf \U$14539 ( \16187 , \16186_nR17f7 );
and \U$14540 ( \16188 , \16167 , \16187 );
xnor \U$14541 ( \16189 , \16145 , \16124 );
and \U$14542 ( \16190 , \16188 , \16189 );
or \U$14543 ( \16191 , \16146 , \16190 );
xnor \U$14544 ( \16192 , \16103 , \16082 );
and \U$14545 ( \16193 , \16191 , \16192 );
or \U$14546 ( \16194 , \16104 , \16193 );
xnor \U$14547 ( \16195 , \16061 , \16040 );
and \U$14548 ( \16196 , \16194 , \16195 );
or \U$14549 ( \16197 , \16062 , \16196 );
xnor \U$14550 ( \16198 , \16019 , \15998 );
and \U$14551 ( \16199 , \16197 , \16198 );
or \U$14552 ( \16200 , \16020 , \16199 );
xnor \U$14553 ( \16201 , \15977 , \15956 );
and \U$14554 ( \16202 , \16200 , \16201 );
or \U$14555 ( \16203 , \15978 , \16202 );
xnor \U$14556 ( \16204 , \15935 , \15914 );
and \U$14557 ( \16205 , \16203 , \16204 );
or \U$14558 ( \16206 , \15936 , \16205 );
xnor \U$14559 ( \16207 , \15893 , \15872 );
and \U$14560 ( \16208 , \16206 , \16207 );
or \U$14561 ( \16209 , \15894 , \16208 );
xnor \U$14562 ( \16210 , \15851 , \15830 );
and \U$14563 ( \16211 , \16209 , \16210 );
or \U$14564 ( \16212 , \15852 , \16211 );
xnor \U$14565 ( \16213 , \15809 , \15788 );
and \U$14566 ( \16214 , \16212 , \16213 );
or \U$14567 ( \16215 , \15810 , \16214 );
xnor \U$14568 ( \16216 , \15767 , \15746 );
and \U$14569 ( \16217 , \16215 , \16216 );
or \U$14570 ( \16218 , \15768 , \16217 );
xnor \U$14571 ( \16219 , \15725 , \15704 );
and \U$14572 ( \16220 , \16218 , \16219 );
or \U$14573 ( \16221 , \15726 , \16220 );
xnor \U$14574 ( \16222 , \15683 , \15637 );
and \U$14575 ( \16223 , \16221 , \16222 );
or \U$14576 ( \16224 , \15684 , \16223 );
buf \U$14577 ( \16225 , \16224 );
and \U$14578 ( \16226 , \15592 , \16225 );
_HMUX r4a2b ( \16227_nR4a2b , \12369 , \15163 , \16226 );
buf \U$14579 ( \16228 , \16227_nR4a2b );
not \U$14580 ( \16229 , \11832 );
nand \U$14581 ( \16230 , \12361 , \16229 );
nor \U$14582 ( \16231 , \12179 , \11015 );
nor \U$14583 ( \16232 , \11090 , \11167 );
nand \U$14584 ( \16233 , \16231 , \16232 );
nor \U$14585 ( \16234 , \11242 , \11319 );
nor \U$14586 ( \16235 , \11395 , \11468 );
nand \U$14587 ( \16236 , \16234 , \16235 );
nor \U$14588 ( \16237 , \16233 , \16236 );
nor \U$14589 ( \16238 , \11537 , \11601 );
nor \U$14590 ( \16239 , \11661 , \11718 );
nand \U$14591 ( \16240 , \16238 , \16239 );
nor \U$14592 ( \16241 , \11756 , \11788 );
nor \U$14593 ( \16242 , \11809 , \11825 );
nand \U$14594 ( \16243 , \16241 , \16242 );
nor \U$14595 ( \16244 , \16240 , \16243 );
nand \U$14596 ( \16245 , \16237 , \16244 );
nor \U$14597 ( \16246 , \12240 , \11944 );
nor \U$14598 ( \16247 , \11989 , \12041 );
nand \U$14599 ( \16248 , \16246 , \16247 );
nor \U$14600 ( \16249 , \12096 , \12135 );
nor \U$14601 ( \16250 , \12156 , \12172 );
nand \U$14602 ( \16251 , \16249 , \16250 );
nor \U$14603 ( \16252 , \16248 , \16251 );
nor \U$14604 ( \16253 , \12260 , \12215 );
nor \U$14605 ( \16254 , \12226 , \12237 );
nand \U$14606 ( \16255 , \16253 , \16254 );
nor \U$14607 ( \16256 , \12265 , \12257 );
not \U$14608 ( \16257 , \12273 );
and \U$14609 ( \16258 , \16256 , \16257 );
or \U$14610 ( \16259 , \12257 , \12275 );
nand \U$14611 ( \16260 , \16259 , \12278 );
nor \U$14612 ( \16261 , \16258 , \16260 );
or \U$14613 ( \16262 , \16255 , \16261 );
or \U$14614 ( \16263 , \12215 , \12280 );
nand \U$14615 ( \16264 , \16263 , \12284 );
and \U$14616 ( \16265 , \16254 , \16264 );
or \U$14617 ( \16266 , \12237 , \12286 );
nand \U$14618 ( \16267 , \16266 , \12289 );
nor \U$14619 ( \16268 , \16265 , \16267 );
nand \U$14620 ( \16269 , \16262 , \16268 );
and \U$14621 ( \16270 , \16252 , \16269 );
or \U$14622 ( \16271 , \11944 , \12291 );
nand \U$14623 ( \16272 , \16271 , \12296 );
and \U$14624 ( \16273 , \16247 , \16272 );
or \U$14625 ( \16274 , \12041 , \12298 );
nand \U$14626 ( \16275 , \16274 , \12301 );
nor \U$14627 ( \16276 , \16273 , \16275 );
or \U$14628 ( \16277 , \16251 , \16276 );
or \U$14629 ( \16278 , \12135 , \12303 );
nand \U$14630 ( \16279 , \16278 , \12307 );
and \U$14631 ( \16280 , \16250 , \16279 );
or \U$14632 ( \16281 , \12172 , \12309 );
nand \U$14633 ( \16282 , \16281 , \12312 );
nor \U$14634 ( \16283 , \16280 , \16282 );
nand \U$14635 ( \16284 , \16277 , \16283 );
nor \U$14636 ( \16285 , \16270 , \16284 );
or \U$14637 ( \16286 , \16245 , \16285 );
or \U$14638 ( \16287 , \11015 , \12314 );
nand \U$14639 ( \16288 , \16287 , \12320 );
and \U$14640 ( \16289 , \16232 , \16288 );
or \U$14641 ( \16290 , \11167 , \12322 );
nand \U$14642 ( \16291 , \16290 , \12325 );
nor \U$14643 ( \16292 , \16289 , \16291 );
or \U$14644 ( \16293 , \16236 , \16292 );
or \U$14645 ( \16294 , \11319 , \12327 );
nand \U$14646 ( \16295 , \16294 , \12331 );
and \U$14647 ( \16296 , \16235 , \16295 );
or \U$14648 ( \16297 , \11468 , \12333 );
nand \U$14649 ( \16298 , \16297 , \12336 );
nor \U$14650 ( \16299 , \16296 , \16298 );
nand \U$14651 ( \16300 , \16293 , \16299 );
and \U$14652 ( \16301 , \16244 , \16300 );
or \U$14653 ( \16302 , \11601 , \12338 );
nand \U$14654 ( \16303 , \16302 , \12343 );
and \U$14655 ( \16304 , \16239 , \16303 );
or \U$14656 ( \16305 , \11718 , \12345 );
nand \U$14657 ( \16306 , \16305 , \12348 );
nor \U$14658 ( \16307 , \16304 , \16306 );
or \U$14659 ( \16308 , \16243 , \16307 );
or \U$14660 ( \16309 , \11788 , \12350 );
nand \U$14661 ( \16310 , \16309 , \12354 );
and \U$14662 ( \16311 , \16242 , \16310 );
or \U$14663 ( \16312 , \11825 , \12356 );
nand \U$14664 ( \16313 , \16312 , \12359 );
nor \U$14665 ( \16314 , \16311 , \16313 );
nand \U$14666 ( \16315 , \16308 , \16314 );
nor \U$14667 ( \16316 , \16301 , \16315 );
nand \U$14668 ( \16317 , \16286 , \16316 );
not \U$14669 ( \16318 , \16317 );
xor \U$14670 ( \16319 , \16230 , \16318 );
buf \U$14671 ( \16320 , \16319 );
not \U$14672 ( \16321 , \14626 );
nand \U$14673 ( \16322 , \15155 , \16321 );
nor \U$14674 ( \16323 , \14973 , \13809 );
nor \U$14675 ( \16324 , \13884 , \13961 );
nand \U$14676 ( \16325 , \16323 , \16324 );
nor \U$14677 ( \16326 , \14036 , \14113 );
nor \U$14678 ( \16327 , \14189 , \14262 );
nand \U$14679 ( \16328 , \16326 , \16327 );
nor \U$14680 ( \16329 , \16325 , \16328 );
nor \U$14681 ( \16330 , \14331 , \14395 );
nor \U$14682 ( \16331 , \14455 , \14512 );
nand \U$14683 ( \16332 , \16330 , \16331 );
nor \U$14684 ( \16333 , \14550 , \14582 );
nor \U$14685 ( \16334 , \14603 , \14619 );
nand \U$14686 ( \16335 , \16333 , \16334 );
nor \U$14687 ( \16336 , \16332 , \16335 );
nand \U$14688 ( \16337 , \16329 , \16336 );
nor \U$14689 ( \16338 , \15034 , \14738 );
nor \U$14690 ( \16339 , \14783 , \14835 );
nand \U$14691 ( \16340 , \16338 , \16339 );
nor \U$14692 ( \16341 , \14890 , \14929 );
nor \U$14693 ( \16342 , \14950 , \14966 );
nand \U$14694 ( \16343 , \16341 , \16342 );
nor \U$14695 ( \16344 , \16340 , \16343 );
nor \U$14696 ( \16345 , \15054 , \15009 );
nor \U$14697 ( \16346 , \15020 , \15031 );
nand \U$14698 ( \16347 , \16345 , \16346 );
nor \U$14699 ( \16348 , \15059 , \15051 );
not \U$14700 ( \16349 , \15067 );
and \U$14701 ( \16350 , \16348 , \16349 );
or \U$14702 ( \16351 , \15051 , \15069 );
nand \U$14703 ( \16352 , \16351 , \15072 );
nor \U$14704 ( \16353 , \16350 , \16352 );
or \U$14705 ( \16354 , \16347 , \16353 );
or \U$14706 ( \16355 , \15009 , \15074 );
nand \U$14707 ( \16356 , \16355 , \15078 );
and \U$14708 ( \16357 , \16346 , \16356 );
or \U$14709 ( \16358 , \15031 , \15080 );
nand \U$14710 ( \16359 , \16358 , \15083 );
nor \U$14711 ( \16360 , \16357 , \16359 );
nand \U$14712 ( \16361 , \16354 , \16360 );
and \U$14713 ( \16362 , \16344 , \16361 );
or \U$14714 ( \16363 , \14738 , \15085 );
nand \U$14715 ( \16364 , \16363 , \15090 );
and \U$14716 ( \16365 , \16339 , \16364 );
or \U$14717 ( \16366 , \14835 , \15092 );
nand \U$14718 ( \16367 , \16366 , \15095 );
nor \U$14719 ( \16368 , \16365 , \16367 );
or \U$14720 ( \16369 , \16343 , \16368 );
or \U$14721 ( \16370 , \14929 , \15097 );
nand \U$14722 ( \16371 , \16370 , \15101 );
and \U$14723 ( \16372 , \16342 , \16371 );
or \U$14724 ( \16373 , \14966 , \15103 );
nand \U$14725 ( \16374 , \16373 , \15106 );
nor \U$14726 ( \16375 , \16372 , \16374 );
nand \U$14727 ( \16376 , \16369 , \16375 );
nor \U$14728 ( \16377 , \16362 , \16376 );
or \U$14729 ( \16378 , \16337 , \16377 );
or \U$14730 ( \16379 , \13809 , \15108 );
nand \U$14731 ( \16380 , \16379 , \15114 );
and \U$14732 ( \16381 , \16324 , \16380 );
or \U$14733 ( \16382 , \13961 , \15116 );
nand \U$14734 ( \16383 , \16382 , \15119 );
nor \U$14735 ( \16384 , \16381 , \16383 );
or \U$14736 ( \16385 , \16328 , \16384 );
or \U$14737 ( \16386 , \14113 , \15121 );
nand \U$14738 ( \16387 , \16386 , \15125 );
and \U$14739 ( \16388 , \16327 , \16387 );
or \U$14740 ( \16389 , \14262 , \15127 );
nand \U$14741 ( \16390 , \16389 , \15130 );
nor \U$14742 ( \16391 , \16388 , \16390 );
nand \U$14743 ( \16392 , \16385 , \16391 );
and \U$14744 ( \16393 , \16336 , \16392 );
or \U$14745 ( \16394 , \14395 , \15132 );
nand \U$14746 ( \16395 , \16394 , \15137 );
and \U$14747 ( \16396 , \16331 , \16395 );
or \U$14748 ( \16397 , \14512 , \15139 );
nand \U$14749 ( \16398 , \16397 , \15142 );
nor \U$14750 ( \16399 , \16396 , \16398 );
or \U$14751 ( \16400 , \16335 , \16399 );
or \U$14752 ( \16401 , \14582 , \15144 );
nand \U$14753 ( \16402 , \16401 , \15148 );
and \U$14754 ( \16403 , \16334 , \16402 );
or \U$14755 ( \16404 , \14619 , \15150 );
nand \U$14756 ( \16405 , \16404 , \15153 );
nor \U$14757 ( \16406 , \16403 , \16405 );
nand \U$14758 ( \16407 , \16400 , \16406 );
nor \U$14759 ( \16408 , \16393 , \16407 );
nand \U$14760 ( \16409 , \16378 , \16408 );
not \U$14761 ( \16410 , \16409 );
xor \U$14762 ( \16411 , \16322 , \16410 );
buf \U$14763 ( \16412 , \16411 );
_HMUX r49ce ( \16413_nR49ce , \16320 , \16412 , \16226 );
buf \U$14764 ( \16414 , \16413_nR49ce );
not \U$14765 ( \16415 , \11825 );
nand \U$14766 ( \16416 , \12359 , \16415 );
nand \U$14767 ( \16417 , \12180 , \11091 );
nand \U$14768 ( \16418 , \11243 , \11396 );
nor \U$14769 ( \16419 , \16417 , \16418 );
nand \U$14770 ( \16420 , \11538 , \11662 );
nand \U$14771 ( \16421 , \11757 , \11810 );
nor \U$14772 ( \16422 , \16420 , \16421 );
nand \U$14773 ( \16423 , \16419 , \16422 );
nand \U$14774 ( \16424 , \12241 , \11990 );
nand \U$14775 ( \16425 , \12097 , \12157 );
nor \U$14776 ( \16426 , \16424 , \16425 );
nand \U$14777 ( \16427 , \12261 , \12227 );
not \U$14778 ( \16428 , \12276 );
or \U$14779 ( \16429 , \16427 , \16428 );
and \U$14780 ( \16430 , \12227 , \12281 );
nor \U$14781 ( \16431 , \16430 , \12287 );
nand \U$14782 ( \16432 , \16429 , \16431 );
and \U$14783 ( \16433 , \16426 , \16432 );
and \U$14784 ( \16434 , \11990 , \12292 );
nor \U$14785 ( \16435 , \16434 , \12299 );
or \U$14786 ( \16436 , \16425 , \16435 );
and \U$14787 ( \16437 , \12157 , \12304 );
nor \U$14788 ( \16438 , \16437 , \12310 );
nand \U$14789 ( \16439 , \16436 , \16438 );
nor \U$14790 ( \16440 , \16433 , \16439 );
or \U$14791 ( \16441 , \16423 , \16440 );
and \U$14792 ( \16442 , \11091 , \12315 );
nor \U$14793 ( \16443 , \16442 , \12323 );
or \U$14794 ( \16444 , \16418 , \16443 );
and \U$14795 ( \16445 , \11396 , \12328 );
nor \U$14796 ( \16446 , \16445 , \12334 );
nand \U$14797 ( \16447 , \16444 , \16446 );
and \U$14798 ( \16448 , \16422 , \16447 );
and \U$14799 ( \16449 , \11662 , \12339 );
nor \U$14800 ( \16450 , \16449 , \12346 );
or \U$14801 ( \16451 , \16421 , \16450 );
and \U$14802 ( \16452 , \11810 , \12351 );
nor \U$14803 ( \16453 , \16452 , \12357 );
nand \U$14804 ( \16454 , \16451 , \16453 );
nor \U$14805 ( \16455 , \16448 , \16454 );
nand \U$14806 ( \16456 , \16441 , \16455 );
not \U$14807 ( \16457 , \16456 );
xor \U$14808 ( \16458 , \16416 , \16457 );
buf \U$14809 ( \16459 , \16458 );
not \U$14810 ( \16460 , \14619 );
nand \U$14811 ( \16461 , \15153 , \16460 );
nand \U$14812 ( \16462 , \14974 , \13885 );
nand \U$14813 ( \16463 , \14037 , \14190 );
nor \U$14814 ( \16464 , \16462 , \16463 );
nand \U$14815 ( \16465 , \14332 , \14456 );
nand \U$14816 ( \16466 , \14551 , \14604 );
nor \U$14817 ( \16467 , \16465 , \16466 );
nand \U$14818 ( \16468 , \16464 , \16467 );
nand \U$14819 ( \16469 , \15035 , \14784 );
nand \U$14820 ( \16470 , \14891 , \14951 );
nor \U$14821 ( \16471 , \16469 , \16470 );
nand \U$14822 ( \16472 , \15055 , \15021 );
not \U$14823 ( \16473 , \15070 );
or \U$14824 ( \16474 , \16472 , \16473 );
and \U$14825 ( \16475 , \15021 , \15075 );
nor \U$14826 ( \16476 , \16475 , \15081 );
nand \U$14827 ( \16477 , \16474 , \16476 );
and \U$14828 ( \16478 , \16471 , \16477 );
and \U$14829 ( \16479 , \14784 , \15086 );
nor \U$14830 ( \16480 , \16479 , \15093 );
or \U$14831 ( \16481 , \16470 , \16480 );
and \U$14832 ( \16482 , \14951 , \15098 );
nor \U$14833 ( \16483 , \16482 , \15104 );
nand \U$14834 ( \16484 , \16481 , \16483 );
nor \U$14835 ( \16485 , \16478 , \16484 );
or \U$14836 ( \16486 , \16468 , \16485 );
and \U$14837 ( \16487 , \13885 , \15109 );
nor \U$14838 ( \16488 , \16487 , \15117 );
or \U$14839 ( \16489 , \16463 , \16488 );
and \U$14840 ( \16490 , \14190 , \15122 );
nor \U$14841 ( \16491 , \16490 , \15128 );
nand \U$14842 ( \16492 , \16489 , \16491 );
and \U$14843 ( \16493 , \16467 , \16492 );
and \U$14844 ( \16494 , \14456 , \15133 );
nor \U$14845 ( \16495 , \16494 , \15140 );
or \U$14846 ( \16496 , \16466 , \16495 );
and \U$14847 ( \16497 , \14604 , \15145 );
nor \U$14848 ( \16498 , \16497 , \15151 );
nand \U$14849 ( \16499 , \16496 , \16498 );
nor \U$14850 ( \16500 , \16493 , \16499 );
nand \U$14851 ( \16501 , \16486 , \16500 );
not \U$14852 ( \16502 , \16501 );
xor \U$14853 ( \16503 , \16461 , \16502 );
buf \U$14854 ( \16504 , \16503 );
_HMUX r4965 ( \16505_nR4965 , \16459 , \16504 , \16226 );
buf \U$14855 ( \16506 , \16505_nR4965 );
not \U$14856 ( \16507 , \11809 );
nand \U$14857 ( \16508 , \12356 , \16507 );
nand \U$14858 ( \16509 , \16250 , \16231 );
nand \U$14859 ( \16510 , \16232 , \16234 );
nor \U$14860 ( \16511 , \16509 , \16510 );
nand \U$14861 ( \16512 , \16235 , \16238 );
nand \U$14862 ( \16513 , \16239 , \16241 );
nor \U$14863 ( \16514 , \16512 , \16513 );
nand \U$14864 ( \16515 , \16511 , \16514 );
nand \U$14865 ( \16516 , \16254 , \16246 );
nand \U$14866 ( \16517 , \16247 , \16249 );
nor \U$14867 ( \16518 , \16516 , \16517 );
nand \U$14868 ( \16519 , \16256 , \16253 );
or \U$14869 ( \16520 , \16519 , \12273 );
and \U$14870 ( \16521 , \16253 , \16260 );
nor \U$14871 ( \16522 , \16521 , \16264 );
nand \U$14872 ( \16523 , \16520 , \16522 );
and \U$14873 ( \16524 , \16518 , \16523 );
and \U$14874 ( \16525 , \16246 , \16267 );
nor \U$14875 ( \16526 , \16525 , \16272 );
or \U$14876 ( \16527 , \16517 , \16526 );
and \U$14877 ( \16528 , \16249 , \16275 );
nor \U$14878 ( \16529 , \16528 , \16279 );
nand \U$14879 ( \16530 , \16527 , \16529 );
nor \U$14880 ( \16531 , \16524 , \16530 );
or \U$14881 ( \16532 , \16515 , \16531 );
and \U$14882 ( \16533 , \16231 , \16282 );
nor \U$14883 ( \16534 , \16533 , \16288 );
or \U$14884 ( \16535 , \16510 , \16534 );
and \U$14885 ( \16536 , \16234 , \16291 );
nor \U$14886 ( \16537 , \16536 , \16295 );
nand \U$14887 ( \16538 , \16535 , \16537 );
and \U$14888 ( \16539 , \16514 , \16538 );
and \U$14889 ( \16540 , \16238 , \16298 );
nor \U$14890 ( \16541 , \16540 , \16303 );
or \U$14891 ( \16542 , \16513 , \16541 );
and \U$14892 ( \16543 , \16241 , \16306 );
nor \U$14893 ( \16544 , \16543 , \16310 );
nand \U$14894 ( \16545 , \16542 , \16544 );
nor \U$14895 ( \16546 , \16539 , \16545 );
nand \U$14896 ( \16547 , \16532 , \16546 );
not \U$14897 ( \16548 , \16547 );
xor \U$14898 ( \16549 , \16508 , \16548 );
buf \U$14899 ( \16550 , \16549 );
not \U$14900 ( \16551 , \14603 );
nand \U$14901 ( \16552 , \15150 , \16551 );
nand \U$14902 ( \16553 , \16342 , \16323 );
nand \U$14903 ( \16554 , \16324 , \16326 );
nor \U$14904 ( \16555 , \16553 , \16554 );
nand \U$14905 ( \16556 , \16327 , \16330 );
nand \U$14906 ( \16557 , \16331 , \16333 );
nor \U$14907 ( \16558 , \16556 , \16557 );
nand \U$14908 ( \16559 , \16555 , \16558 );
nand \U$14909 ( \16560 , \16346 , \16338 );
nand \U$14910 ( \16561 , \16339 , \16341 );
nor \U$14911 ( \16562 , \16560 , \16561 );
nand \U$14912 ( \16563 , \16348 , \16345 );
or \U$14913 ( \16564 , \16563 , \15067 );
and \U$14914 ( \16565 , \16345 , \16352 );
nor \U$14915 ( \16566 , \16565 , \16356 );
nand \U$14916 ( \16567 , \16564 , \16566 );
and \U$14917 ( \16568 , \16562 , \16567 );
and \U$14918 ( \16569 , \16338 , \16359 );
nor \U$14919 ( \16570 , \16569 , \16364 );
or \U$14920 ( \16571 , \16561 , \16570 );
and \U$14921 ( \16572 , \16341 , \16367 );
nor \U$14922 ( \16573 , \16572 , \16371 );
nand \U$14923 ( \16574 , \16571 , \16573 );
nor \U$14924 ( \16575 , \16568 , \16574 );
or \U$14925 ( \16576 , \16559 , \16575 );
and \U$14926 ( \16577 , \16323 , \16374 );
nor \U$14927 ( \16578 , \16577 , \16380 );
or \U$14928 ( \16579 , \16554 , \16578 );
and \U$14929 ( \16580 , \16326 , \16383 );
nor \U$14930 ( \16581 , \16580 , \16387 );
nand \U$14931 ( \16582 , \16579 , \16581 );
and \U$14932 ( \16583 , \16558 , \16582 );
and \U$14933 ( \16584 , \16330 , \16390 );
nor \U$14934 ( \16585 , \16584 , \16395 );
or \U$14935 ( \16586 , \16557 , \16585 );
and \U$14936 ( \16587 , \16333 , \16398 );
nor \U$14937 ( \16588 , \16587 , \16402 );
nand \U$14938 ( \16589 , \16586 , \16588 );
nor \U$14939 ( \16590 , \16583 , \16589 );
nand \U$14940 ( \16591 , \16576 , \16590 );
not \U$14941 ( \16592 , \16591 );
xor \U$14942 ( \16593 , \16552 , \16592 );
buf \U$14943 ( \16594 , \16593 );
_HMUX r48f0 ( \16595_nR48f0 , \16550 , \16594 , \16226 );
buf \U$14944 ( \16596 , \16595_nR48f0 );
not \U$14945 ( \16597 , \11788 );
nand \U$14946 ( \16598 , \12354 , \16597 );
nor \U$14947 ( \16599 , \12181 , \11244 );
nor \U$14948 ( \16600 , \11539 , \11758 );
nand \U$14949 ( \16601 , \16599 , \16600 );
nor \U$14950 ( \16602 , \12242 , \12098 );
not \U$14951 ( \16603 , \12282 );
and \U$14952 ( \16604 , \16602 , \16603 );
or \U$14953 ( \16605 , \12098 , \12293 );
nand \U$14954 ( \16606 , \16605 , \12305 );
nor \U$14955 ( \16607 , \16604 , \16606 );
or \U$14956 ( \16608 , \16601 , \16607 );
or \U$14957 ( \16609 , \11244 , \12316 );
nand \U$14958 ( \16610 , \16609 , \12329 );
and \U$14959 ( \16611 , \16600 , \16610 );
or \U$14960 ( \16612 , \11758 , \12340 );
nand \U$14961 ( \16613 , \16612 , \12352 );
nor \U$14962 ( \16614 , \16611 , \16613 );
nand \U$14963 ( \16615 , \16608 , \16614 );
not \U$14964 ( \16616 , \16615 );
xor \U$14965 ( \16617 , \16598 , \16616 );
buf \U$14966 ( \16618 , \16617 );
not \U$14967 ( \16619 , \14582 );
nand \U$14968 ( \16620 , \15148 , \16619 );
nor \U$14969 ( \16621 , \14975 , \14038 );
nor \U$14970 ( \16622 , \14333 , \14552 );
nand \U$14971 ( \16623 , \16621 , \16622 );
nor \U$14972 ( \16624 , \15036 , \14892 );
not \U$14973 ( \16625 , \15076 );
and \U$14974 ( \16626 , \16624 , \16625 );
or \U$14975 ( \16627 , \14892 , \15087 );
nand \U$14976 ( \16628 , \16627 , \15099 );
nor \U$14977 ( \16629 , \16626 , \16628 );
or \U$14978 ( \16630 , \16623 , \16629 );
or \U$14979 ( \16631 , \14038 , \15110 );
nand \U$14980 ( \16632 , \16631 , \15123 );
and \U$14981 ( \16633 , \16622 , \16632 );
or \U$14982 ( \16634 , \14552 , \15134 );
nand \U$14983 ( \16635 , \16634 , \15146 );
nor \U$14984 ( \16636 , \16633 , \16635 );
nand \U$14985 ( \16637 , \16630 , \16636 );
not \U$14986 ( \16638 , \16637 );
xor \U$14987 ( \16639 , \16620 , \16638 );
buf \U$14988 ( \16640 , \16639 );
_HMUX r486b ( \16641_nR486b , \16618 , \16640 , \16226 );
buf \U$14989 ( \16642 , \16641_nR486b );
not \U$14990 ( \16643 , \11756 );
nand \U$14991 ( \16644 , \12350 , \16643 );
nor \U$14992 ( \16645 , \16251 , \16233 );
nor \U$14993 ( \16646 , \16236 , \16240 );
nand \U$14994 ( \16647 , \16645 , \16646 );
nor \U$14995 ( \16648 , \16255 , \16248 );
not \U$14996 ( \16649 , \16261 );
and \U$14997 ( \16650 , \16648 , \16649 );
or \U$14998 ( \16651 , \16248 , \16268 );
nand \U$14999 ( \16652 , \16651 , \16276 );
nor \U$15000 ( \16653 , \16650 , \16652 );
or \U$15001 ( \16654 , \16647 , \16653 );
or \U$15002 ( \16655 , \16233 , \16283 );
nand \U$15003 ( \16656 , \16655 , \16292 );
and \U$15004 ( \16657 , \16646 , \16656 );
or \U$15005 ( \16658 , \16240 , \16299 );
nand \U$15006 ( \16659 , \16658 , \16307 );
nor \U$15007 ( \16660 , \16657 , \16659 );
nand \U$15008 ( \16661 , \16654 , \16660 );
not \U$15009 ( \16662 , \16661 );
xor \U$15010 ( \16663 , \16644 , \16662 );
buf \U$15011 ( \16664 , \16663 );
not \U$15012 ( \16665 , \14550 );
nand \U$15013 ( \16666 , \15144 , \16665 );
nor \U$15014 ( \16667 , \16343 , \16325 );
nor \U$15015 ( \16668 , \16328 , \16332 );
nand \U$15016 ( \16669 , \16667 , \16668 );
nor \U$15017 ( \16670 , \16347 , \16340 );
not \U$15018 ( \16671 , \16353 );
and \U$15019 ( \16672 , \16670 , \16671 );
or \U$15020 ( \16673 , \16340 , \16360 );
nand \U$15021 ( \16674 , \16673 , \16368 );
nor \U$15022 ( \16675 , \16672 , \16674 );
or \U$15023 ( \16676 , \16669 , \16675 );
or \U$15024 ( \16677 , \16325 , \16375 );
nand \U$15025 ( \16678 , \16677 , \16384 );
and \U$15026 ( \16679 , \16668 , \16678 );
or \U$15027 ( \16680 , \16332 , \16391 );
nand \U$15028 ( \16681 , \16680 , \16399 );
nor \U$15029 ( \16682 , \16679 , \16681 );
nand \U$15030 ( \16683 , \16676 , \16682 );
not \U$15031 ( \16684 , \16683 );
xor \U$15032 ( \16685 , \16666 , \16684 );
buf \U$15033 ( \16686 , \16685 );
_HMUX r47de ( \16687_nR47de , \16664 , \16686 , \16226 );
buf \U$15034 ( \16688 , \16687_nR47de );
not \U$15035 ( \16689 , \11718 );
nand \U$15036 ( \16690 , \12348 , \16689 );
nor \U$15037 ( \16691 , \16425 , \16417 );
nor \U$15038 ( \16692 , \16418 , \16420 );
nand \U$15039 ( \16693 , \16691 , \16692 );
nor \U$15040 ( \16694 , \16427 , \16424 );
and \U$15041 ( \16695 , \16694 , \12276 );
or \U$15042 ( \16696 , \16424 , \16431 );
nand \U$15043 ( \16697 , \16696 , \16435 );
nor \U$15044 ( \16698 , \16695 , \16697 );
or \U$15045 ( \16699 , \16693 , \16698 );
or \U$15046 ( \16700 , \16417 , \16438 );
nand \U$15047 ( \16701 , \16700 , \16443 );
and \U$15048 ( \16702 , \16692 , \16701 );
or \U$15049 ( \16703 , \16420 , \16446 );
nand \U$15050 ( \16704 , \16703 , \16450 );
nor \U$15051 ( \16705 , \16702 , \16704 );
nand \U$15052 ( \16706 , \16699 , \16705 );
not \U$15053 ( \16707 , \16706 );
xor \U$15054 ( \16708 , \16690 , \16707 );
buf \U$15055 ( \16709 , \16708 );
not \U$15056 ( \16710 , \14512 );
nand \U$15057 ( \16711 , \15142 , \16710 );
nor \U$15058 ( \16712 , \16470 , \16462 );
nor \U$15059 ( \16713 , \16463 , \16465 );
nand \U$15060 ( \16714 , \16712 , \16713 );
nor \U$15061 ( \16715 , \16472 , \16469 );
and \U$15062 ( \16716 , \16715 , \15070 );
or \U$15063 ( \16717 , \16469 , \16476 );
nand \U$15064 ( \16718 , \16717 , \16480 );
nor \U$15065 ( \16719 , \16716 , \16718 );
or \U$15066 ( \16720 , \16714 , \16719 );
or \U$15067 ( \16721 , \16462 , \16483 );
nand \U$15068 ( \16722 , \16721 , \16488 );
and \U$15069 ( \16723 , \16713 , \16722 );
or \U$15070 ( \16724 , \16465 , \16491 );
nand \U$15071 ( \16725 , \16724 , \16495 );
nor \U$15072 ( \16726 , \16723 , \16725 );
nand \U$15073 ( \16727 , \16720 , \16726 );
not \U$15074 ( \16728 , \16727 );
xor \U$15075 ( \16729 , \16711 , \16728 );
buf \U$15076 ( \16730 , \16729 );
_HMUX r474d ( \16731_nR474d , \16709 , \16730 , \16226 );
buf \U$15077 ( \16732 , \16731_nR474d );
not \U$15078 ( \16733 , \11661 );
nand \U$15079 ( \16734 , \12345 , \16733 );
nor \U$15080 ( \16735 , \16517 , \16509 );
nor \U$15081 ( \16736 , \16510 , \16512 );
nand \U$15082 ( \16737 , \16735 , \16736 );
nor \U$15083 ( \16738 , \16519 , \16516 );
and \U$15084 ( \16739 , \16738 , \16257 );
or \U$15085 ( \16740 , \16516 , \16522 );
nand \U$15086 ( \16741 , \16740 , \16526 );
nor \U$15087 ( \16742 , \16739 , \16741 );
or \U$15088 ( \16743 , \16737 , \16742 );
or \U$15089 ( \16744 , \16509 , \16529 );
nand \U$15090 ( \16745 , \16744 , \16534 );
and \U$15091 ( \16746 , \16736 , \16745 );
or \U$15092 ( \16747 , \16512 , \16537 );
nand \U$15093 ( \16748 , \16747 , \16541 );
nor \U$15094 ( \16749 , \16746 , \16748 );
nand \U$15095 ( \16750 , \16743 , \16749 );
not \U$15096 ( \16751 , \16750 );
xor \U$15097 ( \16752 , \16734 , \16751 );
buf \U$15098 ( \16753 , \16752 );
not \U$15099 ( \16754 , \14455 );
nand \U$15100 ( \16755 , \15139 , \16754 );
nor \U$15101 ( \16756 , \16561 , \16553 );
nor \U$15102 ( \16757 , \16554 , \16556 );
nand \U$15103 ( \16758 , \16756 , \16757 );
nor \U$15104 ( \16759 , \16563 , \16560 );
and \U$15105 ( \16760 , \16759 , \16349 );
or \U$15106 ( \16761 , \16560 , \16566 );
nand \U$15107 ( \16762 , \16761 , \16570 );
nor \U$15108 ( \16763 , \16760 , \16762 );
or \U$15109 ( \16764 , \16758 , \16763 );
or \U$15110 ( \16765 , \16553 , \16573 );
nand \U$15111 ( \16766 , \16765 , \16578 );
and \U$15112 ( \16767 , \16757 , \16766 );
or \U$15113 ( \16768 , \16556 , \16581 );
nand \U$15114 ( \16769 , \16768 , \16585 );
nor \U$15115 ( \16770 , \16767 , \16769 );
nand \U$15116 ( \16771 , \16764 , \16770 );
not \U$15117 ( \16772 , \16771 );
xor \U$15118 ( \16773 , \16755 , \16772 );
buf \U$15119 ( \16774 , \16773 );
_HMUX r46b4 ( \16775_nR46b4 , \16753 , \16774 , \16226 );
buf \U$15120 ( \16776 , \16775_nR46b4 );
not \U$15121 ( \16777 , \11601 );
nand \U$15122 ( \16778 , \12343 , \16777 );
nand \U$15123 ( \16779 , \12182 , \11540 );
not \U$15124 ( \16780 , \12294 );
or \U$15125 ( \16781 , \16779 , \16780 );
and \U$15126 ( \16782 , \11540 , \12317 );
nor \U$15127 ( \16783 , \16782 , \12341 );
nand \U$15128 ( \16784 , \16781 , \16783 );
not \U$15129 ( \16785 , \16784 );
xor \U$15130 ( \16786 , \16778 , \16785 );
buf \U$15131 ( \16787 , \16786 );
not \U$15132 ( \16788 , \14395 );
nand \U$15133 ( \16789 , \15137 , \16788 );
nand \U$15134 ( \16790 , \14976 , \14334 );
not \U$15135 ( \16791 , \15088 );
or \U$15136 ( \16792 , \16790 , \16791 );
and \U$15137 ( \16793 , \14334 , \15111 );
nor \U$15138 ( \16794 , \16793 , \15135 );
nand \U$15139 ( \16795 , \16792 , \16794 );
not \U$15140 ( \16796 , \16795 );
xor \U$15141 ( \16797 , \16789 , \16796 );
buf \U$15142 ( \16798 , \16797 );
_HMUX r4613 ( \16799_nR4613 , \16787 , \16798 , \16226 );
buf \U$15143 ( \16800 , \16799_nR4613 );
not \U$15144 ( \16801 , \11537 );
nand \U$15145 ( \16802 , \12338 , \16801 );
nand \U$15146 ( \16803 , \16252 , \16237 );
not \U$15147 ( \16804 , \16269 );
or \U$15148 ( \16805 , \16803 , \16804 );
and \U$15149 ( \16806 , \16237 , \16284 );
nor \U$15150 ( \16807 , \16806 , \16300 );
nand \U$15151 ( \16808 , \16805 , \16807 );
not \U$15152 ( \16809 , \16808 );
xor \U$15153 ( \16810 , \16802 , \16809 );
buf \U$15154 ( \16811 , \16810 );
not \U$15155 ( \16812 , \14331 );
nand \U$15156 ( \16813 , \15132 , \16812 );
nand \U$15157 ( \16814 , \16344 , \16329 );
not \U$15158 ( \16815 , \16361 );
or \U$15159 ( \16816 , \16814 , \16815 );
and \U$15160 ( \16817 , \16329 , \16376 );
nor \U$15161 ( \16818 , \16817 , \16392 );
nand \U$15162 ( \16819 , \16816 , \16818 );
not \U$15163 ( \16820 , \16819 );
xor \U$15164 ( \16821 , \16813 , \16820 );
buf \U$15165 ( \16822 , \16821 );
_HMUX r4570 ( \16823_nR4570 , \16811 , \16822 , \16226 );
buf \U$15166 ( \16824 , \16823_nR4570 );
not \U$15167 ( \16825 , \11468 );
nand \U$15168 ( \16826 , \12336 , \16825 );
nand \U$15169 ( \16827 , \16426 , \16419 );
not \U$15170 ( \16828 , \16432 );
or \U$15171 ( \16829 , \16827 , \16828 );
and \U$15172 ( \16830 , \16419 , \16439 );
nor \U$15173 ( \16831 , \16830 , \16447 );
nand \U$15174 ( \16832 , \16829 , \16831 );
not \U$15175 ( \16833 , \16832 );
xor \U$15176 ( \16834 , \16826 , \16833 );
buf \U$15177 ( \16835 , \16834 );
not \U$15178 ( \16836 , \14262 );
nand \U$15179 ( \16837 , \15130 , \16836 );
nand \U$15180 ( \16838 , \16471 , \16464 );
not \U$15181 ( \16839 , \16477 );
or \U$15182 ( \16840 , \16838 , \16839 );
and \U$15183 ( \16841 , \16464 , \16484 );
nor \U$15184 ( \16842 , \16841 , \16492 );
nand \U$15185 ( \16843 , \16840 , \16842 );
not \U$15186 ( \16844 , \16843 );
xor \U$15187 ( \16845 , \16837 , \16844 );
buf \U$15188 ( \16846 , \16845 );
_HMUX r44bd ( \16847_nR44bd , \16835 , \16846 , \16226 );
buf \U$15189 ( \16848 , \16847_nR44bd );
not \U$15190 ( \16849 , \11395 );
nand \U$15191 ( \16850 , \12333 , \16849 );
nand \U$15192 ( \16851 , \16518 , \16511 );
not \U$15193 ( \16852 , \16523 );
or \U$15194 ( \16853 , \16851 , \16852 );
and \U$15195 ( \16854 , \16511 , \16530 );
nor \U$15196 ( \16855 , \16854 , \16538 );
nand \U$15197 ( \16856 , \16853 , \16855 );
not \U$15198 ( \16857 , \16856 );
xor \U$15199 ( \16858 , \16850 , \16857 );
buf \U$15200 ( \16859 , \16858 );
not \U$15201 ( \16860 , \14189 );
nand \U$15202 ( \16861 , \15127 , \16860 );
nand \U$15203 ( \16862 , \16562 , \16555 );
not \U$15204 ( \16863 , \16567 );
or \U$15205 ( \16864 , \16862 , \16863 );
and \U$15206 ( \16865 , \16555 , \16574 );
nor \U$15207 ( \16866 , \16865 , \16582 );
nand \U$15208 ( \16867 , \16864 , \16866 );
not \U$15209 ( \16868 , \16867 );
xor \U$15210 ( \16869 , \16861 , \16868 );
buf \U$15211 ( \16870 , \16869 );
_HMUX r4404 ( \16871_nR4404 , \16859 , \16870 , \16226 );
buf \U$15212 ( \16872 , \16871_nR4404 );
not \U$15213 ( \16873 , \11319 );
nand \U$15214 ( \16874 , \12331 , \16873 );
nand \U$15215 ( \16875 , \16602 , \16599 );
or \U$15216 ( \16876 , \16875 , \12282 );
and \U$15217 ( \16877 , \16599 , \16606 );
nor \U$15218 ( \16878 , \16877 , \16610 );
nand \U$15219 ( \16879 , \16876 , \16878 );
not \U$15220 ( \16880 , \16879 );
xor \U$15221 ( \16881 , \16874 , \16880 );
buf \U$15222 ( \16882 , \16881 );
not \U$15223 ( \16883 , \14113 );
nand \U$15224 ( \16884 , \15125 , \16883 );
nand \U$15225 ( \16885 , \16624 , \16621 );
or \U$15226 ( \16886 , \16885 , \15076 );
and \U$15227 ( \16887 , \16621 , \16628 );
nor \U$15228 ( \16888 , \16887 , \16632 );
nand \U$15229 ( \16889 , \16886 , \16888 );
not \U$15230 ( \16890 , \16889 );
xor \U$15231 ( \16891 , \16884 , \16890 );
buf \U$15232 ( \16892 , \16891 );
_HMUX r4343 ( \16893_nR4343 , \16882 , \16892 , \16226 );
buf \U$15233 ( \16894 , \16893_nR4343 );
not \U$15234 ( \16895 , \11242 );
nand \U$15235 ( \16896 , \12327 , \16895 );
nand \U$15236 ( \16897 , \16648 , \16645 );
or \U$15237 ( \16898 , \16897 , \16261 );
and \U$15238 ( \16899 , \16645 , \16652 );
nor \U$15239 ( \16900 , \16899 , \16656 );
nand \U$15240 ( \16901 , \16898 , \16900 );
not \U$15241 ( \16902 , \16901 );
xor \U$15242 ( \16903 , \16896 , \16902 );
buf \U$15243 ( \16904 , \16903 );
not \U$15244 ( \16905 , \14036 );
nand \U$15245 ( \16906 , \15121 , \16905 );
nand \U$15246 ( \16907 , \16670 , \16667 );
or \U$15247 ( \16908 , \16907 , \16353 );
and \U$15248 ( \16909 , \16667 , \16674 );
nor \U$15249 ( \16910 , \16909 , \16678 );
nand \U$15250 ( \16911 , \16908 , \16910 );
not \U$15251 ( \16912 , \16911 );
xor \U$15252 ( \16913 , \16906 , \16912 );
buf \U$15253 ( \16914 , \16913 );
_HMUX r4284 ( \16915_nR4284 , \16904 , \16914 , \16226 );
buf \U$15254 ( \16916 , \16915_nR4284 );
not \U$15255 ( \16917 , \11167 );
nand \U$15256 ( \16918 , \12325 , \16917 );
nand \U$15257 ( \16919 , \16694 , \16691 );
or \U$15258 ( \16920 , \16919 , \16428 );
and \U$15259 ( \16921 , \16691 , \16697 );
nor \U$15260 ( \16922 , \16921 , \16701 );
nand \U$15261 ( \16923 , \16920 , \16922 );
not \U$15262 ( \16924 , \16923 );
xor \U$15263 ( \16925 , \16918 , \16924 );
buf \U$15264 ( \16926 , \16925 );
not \U$15265 ( \16927 , \13961 );
nand \U$15266 ( \16928 , \15119 , \16927 );
nand \U$15267 ( \16929 , \16715 , \16712 );
or \U$15268 ( \16930 , \16929 , \16473 );
and \U$15269 ( \16931 , \16712 , \16718 );
nor \U$15270 ( \16932 , \16931 , \16722 );
nand \U$15271 ( \16933 , \16930 , \16932 );
not \U$15272 ( \16934 , \16933 );
xor \U$15273 ( \16935 , \16928 , \16934 );
buf \U$15274 ( \16936 , \16935 );
_HMUX r41c5 ( \16937_nR41c5 , \16926 , \16936 , \16226 );
buf \U$15275 ( \16938 , \16937_nR41c5 );
not \U$15276 ( \16939 , \11090 );
nand \U$15277 ( \16940 , \12322 , \16939 );
nand \U$15278 ( \16941 , \16738 , \16735 );
or \U$15279 ( \16942 , \16941 , \12273 );
and \U$15280 ( \16943 , \16735 , \16741 );
nor \U$15281 ( \16944 , \16943 , \16745 );
nand \U$15282 ( \16945 , \16942 , \16944 );
not \U$15283 ( \16946 , \16945 );
xor \U$15284 ( \16947 , \16940 , \16946 );
buf \U$15285 ( \16948 , \16947 );
not \U$15286 ( \16949 , \13884 );
nand \U$15287 ( \16950 , \15116 , \16949 );
nand \U$15288 ( \16951 , \16759 , \16756 );
or \U$15289 ( \16952 , \16951 , \15067 );
and \U$15290 ( \16953 , \16756 , \16762 );
nor \U$15291 ( \16954 , \16953 , \16766 );
nand \U$15292 ( \16955 , \16952 , \16954 );
not \U$15293 ( \16956 , \16955 );
xor \U$15294 ( \16957 , \16950 , \16956 );
buf \U$15295 ( \16958 , \16957 );
_HMUX r40dc ( \16959_nR40dc , \16948 , \16958 , \16226 );
buf \U$15296 ( \16960 , \16959_nR40dc );
not \U$15297 ( \16961 , \11015 );
nand \U$15298 ( \16962 , \12320 , \16961 );
xor \U$15299 ( \16963 , \16962 , \12318 );
buf \U$15300 ( \16964 , \16963 );
not \U$15301 ( \16965 , \13809 );
nand \U$15302 ( \16966 , \15114 , \16965 );
xor \U$15303 ( \16967 , \16966 , \15112 );
buf \U$15304 ( \16968 , \16967 );
_HMUX r3ff5 ( \16969_nR3ff5 , \16964 , \16968 , \16226 );
buf \U$15305 ( \16970 , \16969_nR3ff5 );
not \U$15306 ( \16971 , \12179 );
nand \U$15307 ( \16972 , \12314 , \16971 );
xor \U$15308 ( \16973 , \16972 , \16285 );
buf \U$15309 ( \16974 , \16973 );
not \U$15310 ( \16975 , \14973 );
nand \U$15311 ( \16976 , \15108 , \16975 );
xor \U$15312 ( \16977 , \16976 , \16377 );
buf \U$15313 ( \16978 , \16977 );
_HMUX r3f1c ( \16979_nR3f1c , \16974 , \16978 , \16226 );
buf \U$15314 ( \16980 , \16979_nR3f1c );
not \U$15315 ( \16981 , \12172 );
nand \U$15316 ( \16982 , \12312 , \16981 );
xor \U$15317 ( \16983 , \16982 , \16440 );
buf \U$15318 ( \16984 , \16983 );
not \U$15319 ( \16985 , \14966 );
nand \U$15320 ( \16986 , \15106 , \16985 );
xor \U$15321 ( \16987 , \16986 , \16485 );
buf \U$15322 ( \16988 , \16987 );
_HMUX r3e43 ( \16989_nR3e43 , \16984 , \16988 , \16226 );
buf \U$15323 ( \16990 , \16989_nR3e43 );
not \U$15324 ( \16991 , \12156 );
nand \U$15325 ( \16992 , \12309 , \16991 );
xor \U$15326 ( \16993 , \16992 , \16531 );
buf \U$15327 ( \16994 , \16993 );
not \U$15328 ( \16995 , \14950 );
nand \U$15329 ( \16996 , \15103 , \16995 );
xor \U$15330 ( \16997 , \16996 , \16575 );
buf \U$15331 ( \16998 , \16997 );
_HMUX r3d72 ( \16999_nR3d72 , \16994 , \16998 , \16226 );
buf \U$15332 ( \17000 , \16999_nR3d72 );
not \U$15333 ( \17001 , \12135 );
nand \U$15334 ( \17002 , \12307 , \17001 );
xor \U$15335 ( \17003 , \17002 , \16607 );
buf \U$15336 ( \17004 , \17003 );
not \U$15337 ( \17005 , \14929 );
nand \U$15338 ( \17006 , \15101 , \17005 );
xor \U$15339 ( \17007 , \17006 , \16629 );
buf \U$15340 ( \17008 , \17007 );
_HMUX r3c9d ( \17009_nR3c9d , \17004 , \17008 , \16226 );
buf \U$15341 ( \17010 , \17009_nR3c9d );
not \U$15342 ( \17011 , \12096 );
nand \U$15343 ( \17012 , \12303 , \17011 );
xor \U$15344 ( \17013 , \17012 , \16653 );
buf \U$15345 ( \17014 , \17013 );
not \U$15346 ( \17015 , \14890 );
nand \U$15347 ( \17016 , \15097 , \17015 );
xor \U$15348 ( \17017 , \17016 , \16675 );
buf \U$15349 ( \17018 , \17017 );
_HMUX r3bd2 ( \17019_nR3bd2 , \17014 , \17018 , \16226 );
buf \U$15350 ( \17020 , \17019_nR3bd2 );
not \U$15351 ( \17021 , \12041 );
nand \U$15352 ( \17022 , \12301 , \17021 );
xor \U$15353 ( \17023 , \17022 , \16698 );
buf \U$15354 ( \17024 , \17023 );
not \U$15355 ( \17025 , \14835 );
nand \U$15356 ( \17026 , \15095 , \17025 );
xor \U$15357 ( \17027 , \17026 , \16719 );
buf \U$15358 ( \17028 , \17027 );
_HMUX r3ab9 ( \17029_nR3ab9 , \17024 , \17028 , \16226 );
buf \U$15359 ( \17030 , \17029_nR3ab9 );
not \U$15360 ( \17031 , \11989 );
nand \U$15361 ( \17032 , \12298 , \17031 );
xor \U$15362 ( \17033 , \17032 , \16742 );
buf \U$15363 ( \17034 , \17033 );
not \U$15364 ( \17035 , \14783 );
nand \U$15365 ( \17036 , \15092 , \17035 );
xor \U$15366 ( \17037 , \17036 , \16763 );
buf \U$15367 ( \17038 , \17037 );
_HMUX r3a04 ( \17039_nR3a04 , \17034 , \17038 , \16226 );
buf \U$15368 ( \17040 , \17039_nR3a04 );
not \U$15369 ( \17041 , \11944 );
nand \U$15370 ( \17042 , \12296 , \17041 );
xor \U$15371 ( \17043 , \17042 , \16780 );
buf \U$15372 ( \17044 , \17043 );
not \U$15373 ( \17045 , \14738 );
nand \U$15374 ( \17046 , \15090 , \17045 );
xor \U$15375 ( \17047 , \17046 , \16791 );
buf \U$15376 ( \17048 , \17047 );
_HMUX r38d1 ( \17049_nR38d1 , \17044 , \17048 , \16226 );
buf \U$15377 ( \17050 , \17049_nR38d1 );
not \U$15378 ( \17051 , \12240 );
nand \U$15379 ( \17052 , \12291 , \17051 );
xor \U$15380 ( \17053 , \17052 , \16804 );
buf \U$15381 ( \17054 , \17053 );
not \U$15382 ( \17055 , \15034 );
nand \U$15383 ( \17056 , \15085 , \17055 );
xor \U$15384 ( \17057 , \17056 , \16815 );
buf \U$15385 ( \17058 , \17057 );
_HMUX r3834 ( \17059_nR3834 , \17054 , \17058 , \16226 );
buf \U$15386 ( \17060 , \17059_nR3834 );
not \U$15387 ( \17061 , \12237 );
nand \U$15388 ( \17062 , \12289 , \17061 );
xor \U$15389 ( \17063 , \17062 , \16828 );
buf \U$15390 ( \17064 , \17063 );
not \U$15391 ( \17065 , \15031 );
nand \U$15392 ( \17066 , \15083 , \17065 );
xor \U$15393 ( \17067 , \17066 , \16839 );
buf \U$15394 ( \17068 , \17067 );
_HMUX r3719 ( \17069_nR3719 , \17064 , \17068 , \16226 );
buf \U$15395 ( \17070 , \17069_nR3719 );
not \U$15396 ( \17071 , \12226 );
nand \U$15397 ( \17072 , \12286 , \17071 );
xor \U$15398 ( \17073 , \17072 , \16852 );
buf \U$15399 ( \17074 , \17073 );
not \U$15400 ( \17075 , \15020 );
nand \U$15401 ( \17076 , \15080 , \17075 );
xor \U$15402 ( \17077 , \17076 , \16863 );
buf \U$15403 ( \17078 , \17077 );
_HMUX r3690 ( \17079_nR3690 , \17074 , \17078 , \16226 );
buf \U$15404 ( \17080 , \17079_nR3690 );
not \U$15405 ( \17081 , \12215 );
nand \U$15406 ( \17082 , \12284 , \17081 );
xor \U$15407 ( \17083 , \17082 , \12282 );
buf \U$15408 ( \17084 , \17083 );
not \U$15409 ( \17085 , \15009 );
nand \U$15410 ( \17086 , \15078 , \17085 );
xor \U$15411 ( \17087 , \17086 , \15076 );
buf \U$15412 ( \17088 , \17087 );
_HMUX r3589 ( \17089_nR3589 , \17084 , \17088 , \16226 );
buf \U$15413 ( \17090 , \17089_nR3589 );
not \U$15414 ( \17091 , \12260 );
nand \U$15415 ( \17092 , \12280 , \17091 );
xor \U$15416 ( \17093 , \17092 , \16261 );
buf \U$15417 ( \17094 , \17093 );
not \U$15418 ( \17095 , \15054 );
nand \U$15419 ( \17096 , \15074 , \17095 );
xor \U$15420 ( \17097 , \17096 , \16353 );
buf \U$15421 ( \17098 , \17097 );
_HMUX r351c ( \17099_nR351c , \17094 , \17098 , \16226 );
buf \U$15422 ( \17100 , \17099_nR351c );
not \U$15423 ( \17101 , \12257 );
nand \U$15424 ( \17102 , \12278 , \17101 );
xor \U$15425 ( \17103 , \17102 , \16428 );
buf \U$15426 ( \17104 , \17103 );
not \U$15427 ( \17105 , \15051 );
nand \U$15428 ( \17106 , \15072 , \17105 );
xor \U$15429 ( \17107 , \17106 , \16473 );
buf \U$15430 ( \17108 , \17107 );
_HMUX r342f ( \17109_nR342f , \17104 , \17108 , \16226 );
buf \U$15431 ( \17110 , \17109_nR342f );
not \U$15432 ( \17111 , \12265 );
nand \U$15433 ( \17112 , \12275 , \17111 );
xor \U$15434 ( \17113 , \17112 , \12273 );
buf \U$15435 ( \17114 , \17113 );
not \U$15436 ( \17115 , \15059 );
nand \U$15437 ( \17116 , \15069 , \17115 );
xor \U$15438 ( \17117 , \17116 , \15067 );
buf \U$15439 ( \17118 , \17117 );
_HMUX r33da ( \17119_nR33da , \17114 , \17118 , \16226 );
buf \U$15440 ( \17120 , \17119_nR33da );
nor \U$15441 ( \17121 , \12269 , \12272 );
not \U$15442 ( \17122 , \17121 );
nand \U$15443 ( \17123 , \12273 , \17122 );
not \U$15444 ( \17124 , \17123 );
buf \U$15445 ( \17125 , \17124 );
nor \U$15446 ( \17126 , \15063 , \15066 );
not \U$15447 ( \17127 , \17126 );
nand \U$15448 ( \17128 , \15067 , \17127 );
not \U$15449 ( \17129 , \17128 );
buf \U$15450 ( \17130 , \17129 );
_HMUX r3309 ( \17131_nR3309 , \17125 , \17130 , \16226 );
buf \U$15451 ( \17132 , \17131_nR3309 );
xor \U$15452 ( \17133 , \12271 , \10430 );
buf \U$15453 ( \17134 , \17133 );
xor \U$15454 ( \17135 , \15065 , \13224 );
buf \U$15455 ( \17136 , \17135 );
_HMUX r32c4 ( \17137_nR32c4 , \17134 , \17136 , \16226 );
buf \U$15456 ( \17138 , \17137_nR32c4 );
endmodule

